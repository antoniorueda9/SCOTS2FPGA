// Benchmark "DD" written by ABC on Sun Jun  9 18:29:03 2019

module DD ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29,
    po0  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29;
  output po0;
  wire n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
    n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
    n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
    n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
    n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
    n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
    n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
    n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
    n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
    n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
    n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
    n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
    n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
    n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
    n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
    n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
    n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
    n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
    n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
    n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
    n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
    n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
    n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
    n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
    n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
    n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
    n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
    n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
    n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
    n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
    n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
    n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
    n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
    n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
    n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
    n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
    n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
    n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
    n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
    n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
    n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
    n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
    n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
    n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
    n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
    n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
    n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
    n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
    n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
    n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
    n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
    n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
    n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
    n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
    n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
    n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
    n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
    n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
    n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
    n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
    n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
    n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
    n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
    n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
    n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
    n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
    n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
    n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
    n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
    n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
    n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
    n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
    n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
    n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
    n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
    n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
    n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
    n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
    n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
    n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
    n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
    n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
    n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
    n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
    n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
    n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
    n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
    n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
    n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
    n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
    n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
    n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
    n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
    n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
    n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
    n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
    n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
    n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
    n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
    n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
    n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
    n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
    n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
    n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
    n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
    n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
    n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
    n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
    n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
    n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
    n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
    n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
    n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
    n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
    n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
    n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
    n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
    n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
    n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
    n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
    n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
    n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
    n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
    n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
    n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
    n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
    n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
    n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
    n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
    n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
    n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
    n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
    n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
    n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
    n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
    n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
    n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
    n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
    n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
    n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
    n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
    n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
    n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
    n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
    n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
    n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
    n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
    n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
    n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
    n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
    n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
    n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
    n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
    n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
    n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
    n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
    n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
    n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
    n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
    n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
    n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
    n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
    n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
    n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
    n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
    n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
    n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
    n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
    n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
    n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
    n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
    n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
    n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
    n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
    n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
    n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
    n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
    n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
    n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
    n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
    n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
    n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
    n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
    n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
    n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
    n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
    n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
    n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
    n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
    n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
    n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
    n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
    n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
    n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
    n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
    n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
    n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
    n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
    n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
    n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
    n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
    n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
    n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
    n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
    n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
    n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
    n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
    n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
    n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
    n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
    n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
    n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
    n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
    n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
    n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
    n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
    n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
    n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
    n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
    n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
    n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
    n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
    n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
    n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
    n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
    n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
    n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
    n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
    n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
    n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
    n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
    n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
    n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
    n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
    n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
    n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
    n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
    n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
    n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
    n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
    n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
    n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
    n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
    n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
    n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
    n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
    n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
    n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
    n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
    n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
    n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
    n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
    n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
    n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
    n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
    n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
    n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
    n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
    n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
    n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
    n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
    n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
    n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
    n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
    n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
    n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
    n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
    n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
    n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
    n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
    n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
    n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
    n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
    n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
    n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
    n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
    n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
    n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
    n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
    n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
    n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
    n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
    n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
    n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
    n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
    n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
    n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
    n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
    n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
    n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
    n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
    n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
    n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
    n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
    n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
    n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
    n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
    n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
    n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
    n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
    n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
    n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
    n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
    n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
    n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
    n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
    n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
    n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
    n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
    n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
    n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
    n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
    n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
    n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
    n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
    n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
    n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
    n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
    n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
    n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
    n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
    n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
    n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
    n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
    n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
    n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
    n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
    n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
    n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
    n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
    n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
    n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
    n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
    n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
    n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
    n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
    n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
    n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
    n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
    n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
    n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
    n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
    n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
    n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
    n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
    n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
    n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
    n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
    n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
    n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
    n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
    n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
    n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
    n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
    n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
    n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
    n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
    n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
    n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
    n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
    n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
    n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
    n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
    n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
    n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
    n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
    n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
    n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
    n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
    n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
    n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
    n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
    n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
    n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
    n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
    n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
    n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
    n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
    n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
    n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
    n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
    n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
    n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
    n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
    n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
    n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
    n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
    n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
    n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
    n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
    n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
    n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
    n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
    n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
    n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
    n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
    n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
    n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
    n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
    n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
    n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
    n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
    n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
    n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
    n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
    n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
    n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
    n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
    n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
    n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
    n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
    n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
    n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
    n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
    n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
    n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
    n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
    n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
    n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
    n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
    n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
    n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
    n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
    n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
    n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
    n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
    n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
    n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
    n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
    n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
    n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
    n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
    n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
    n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
    n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
    n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
    n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
    n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
    n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
    n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
    n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
    n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
    n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
    n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
    n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
    n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
    n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
    n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
    n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
    n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
    n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
    n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
    n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
    n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
    n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
    n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
    n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
    n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
    n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
    n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
    n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
    n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
    n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
    n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
    n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
    n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
    n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
    n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
    n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
    n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
    n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
    n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
    n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
    n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
    n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
    n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
    n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
    n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
    n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
    n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
    n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
    n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
    n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
    n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
    n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
    n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
    n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
    n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
    n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
    n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
    n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
    n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
    n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
    n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
    n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
    n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
    n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
    n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
    n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
    n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
    n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
    n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
    n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
    n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
    n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
    n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
    n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
    n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
    n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
    n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
    n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
    n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
    n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
    n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
    n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
    n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
    n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
    n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
    n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
    n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
    n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
    n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
    n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
    n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
    n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
    n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
    n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
    n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
    n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
    n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
    n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
    n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
    n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
    n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
    n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
    n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
    n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
    n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
    n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
    n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
    n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
    n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
    n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
    n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
    n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
    n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
    n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
    n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
    n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
    n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
    n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
    n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
    n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
    n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
    n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
    n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
    n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
    n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
    n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
    n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
    n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
    n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
    n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
    n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
    n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
    n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
    n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
    n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
    n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
    n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
    n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
    n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
    n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
    n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
    n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
    n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
    n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
    n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
    n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
    n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
    n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
    n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
    n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
    n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
    n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
    n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
    n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
    n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
    n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
    n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
    n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
    n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
    n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
    n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
    n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
    n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
    n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
    n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
    n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
    n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
    n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
    n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
    n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
    n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
    n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
    n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
    n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
    n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
    n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
    n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
    n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
    n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
    n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
    n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
    n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
    n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
    n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
    n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
    n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
    n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
    n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
    n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
    n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
    n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
    n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
    n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
    n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
    n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
    n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
    n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
    n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
    n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
    n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
    n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
    n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
    n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
    n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
    n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
    n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
    n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
    n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
    n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
    n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
    n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
    n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
    n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
    n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
    n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
    n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
    n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
    n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
    n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
    n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
    n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
    n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
    n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
    n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
    n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
    n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
    n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
    n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
    n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
    n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
    n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
    n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
    n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
    n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
    n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
    n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
    n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
    n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
    n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
    n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
    n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
    n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
    n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
    n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
    n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
    n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
    n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
    n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
    n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
    n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
    n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
    n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
    n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
    n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
    n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
    n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
    n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
    n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
    n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
    n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
    n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
    n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
    n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
    n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
    n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429,
    n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
    n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
    n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
    n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
    n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
    n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
    n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
    n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
    n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
    n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
    n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
    n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
    n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
    n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
    n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
    n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
    n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
    n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
    n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
    n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726,
    n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
    n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
    n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
    n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798,
    n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
    n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
    n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852,
    n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870,
    n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
    n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
    n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
    n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942,
    n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
    n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
    n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
    n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
    n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
    n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014,
    n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
    n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
    n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
    n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
    n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
    n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
    n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
    n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086,
    n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
    n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
    n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
    n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
    n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
    n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
    n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
    n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
    n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
    n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
    n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212,
    n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230,
    n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
    n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
    n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
    n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
    n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
    n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
    n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
    n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
    n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
    n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
    n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
    n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
    n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
    n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
    n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
    n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
    n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
    n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
    n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
    n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
    n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
    n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
    n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
    n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
    n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
    n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
    n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
    n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
    n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716,
    n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
    n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
    n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
    n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
    n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
    n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
    n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
    n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788,
    n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
    n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
    n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
    n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
    n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
    n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
    n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
    n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
    n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
    n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
    n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
    n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
    n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
    n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
    n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932,
    n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950,
    n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
    n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
    n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
    n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
    n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
    n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
    n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
    n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
    n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
    n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
    n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
    n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
    n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
    n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
    n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
    n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
    n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
    n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
    n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
    n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
    n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
    n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
    n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
    n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238,
    n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
    n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
    n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292,
    n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310,
    n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
    n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
    n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
    n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
    n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
    n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364,
    n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
    n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382,
    n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
    n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
    n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
    n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
    n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
    n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
    n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
    n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454,
    n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
    n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
    n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
    n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
    n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
    n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
    n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
    n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
    n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
    n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
    n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
    n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
    n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
    n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
    n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598,
    n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
    n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
    n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
    n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
    n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
    n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
    n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
    n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
    n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
    n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
    n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
    n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
    n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
    n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
    n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
    n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
    n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
    n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
    n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
    n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
    n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
    n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
    n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
    n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
    n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
    n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
    n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
    n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
    n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
    n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
    n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
    n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
    n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
    n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
    n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102,
    n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
    n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
    n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
    n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
    n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
    n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
    n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
    n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
    n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
    n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
    n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
    n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
    n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
    n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
    n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
    n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
    n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
    n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
    n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
    n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
    n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
    n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
    n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
    n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
    n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
    n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
    n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
    n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
    n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
    n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
    n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
    n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
    n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
    n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
    n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
    n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
    n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
    n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
    n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
    n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
    n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
    n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
    n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
    n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
    n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
    n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
    n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
    n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
    n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
    n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
    n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
    n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
    n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
    n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
    n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
    n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
    n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
    n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
    n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
    n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
    n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
    n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
    n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
    n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
    n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
    n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
    n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
    n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
    n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
    n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
    n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
    n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
    n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
    n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
    n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
    n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
    n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
    n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
    n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
    n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542,
    n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
    n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
    n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
    n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614,
    n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
    n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
    n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
    n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686,
    n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
    n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
    n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
    n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758,
    n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
    n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
    n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
    n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
    n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
    n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
    n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
    n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
    n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
    n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
    n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
    n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
    n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
    n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
    n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
    n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
    n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
    n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
    n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
    n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
    n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
    n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
    n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
    n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
    n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
    n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
    n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
    n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
    n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
    n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
    n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
    n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
    n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
    n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
    n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
    n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
    n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
    n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
    n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334,
    n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
    n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
    n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
    n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
    n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
    n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
    n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
    n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406,
    n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
    n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
    n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
    n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
    n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
    n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
    n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
    n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
    n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550,
    n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559,
    n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
    n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
    n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
    n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
    n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
    n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
    n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
    n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
    n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
    n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
    n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
    n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
    n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
    n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
    n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784,
    n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
    n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
    n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838,
    n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856,
    n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
    n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
    n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
    n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928,
    n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
    n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
    n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
    n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000,
    n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
    n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
    n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054,
    n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072,
    n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
    n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
    n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
    n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
    n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
    n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
    n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198,
    n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216,
    n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
    n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
    n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
    n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
    n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
    n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
    n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
    n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
    n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
    n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
    n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
    n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
    n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
    n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
    n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
    n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486,
    n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
    n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504,
    n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
    n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
    n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558,
    n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
    n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
    n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
    n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
    n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630,
    n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
    n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648,
    n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
    n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
    n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
    n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
    n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
    n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
    n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720,
    n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
    n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
    n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
    n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
    n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
    n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
    n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846,
    n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864,
    n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
    n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
    n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
    n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936,
    n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
    n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
    n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990,
    n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
    n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
    n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
    n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
    n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
    n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
    n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
    n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
    n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
    n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
    n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
    n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
    n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
    n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
    n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
    n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
    n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
    n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
    n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
    n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
    n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
    n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
    n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764,
    n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
    n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
    n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
    n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
    n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
    n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
    n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
    n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980,
    n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989,
    n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
    n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
    n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
    n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
    n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
    n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
    n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
    n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061,
    n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
    n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
    n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
    n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
    n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
    n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
    n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
    n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
    n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
    n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
    n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
    n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
    n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
    n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
    n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
    n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412,
    n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
    n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
    n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
    n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
    n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
    n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
    n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
    n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
    n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
    n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
    n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
    n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
    n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
    n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
    n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
    n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
    n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
    n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
    n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
    n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628,
    n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637,
    n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
    n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
    n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
    n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
    n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
    n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
    n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709,
    n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
    n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
    n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
    n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
    n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
    n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
    n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
    n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
    n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
    n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
    n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
    n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
    n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
    n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853,
    n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
    n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
    n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
    n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916,
    n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925,
    n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
    n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
    n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
    n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
    n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
    n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
    n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997,
    n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
    n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
    n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
    n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
    n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
    n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
    n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060,
    n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
    n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
    n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
    n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
    n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114,
    n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
    n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132,
    n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141,
    n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
    n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
    n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
    n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
    n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204,
    n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213,
    n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
    n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
    n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
    n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
    n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258,
    n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
    n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
    n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285,
    n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
    n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
    n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
    n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
    n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
    n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
    n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348,
    n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357,
    n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
    n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
    n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
    n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
    n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
    n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
    n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
    n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
    n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
    n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
    n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
    n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
    n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
    n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
    n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501,
    n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
    n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
    n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
    n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
    n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
    n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
    n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564,
    n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573,
    n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
    n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
    n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
    n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
    n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
    n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
    n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
    n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
    n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
    n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
    n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
    n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
    n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
    n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
    n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
    n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789,
    n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
    n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
    n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816,
    n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
    n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
    n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
    n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
    n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861,
    n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
    n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
    n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888,
    n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
    n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906,
    n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
    n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
    n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933,
    n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
    n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
    n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960,
    n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
    n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
    n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
    n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
    n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005,
    n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
    n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023,
    n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
    n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
    n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
    n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077,
    n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
    n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095,
    n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
    n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
    n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
    n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
    n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
    n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149,
    n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
    n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167,
    n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176,
    n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
    n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
    n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
    n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
    n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221,
    n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
    n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239,
    n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248,
    n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
    n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
    n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
    n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
    n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293,
    n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
    n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320,
    n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
    n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
    n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
    n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
    n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
    n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
    n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
    n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
    n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437,
    n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
    n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455,
    n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
    n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
    n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
    n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
    n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
    n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509,
    n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
    n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
    n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
    n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
    n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
    n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
    n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
    n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581,
    n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
    n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599,
    n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608,
    n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
    n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
    n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
    n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644,
    n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653,
    n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
    n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
    n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680,
    n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
    n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
    n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
    n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
    n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725,
    n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
    n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743,
    n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752,
    n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
    n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
    n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
    n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788,
    n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797,
    n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
    n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815,
    n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824,
    n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
    n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
    n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
    n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
    n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
    n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887,
    n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
    n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
    n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
    n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
    n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
    n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941,
    n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
    n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959,
    n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968,
    n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
    n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
    n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
    n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013,
    n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
    n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040,
    n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
    n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
    n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
    n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076,
    n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085,
    n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
    n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103,
    n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
    n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
    n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
    n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
    n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148,
    n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157,
    n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
    n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
    n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184,
    n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
    n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202,
    n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
    n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
    n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229,
    n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
    n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
    n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
    n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
    n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
    n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328,
    n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
    n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
    n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
    n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400,
    n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
    n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
    n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
    n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
    n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445,
    n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
    n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463,
    n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472,
    n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
    n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
    n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
    n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
    n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535,
    n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544,
    n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
    n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562,
    n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
    n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
    n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589,
    n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
    n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616,
    n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
    n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634,
    n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
    n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652,
    n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661,
    n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
    n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679,
    n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688,
    n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
    n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
    n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
    n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
    n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
    n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
    n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
    n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805,
    n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
    n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823,
    n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832,
    n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
    n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850,
    n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
    n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868,
    n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877,
    n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
    n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895,
    n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904,
    n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
    n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922,
    n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
    n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940,
    n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949,
    n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
    n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
    n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976,
    n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
    n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994,
    n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
    n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
    n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021,
    n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
    n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039,
    n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048,
    n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
    n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
    n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
    n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084,
    n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093,
    n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
    n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111,
    n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120,
    n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
    n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
    n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156,
    n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165,
    n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
    n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183,
    n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192,
    n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
    n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
    n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
    n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228,
    n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237,
    n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
    n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255,
    n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264,
    n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
    n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282,
    n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
    n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300,
    n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309,
    n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
    n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
    n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
    n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
    n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
    n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
    n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
    n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381,
    n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
    n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
    n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
    n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
    n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426,
    n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
    n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444,
    n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453,
    n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
    n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
    n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
    n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
    n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
    n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
    n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516,
    n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525,
    n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
    n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
    n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552,
    n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
    n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
    n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
    n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588,
    n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597,
    n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
    n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
    n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624,
    n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
    n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642,
    n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
    n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660,
    n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669,
    n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
    n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
    n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696,
    n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
    n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714,
    n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
    n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732,
    n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741,
    n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
    n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
    n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
    n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786,
    n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
    n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804,
    n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813,
    n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
    n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831,
    n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840,
    n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
    n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
    n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
    n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876,
    n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885,
    n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
    n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903,
    n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912,
    n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
    n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
    n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
    n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948,
    n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957,
    n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
    n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975,
    n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984,
    n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
    n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002,
    n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
    n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020,
    n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029,
    n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
    n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047,
    n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056,
    n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
    n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
    n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092,
    n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101,
    n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
    n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119,
    n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
    n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173,
    n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191,
    n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200,
    n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
    n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
    n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236,
    n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
    n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
    n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
    n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308,
    n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317,
    n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
    n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
    n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
    n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
    n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
    n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
    n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
    n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389,
    n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
    n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
    n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
    n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
    n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452,
    n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
    n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
    n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
    n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524,
    n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
    n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
    n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
    n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
    n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
    n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632,
    n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650,
    n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
    n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668,
    n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677,
    n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
    n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704,
    n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
    n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722,
    n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740,
    n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749,
    n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
    n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776,
    n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
    n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794,
    n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
    n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812,
    n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821,
    n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
    n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839,
    n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
    n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
    n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866,
    n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
    n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884,
    n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893,
    n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
    n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911,
    n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920,
    n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
    n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938,
    n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956,
    n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965,
    n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
    n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983,
    n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992,
    n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
    n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010,
    n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
    n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028,
    n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037,
    n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
    n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
    n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064,
    n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
    n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082,
    n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
    n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100,
    n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109,
    n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
    n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127,
    n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
    n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
    n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
    n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
    n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172,
    n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181,
    n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
    n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199,
    n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
    n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
    n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226,
    n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
    n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244,
    n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253,
    n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
    n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271,
    n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280,
    n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
    n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298,
    n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
    n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316,
    n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325,
    n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
    n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
    n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
    n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
    n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388,
    n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397,
    n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
    n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415,
    n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424,
    n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
    n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442,
    n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
    n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460,
    n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
    n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487,
    n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496,
    n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
    n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514,
    n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
    n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532,
    n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541,
    n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
    n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568,
    n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
    n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
    n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
    n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604,
    n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613,
    n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
    n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
    n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640,
    n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
    n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
    n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
    n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676,
    n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685,
    n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
    n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703,
    n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712,
    n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
    n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
    n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
    n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748,
    n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757,
    n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
    n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775,
    n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784,
    n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
    n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
    n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829,
    n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847,
    n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
    n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
    n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
    n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892,
    n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901,
    n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
    n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919,
    n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
    n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
    n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
    n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
    n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964,
    n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973,
    n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
    n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991,
    n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
    n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
    n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
    n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
    n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036,
    n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045,
    n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
    n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063,
    n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
    n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
    n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
    n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117,
    n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
    n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
    n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
    n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
    n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
    n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
    n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180,
    n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189,
    n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
    n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207,
    n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
    n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
    n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
    n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
    n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252,
    n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261,
    n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
    n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
    n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
    n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
    n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
    n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
    n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324,
    n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333,
    n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
    n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351,
    n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
    n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
    n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
    n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
    n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396,
    n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405,
    n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
    n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423,
    n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
    n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
    n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
    n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
    n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468,
    n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477,
    n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
    n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495,
    n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
    n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
    n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
    n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531,
    n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540,
    n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549,
    n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
    n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567,
    n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
    n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
    n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594,
    n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603,
    n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612,
    n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621,
    n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
    n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639,
    n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
    n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
    n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666,
    n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675,
    n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684,
    n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693,
    n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
    n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711,
    n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720,
    n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
    n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738,
    n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747,
    n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756,
    n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765,
    n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
    n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783,
    n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
    n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
    n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
    n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819,
    n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828,
    n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837,
    n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
    n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
    n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
    n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
    n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
    n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
    n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900,
    n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909,
    n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
    n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927,
    n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936,
    n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
    n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954,
    n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963,
    n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972,
    n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981,
    n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
    n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999,
    n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008,
    n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
    n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026,
    n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035,
    n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044,
    n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053,
    n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
    n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071,
    n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080,
    n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
    n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
    n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
    n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116,
    n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125,
    n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
    n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143,
    n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
    n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
    n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170,
    n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179,
    n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188,
    n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197,
    n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
    n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215,
    n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
    n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
    n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242,
    n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251,
    n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260,
    n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269,
    n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
    n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287,
    n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
    n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
    n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
    n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
    n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332,
    n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341,
    n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
    n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359,
    n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368,
    n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
    n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
    n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395,
    n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404,
    n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413,
    n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
    n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431,
    n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
    n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
    n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
    n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467,
    n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476,
    n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485,
    n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
    n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
    n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
    n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
    n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
    n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
    n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
    n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
    n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
    n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
    n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
    n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
    n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620,
    n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629,
    n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
    n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647,
    n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
    n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
    n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
    n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683,
    n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692,
    n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701,
    n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
    n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
    n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
    n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
    n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
    n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
    n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764,
    n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773,
    n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
    n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
    n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
    n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
    n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
    n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
    n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836,
    n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845,
    n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
    n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863,
    n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
    n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
    n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
    n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
    n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908,
    n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917,
    n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
    n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
    n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
    n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
    n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980,
    n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989,
    n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
    n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
    n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
    n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
    n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
    n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
    n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052,
    n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061,
    n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
    n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079,
    n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
    n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
    n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
    n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124,
    n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133,
    n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
    n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151,
    n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160,
    n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
    n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
    n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196,
    n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
    n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223,
    n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
    n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
    n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
    n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259,
    n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268,
    n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277,
    n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
    n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295,
    n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
    n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
    n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
    n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331,
    n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340,
    n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349,
    n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
    n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367,
    n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
    n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
    n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
    n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403,
    n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412,
    n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421,
    n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
    n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439,
    n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
    n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
    n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
    n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475,
    n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484,
    n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493,
    n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502,
    n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511,
    n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
    n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
    n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
    n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
    n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556,
    n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565,
    n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574,
    n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583,
    n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
    n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
    n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
    n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
    n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628,
    n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637,
    n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646,
    n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
    n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
    n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700,
    n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
    n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727,
    n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
    n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
    n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
    n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763,
    n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772,
    n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, n39781,
    n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
    n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799,
    n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
    n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
    n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
    n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
    n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844,
    n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852, n39853,
    n39854, n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
    n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871,
    n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
    n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
    n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
    n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
    n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916,
    n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924, n39925,
    n39926, n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
    n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943,
    n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
    n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
    n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
    n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979,
    n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988,
    n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996, n39997,
    n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006,
    n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015,
    n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
    n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
    n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
    n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051,
    n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060,
    n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068, n40069,
    n40070, n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078,
    n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087,
    n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
    n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
    n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
    n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123,
    n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132,
    n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141,
    n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
    n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159,
    n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
    n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
    n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
    n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
    n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204,
    n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212, n40213,
    n40214, n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222,
    n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
    n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
    n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
    n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
    n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276,
    n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284, n40285,
    n40286, n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294,
    n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303,
    n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
    n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
    n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
    n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339,
    n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348,
    n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356, n40357,
    n40358, n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
    n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375,
    n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
    n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
    n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
    n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411,
    n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420,
    n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428, n40429,
    n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438,
    n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447,
    n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
    n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
    n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
    n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
    n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492,
    n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501,
    n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
    n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
    n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
    n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
    n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
    n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
    n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564,
    n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573,
    n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582,
    n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591,
    n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
    n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
    n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
    n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
    n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636,
    n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645,
    n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654,
    n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663,
    n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
    n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
    n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
    n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
    n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708,
    n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717,
    n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
    n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
    n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
    n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
    n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
    n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
    n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780,
    n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789,
    n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
    n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807,
    n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
    n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
    n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
    n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
    n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852,
    n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861,
    n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
    n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879,
    n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888,
    n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
    n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
    n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
    n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924,
    n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933,
    n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942,
    n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951,
    n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960,
    n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
    n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
    n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
    n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996,
    n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005,
    n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014,
    n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023,
    n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032,
    n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
    n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
    n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
    n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068,
    n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077,
    n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086,
    n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095,
    n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104,
    n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
    n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
    n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
    n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
    n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149,
    n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158,
    n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167,
    n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
    n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
    n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
    n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
    n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212,
    n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221,
    n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230,
    n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
    n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
    n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
    n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284,
    n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293,
    n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302,
    n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311,
    n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320,
    n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
    n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
    n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
    n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356,
    n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365,
    n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374,
    n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383,
    n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392,
    n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
    n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
    n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419,
    n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428,
    n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437,
    n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446,
    n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455,
    n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464,
    n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
    n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
    n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491,
    n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500,
    n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509,
    n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518,
    n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
    n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536,
    n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
    n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
    n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563,
    n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572,
    n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581,
    n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590,
    n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
    n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
    n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
    n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
    n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644,
    n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653,
    n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662,
    n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671,
    n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
    n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
    n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
    n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707,
    n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716,
    n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724, n41725,
    n41726, n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734,
    n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743,
    n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752,
    n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
    n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
    n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779,
    n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788,
    n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796, n41797,
    n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806,
    n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815,
    n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824,
    n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
    n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
    n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851,
    n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860,
    n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868, n41869,
    n41870, n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878,
    n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887,
    n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896,
    n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
    n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
    n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
    n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932,
    n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940, n41941,
    n41942, n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950,
    n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959,
    n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968,
    n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
    n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
    n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995,
    n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004,
    n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42013,
    n42014, n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022,
    n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031,
    n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
    n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
    n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
    n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
    n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076,
    n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085,
    n42086, n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
    n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103,
    n42104, n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112,
    n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
    n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
    n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139,
    n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148,
    n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157,
    n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
    n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174, n42175,
    n42176, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
    n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
    n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
    n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211,
    n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220,
    n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229,
    n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
    n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246, n42247,
    n42248, n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256,
    n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
    n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
    n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283,
    n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292,
    n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301,
    n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310,
    n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318, n42319,
    n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328,
    n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337,
    n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
    n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
    n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364,
    n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373,
    n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382,
    n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390, n42391,
    n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400,
    n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409,
    n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
    n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427,
    n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436,
    n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444, n42445,
    n42446, n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
    n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462, n42463,
    n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472,
    n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481,
    n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
    n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
    n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508,
    n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517,
    n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526,
    n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535,
    n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544,
    n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553,
    n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
    n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
    n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580,
    n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589,
    n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
    n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607,
    n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616,
    n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625,
    n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
    n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643,
    n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652,
    n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42661,
    n42662, n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
    n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679,
    n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688,
    n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697,
    n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
    n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715,
    n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724,
    n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732, n42733,
    n42734, n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
    n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751,
    n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760,
    n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769,
    n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
    n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787,
    n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796,
    n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804, n42805,
    n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814,
    n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823,
    n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
    n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
    n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
    n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859,
    n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868,
    n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876, n42877,
    n42878, n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886,
    n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895,
    n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904,
    n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
    n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
    n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931,
    n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940,
    n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949,
    n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
    n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967,
    n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976,
    n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985,
    n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
    n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
    n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012,
    n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020, n43021,
    n43022, n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030,
    n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039,
    n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048,
    n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057,
    n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
    n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
    n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084,
    n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092, n43093,
    n43094, n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
    n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111,
    n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120,
    n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
    n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
    n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156,
    n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165,
    n43166, n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174,
    n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182, n43183,
    n43184, n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192,
    n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201,
    n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
    n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
    n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228,
    n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237,
    n43238, n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246,
    n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255,
    n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264,
    n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273,
    n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
    n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
    n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300,
    n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308, n43309,
    n43310, n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318,
    n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326, n43327,
    n43328, n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336,
    n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
    n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
    n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
    n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372,
    n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381,
    n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
    n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399,
    n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
    n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
    n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
    n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
    n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444,
    n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453,
    n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
    n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471,
    n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
    n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
    n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
    n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
    n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516,
    n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525,
    n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
    n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543,
    n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552,
    n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
    n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
    n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588,
    n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597,
    n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
    n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615,
    n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624,
    n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
    n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
    n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
    n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660,
    n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669,
    n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
    n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687,
    n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
    n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
    n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
    n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
    n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732,
    n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741,
    n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
    n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759,
    n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768,
    n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
    n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
    n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
    n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804,
    n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813,
    n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
    n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831,
    n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840,
    n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
    n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
    n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
    n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876,
    n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885,
    n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
    n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903,
    n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
    n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
    n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
    n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
    n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948,
    n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957,
    n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
    n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975,
    n43976, n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984,
    n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993,
    n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
    n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
    n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020,
    n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029,
    n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038,
    n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047,
    n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056,
    n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065,
    n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
    n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
    n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092,
    n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100, n44101,
    n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110,
    n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119,
    n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128,
    n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137,
    n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
    n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
    n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164,
    n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173,
    n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
    n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191,
    n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200,
    n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209,
    n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
    n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
    n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236,
    n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245,
    n44246, n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254,
    n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263,
    n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272,
    n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281,
    n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
    n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
    n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308,
    n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316, n44317,
    n44318, n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326,
    n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335,
    n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344,
    n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353,
    n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
    n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
    n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380,
    n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388, n44389,
    n44390, n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398,
    n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406, n44407,
    n44408, n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416,
    n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425,
    n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
    n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
    n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452,
    n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460, n44461,
    n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
    n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478, n44479,
    n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488,
    n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497,
    n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
    n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
    n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524,
    n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532, n44533,
    n44534, n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542,
    n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551,
    n44552, n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560,
    n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
    n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
    n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
    n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596,
    n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604, n44605,
    n44606, n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614,
    n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622, n44623,
    n44624, n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632,
    n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
    n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
    n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
    n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668,
    n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676, n44677,
    n44678, n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686,
    n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694, n44695,
    n44696, n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704,
    n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713,
    n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
    n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
    n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740,
    n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748, n44749,
    n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758,
    n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766, n44767,
    n44768, n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776,
    n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785,
    n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
    n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
    n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812,
    n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821,
    n44822, n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
    n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838, n44839,
    n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848,
    n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857,
    n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
    n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
    n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884,
    n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892, n44893,
    n44894, n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
    n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910, n44911,
    n44912, n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920,
    n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929,
    n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
    n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
    n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956,
    n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965,
    n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
    n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983,
    n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
    n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
    n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
    n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
    n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028,
    n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037,
    n45038, n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046,
    n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055,
    n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064,
    n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073,
    n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
    n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
    n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100,
    n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109,
    n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118,
    n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127,
    n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136,
    n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145,
    n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
    n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
    n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172,
    n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180, n45181,
    n45182, n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190,
    n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199,
    n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208,
    n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217,
    n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
    n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
    n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244,
    n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252, n45253,
    n45254, n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262,
    n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271,
    n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280,
    n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289,
    n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
    n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307,
    n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316,
    n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324, n45325,
    n45326, n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334,
    n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343,
    n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
    n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361,
    n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
    n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379,
    n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388,
    n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397,
    n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
    n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415,
    n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424,
    n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
    n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
    n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
    n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460,
    n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469,
    n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
    n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487,
    n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496,
    n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505,
    n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
    n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523,
    n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532,
    n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541,
    n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550,
    n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559,
    n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568,
    n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577,
    n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
    n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595,
    n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604,
    n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613,
    n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622,
    n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631,
    n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640,
    n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649,
    n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
    n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667,
    n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676,
    n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685,
    n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
    n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703,
    n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712,
    n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721,
    n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
    n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739,
    n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748,
    n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756, n45757,
    n45758, n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
    n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775,
    n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784,
    n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793,
    n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
    n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811,
    n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820,
    n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828, n45829,
    n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838,
    n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847,
    n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
    n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865,
    n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
    n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883,
    n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892,
    n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900, n45901,
    n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910,
    n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919,
    n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928,
    n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
    n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
    n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955,
    n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964,
    n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973,
    n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
    n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991,
    n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000,
    n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009,
    n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
    n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027,
    n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036,
    n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045,
    n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054,
    n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063,
    n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072,
    n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081,
    n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
    n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099,
    n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108,
    n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116, n46117,
    n46118, n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
    n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135,
    n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144,
    n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153,
    n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
    n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171,
    n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180,
    n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188, n46189,
    n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198,
    n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207,
    n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216,
    n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225,
    n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
    n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243,
    n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252,
    n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261,
    n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270,
    n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279,
    n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288,
    n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297,
    n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
    n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315,
    n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324,
    n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333,
    n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342,
    n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351,
    n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360,
    n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369,
    n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
    n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387,
    n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396,
    n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405,
    n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414,
    n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423,
    n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432,
    n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441,
    n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
    n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459,
    n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468,
    n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477,
    n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486,
    n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495,
    n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504,
    n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513,
    n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
    n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531,
    n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540,
    n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549,
    n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558,
    n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567,
    n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576,
    n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585,
    n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
    n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603,
    n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612,
    n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621,
    n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630,
    n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639,
    n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648,
    n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657,
    n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
    n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675,
    n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684,
    n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693,
    n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702,
    n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711,
    n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720,
    n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729,
    n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
    n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747,
    n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756,
    n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765,
    n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774,
    n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783,
    n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792,
    n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801,
    n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
    n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
    n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828,
    n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837,
    n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846,
    n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855,
    n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864,
    n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873,
    n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
    n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891,
    n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900,
    n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909,
    n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918,
    n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927,
    n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936,
    n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945,
    n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
    n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
    n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972,
    n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981,
    n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990,
    n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999,
    n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008,
    n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017,
    n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
    n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035,
    n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044,
    n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052, n47053,
    n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062,
    n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071,
    n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080,
    n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
    n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
    n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107,
    n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116,
    n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125,
    n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
    n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143,
    n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152,
    n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
    n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
    n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179,
    n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188,
    n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197,
    n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206,
    n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215,
    n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224,
    n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233,
    n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
    n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251,
    n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260,
    n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269,
    n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
    n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287,
    n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296,
    n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305,
    n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
    n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323,
    n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332,
    n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340, n47341,
    n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350,
    n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359,
    n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
    n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
    n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
    n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395,
    n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404,
    n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413,
    n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422,
    n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431,
    n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440,
    n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449,
    n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
    n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467,
    n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476,
    n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484, n47485,
    n47486, n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494,
    n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503,
    n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512,
    n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521,
    n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
    n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539,
    n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548,
    n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557,
    n47558, n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566,
    n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575,
    n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584,
    n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593,
    n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
    n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611,
    n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620,
    n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629,
    n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638,
    n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647,
    n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656,
    n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
    n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
    n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683,
    n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692,
    n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701,
    n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710,
    n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719,
    n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728,
    n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737,
    n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
    n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755,
    n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764,
    n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773,
    n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782,
    n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791,
    n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800,
    n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809,
    n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
    n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827,
    n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836,
    n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845,
    n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
    n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863,
    n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872,
    n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881,
    n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
    n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899,
    n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908,
    n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917,
    n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926,
    n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935,
    n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944,
    n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953,
    n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
    n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971,
    n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980,
    n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989,
    n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998,
    n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007,
    n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016,
    n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025,
    n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
    n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043,
    n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052,
    n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061,
    n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070,
    n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079,
    n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088,
    n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097,
    n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
    n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115,
    n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124,
    n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133,
    n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
    n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151,
    n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
    n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169,
    n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
    n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187,
    n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196,
    n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205,
    n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214,
    n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223,
    n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232,
    n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241,
    n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
    n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259,
    n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268,
    n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277,
    n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286,
    n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295,
    n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304,
    n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313,
    n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
    n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331,
    n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340,
    n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349,
    n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358,
    n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367,
    n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376,
    n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385,
    n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
    n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403,
    n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412,
    n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421,
    n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430,
    n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439,
    n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448,
    n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457,
    n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
    n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475,
    n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484,
    n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493,
    n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502,
    n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511,
    n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520,
    n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529,
    n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
    n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547,
    n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556,
    n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565,
    n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574,
    n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583,
    n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592,
    n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601,
    n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
    n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619,
    n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628,
    n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637,
    n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646,
    n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655,
    n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664,
    n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673,
    n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
    n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691,
    n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700,
    n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709,
    n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718,
    n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727,
    n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
    n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745,
    n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
    n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763,
    n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772,
    n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781,
    n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790,
    n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799,
    n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808,
    n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817,
    n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
    n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835,
    n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844,
    n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853,
    n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862,
    n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871,
    n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880,
    n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889,
    n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
    n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907,
    n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916,
    n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925,
    n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934,
    n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943,
    n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952,
    n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961,
    n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
    n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979,
    n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988,
    n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997,
    n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006,
    n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015,
    n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024,
    n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033,
    n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
    n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051,
    n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060,
    n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069,
    n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078,
    n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087,
    n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096,
    n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105,
    n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
    n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123,
    n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132,
    n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141,
    n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150,
    n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159,
    n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168,
    n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177,
    n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
    n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195,
    n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204,
    n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213,
    n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222,
    n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231,
    n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240,
    n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249,
    n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
    n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267,
    n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276,
    n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285,
    n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294,
    n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303,
    n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312,
    n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321,
    n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
    n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339,
    n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348,
    n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357,
    n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366,
    n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375,
    n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384,
    n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393,
    n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
    n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411,
    n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420,
    n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429,
    n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438,
    n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447,
    n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456,
    n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465,
    n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
    n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483,
    n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492,
    n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500, n49501,
    n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510,
    n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519,
    n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528,
    n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537,
    n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
    n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555,
    n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564,
    n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573,
    n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582,
    n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591,
    n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600,
    n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609,
    n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
    n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627,
    n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636,
    n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645,
    n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654,
    n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663,
    n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672,
    n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681,
    n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
    n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699,
    n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708,
    n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716, n49717,
    n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726,
    n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735,
    n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744,
    n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753,
    n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
    n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771,
    n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780,
    n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789,
    n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
    n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807,
    n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816,
    n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825,
    n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
    n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843,
    n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852,
    n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860, n49861,
    n49862, n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870,
    n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879,
    n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888,
    n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897,
    n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
    n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915,
    n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924,
    n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933,
    n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942,
    n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951,
    n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960,
    n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969,
    n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
    n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987,
    n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996,
    n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004, n50005,
    n50006, n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
    n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023,
    n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032,
    n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041,
    n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
    n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059,
    n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068,
    n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076, n50077,
    n50078, n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086,
    n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095,
    n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104,
    n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113,
    n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
    n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131,
    n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140,
    n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148, n50149,
    n50150, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158,
    n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167,
    n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
    n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185,
    n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
    n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203,
    n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212,
    n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221,
    n50222, n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230,
    n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239,
    n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248,
    n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257,
    n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
    n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275,
    n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284,
    n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292, n50293,
    n50294, n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302,
    n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311,
    n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
    n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329,
    n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
    n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347,
    n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356,
    n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365,
    n50366, n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374,
    n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383,
    n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
    n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401,
    n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
    n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419,
    n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428,
    n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437,
    n50438, n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446,
    n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455,
    n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464,
    n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473,
    n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
    n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491,
    n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500,
    n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508, n50509,
    n50510, n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518,
    n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527,
    n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536,
    n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545,
    n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
    n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
    n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572,
    n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581,
    n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590,
    n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599,
    n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
    n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617,
    n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
    n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635,
    n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644,
    n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652, n50653,
    n50654, n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662,
    n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671,
    n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680,
    n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689,
    n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
    n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
    n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716,
    n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724, n50725,
    n50726, n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734,
    n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743,
    n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752,
    n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761,
    n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
    n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779,
    n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788,
    n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797,
    n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806,
    n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815,
    n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824,
    n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833,
    n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
    n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851,
    n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860,
    n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868, n50869,
    n50870, n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878,
    n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887,
    n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896,
    n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905,
    n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
    n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923,
    n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932,
    n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940, n50941,
    n50942, n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950,
    n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959,
    n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968,
    n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977,
    n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
    n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995,
    n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004,
    n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012, n51013,
    n51014, n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022,
    n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031,
    n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040,
    n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049,
    n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
    n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067,
    n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076,
    n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51085,
    n51086, n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094,
    n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103,
    n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112,
    n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121,
    n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
    n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139,
    n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148,
    n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157,
    n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166,
    n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175,
    n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184,
    n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193,
    n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
    n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211,
    n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220,
    n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228, n51229,
    n51230, n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238,
    n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247,
    n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256,
    n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265,
    n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
    n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283,
    n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292,
    n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301,
    n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310,
    n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319,
    n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328,
    n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337,
    n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
    n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355,
    n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364,
    n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373,
    n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382,
    n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391,
    n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400,
    n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409,
    n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
    n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427,
    n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436,
    n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445,
    n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454,
    n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463,
    n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472,
    n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481,
    n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
    n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499,
    n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508,
    n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517,
    n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526,
    n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535,
    n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544,
    n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553,
    n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
    n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571,
    n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580,
    n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589,
    n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598,
    n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607,
    n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616,
    n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625,
    n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
    n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643,
    n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652,
    n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661,
    n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670,
    n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679,
    n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688,
    n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697,
    n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
    n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715,
    n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724,
    n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733,
    n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742,
    n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751,
    n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760,
    n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769,
    n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
    n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787,
    n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796,
    n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805,
    n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814,
    n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823,
    n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832,
    n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841,
    n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
    n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859,
    n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868,
    n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877,
    n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886,
    n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895,
    n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904,
    n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913,
    n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
    n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931,
    n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940,
    n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949,
    n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958,
    n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967,
    n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976,
    n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985,
    n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
    n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003,
    n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012,
    n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021,
    n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030,
    n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039,
    n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048,
    n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057,
    n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
    n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075,
    n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084,
    n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093,
    n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102,
    n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111,
    n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120,
    n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129,
    n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
    n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147,
    n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156,
    n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165,
    n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174,
    n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183,
    n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192,
    n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201,
    n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
    n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219,
    n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228,
    n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237,
    n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246,
    n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255,
    n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264,
    n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273,
    n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
    n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291,
    n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
    n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309,
    n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318,
    n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327,
    n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336,
    n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345,
    n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
    n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363,
    n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372,
    n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381,
    n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390,
    n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399,
    n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408,
    n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417,
    n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
    n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435,
    n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444,
    n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453,
    n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462,
    n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471,
    n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480,
    n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489,
    n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
    n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507,
    n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
    n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525,
    n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534,
    n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543,
    n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552,
    n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561,
    n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
    n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579,
    n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
    n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597,
    n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606,
    n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615,
    n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624,
    n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633,
    n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
    n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651,
    n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660,
    n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669,
    n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678,
    n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687,
    n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696,
    n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705,
    n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
    n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723,
    n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732,
    n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741,
    n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750,
    n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759,
    n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768,
    n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777,
    n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
    n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795,
    n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804,
    n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813,
    n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822,
    n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831,
    n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840,
    n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849,
    n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
    n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867,
    n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876,
    n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885,
    n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894,
    n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903,
    n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912,
    n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921,
    n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
    n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939,
    n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948,
    n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957,
    n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966,
    n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975,
    n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984,
    n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993,
    n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
    n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011,
    n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020,
    n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029,
    n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038,
    n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047,
    n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056,
    n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065,
    n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
    n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083,
    n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
    n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101,
    n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110,
    n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119,
    n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128,
    n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137,
    n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
    n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155,
    n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164,
    n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173,
    n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182,
    n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191,
    n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200,
    n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
    n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
    n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227,
    n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
    n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245,
    n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254,
    n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263,
    n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272,
    n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281,
    n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
    n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299,
    n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308,
    n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317,
    n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326,
    n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335,
    n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344,
    n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353,
    n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
    n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371,
    n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380,
    n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389,
    n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398,
    n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407,
    n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416,
    n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425,
    n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
    n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443,
    n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452,
    n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461,
    n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470,
    n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479,
    n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488,
    n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497,
    n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
    n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515,
    n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524,
    n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533,
    n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542,
    n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550, n53551,
    n53552, n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560,
    n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569,
    n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
    n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587,
    n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596,
    n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605,
    n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614,
    n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623,
    n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632,
    n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641,
    n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
    n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659,
    n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668,
    n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677,
    n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686,
    n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695,
    n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704,
    n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713,
    n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
    n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731,
    n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740,
    n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749,
    n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758,
    n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766, n53767,
    n53768, n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776,
    n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785,
    n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
    n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803,
    n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812,
    n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821,
    n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830,
    n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838, n53839,
    n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848,
    n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857,
    n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
    n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875,
    n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884,
    n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893,
    n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902,
    n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911,
    n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920,
    n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929,
    n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
    n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947,
    n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956,
    n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965,
    n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974,
    n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983,
    n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992,
    n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001,
    n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
    n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019,
    n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028,
    n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037,
    n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046,
    n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055,
    n54056, n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064,
    n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073,
    n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
    n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091,
    n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100,
    n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108, n54109,
    n54110, n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118,
    n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127,
    n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136,
    n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145,
    n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
    n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163,
    n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172,
    n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181,
    n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190,
    n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199,
    n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208,
    n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217,
    n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
    n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235,
    n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244,
    n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, n54253,
    n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262,
    n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271,
    n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280,
    n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289,
    n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
    n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307,
    n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316,
    n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324, n54325,
    n54326, n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334,
    n54335, n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343,
    n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352,
    n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361,
    n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
    n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379,
    n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388,
    n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396, n54397,
    n54398, n54399, n54400, n54401, n54402, n54403, n54404, n54405, n54406,
    n54407, n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415,
    n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424,
    n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433,
    n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
    n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451,
    n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460,
    n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468, n54469,
    n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478,
    n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487,
    n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496,
    n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505,
    n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
    n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523,
    n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532,
    n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541,
    n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550,
    n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559,
    n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568,
    n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
    n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
    n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595,
    n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604,
    n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613,
    n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622,
    n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631,
    n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640,
    n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649,
    n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
    n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667,
    n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676,
    n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685,
    n54686, n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694,
    n54695, n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703,
    n54704, n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712,
    n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721,
    n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
    n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739,
    n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748,
    n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756, n54757,
    n54758, n54759, n54760, n54761, n54762, n54763, n54764, n54765, n54766,
    n54767, n54768, n54769, n54770, n54771, n54772, n54773, n54774, n54775,
    n54776, n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784,
    n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793,
    n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
    n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811,
    n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820,
    n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828, n54829,
    n54830, n54831, n54832, n54833, n54834, n54835, n54836, n54837, n54838,
    n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846, n54847,
    n54848, n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856,
    n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865,
    n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
    n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883,
    n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892,
    n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900, n54901,
    n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54910,
    n54911, n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919,
    n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928,
    n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937,
    n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
    n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955,
    n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964,
    n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972, n54973,
    n54974, n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982,
    n54983, n54984, n54985, n54986, n54987, n54988, n54989, n54990, n54991,
    n54992, n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000,
    n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009,
    n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
    n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027,
    n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036,
    n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044, n55045,
    n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053, n55054,
    n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062, n55063,
    n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072,
    n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081,
    n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090,
    n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099,
    n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108,
    n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116, n55117,
    n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125, n55126,
    n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135,
    n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144,
    n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153,
    n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162,
    n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171,
    n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180,
    n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189,
    n55190, n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198,
    n55199, n55200, n55201, n55202, n55203, n55204, n55205, n55206, n55207,
    n55208, n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216,
    n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225,
    n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234,
    n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243,
    n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252,
    n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261,
    n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269, n55270,
    n55271, n55272, n55273, n55274, n55275, n55276, n55277, n55278, n55279,
    n55280, n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288,
    n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297,
    n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
    n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315,
    n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324,
    n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333,
    n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342,
    n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351,
    n55352, n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360,
    n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369,
    n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
    n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387,
    n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396,
    n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404, n55405,
    n55406, n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414,
    n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422, n55423,
    n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432,
    n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441,
    n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450,
    n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459,
    n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468,
    n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476, n55477,
    n55478, n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486,
    n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494, n55495,
    n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504,
    n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513,
    n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522,
    n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531,
    n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540,
    n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549,
    n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558,
    n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567,
    n55568, n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576,
    n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585,
    n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594,
    n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603,
    n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612,
    n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620, n55621,
    n55622, n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630,
    n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639,
    n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648,
    n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657,
    n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666,
    n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675,
    n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684,
    n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692, n55693,
    n55694, n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702,
    n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711,
    n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720,
    n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729,
    n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738,
    n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747,
    n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756,
    n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764, n55765,
    n55766, n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774,
    n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782, n55783,
    n55784, n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792,
    n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801,
    n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810,
    n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819,
    n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828,
    n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836, n55837,
    n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845, n55846,
    n55847, n55848, n55849, n55850, n55851, n55852, n55853, n55854, n55855,
    n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864,
    n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873,
    n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
    n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891,
    n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900,
    n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909,
    n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918,
    n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927,
    n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936,
    n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945,
    n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954,
    n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963,
    n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972,
    n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981,
    n55982, n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990,
    n55991, n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999,
    n56000, n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008,
    n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017,
    n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026,
    n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035,
    n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044,
    n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053,
    n56054, n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062,
    n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071,
    n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080,
    n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089,
    n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098,
    n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107,
    n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116,
    n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125,
    n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134,
    n56135, n56136, n56137, n56138, n56139, n56140, n56141, n56142, n56143,
    n56144, n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152,
    n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161,
    n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170,
    n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179,
    n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188,
    n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196, n56197,
    n56198, n56199, n56200, n56201, n56202, n56203, n56204, n56205, n56206,
    n56207, n56208, n56209, n56210, n56211, n56212, n56213, n56214, n56215,
    n56216, n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224,
    n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233,
    n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
    n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251,
    n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260,
    n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268, n56269,
    n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277, n56278,
    n56279, n56280, n56281, n56282, n56283, n56284, n56285, n56286, n56287,
    n56288, n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296,
    n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305,
    n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314,
    n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323,
    n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332,
    n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340, n56341,
    n56342, n56343, n56344, n56345, n56346, n56347, n56348, n56349, n56350,
    n56351, n56352, n56353, n56354, n56355, n56356, n56357, n56358, n56359,
    n56360, n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368,
    n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377,
    n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386,
    n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394, n56395,
    n56396, n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404,
    n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412, n56413,
    n56414, n56415, n56416, n56417, n56418, n56419, n56420, n56421, n56422,
    n56423, n56424, n56425, n56426, n56427, n56428, n56429, n56430, n56431,
    n56432, n56433, n56434, n56435, n56436, n56437, n56438, n56439, n56440,
    n56441, n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449,
    n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458,
    n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466, n56467,
    n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476,
    n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484, n56485,
    n56486, n56487, n56488, n56489, n56490, n56491, n56492, n56493, n56494,
    n56495, n56496, n56497, n56498, n56499, n56500, n56501, n56502, n56503,
    n56504, n56505, n56506, n56507, n56508, n56509, n56510, n56511, n56512,
    n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521,
    n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
    n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539,
    n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548,
    n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556, n56557,
    n56558, n56559, n56560, n56561, n56562, n56563, n56564, n56565, n56566,
    n56567, n56568, n56569, n56570, n56571, n56572, n56573, n56574, n56575,
    n56576, n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584,
    n56585, n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593,
    n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
    n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611,
    n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620,
    n56621, n56622, n56623, n56624, n56625, n56626, n56627, n56628, n56629,
    n56630, n56631, n56632, n56633, n56634, n56635, n56636, n56637, n56638,
    n56639, n56640, n56641, n56642, n56643, n56644, n56645, n56646, n56647,
    n56648, n56649, n56650, n56651, n56652, n56653, n56654, n56655, n56656,
    n56657, n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665,
    n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674,
    n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683,
    n56684, n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692,
    n56693, n56694, n56695, n56696, n56697, n56698, n56699, n56700, n56701,
    n56702, n56703, n56704, n56705, n56706, n56707, n56708, n56709, n56710,
    n56711, n56712, n56713, n56714, n56715, n56716, n56717, n56718, n56719,
    n56720, n56721, n56722, n56723, n56724, n56725, n56726, n56727, n56728,
    n56729, n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737,
    n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746,
    n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754, n56755,
    n56756, n56757, n56758, n56759, n56760, n56761, n56762, n56763, n56764,
    n56765, n56766, n56767, n56768, n56769, n56770, n56771, n56772, n56773,
    n56774, n56775, n56776, n56777, n56778, n56779, n56780, n56781, n56782,
    n56783, n56784, n56785, n56786, n56787, n56788, n56789, n56790, n56791,
    n56792, n56793, n56794, n56795, n56796, n56797, n56798, n56799, n56800,
    n56801, n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809,
    n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818,
    n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826, n56827,
    n56828, n56829, n56830, n56831, n56832, n56833, n56834, n56835, n56836,
    n56837, n56838, n56839, n56840, n56841, n56842, n56843, n56844, n56845,
    n56846, n56847, n56848, n56849, n56850, n56851, n56852, n56853, n56854,
    n56855, n56856, n56857, n56858, n56859, n56860, n56861, n56862, n56863,
    n56864, n56865, n56866, n56867, n56868, n56869, n56870, n56871, n56872,
    n56873, n56874, n56875, n56876, n56877, n56878, n56879, n56880, n56881,
    n56882, n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890,
    n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898, n56899,
    n56900, n56901, n56902, n56903, n56904, n56905, n56906, n56907, n56908,
    n56909, n56910, n56911, n56912, n56913, n56914, n56915, n56916, n56917,
    n56918, n56919, n56920, n56921, n56922, n56923, n56924, n56925, n56926,
    n56927, n56928, n56929, n56930, n56931, n56932, n56933, n56934, n56935,
    n56936, n56937, n56938, n56939, n56940, n56941, n56942, n56943, n56944,
    n56945, n56946, n56947, n56948, n56949, n56950, n56951, n56952, n56953,
    n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962,
    n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970, n56971,
    n56972, n56973, n56974, n56975, n56976, n56977, n56978, n56979, n56980,
    n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988, n56989,
    n56990, n56991, n56992, n56993, n56994, n56995, n56996, n56997, n56998,
    n56999, n57000, n57001, n57002, n57003, n57004, n57005, n57006, n57007,
    n57008, n57009, n57010, n57011, n57012, n57013, n57014, n57015, n57016,
    n57017, n57018, n57019, n57020, n57021, n57022, n57023, n57024, n57025,
    n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034,
    n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042, n57043,
    n57044, n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052,
    n57053, n57054, n57055, n57056, n57057, n57058, n57059, n57060, n57061,
    n57062, n57063, n57064, n57065, n57066, n57067, n57068, n57069, n57070,
    n57071, n57072, n57073, n57074, n57075, n57076, n57077, n57078, n57079,
    n57080, n57081, n57082, n57083, n57084, n57085, n57086, n57087, n57088,
    n57089, n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097,
    n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
    n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115,
    n57116, n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124,
    n57125, n57126, n57127, n57128, n57129, n57130, n57131, n57132, n57133,
    n57134, n57135, n57136, n57137, n57138, n57139, n57140, n57141, n57142,
    n57143, n57144, n57145, n57146, n57147, n57148, n57149, n57150, n57151,
    n57152, n57153, n57154, n57155, n57156, n57157, n57158, n57159, n57160,
    n57161, n57162, n57163, n57164, n57165, n57166, n57167, n57168, n57169,
    n57170, n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178,
    n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186, n57187,
    n57188, n57189, n57190, n57191, n57192, n57193, n57194, n57195, n57196,
    n57197, n57198, n57199, n57200, n57201, n57202, n57203, n57204, n57205,
    n57206, n57207, n57208, n57209, n57210, n57211, n57212, n57213, n57214,
    n57215, n57216, n57217, n57218, n57219, n57220, n57221, n57222, n57223,
    n57224, n57225, n57226, n57227, n57228, n57229, n57230, n57231, n57232,
    n57233, n57234, n57235, n57236, n57237, n57238, n57239, n57240, n57241,
    n57242, n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250,
    n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258, n57259,
    n57260, n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268,
    n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276, n57277,
    n57278, n57279, n57280, n57281, n57282, n57283, n57284, n57285, n57286,
    n57287, n57288, n57289, n57290, n57291, n57292, n57293, n57294, n57295,
    n57296, n57297, n57298, n57299, n57300, n57301, n57302, n57303, n57304,
    n57305, n57306, n57307, n57308, n57309, n57310, n57311, n57312, n57313,
    n57314, n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322,
    n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330, n57331,
    n57332, n57333, n57334, n57335, n57336, n57337, n57338, n57339, n57340,
    n57341, n57342, n57343, n57344, n57345, n57346, n57347, n57348, n57349,
    n57350, n57351, n57352, n57353, n57354, n57355, n57356, n57357, n57358,
    n57359, n57360, n57361, n57362, n57363, n57364, n57365, n57366, n57367,
    n57368, n57369, n57370, n57371, n57372, n57373, n57374, n57375, n57376,
    n57377, n57378, n57379, n57380, n57381, n57382, n57383, n57384, n57385,
    n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394,
    n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402, n57403,
    n57404, n57405, n57406, n57407, n57408, n57409, n57410, n57411, n57412,
    n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420, n57421,
    n57422, n57423, n57424, n57425, n57426, n57427, n57428, n57429, n57430,
    n57431, n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439,
    n57440, n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448,
    n57449, n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457,
    n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
    n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474, n57475,
    n57476, n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484,
    n57485, n57486, n57487, n57488, n57489, n57490, n57491, n57492, n57493,
    n57494, n57495, n57496, n57497, n57498, n57499, n57500, n57501, n57502,
    n57503, n57504, n57505, n57506, n57507, n57508, n57509, n57510, n57511,
    n57512, n57513, n57514, n57515, n57516, n57517, n57518, n57519, n57520,
    n57521, n57522, n57523, n57524, n57525, n57526, n57527, n57528, n57529,
    n57530, n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538,
    n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546, n57547,
    n57548, n57549, n57550, n57551, n57552, n57553, n57554, n57555, n57556,
    n57557, n57558, n57559, n57560, n57561, n57562, n57563, n57564, n57565,
    n57566, n57567, n57568, n57569, n57570, n57571, n57572, n57573, n57574,
    n57575, n57576, n57577, n57578, n57579, n57580, n57581, n57582, n57583,
    n57584, n57585, n57586, n57587, n57588, n57589, n57590, n57591, n57592,
    n57593, n57594, n57595, n57596, n57597, n57598, n57599, n57600, n57601,
    n57602, n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610,
    n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618, n57619,
    n57620, n57621, n57622, n57623, n57624, n57625, n57626, n57627, n57628,
    n57629, n57630, n57631, n57632, n57633, n57634, n57635, n57636, n57637,
    n57638, n57639, n57640, n57641, n57642, n57643, n57644, n57645, n57646,
    n57647, n57648, n57649, n57650, n57651, n57652, n57653, n57654, n57655,
    n57656, n57657, n57658, n57659, n57660, n57661, n57662, n57663, n57664,
    n57665, n57666, n57667, n57668, n57669, n57670, n57671, n57672, n57673,
    n57674, n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682,
    n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690, n57691,
    n57692, n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700,
    n57701, n57702, n57703, n57704, n57705, n57706, n57707, n57708, n57709,
    n57710, n57711, n57712, n57713, n57714, n57715, n57716, n57717, n57718,
    n57719, n57720, n57721, n57722, n57723, n57724, n57725, n57726, n57727,
    n57728, n57729, n57730, n57731, n57732, n57733, n57734, n57735, n57736,
    n57737, n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745,
    n57746, n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
    n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762, n57763,
    n57764, n57765, n57766, n57767, n57768, n57769, n57770, n57771, n57772,
    n57773, n57774, n57775, n57776, n57777, n57778, n57779, n57780, n57781,
    n57782, n57783, n57784, n57785, n57786, n57787, n57788, n57789, n57790,
    n57791, n57792, n57793, n57794, n57795, n57796, n57797, n57798, n57799,
    n57800, n57801, n57802, n57803, n57804, n57805, n57806, n57807, n57808,
    n57809, n57810, n57811, n57812, n57813, n57814, n57815, n57816, n57817,
    n57818, n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826,
    n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834, n57835,
    n57836, n57837, n57838, n57839, n57840, n57841, n57842, n57843, n57844,
    n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852, n57853,
    n57854, n57855, n57856, n57857, n57858, n57859, n57860, n57861, n57862,
    n57863, n57864, n57865, n57866, n57867, n57868, n57869, n57870, n57871,
    n57872, n57873, n57874, n57875, n57876, n57877, n57878, n57879, n57880,
    n57881, n57882, n57883, n57884, n57885, n57886, n57887, n57888, n57889,
    n57890, n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
    n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906, n57907,
    n57908, n57909, n57910, n57911, n57912, n57913, n57914, n57915, n57916,
    n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924, n57925,
    n57926, n57927, n57928, n57929, n57930, n57931, n57932, n57933, n57934,
    n57935, n57936, n57937, n57938, n57939, n57940, n57941, n57942, n57943,
    n57944, n57945, n57946, n57947, n57948, n57949, n57950, n57951, n57952,
    n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961,
    n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
    n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978, n57979,
    n57980, n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988,
    n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997,
    n57998, n57999, n58000, n58001, n58002, n58003, n58004, n58005, n58006,
    n58007, n58008, n58009, n58010, n58011, n58012, n58013, n58014, n58015,
    n58016, n58017, n58018, n58019, n58020, n58021, n58022, n58023, n58024,
    n58025, n58026, n58027, n58028, n58029, n58030, n58031, n58032, n58033,
    n58034, n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042,
    n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050, n58051,
    n58052, n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060,
    n58061, n58062, n58063, n58064, n58065, n58066, n58067, n58068, n58069,
    n58070, n58071, n58072, n58073, n58074, n58075, n58076, n58077, n58078,
    n58079, n58080, n58081, n58082, n58083, n58084, n58085, n58086, n58087,
    n58088, n58089, n58090, n58091, n58092, n58093, n58094, n58095, n58096,
    n58097, n58098, n58099, n58100, n58101, n58102, n58103, n58104, n58105,
    n58106, n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114,
    n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122, n58123,
    n58124, n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132,
    n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140, n58141,
    n58142, n58143, n58144, n58145, n58146, n58147, n58148, n58149, n58150,
    n58151, n58152, n58153, n58154, n58155, n58156, n58157, n58158, n58159,
    n58160, n58161, n58162, n58163, n58164, n58165, n58166, n58167, n58168,
    n58169, n58170, n58171, n58172, n58173, n58174, n58175, n58176, n58177,
    n58178, n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186,
    n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194, n58195,
    n58196, n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204,
    n58205, n58206, n58207, n58208, n58209, n58210, n58211, n58212, n58213,
    n58214, n58215, n58216, n58217, n58218, n58219, n58220, n58221, n58222,
    n58223, n58224, n58225, n58226, n58227, n58228, n58229, n58230, n58231,
    n58232, n58233, n58234, n58235, n58236, n58237, n58238, n58239, n58240,
    n58241, n58242, n58243, n58244, n58245, n58246, n58247, n58248, n58249,
    n58250, n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258,
    n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266, n58267,
    n58268, n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276,
    n58277, n58278, n58279, n58280, n58281, n58282, n58283, n58284, n58285,
    n58286, n58287, n58288, n58289, n58290, n58291, n58292, n58293, n58294,
    n58295, n58296, n58297, n58298, n58299, n58300, n58301, n58302, n58303,
    n58304, n58305, n58306, n58307, n58308, n58309, n58310, n58311, n58312,
    n58313, n58314, n58315, n58316, n58317, n58318, n58319, n58320, n58321,
    n58322, n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330,
    n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338, n58339,
    n58340, n58341, n58342, n58343, n58344, n58345, n58346, n58347, n58348,
    n58349, n58350, n58351, n58352, n58353, n58354, n58355, n58356, n58357,
    n58358, n58359, n58360, n58361, n58362, n58363, n58364, n58365, n58366,
    n58367, n58368, n58369, n58370, n58371, n58372, n58373, n58374, n58375,
    n58376, n58377, n58378, n58379, n58380, n58381, n58382, n58383, n58384,
    n58385, n58386, n58387, n58388, n58389, n58390, n58391, n58392, n58393,
    n58394, n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402,
    n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410, n58411,
    n58412, n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420,
    n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428, n58429,
    n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437, n58438,
    n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446, n58447,
    n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455, n58456,
    n58457, n58458, n58459, n58460, n58461, n58462, n58463, n58464, n58465,
    n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
    n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482, n58483,
    n58484, n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492,
    n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500, n58501,
    n58502, n58503, n58504, n58505, n58506, n58507, n58508, n58509, n58510,
    n58511, n58512, n58513, n58514, n58515, n58516, n58517, n58518, n58519,
    n58520, n58521, n58522, n58523, n58524, n58525, n58526, n58527, n58528,
    n58529, n58530, n58531, n58532, n58533, n58534, n58535, n58536, n58537,
    n58538, n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
    n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554, n58555,
    n58556, n58557, n58558, n58559, n58560, n58561, n58562, n58563, n58564,
    n58565, n58566, n58567, n58568, n58569, n58570, n58571, n58572, n58573,
    n58574, n58575, n58576, n58577, n58578, n58579, n58580, n58581, n58582,
    n58583, n58584, n58585, n58586, n58587, n58588, n58589, n58590, n58591,
    n58592, n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600,
    n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608, n58609,
    n58610, n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618,
    n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626, n58627,
    n58628, n58629, n58630, n58631, n58632, n58633, n58634, n58635, n58636,
    n58637, n58638, n58639, n58640, n58641, n58642, n58643, n58644, n58645,
    n58646, n58647, n58648, n58649, n58650, n58651, n58652, n58653, n58654,
    n58655, n58656, n58657, n58658, n58659, n58660, n58661, n58662, n58663,
    n58664, n58665, n58666, n58667, n58668, n58669, n58670, n58671, n58672,
    n58673, n58674, n58675, n58676, n58677, n58678, n58679, n58680, n58681,
    n58682, n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690,
    n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698, n58699,
    n58700, n58701, n58702, n58703, n58704, n58705, n58706, n58707, n58708,
    n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716, n58717,
    n58718, n58719, n58720, n58721, n58722, n58723, n58724, n58725, n58726,
    n58727, n58728, n58729, n58730, n58731, n58732, n58733, n58734, n58735,
    n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58743, n58744,
    n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752, n58753,
    n58754, n58755, n58756, n58757, n58758, n58759, n58760, n58761, n58762,
    n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770, n58771,
    n58772, n58773, n58774, n58775, n58776, n58777, n58778, n58779, n58780,
    n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788, n58789,
    n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797, n58798,
    n58799, n58800, n58801, n58802, n58803, n58804, n58805, n58806, n58807,
    n58808, n58809, n58810, n58811, n58812, n58813, n58814, n58815, n58816,
    n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824, n58825,
    n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833, n58834,
    n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842, n58843,
    n58844, n58845, n58846, n58847, n58848, n58849, n58850, n58851, n58852,
    n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860, n58861,
    n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869, n58870,
    n58871, n58872, n58873, n58874, n58875, n58876, n58877, n58878, n58879,
    n58880, n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888,
    n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896, n58897,
    n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906,
    n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914, n58915,
    n58916, n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924,
    n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932, n58933,
    n58934, n58935, n58936, n58937, n58938, n58939, n58940, n58941, n58942,
    n58943, n58944, n58945, n58946, n58947, n58948, n58949, n58950, n58951,
    n58952, n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960,
    n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968, n58969,
    n58970, n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978,
    n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986, n58987,
    n58988, n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996,
    n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004, n59005,
    n59006, n59007, n59008, n59009, n59010, n59011, n59012, n59013, n59014,
    n59015, n59016, n59017, n59018, n59019, n59020, n59021, n59022, n59023,
    n59024, n59025, n59026, n59027, n59028, n59029, n59030, n59031, n59032,
    n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040, n59041,
    n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049, n59050,
    n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058, n59059,
    n59060, n59061, n59062, n59063, n59064, n59065, n59066, n59067, n59068,
    n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076, n59077,
    n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085, n59086,
    n59087, n59088, n59089, n59090, n59091, n59092, n59093, n59094, n59095,
    n59096, n59097, n59098, n59099, n59100, n59101, n59102, n59103, n59104,
    n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112, n59113,
    n59114, n59115, n59116, n59117, n59118, n59119, n59120, n59121, n59122,
    n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130, n59131,
    n59132, n59133, n59134, n59135, n59136, n59137, n59138, n59139, n59140,
    n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148, n59149,
    n59150, n59151, n59152, n59153, n59154, n59155, n59156, n59157, n59158,
    n59159, n59160, n59161, n59162, n59163, n59164, n59165, n59166, n59167,
    n59168, n59169, n59170, n59171, n59172, n59173, n59174, n59175, n59176,
    n59177, n59178, n59179, n59180, n59181, n59182, n59183, n59184, n59185,
    n59186, n59187, n59188, n59189, n59190, n59191, n59192, n59193, n59194,
    n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202, n59203,
    n59204, n59205, n59206, n59207, n59208, n59209, n59210, n59211, n59212,
    n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220, n59221,
    n59222, n59223, n59224, n59225, n59226, n59227, n59228, n59229, n59230,
    n59231, n59232, n59233, n59234, n59235, n59236, n59237, n59238, n59239,
    n59240, n59241, n59242, n59243, n59244, n59245, n59246, n59247, n59248,
    n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256, n59257,
    n59258, n59259, n59260, n59261, n59262, n59263, n59264, n59265, n59266,
    n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274, n59275,
    n59276, n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284,
    n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292, n59293,
    n59294, n59295, n59296, n59297, n59298, n59299, n59300, n59301, n59302,
    n59303, n59304, n59305, n59306, n59307, n59308, n59309, n59310, n59311,
    n59312, n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59320,
    n59321, n59322, n59323, n59324, n59325, n59326, n59327, n59328, n59329,
    n59330, n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338,
    n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346, n59347,
    n59348, n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356,
    n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364, n59365,
    n59366, n59367, n59368, n59369, n59370, n59371, n59372, n59373, n59374,
    n59375, n59376, n59377, n59378, n59379, n59380, n59381, n59382, n59383,
    n59384, n59385, n59386, n59387, n59388, n59389, n59390, n59391, n59392,
    n59393, n59394, n59395, n59396, n59397, n59398, n59399, n59400, n59401,
    n59402, n59403, n59404, n59405, n59406, n59407, n59408, n59409, n59410,
    n59411, n59412, n59413, n59414, n59415, n59416, n59417, n59418, n59419,
    n59420, n59421, n59422, n59423, n59424, n59425, n59426, n59427, n59428,
    n59429, n59430, n59431, n59432, n59433, n59434, n59435, n59436, n59437,
    n59438, n59439, n59440, n59441, n59442, n59443, n59444, n59445, n59446,
    n59447, n59448, n59449, n59450, n59451, n59452, n59453, n59454, n59455,
    n59456, n59457, n59458, n59459, n59460, n59461, n59462, n59463, n59464,
    n59465, n59466, n59467, n59468, n59469, n59470, n59471, n59472, n59473,
    n59474, n59475, n59476, n59477, n59478, n59479, n59480, n59481, n59482,
    n59483, n59484, n59485, n59486, n59487, n59488, n59489, n59490, n59491,
    n59492, n59493, n59494, n59495, n59496, n59497, n59498, n59499, n59500,
    n59501, n59502, n59503, n59504, n59505, n59506, n59507, n59508, n59509,
    n59510, n59511, n59512, n59513, n59514, n59515, n59516, n59517, n59518,
    n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526, n59527,
    n59528, n59529, n59530, n59531, n59532, n59533, n59534, n59535, n59536,
    n59537, n59538, n59539, n59540, n59541, n59542, n59543, n59544, n59545,
    n59546, n59547, n59548, n59549, n59550, n59551, n59552, n59553, n59554,
    n59555, n59556, n59557, n59558, n59559, n59560, n59561, n59562, n59563,
    n59564, n59565, n59566, n59567, n59568, n59569, n59570, n59571, n59572,
    n59573, n59574, n59575, n59576, n59577, n59578, n59579, n59580, n59581,
    n59582, n59583, n59584, n59585, n59586, n59587, n59588, n59589, n59590,
    n59591, n59592, n59593, n59594, n59595, n59596, n59597, n59598, n59599,
    n59600, n59601, n59602, n59603, n59604, n59605, n59606, n59607, n59608,
    n59609, n59610, n59611, n59612, n59613, n59614, n59615, n59616, n59617,
    n59618, n59619, n59620, n59621, n59622, n59623, n59624, n59625, n59626,
    n59627, n59628, n59629, n59630, n59631, n59632, n59633, n59634, n59635,
    n59636, n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644,
    n59645, n59646, n59647, n59648, n59649, n59650, n59651, n59652, n59653,
    n59654, n59655, n59656, n59657, n59658, n59659, n59660, n59661, n59662,
    n59663, n59664, n59665, n59666, n59667, n59668, n59669, n59670, n59671,
    n59672, n59673, n59674, n59675, n59676, n59677, n59678, n59679, n59680,
    n59681, n59682, n59683, n59684, n59685, n59686, n59687, n59688, n59689,
    n59690, n59691, n59692, n59693, n59694, n59695, n59696, n59697, n59698,
    n59699, n59700, n59701, n59702, n59703, n59704, n59705, n59706, n59707,
    n59708, n59709, n59710, n59711, n59712, n59713, n59714, n59715, n59716,
    n59717, n59718, n59719, n59720, n59721, n59722, n59723, n59724, n59725,
    n59726, n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734,
    n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742, n59743,
    n59744, n59745, n59746, n59747, n59748, n59749, n59750, n59751, n59752,
    n59753, n59754, n59755, n59756, n59757, n59758, n59759, n59760, n59761,
    n59762, n59763, n59764, n59765, n59766, n59767, n59768, n59769, n59770,
    n59771, n59772, n59773, n59774, n59775, n59776, n59777, n59778, n59779,
    n59780, n59781, n59782, n59783, n59784, n59785, n59786, n59787, n59788,
    n59789, n59790, n59791, n59792, n59793, n59794, n59795, n59796, n59797,
    n59798, n59799, n59800, n59801, n59802, n59803, n59804, n59805, n59806,
    n59807, n59808, n59809, n59810, n59811, n59812, n59813, n59814, n59815,
    n59816, n59817, n59818, n59819, n59820, n59821, n59822, n59823, n59824,
    n59825, n59826, n59827, n59828, n59829, n59830, n59831, n59832, n59833,
    n59834, n59835, n59836, n59837, n59838, n59839, n59840, n59841, n59842,
    n59843, n59844, n59845, n59846, n59847, n59848, n59849, n59850, n59851,
    n59852, n59853, n59854, n59855, n59856, n59857, n59858, n59859, n59860,
    n59861, n59862, n59863, n59864, n59865, n59866, n59867, n59868, n59869,
    n59870, n59871, n59872, n59873, n59874, n59875, n59876, n59877, n59878,
    n59879, n59880, n59881, n59882, n59883, n59884, n59885, n59886, n59887,
    n59888, n59889, n59890, n59891, n59892, n59893, n59894, n59895, n59896,
    n59897, n59898, n59899, n59900, n59901, n59902, n59903, n59904, n59905,
    n59906, n59907, n59908, n59909, n59910, n59911, n59912, n59913, n59914,
    n59915, n59916, n59917, n59918, n59919, n59920, n59921, n59922, n59923,
    n59924, n59925, n59926, n59927, n59928, n59929, n59930, n59931, n59932,
    n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59940, n59941,
    n59942, n59943, n59944, n59945, n59946, n59947, n59948, n59949, n59950,
    n59951, n59952, n59953, n59954, n59955, n59956, n59957, n59958, n59959,
    n59960, n59961, n59962, n59963, n59964, n59965, n59966, n59967, n59968,
    n59969, n59970, n59971, n59972, n59973, n59974, n59975, n59976, n59977,
    n59978, n59979, n59980, n59981, n59982, n59983, n59984, n59985, n59986,
    n59987, n59988, n59989, n59990, n59991, n59992, n59993, n59994, n59995,
    n59996, n59997, n59998, n59999, n60000, n60001, n60002, n60003, n60004,
    n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012, n60013,
    n60014, n60015, n60016, n60017, n60018, n60019, n60020, n60021, n60022,
    n60023, n60024, n60025, n60026, n60027, n60028, n60029, n60030, n60031,
    n60032, n60033, n60034, n60035, n60036, n60037, n60038, n60039, n60040,
    n60041, n60042, n60043, n60044, n60045, n60046, n60047, n60048, n60049,
    n60050, n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058,
    n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066, n60067,
    n60068, n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076,
    n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084, n60085,
    n60086, n60087, n60088, n60089, n60090, n60091, n60092, n60093, n60094,
    n60095, n60096, n60097, n60098, n60099, n60100, n60101, n60102, n60103,
    n60104, n60105, n60106, n60107, n60108, n60109, n60110, n60111, n60112,
    n60113, n60114, n60115, n60116, n60117, n60118, n60119, n60120, n60121,
    n60122, n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130,
    n60131, n60132, n60133, n60134, n60135, n60136, n60137, n60138, n60139,
    n60140, n60141, n60142, n60143, n60144, n60145, n60146, n60147, n60148,
    n60149, n60150, n60151, n60152, n60153, n60154, n60155, n60156, n60157,
    n60158, n60159, n60160, n60161, n60162, n60163, n60164, n60165, n60166,
    n60167, n60168, n60169, n60170, n60171, n60172, n60173, n60174, n60175,
    n60176, n60177, n60178, n60179, n60180, n60181, n60182, n60183, n60184,
    n60185, n60186, n60187, n60188, n60189, n60190, n60191, n60192, n60193,
    n60194, n60195, n60196, n60197, n60198, n60199, n60200, n60201, n60202,
    n60203, n60204, n60205, n60206, n60207, n60208, n60209, n60210, n60211,
    n60212, n60213, n60214, n60215, n60216, n60217, n60218, n60219, n60220,
    n60221, n60222, n60223, n60224, n60225, n60226, n60227, n60228, n60229,
    n60230, n60231, n60232, n60233, n60234, n60235, n60236, n60237, n60238,
    n60239, n60240, n60241, n60242, n60243, n60244, n60245, n60246, n60247,
    n60248, n60249, n60250, n60251, n60252, n60253, n60254, n60255, n60256,
    n60257, n60258, n60259, n60260, n60261, n60262, n60263, n60264, n60265,
    n60266, n60267, n60268, n60269, n60270, n60271, n60272, n60273, n60274,
    n60275, n60276, n60277, n60278, n60279, n60280, n60281, n60282, n60283,
    n60284, n60285, n60286, n60287, n60288, n60289, n60290, n60291, n60292,
    n60293, n60294, n60295, n60296, n60297, n60298, n60299, n60300, n60301,
    n60302, n60303, n60304, n60305, n60306, n60307, n60308, n60309, n60310,
    n60311, n60312, n60313, n60314, n60315, n60316, n60317, n60318, n60319,
    n60320, n60321, n60322, n60323, n60324, n60325, n60326, n60327, n60328,
    n60329, n60330, n60331, n60332, n60333, n60334, n60335, n60336, n60337,
    n60338, n60339, n60340, n60341, n60342, n60343, n60344, n60345, n60346,
    n60347, n60348, n60349, n60350, n60351, n60352, n60353, n60354, n60355,
    n60356, n60357, n60358, n60359, n60360, n60361, n60362, n60363, n60364,
    n60365, n60366, n60367, n60368, n60369, n60370, n60371, n60372, n60373,
    n60374, n60375, n60376, n60377, n60378, n60379, n60380, n60381, n60382,
    n60383, n60384, n60385, n60386, n60387, n60388, n60389, n60390, n60391,
    n60392, n60393, n60394, n60395, n60396, n60397, n60398, n60399, n60400,
    n60401, n60402, n60403, n60404, n60405, n60406, n60407, n60408, n60409,
    n60410, n60411, n60412, n60413, n60414, n60415, n60416, n60417, n60418,
    n60419, n60420, n60421, n60422, n60423, n60424, n60425, n60426, n60427,
    n60428, n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60436,
    n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444, n60445,
    n60446, n60447, n60448, n60449, n60450, n60451, n60452, n60453, n60454,
    n60455, n60456, n60457, n60458, n60459, n60460, n60461, n60462, n60463,
    n60464, n60465, n60466, n60467, n60468, n60469, n60470, n60471, n60472,
    n60473, n60474, n60475, n60476, n60477, n60478, n60479, n60480, n60481,
    n60482, n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490,
    n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498, n60499,
    n60500, n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508,
    n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516, n60517,
    n60518, n60519, n60520, n60521, n60522, n60523, n60524, n60525, n60526,
    n60527, n60528, n60529, n60530, n60531, n60532, n60533, n60534, n60535,
    n60536, n60537, n60538, n60539, n60540, n60541, n60542, n60543, n60544,
    n60545, n60546, n60547, n60548, n60549, n60550, n60551, n60552, n60553,
    n60554, n60555, n60556, n60557, n60558, n60559, n60560, n60561, n60562,
    n60563, n60564, n60565, n60566, n60567, n60568, n60569, n60570, n60571,
    n60572, n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580,
    n60581, n60582, n60583, n60584, n60585, n60586, n60587, n60588, n60589,
    n60590, n60591, n60592, n60593, n60594, n60595, n60596, n60597, n60598,
    n60599, n60600, n60601, n60602, n60603, n60604, n60605, n60606, n60607,
    n60608, n60609, n60610, n60611, n60612, n60613, n60614, n60615, n60616,
    n60617, n60618, n60619, n60620, n60621, n60622, n60623, n60624, n60625,
    n60626, n60627, n60628, n60629, n60630, n60631, n60632, n60633, n60634,
    n60635, n60636, n60637, n60638, n60639, n60640, n60641, n60642, n60643,
    n60644, n60645, n60646, n60647, n60648, n60649, n60650, n60651, n60652,
    n60653, n60654, n60655, n60656, n60657, n60658, n60659, n60660, n60661,
    n60662, n60663, n60664, n60665, n60666, n60667, n60668, n60669, n60670,
    n60671, n60672, n60673, n60674, n60675, n60676, n60677, n60678, n60679,
    n60680, n60681, n60682, n60683, n60684, n60685, n60686, n60687, n60688,
    n60689, n60690, n60691, n60692, n60693, n60694, n60695, n60696, n60697,
    n60698, n60699, n60700, n60701, n60702, n60703, n60704, n60705, n60706,
    n60707, n60708, n60709, n60710, n60711, n60712, n60713, n60714, n60715,
    n60716, n60717, n60718, n60719, n60720, n60721, n60722, n60723, n60724,
    n60725, n60726, n60727, n60728, n60729, n60730, n60731, n60732, n60733,
    n60734, n60735, n60736, n60737, n60738, n60739, n60740, n60741, n60742,
    n60743, n60744, n60745, n60746, n60747, n60748, n60749, n60750, n60751,
    n60752, n60753, n60754, n60755, n60756, n60757, n60758, n60759, n60760,
    n60761, n60762, n60763, n60764, n60765, n60766, n60767, n60768, n60769,
    n60770, n60771, n60772, n60773, n60774, n60775, n60776, n60777, n60778,
    n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786, n60787,
    n60788, n60789, n60790, n60791, n60792, n60793, n60794, n60795, n60796,
    n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60804, n60805,
    n60806, n60807, n60808, n60809, n60810, n60811, n60812, n60813, n60814,
    n60815, n60816, n60817, n60818, n60819, n60820, n60821, n60822, n60823,
    n60824, n60825, n60826, n60827, n60828, n60829, n60830, n60831, n60832,
    n60833, n60834, n60835, n60836, n60837, n60838, n60839, n60840, n60841,
    n60842, n60843, n60844, n60845, n60846, n60847, n60848, n60849, n60850,
    n60851, n60852, n60853, n60854, n60855, n60856, n60857, n60858, n60859,
    n60860, n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868,
    n60869, n60870, n60871, n60872, n60873, n60874, n60875, n60876, n60877,
    n60878, n60879, n60880, n60881, n60882, n60883, n60884, n60885, n60886,
    n60887, n60888, n60889, n60890, n60891, n60892, n60893, n60894, n60895,
    n60896, n60897, n60898, n60899, n60900, n60901, n60902, n60903, n60904,
    n60905, n60906, n60907, n60908, n60909, n60910, n60911, n60912, n60913,
    n60914, n60915, n60916, n60917, n60918, n60919, n60920, n60921, n60922,
    n60923, n60924, n60925, n60926, n60927, n60928, n60929, n60930, n60931,
    n60932, n60933, n60934, n60935, n60936, n60937, n60938, n60939, n60940,
    n60941, n60942, n60943, n60944, n60945, n60946, n60947, n60948, n60949,
    n60950, n60951, n60952, n60953, n60954, n60955, n60956, n60957, n60958,
    n60959, n60960, n60961, n60962, n60963, n60964, n60965, n60966, n60967,
    n60968, n60969, n60970, n60971, n60972, n60973, n60974, n60975, n60976,
    n60977, n60978, n60979, n60980, n60981, n60982, n60983, n60984, n60985,
    n60986, n60987, n60988, n60989, n60990, n60991, n60992, n60993, n60994,
    n60995, n60996, n60997, n60998, n60999, n61000, n61001, n61002, n61003,
    n61004, n61005, n61006, n61007, n61008, n61009, n61010, n61011, n61012,
    n61013, n61014, n61015, n61016, n61017, n61018, n61019, n61020, n61021,
    n61022, n61023, n61024, n61025, n61026, n61027, n61028, n61029, n61030,
    n61031, n61032, n61033, n61034, n61035, n61036, n61037, n61038, n61039,
    n61040, n61041, n61042, n61043, n61044, n61045, n61046, n61047, n61048,
    n61049, n61050, n61051, n61052, n61053, n61054, n61055, n61056, n61057,
    n61058, n61059, n61060, n61061, n61062, n61063, n61064, n61065, n61066,
    n61067, n61068, n61069, n61070, n61071, n61072, n61073, n61074, n61075,
    n61076, n61077, n61078, n61079, n61080, n61081, n61082, n61083, n61084,
    n61085, n61086, n61087, n61088, n61089, n61090, n61091, n61092, n61093,
    n61094, n61095, n61096, n61097, n61098, n61099, n61100, n61101, n61102,
    n61103, n61104, n61105, n61106, n61107, n61108, n61109, n61110, n61111,
    n61112, n61113, n61114, n61115, n61116, n61117, n61118, n61119, n61120,
    n61121, n61122, n61123, n61124, n61125, n61126, n61127, n61128, n61129,
    n61130, n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138,
    n61139, n61140, n61141, n61142, n61143, n61144, n61145, n61146, n61147,
    n61148, n61149, n61150, n61151, n61152, n61153, n61154, n61155, n61156,
    n61157, n61158, n61159, n61160, n61161, n61162, n61163, n61164, n61165,
    n61166, n61167, n61168, n61169, n61170, n61171, n61172, n61173, n61174,
    n61175, n61176, n61177, n61178, n61179, n61180, n61181, n61182, n61183,
    n61184, n61185, n61186, n61187, n61188, n61189, n61190, n61191, n61192,
    n61193, n61194, n61195, n61196, n61197, n61198, n61199, n61200, n61201,
    n61202, n61203, n61204, n61205, n61206, n61207, n61208, n61209, n61210,
    n61211, n61212, n61213, n61214, n61215, n61216, n61217, n61218, n61219,
    n61220, n61221, n61222, n61223, n61224, n61225, n61226, n61227, n61228,
    n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236, n61237,
    n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61245, n61246,
    n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61254, n61255,
    n61256, n61257, n61258, n61259, n61260, n61261, n61262, n61263, n61264,
    n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272, n61273,
    n61274, n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282,
    n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290, n61291,
    n61292, n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300,
    n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308, n61309,
    n61310, n61311, n61312, n61313, n61314, n61315, n61316, n61317, n61318,
    n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326, n61327,
    n61328, n61329, n61330, n61331, n61332, n61333, n61334, n61335, n61336,
    n61337, n61338, n61339, n61340, n61341, n61342, n61343, n61344, n61345,
    n61346, n61347, n61348, n61349, n61350, n61351, n61352, n61353, n61354,
    n61355, n61356, n61357, n61358, n61359, n61360, n61361, n61362, n61363,
    n61364, n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372,
    n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380, n61381,
    n61382, n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390,
    n61391, n61392, n61393, n61394, n61395, n61396, n61397, n61398, n61399,
    n61400, n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408,
    n61409, n61410, n61411, n61412, n61413, n61414, n61415, n61416, n61417,
    n61418, n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426,
    n61427, n61428, n61429, n61430, n61431, n61432, n61433, n61434, n61435,
    n61436, n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444,
    n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452, n61453,
    n61454, n61455, n61456, n61457, n61458, n61459, n61460, n61461, n61462,
    n61463, n61464, n61465, n61466, n61467, n61468, n61469, n61470, n61471,
    n61472, n61473, n61474, n61475, n61476, n61477, n61478, n61479, n61480,
    n61481, n61482, n61483, n61484, n61485, n61486, n61487, n61488, n61489,
    n61490, n61491, n61492, n61493, n61494, n61495, n61496, n61497, n61498,
    n61499, n61500, n61501, n61502, n61503, n61504, n61505, n61506, n61507,
    n61508, n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516,
    n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524, n61525,
    n61526, n61527, n61528, n61529, n61530, n61531, n61532, n61533, n61534,
    n61535, n61536, n61537, n61538, n61539, n61540, n61541, n61542, n61543,
    n61544, n61545, n61546, n61547, n61548, n61549, n61550, n61551, n61552,
    n61553, n61554, n61555, n61556, n61557, n61558, n61559, n61560, n61561,
    n61562, n61563, n61564, n61565, n61566, n61567, n61568, n61569, n61570,
    n61571, n61572, n61573, n61574, n61575, n61576, n61577, n61578, n61579,
    n61580, n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588,
    n61589, n61590, n61591, n61592, n61593, n61594, n61595, n61596, n61597,
    n61598, n61599, n61600, n61601, n61602, n61603, n61604, n61605, n61606,
    n61607, n61608, n61609, n61610, n61611, n61612, n61613, n61614, n61615,
    n61616, n61617, n61618, n61619, n61620, n61621, n61622, n61623, n61624,
    n61625, n61626, n61627, n61628, n61629, n61630, n61631, n61632, n61633,
    n61634, n61635, n61636, n61637, n61638, n61639, n61640, n61641, n61642,
    n61643, n61644, n61645, n61646, n61647, n61648, n61649, n61650, n61651,
    n61652, n61653, n61654, n61655, n61656, n61657, n61658, n61659, n61660,
    n61661, n61662, n61663, n61664, n61665, n61666, n61667, n61668, n61669,
    n61670, n61671, n61672, n61673, n61674, n61675, n61676, n61677, n61678,
    n61679, n61680, n61681, n61682, n61683, n61684, n61685, n61686, n61687,
    n61688, n61689, n61690, n61691, n61692, n61693, n61694, n61695, n61696,
    n61697, n61698, n61699, n61700, n61701, n61702, n61703, n61704, n61705,
    n61706, n61707, n61708, n61709, n61710, n61711, n61712, n61713, n61714,
    n61715, n61716, n61717, n61718, n61719, n61720, n61721, n61722, n61723,
    n61724, n61725, n61726, n61727, n61728, n61729, n61730, n61731, n61732,
    n61733, n61734, n61735, n61736, n61737, n61738, n61739, n61740, n61741,
    n61742, n61743, n61744, n61745, n61746, n61747, n61748, n61749, n61750,
    n61751, n61752, n61753, n61754, n61755, n61756, n61757, n61758, n61759,
    n61760, n61761, n61762, n61763, n61764, n61765, n61766, n61767, n61768,
    n61769, n61770, n61771, n61772, n61773, n61774, n61775, n61776, n61777,
    n61778, n61779, n61780, n61781, n61782, n61783, n61784, n61785, n61786,
    n61787, n61788, n61789, n61790, n61791, n61792, n61793, n61794, n61795,
    n61796, n61797, n61798, n61799, n61800, n61801, n61802, n61803, n61804,
    n61805, n61806, n61807, n61808, n61809, n61810, n61811, n61812, n61813,
    n61814, n61815, n61816, n61817, n61818, n61819, n61820, n61821, n61822,
    n61823, n61824, n61825, n61826, n61827, n61828, n61829, n61830, n61831,
    n61832, n61833, n61834, n61835, n61836, n61837, n61838, n61839, n61840,
    n61841, n61842, n61843, n61844, n61845, n61846, n61847, n61848, n61849,
    n61850, n61851, n61852, n61853, n61854, n61855, n61856, n61857, n61858,
    n61859, n61860, n61861, n61862, n61863, n61864, n61865, n61866, n61867,
    n61868, n61869, n61870, n61871, n61872, n61873, n61874, n61875, n61876,
    n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884, n61885,
    n61886, n61887, n61888, n61889, n61890, n61891, n61892, n61893, n61894,
    n61895, n61896, n61897, n61898, n61899, n61900, n61901, n61902, n61903,
    n61904, n61905, n61906, n61907, n61908, n61909, n61910, n61911, n61912,
    n61913, n61914, n61915, n61916, n61917, n61918, n61919, n61920, n61921,
    n61922, n61923, n61924, n61925, n61926, n61927, n61928, n61929, n61930,
    n61931, n61932, n61933, n61934, n61935, n61936, n61937, n61938, n61939,
    n61940, n61941, n61942, n61943, n61944, n61945, n61946, n61947, n61948,
    n61949, n61950, n61951, n61952, n61953, n61954, n61955, n61956, n61957,
    n61958, n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966,
    n61967, n61968, n61969, n61970, n61971, n61972, n61973, n61974, n61975,
    n61976, n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984,
    n61985, n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993,
    n61994, n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62002,
    n62003, n62004, n62005, n62006, n62007, n62008, n62009, n62010, n62011,
    n62012, n62013, n62014, n62015, n62016, n62017, n62018, n62019, n62020,
    n62021, n62022, n62023, n62024, n62025, n62026, n62027, n62028, n62029,
    n62030, n62031, n62032, n62033, n62034, n62035, n62036, n62037, n62038,
    n62039, n62040, n62041, n62042, n62043, n62044, n62045, n62046, n62047,
    n62048, n62049, n62050, n62051, n62052, n62053, n62054, n62055, n62056,
    n62057, n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065,
    n62066, n62067, n62068, n62069, n62070, n62071, n62072, n62073, n62074,
    n62075, n62076, n62077, n62078, n62079, n62080, n62081, n62082, n62083,
    n62084, n62085, n62086, n62087, n62088, n62089, n62090, n62091, n62092,
    n62093, n62094, n62095, n62096, n62097, n62098, n62099, n62100, n62101,
    n62102, n62103, n62104, n62105, n62106, n62107, n62108, n62109, n62110,
    n62111, n62112, n62113, n62114, n62115, n62116, n62117, n62118, n62119,
    n62120, n62121, n62122, n62123, n62124, n62125, n62126, n62127, n62128,
    n62129, n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137,
    n62138, n62139, n62140, n62141, n62142, n62143, n62144, n62145, n62146,
    n62147, n62148, n62149, n62150, n62151, n62152, n62153, n62154, n62155,
    n62156, n62157, n62158, n62159, n62160, n62161, n62162, n62163, n62164,
    n62165, n62166, n62167, n62168, n62169, n62170, n62171, n62172, n62173,
    n62174, n62175, n62176, n62177, n62178, n62179, n62180, n62181, n62182,
    n62183, n62184, n62185, n62186, n62187, n62188, n62189, n62190, n62191,
    n62192, n62193, n62194, n62195, n62196, n62197, n62198, n62199, n62200,
    n62201, n62202, n62203, n62204, n62205, n62206, n62207, n62208, n62209,
    n62210, n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218,
    n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226, n62227,
    n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235, n62236,
    n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244, n62245,
    n62246, n62247, n62248, n62249, n62250, n62251, n62252, n62253, n62254,
    n62255, n62256, n62257, n62258, n62259, n62260, n62261, n62262, n62263,
    n62264, n62265, n62266, n62267, n62268, n62269, n62270, n62271, n62272,
    n62273, n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281,
    n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290,
    n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299,
    n62300, n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308,
    n62309, n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317,
    n62318, n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326,
    n62327, n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335,
    n62336, n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344,
    n62345, n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353,
    n62354, n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362,
    n62363, n62364, n62365, n62366, n62367, n62368, n62369, n62370, n62371,
    n62372, n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380,
    n62381, n62382, n62383, n62384, n62385, n62386, n62387, n62388, n62389,
    n62390, n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398,
    n62399, n62400, n62401, n62402, n62403, n62404, n62405, n62406, n62407,
    n62408, n62409, n62410, n62411, n62412, n62413, n62414, n62415, n62416,
    n62417, n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425,
    n62426, n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434,
    n62435, n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443,
    n62444, n62445, n62446, n62447, n62448, n62449, n62450, n62451, n62452,
    n62453, n62454, n62455, n62456, n62457, n62458, n62459, n62460, n62461,
    n62462, n62463, n62464, n62465, n62466, n62467, n62468, n62469, n62470,
    n62471, n62472, n62473, n62474, n62475, n62476, n62477, n62478, n62479,
    n62480, n62481, n62482, n62483, n62484, n62485, n62486, n62487, n62488,
    n62489, n62490, n62491, n62492, n62493, n62494, n62495, n62496, n62497,
    n62498, n62499, n62500, n62501, n62502, n62503, n62504, n62505, n62506,
    n62507, n62508, n62509, n62510, n62511, n62512, n62513, n62514, n62515,
    n62516, n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524,
    n62525, n62526, n62527, n62528, n62529, n62530, n62531, n62532, n62533,
    n62534, n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542,
    n62543, n62544, n62545, n62546, n62547, n62548, n62549, n62550, n62551,
    n62552, n62553, n62554, n62555, n62556, n62557, n62558, n62559, n62560,
    n62561, n62562, n62563, n62564, n62565, n62566, n62567, n62568, n62569,
    n62570, n62571, n62572, n62573, n62574, n62575, n62576, n62577, n62578,
    n62579, n62580, n62581, n62582, n62583, n62584, n62585, n62586, n62587,
    n62588, n62589, n62590, n62591, n62592, n62593, n62594, n62595, n62596,
    n62597, n62598, n62599, n62600, n62601, n62602, n62603, n62604, n62605,
    n62606, n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614,
    n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622, n62623,
    n62624, n62625, n62626, n62627, n62628, n62629, n62630, n62631, n62632,
    n62633, n62634, n62635, n62636, n62637, n62638, n62639, n62640, n62641,
    n62642, n62643, n62644, n62645, n62646, n62647, n62648, n62649, n62650,
    n62651, n62652, n62653, n62654, n62655, n62656, n62657, n62658, n62659,
    n62660, n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668,
    n62669, n62670, n62671, n62672, n62673, n62674, n62675, n62676, n62677,
    n62678, n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686,
    n62687, n62688, n62689, n62690, n62691, n62692, n62693, n62694, n62695,
    n62696, n62697, n62698, n62699, n62700, n62701, n62702, n62703, n62704,
    n62705, n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713,
    n62714, n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722,
    n62723, n62724, n62725, n62726, n62727, n62728, n62729, n62730, n62731,
    n62732, n62733, n62734, n62735, n62736, n62737, n62738, n62739, n62740,
    n62741, n62742, n62743, n62744, n62745, n62746, n62747, n62748, n62749,
    n62750, n62751, n62752, n62753, n62754, n62755, n62756, n62757, n62758,
    n62759, n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767,
    n62768, n62769, n62770, n62771, n62772, n62773, n62774, n62775, n62776,
    n62777, n62778, n62779, n62780, n62781, n62782, n62783, n62784, n62785,
    n62786, n62787, n62788, n62789, n62790, n62791, n62792, n62793, n62794,
    n62795, n62796, n62797, n62798, n62799, n62800, n62801, n62802, n62803,
    n62804, n62805, n62806, n62807, n62808, n62809, n62810, n62811, n62812,
    n62813, n62814, n62815, n62816, n62817, n62818, n62819, n62820, n62821,
    n62822, n62823, n62824, n62825, n62826, n62827, n62828, n62829, n62830,
    n62831, n62832, n62833, n62834, n62835, n62836, n62837, n62838, n62839,
    n62840, n62841, n62842, n62843, n62844, n62845, n62846, n62847, n62848,
    n62849, n62850, n62851, n62852, n62853, n62854, n62855, n62856, n62857,
    n62858, n62859, n62860, n62861, n62862, n62863, n62864, n62865, n62866,
    n62867, n62868, n62869, n62870, n62871, n62872, n62873, n62874, n62875,
    n62876, n62877, n62878, n62879, n62880, n62881, n62882, n62883, n62884,
    n62885, n62886, n62887, n62888, n62889, n62890, n62891, n62892, n62893,
    n62894, n62895, n62896, n62897, n62898, n62899, n62900, n62901, n62902,
    n62903, n62904, n62905, n62906, n62907, n62908, n62909, n62910, n62911,
    n62912, n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920,
    n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928, n62929,
    n62930, n62931, n62932, n62933, n62934, n62935, n62936, n62937, n62938,
    n62939, n62940, n62941, n62942, n62943, n62944, n62945, n62946, n62947,
    n62948, n62949, n62950, n62951, n62952, n62953, n62954, n62955, n62956,
    n62957, n62958, n62959, n62960, n62961, n62962, n62963, n62964, n62965,
    n62966, n62967, n62968, n62969, n62970, n62971, n62972, n62973, n62974,
    n62975, n62976, n62977, n62978, n62979, n62980, n62981, n62982, n62983,
    n62984, n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992,
    n62993, n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001,
    n63002, n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010,
    n63011, n63012, n63013, n63014, n63015, n63016, n63017, n63018, n63019,
    n63020, n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028,
    n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036, n63037,
    n63038, n63039, n63040, n63041, n63042, n63043, n63044, n63045, n63046,
    n63047, n63048, n63049, n63050, n63051, n63052, n63053, n63054, n63055,
    n63056, n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064,
    n63065, n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073,
    n63074, n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082,
    n63083, n63084, n63085, n63086, n63087, n63088, n63089, n63090, n63091,
    n63092, n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100,
    n63101, n63102, n63103, n63104, n63105, n63106, n63107, n63108, n63109,
    n63110, n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63118,
    n63119, n63120, n63121, n63122, n63123, n63124, n63125, n63126, n63127,
    n63128, n63129, n63130, n63131, n63132, n63133, n63134, n63135, n63136,
    n63137, n63138, n63139, n63140, n63141, n63142, n63143, n63144, n63145,
    n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153, n63154,
    n63155, n63156, n63157, n63158, n63159, n63160, n63161, n63162, n63163,
    n63164, n63165, n63166, n63167, n63168, n63169, n63170, n63171, n63172,
    n63173, n63174, n63175, n63176, n63177, n63178, n63179, n63180, n63181,
    n63182, n63183, n63184, n63185, n63186, n63187, n63188, n63189, n63190,
    n63191, n63192, n63193, n63194, n63195, n63196, n63197, n63198, n63199,
    n63200, n63201, n63202, n63203, n63204, n63205, n63206, n63207, n63208,
    n63209, n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217,
    n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225, n63226,
    n63227, n63228, n63229, n63230, n63231, n63232, n63233, n63234, n63235,
    n63236, n63237, n63238, n63239, n63240, n63241, n63242, n63243, n63244,
    n63245, n63246, n63247, n63248, n63249, n63250, n63251, n63252, n63253,
    n63254, n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262,
    n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270, n63271,
    n63272, n63273, n63274, n63275, n63276, n63277, n63278, n63279, n63280,
    n63281, n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289,
    n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298,
    n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306, n63307,
    n63308, n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316,
    n63317, n63318, n63319, n63320, n63321, n63322, n63323, n63324, n63325,
    n63326, n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63334,
    n63335, n63336, n63337, n63338, n63339, n63340, n63341, n63342, n63343,
    n63344, n63345, n63346, n63347, n63348, n63349, n63350, n63351, n63352,
    n63353, n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361,
    n63362, n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370,
    n63371, n63372, n63373, n63374, n63375, n63376, n63377, n63378, n63379,
    n63380, n63381, n63382, n63383, n63384, n63385, n63386, n63387, n63388,
    n63389, n63390, n63391, n63392, n63393, n63394, n63395, n63396, n63397,
    n63398, n63399, n63400, n63401, n63402, n63403, n63404, n63405, n63406,
    n63407, n63408, n63409, n63410, n63411, n63412, n63413, n63414, n63415,
    n63416, n63417, n63418, n63419, n63420, n63421, n63422, n63423, n63424,
    n63425, n63426, n63427, n63428, n63429, n63430, n63431, n63432, n63433,
    n63434, n63435, n63436, n63437, n63438, n63439, n63440, n63441, n63442,
    n63443, n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451,
    n63452, n63453, n63454, n63455, n63456, n63457, n63458, n63459, n63460,
    n63461, n63462, n63463, n63464, n63465, n63466, n63467, n63468, n63469,
    n63470, n63471, n63472, n63473, n63474, n63475, n63476, n63477, n63478,
    n63479, n63480, n63481, n63482, n63483, n63484, n63485, n63486, n63487,
    n63488, n63489, n63490, n63491, n63492, n63493, n63494, n63495, n63496,
    n63497, n63498, n63499, n63500, n63501, n63502, n63503, n63504, n63505,
    n63506, n63507, n63508, n63509, n63510, n63511, n63512, n63513, n63514,
    n63515, n63516, n63517, n63518, n63519, n63520, n63521, n63522, n63523,
    n63524, n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532,
    n63533, n63534, n63535, n63536, n63537, n63538, n63539, n63540, n63541,
    n63542, n63543, n63544, n63545, n63546, n63547, n63548, n63549, n63550,
    n63551, n63552, n63553, n63554, n63555, n63556, n63557, n63558, n63559,
    n63560, n63561, n63562, n63563, n63564, n63565, n63566, n63567, n63568,
    n63569, n63570, n63571, n63572, n63573, n63574, n63575, n63576, n63577,
    n63578, n63579, n63580, n63581, n63582, n63583, n63584, n63585, n63586,
    n63587, n63588, n63589, n63590, n63591, n63592, n63593, n63594, n63595,
    n63596, n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604,
    n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612, n63613,
    n63614, n63615, n63616, n63617, n63618, n63619, n63620, n63621, n63622,
    n63623, n63624, n63625, n63626, n63627, n63628, n63629, n63630, n63631,
    n63632, n63633, n63634, n63635, n63636, n63637, n63638, n63639, n63640,
    n63641, n63642, n63643, n63644, n63645, n63646, n63647, n63648, n63649,
    n63650, n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658,
    n63659, n63660, n63661, n63662, n63663, n63664, n63665, n63666, n63667,
    n63668, n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676,
    n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684, n63685,
    n63686, n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694,
    n63695, n63696, n63697, n63698, n63699, n63700, n63701, n63702, n63703,
    n63704, n63705, n63706, n63707, n63708, n63709, n63710, n63711, n63712,
    n63713, n63714, n63715, n63716, n63717, n63718, n63719, n63720, n63721,
    n63722, n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730,
    n63731, n63732, n63733, n63734, n63735, n63736, n63737, n63738, n63739,
    n63740, n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748,
    n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756, n63757,
    n63758, n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766,
    n63767, n63768, n63769, n63770, n63771, n63772, n63773, n63774, n63775,
    n63776, n63777, n63778, n63779, n63780, n63781, n63782, n63783, n63784,
    n63785, n63786, n63787, n63788, n63789, n63790, n63791, n63792, n63793,
    n63794, n63795, n63796, n63797, n63798, n63799, n63800, n63801, n63802,
    n63803, n63804, n63805, n63806, n63807, n63808, n63809, n63810, n63811,
    n63812, n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
    n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828, n63829,
    n63830, n63831, n63832, n63833, n63834, n63835, n63836, n63837, n63838,
    n63839, n63840, n63841, n63842, n63843, n63844, n63845, n63846, n63847,
    n63848, n63849, n63850, n63851, n63852, n63853, n63854, n63855, n63856,
    n63857, n63858, n63859, n63860, n63861, n63862, n63863, n63864, n63865,
    n63866, n63867, n63868, n63869, n63870, n63871, n63872, n63873, n63874,
    n63875, n63876, n63877, n63878, n63879, n63880, n63881, n63882, n63883,
    n63884, n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892,
    n63893, n63894, n63895, n63896, n63897, n63898, n63899, n63900, n63901,
    n63902, n63903, n63904, n63905, n63906, n63907, n63908, n63909, n63910,
    n63911, n63912, n63913, n63914, n63915, n63916, n63917, n63918, n63919,
    n63920, n63921, n63922, n63923, n63924, n63925, n63926, n63927, n63928,
    n63929, n63930, n63931, n63932, n63933, n63934, n63935, n63936, n63937,
    n63938, n63939, n63940, n63941, n63942, n63943, n63944, n63945, n63946,
    n63947, n63948, n63949, n63950, n63951, n63952, n63953, n63954, n63955,
    n63956, n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964,
    n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972, n63973,
    n63974, n63975, n63976, n63977, n63978, n63979, n63980, n63981, n63982,
    n63983, n63984, n63985, n63986, n63987, n63988, n63989, n63990, n63991,
    n63992, n63993, n63994, n63995, n63996, n63997, n63998, n63999, n64000,
    n64001, n64002, n64003, n64004, n64005, n64006, n64007, n64008, n64009,
    n64010, n64011, n64012, n64013, n64014, n64015, n64016, n64017, n64018,
    n64019, n64020, n64021, n64022, n64023, n64024, n64025, n64026, n64027,
    n64028, n64029, n64030, n64031, n64032, n64033, n64034, n64035, n64036,
    n64037, n64038, n64039, n64040, n64041, n64042, n64043, n64044, n64045,
    n64046, n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054,
    n64055, n64056, n64057, n64058, n64059, n64060, n64061, n64062, n64063,
    n64064, n64065, n64066, n64067, n64068, n64069, n64070, n64071, n64072,
    n64073, n64074, n64075, n64076, n64077, n64078, n64079, n64080, n64081,
    n64082, n64083, n64084, n64085, n64086, n64087, n64088, n64089, n64090,
    n64091, n64092, n64093, n64094, n64095, n64096, n64097, n64098, n64099,
    n64100, n64101, n64102, n64103, n64104, n64105, n64106, n64107, n64108,
    n64109, n64110, n64111, n64112, n64113, n64114, n64115, n64116, n64117,
    n64118, n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64126,
    n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134, n64135,
    n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143, n64144,
    n64145, n64146, n64147, n64148, n64149, n64150, n64151, n64152, n64153,
    n64154, n64155, n64156, n64157, n64158, n64159, n64160, n64161, n64162,
    n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170, n64171,
    n64172, n64173, n64174, n64175, n64176, n64177, n64178, n64179, n64180,
    n64181, n64182, n64183, n64184, n64185, n64186, n64187, n64188, n64189,
    n64190, n64191, n64192, n64193, n64194, n64195, n64196, n64197, n64198,
    n64199, n64200, n64201, n64202, n64203, n64204, n64205, n64206, n64207,
    n64208, n64209, n64210, n64211, n64212, n64213, n64214, n64215, n64216,
    n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224, n64225,
    n64226, n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234,
    n64235, n64236, n64237, n64238, n64239, n64240, n64241, n64242, n64243,
    n64244, n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252,
    n64253, n64254, n64255, n64256, n64257, n64258, n64259, n64260, n64261,
    n64262, n64263, n64264, n64265, n64266, n64267, n64268, n64269, n64270,
    n64271, n64272, n64273, n64274, n64275, n64276, n64277, n64278, n64279,
    n64280, n64281, n64282, n64283, n64284, n64285, n64286, n64287, n64288,
    n64289, n64290, n64291, n64292, n64293, n64294, n64295, n64296, n64297,
    n64298, n64299, n64300, n64301, n64302, n64303, n64304, n64305, n64306,
    n64307, n64308, n64309, n64310, n64311, n64312, n64313, n64314, n64315,
    n64316, n64317, n64318, n64319, n64320, n64321, n64322, n64323, n64324,
    n64325, n64326, n64327, n64328, n64329, n64330, n64331, n64332, n64333,
    n64334, n64335, n64336, n64337, n64338, n64339, n64340, n64341, n64342,
    n64343, n64344, n64345, n64346, n64347, n64348, n64349, n64350, n64351,
    n64352, n64353, n64354, n64355, n64356, n64357, n64358, n64359, n64360,
    n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368, n64369,
    n64370, n64371, n64372, n64373, n64374, n64375, n64376, n64377, n64378,
    n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386, n64387,
    n64388, n64389, n64390, n64391, n64392, n64393, n64394, n64395, n64396,
    n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404, n64405,
    n64406, n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414,
    n64415, n64416, n64417, n64418, n64419, n64420, n64421, n64422, n64423,
    n64424, n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432,
    n64433, n64434, n64435, n64436, n64437, n64438, n64439, n64440, n64441,
    n64442, n64443, n64444, n64445, n64446, n64447, n64448, n64449, n64450,
    n64451, n64452, n64453, n64454, n64455, n64456, n64457, n64458, n64459,
    n64460, n64461, n64462, n64463, n64464, n64465, n64466, n64467, n64468,
    n64469, n64470, n64471, n64472, n64473, n64474, n64475, n64476, n64477,
    n64478, n64479, n64480, n64481, n64482, n64483, n64484, n64485, n64486,
    n64487, n64488, n64489, n64490, n64491, n64492, n64493, n64494, n64495,
    n64496, n64497, n64498, n64499, n64500, n64501, n64502, n64503, n64504,
    n64505, n64506, n64507, n64508, n64509, n64510, n64511, n64512, n64513,
    n64514, n64515, n64516, n64517, n64518, n64519, n64520, n64521, n64522,
    n64523, n64524, n64525, n64526, n64527, n64528, n64529, n64530, n64531,
    n64532, n64533, n64534, n64535, n64536, n64537, n64538, n64539, n64540,
    n64541, n64542, n64543, n64544, n64545, n64546, n64547, n64548, n64549,
    n64550, n64551, n64552, n64553, n64554, n64555, n64556, n64557, n64558,
    n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566, n64567,
    n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64575, n64576,
    n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64584, n64585,
    n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593, n64594,
    n64595, n64596, n64597, n64598, n64599, n64600, n64601, n64602, n64603,
    n64604, n64605, n64606, n64607, n64608, n64609, n64610, n64611, n64612,
    n64613, n64614, n64615, n64616, n64617, n64618, n64619, n64620, n64621,
    n64622, n64623, n64624, n64625, n64626, n64627, n64628, n64629, n64630,
    n64631, n64632, n64633, n64634, n64635, n64636, n64637, n64638, n64639,
    n64640, n64641, n64642, n64643, n64644, n64645, n64646, n64647, n64648,
    n64649, n64650, n64651, n64652, n64653, n64654, n64655, n64656, n64657,
    n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665, n64666,
    n64667, n64668, n64669, n64670, n64671, n64672, n64673, n64674, n64675,
    n64676, n64677, n64678, n64679, n64680, n64681, n64682, n64683, n64684,
    n64685, n64686, n64687, n64688, n64689, n64690, n64691, n64692, n64693,
    n64694, n64695, n64696, n64697, n64698, n64699, n64700, n64701, n64702,
    n64703, n64704, n64705, n64706, n64707, n64708, n64709, n64710, n64711,
    n64712, n64713, n64714, n64715, n64716, n64717, n64718, n64719, n64720,
    n64721, n64722, n64723, n64724, n64725, n64726, n64727, n64728, n64729,
    n64730, n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738,
    n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746, n64747,
    n64748, n64749, n64750, n64751, n64752, n64753, n64754, n64755, n64756,
    n64757, n64758, n64759, n64760, n64761, n64762, n64763, n64764, n64765,
    n64766, n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774,
    n64775, n64776, n64777, n64778, n64779, n64780, n64781, n64782, n64783,
    n64784, n64785, n64786, n64787, n64788, n64789, n64790, n64791, n64792,
    n64793, n64794, n64795, n64796, n64797, n64798, n64799, n64800, n64801,
    n64802, n64803, n64804, n64805, n64806, n64807, n64808, n64809, n64810,
    n64811, n64812, n64813, n64814, n64815, n64816, n64817, n64818, n64819,
    n64820, n64821, n64822, n64823, n64824, n64825, n64826, n64827, n64828,
    n64829, n64830, n64831, n64832, n64833, n64834, n64835, n64836, n64837,
    n64838, n64839, n64840, n64841, n64842, n64843, n64844, n64845, n64846,
    n64847, n64848, n64849, n64850, n64851, n64852, n64853, n64854, n64855,
    n64856, n64857, n64858, n64859, n64860, n64861, n64862, n64863, n64864,
    n64865, n64866, n64867, n64868, n64869, n64870, n64871, n64872, n64873,
    n64874, n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882,
    n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890, n64891,
    n64892, n64893, n64894, n64895, n64896, n64897, n64898, n64899, n64900,
    n64901, n64902, n64903, n64904, n64905, n64906, n64907, n64908, n64909,
    n64910, n64911, n64912, n64913, n64914, n64915, n64916, n64917, n64918,
    n64919, n64920, n64921, n64922, n64923, n64924, n64925, n64926, n64927,
    n64928, n64929, n64930, n64931, n64932, n64933, n64934, n64935, n64936,
    n64937, n64938, n64939, n64940, n64941, n64942, n64943, n64944, n64945,
    n64946, n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954,
    n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962, n64963,
    n64964, n64965, n64966, n64967, n64968, n64969, n64970, n64971, n64972,
    n64973, n64974, n64975, n64976, n64977, n64978, n64979, n64980, n64981,
    n64982, n64983, n64984, n64985, n64986, n64987, n64988, n64989, n64990,
    n64991, n64992, n64993, n64994, n64995, n64996, n64997, n64998, n64999,
    n65000, n65001, n65002, n65003, n65004, n65005, n65006, n65007, n65008,
    n65009, n65010, n65011, n65012, n65013, n65014, n65015, n65016, n65017,
    n65018, n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026,
    n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034, n65035,
    n65036, n65037, n65038, n65039, n65040, n65041, n65042, n65043, n65044,
    n65045, n65046, n65047, n65048, n65049, n65050, n65051, n65052, n65053,
    n65054, n65055, n65056, n65057, n65058, n65059, n65060, n65061, n65062,
    n65063, n65064, n65065, n65066, n65067, n65068, n65069, n65070, n65071,
    n65072, n65073, n65074, n65075, n65076, n65077, n65078, n65079, n65080,
    n65081, n65082, n65083, n65084, n65085, n65086, n65087, n65088, n65089,
    n65090, n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098,
    n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106, n65107,
    n65108, n65109, n65110, n65111, n65112, n65113, n65114, n65115, n65116,
    n65117, n65118, n65119, n65120, n65121, n65122, n65123, n65124, n65125,
    n65126, n65127, n65128, n65129, n65130, n65131, n65132, n65133, n65134,
    n65135, n65136, n65137, n65138, n65139, n65140, n65141, n65142, n65143,
    n65144, n65145, n65146, n65147, n65148, n65149, n65150, n65151, n65152,
    n65153, n65154, n65155, n65156, n65157, n65158, n65159, n65160, n65161,
    n65162, n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170,
    n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178, n65179,
    n65180, n65181, n65182, n65183, n65184, n65185, n65186, n65187, n65188,
    n65189, n65190, n65191, n65192, n65193, n65194, n65195, n65196, n65197,
    n65198, n65199, n65200, n65201, n65202, n65203, n65204, n65205, n65206,
    n65207, n65208, n65209, n65210, n65211, n65212, n65213, n65214, n65215,
    n65216, n65217, n65218, n65219, n65220, n65221, n65222, n65223, n65224,
    n65225, n65226, n65227, n65228, n65229, n65230, n65231, n65232, n65233,
    n65234, n65235, n65236, n65237, n65238, n65239, n65240, n65241, n65242,
    n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250, n65251,
    n65252, n65253, n65254, n65255, n65256, n65257, n65258, n65259, n65260,
    n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268, n65269,
    n65270, n65271, n65272, n65273, n65274, n65275, n65276, n65277, n65278,
    n65279, n65280, n65281, n65282, n65283, n65284, n65285, n65286, n65287,
    n65288, n65289, n65290, n65291, n65292, n65293, n65294, n65295, n65296,
    n65297, n65298, n65299, n65300, n65301, n65302, n65303, n65304, n65305,
    n65306, n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314,
    n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322, n65323,
    n65324, n65325, n65326, n65327, n65328, n65329, n65330, n65331, n65332,
    n65333, n65334, n65335, n65336, n65337, n65338, n65339, n65340, n65341,
    n65342, n65343, n65344, n65345, n65346, n65347, n65348, n65349, n65350,
    n65351, n65352, n65353, n65354, n65355, n65356, n65357, n65358, n65359,
    n65360, n65361, n65362, n65363, n65364, n65365, n65366, n65367, n65368,
    n65369, n65370, n65371, n65372, n65373, n65374, n65375, n65376, n65377,
    n65378, n65379, n65380, n65381, n65382, n65383, n65384, n65385, n65386,
    n65387, n65388, n65389, n65390, n65391, n65392, n65393, n65394, n65395,
    n65396, n65397, n65398, n65399, n65400, n65401, n65402, n65403, n65404,
    n65405, n65406, n65407, n65408, n65409, n65410, n65411, n65412, n65413,
    n65414, n65415, n65416, n65417, n65418, n65419, n65420, n65421, n65422,
    n65423, n65424, n65425, n65426, n65427, n65428, n65429, n65430, n65431,
    n65432, n65433, n65434, n65435, n65436, n65437, n65438, n65439, n65440,
    n65441, n65442, n65443, n65444, n65445, n65446, n65447, n65448, n65449,
    n65450, n65451, n65452, n65453, n65454, n65455, n65456, n65457, n65458,
    n65459, n65460, n65461, n65462, n65463, n65464, n65465, n65466, n65467,
    n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475, n65476,
    n65477, n65478, n65479, n65480, n65481, n65482, n65483, n65484, n65485,
    n65486, n65487, n65488, n65489, n65490, n65491, n65492, n65493, n65494,
    n65495, n65496, n65497, n65498, n65499, n65500, n65501, n65502, n65503,
    n65504, n65505, n65506, n65507, n65508, n65509, n65510, n65511, n65512,
    n65513, n65514, n65515, n65516, n65517, n65518, n65519, n65520, n65521,
    n65522, n65523, n65524, n65525, n65526, n65527, n65528, n65529, n65530,
    n65531, n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539,
    n65540, n65541, n65542, n65543, n65544, n65545, n65546, n65547, n65548,
    n65549, n65550, n65551, n65552, n65553, n65554, n65555, n65556, n65557,
    n65558, n65559, n65560, n65561, n65562, n65563, n65564, n65565, n65566,
    n65567, n65568, n65569, n65570, n65571, n65572, n65573, n65574, n65575,
    n65576, n65577, n65578, n65579, n65580, n65581, n65582, n65583, n65584,
    n65585, n65586, n65587, n65588, n65589, n65590, n65591, n65592, n65593,
    n65594, n65595, n65596, n65597, n65598, n65599, n65600, n65601, n65602,
    n65603, n65604, n65605, n65606, n65607, n65608, n65609, n65610, n65611,
    n65612, n65613, n65614, n65615, n65616, n65617, n65618, n65619, n65620,
    n65621, n65622, n65623, n65624, n65625, n65626, n65627, n65628, n65629,
    n65630, n65631, n65632, n65633, n65634, n65635, n65636, n65637, n65638,
    n65639, n65640, n65641, n65642, n65643, n65644, n65645, n65646, n65647,
    n65648, n65649, n65650, n65651, n65652, n65653, n65654, n65655, n65656,
    n65657, n65658, n65659, n65660, n65661, n65662, n65663, n65664, n65665,
    n65666, n65667, n65668, n65669, n65670, n65671, n65672, n65673, n65674,
    n65675, n65676, n65677, n65678, n65679, n65680, n65681, n65682, n65683,
    n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691, n65692,
    n65693, n65694, n65695, n65696, n65697, n65698, n65699, n65700, n65701,
    n65702, n65703, n65704, n65705, n65706, n65707, n65708, n65709, n65710,
    n65711, n65712, n65713, n65714, n65715, n65716, n65717, n65718, n65719,
    n65720, n65721, n65722, n65723, n65724, n65725, n65726, n65727, n65728,
    n65729, n65730, n65731, n65732, n65733, n65734, n65735, n65736, n65737,
    n65738, n65739, n65740, n65741, n65742, n65743, n65744, n65745, n65746,
    n65747, n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755,
    n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763, n65764,
    n65765, n65766, n65767, n65768, n65769, n65770, n65771, n65772, n65773,
    n65774, n65775, n65776, n65777, n65778, n65779, n65780, n65781, n65782,
    n65783, n65784, n65785, n65786, n65787, n65788, n65789, n65790, n65791,
    n65792, n65793, n65794, n65795, n65796, n65797, n65798, n65799, n65800,
    n65801, n65802, n65803, n65804, n65805, n65806, n65807, n65808, n65809,
    n65810, n65811, n65812, n65813, n65814, n65815, n65816, n65817, n65818,
    n65819, n65820, n65821, n65822, n65823, n65824, n65825, n65826, n65827,
    n65828, n65829, n65830, n65831, n65832, n65833, n65834, n65835, n65836,
    n65837, n65838, n65839, n65840, n65841, n65842, n65843, n65844, n65845,
    n65846, n65847, n65848, n65849, n65850, n65851, n65852, n65853, n65854,
    n65855, n65856, n65857, n65858, n65859, n65860, n65861, n65862, n65863,
    n65864, n65865, n65866, n65867, n65868, n65869, n65870, n65871, n65872,
    n65873, n65874, n65875, n65876, n65877, n65878, n65879, n65880, n65881,
    n65882, n65883, n65884, n65885, n65886, n65887, n65888, n65889, n65890,
    n65891, n65892, n65893, n65894, n65895, n65896, n65897, n65898, n65899,
    n65900, n65901, n65902, n65903, n65904, n65905, n65906, n65907, n65908,
    n65909, n65910, n65911, n65912, n65913, n65914, n65915, n65916, n65917,
    n65918, n65919, n65920, n65921, n65922, n65923, n65924, n65925, n65926,
    n65927, n65928, n65929, n65930, n65931, n65932, n65933, n65934, n65935,
    n65936, n65937, n65938, n65939, n65940, n65941, n65942, n65943, n65944,
    n65945, n65946, n65947, n65948, n65949, n65950, n65951, n65952, n65953,
    n65954, n65955, n65956, n65957, n65958, n65959, n65960, n65961, n65962,
    n65963, n65964, n65965, n65966, n65967, n65968, n65969, n65970, n65971,
    n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979, n65980,
    n65981, n65982, n65983, n65984, n65985, n65986, n65987, n65988, n65989,
    n65990, n65991, n65992, n65993, n65994, n65995, n65996, n65997, n65998,
    n65999, n66000, n66001, n66002, n66003, n66004, n66005, n66006, n66007,
    n66008, n66009, n66010, n66011, n66012, n66013, n66014, n66015, n66016,
    n66017, n66018, n66019, n66020, n66021, n66022, n66023, n66024, n66025,
    n66026, n66027, n66028, n66029, n66030, n66031, n66032, n66033, n66034,
    n66035, n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043,
    n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051, n66052,
    n66053, n66054, n66055, n66056, n66057, n66058, n66059, n66060, n66061,
    n66062, n66063, n66064, n66065, n66066, n66067, n66068, n66069, n66070,
    n66071, n66072, n66073, n66074, n66075, n66076, n66077, n66078, n66079,
    n66080, n66081, n66082, n66083, n66084, n66085, n66086, n66087, n66088,
    n66089, n66090, n66091, n66092, n66093, n66094, n66095, n66096, n66097,
    n66098, n66099, n66100, n66101, n66102, n66103, n66104, n66105, n66106,
    n66107, n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115,
    n66116, n66117, n66118, n66119, n66120, n66121, n66122, n66123, n66124,
    n66125, n66126, n66127, n66128, n66129, n66130, n66131, n66132, n66133,
    n66134, n66135, n66136, n66137, n66138, n66139, n66140, n66141, n66142,
    n66143, n66144, n66145, n66146, n66147, n66148, n66149, n66150, n66151,
    n66152, n66153, n66154, n66155, n66156, n66157, n66158, n66159, n66160,
    n66161, n66162, n66163, n66164, n66165, n66166, n66167, n66168, n66169,
    n66170, n66171, n66172, n66173, n66174, n66175, n66176, n66177, n66178,
    n66179, n66180, n66181, n66182, n66183, n66184, n66185, n66186, n66187,
    n66188, n66189, n66190, n66191, n66192, n66193, n66194, n66195, n66196,
    n66197, n66198, n66199, n66200, n66201, n66202, n66203, n66204, n66205,
    n66206, n66207, n66208, n66209, n66210, n66211, n66212, n66213, n66214,
    n66215, n66216, n66217, n66218, n66219, n66220, n66221, n66222, n66223,
    n66224, n66225, n66226, n66227, n66228, n66229, n66230, n66231, n66232,
    n66233, n66234, n66235, n66236, n66237, n66238, n66239, n66240, n66241,
    n66242, n66243, n66244, n66245, n66246, n66247, n66248, n66249, n66250,
    n66251, n66252, n66253, n66254, n66255, n66256, n66257, n66258, n66259,
    n66260, n66261, n66262, n66263, n66264, n66265, n66266, n66267, n66268,
    n66269, n66270, n66271, n66272, n66273, n66274, n66275, n66276, n66277,
    n66278, n66279, n66280, n66281, n66282, n66283, n66284, n66285, n66286,
    n66287, n66288, n66289, n66290, n66291, n66292, n66293, n66294, n66295,
    n66296, n66297, n66298, n66299, n66300, n66301, n66302, n66303, n66304,
    n66305, n66306, n66307, n66308, n66309, n66310, n66311, n66312, n66313,
    n66314, n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66322,
    n66323, n66324, n66325, n66326, n66327, n66328, n66329, n66330, n66331,
    n66332, n66333, n66334, n66335, n66336, n66337, n66338, n66339, n66340,
    n66341, n66342, n66343, n66344, n66345, n66346, n66347, n66348, n66349,
    n66350, n66351, n66352, n66353, n66354, n66355, n66356, n66357, n66358,
    n66359, n66360, n66361, n66362, n66363, n66364, n66365, n66366, n66367,
    n66368, n66369, n66370, n66371, n66372, n66373, n66374, n66375, n66376,
    n66377, n66378, n66379, n66380, n66381, n66382, n66383, n66384, n66385,
    n66386, n66387, n66388, n66389, n66390, n66391, n66392, n66393, n66394,
    n66395, n66396, n66397, n66398, n66399, n66400, n66401, n66402, n66403,
    n66404, n66405, n66406, n66407, n66408, n66409, n66410, n66411, n66412,
    n66413, n66414, n66415, n66416, n66417, n66418, n66419, n66420, n66421,
    n66422, n66423, n66424, n66425, n66426, n66427, n66428, n66429, n66430,
    n66431, n66432, n66433, n66434, n66435, n66436, n66437, n66438, n66439,
    n66440, n66441, n66442, n66443, n66444, n66445, n66446, n66447, n66448,
    n66449, n66450, n66451, n66452, n66453, n66454, n66455, n66456, n66457,
    n66458, n66459, n66460, n66461, n66462, n66463, n66464, n66465, n66466,
    n66467, n66468, n66469, n66470, n66471, n66472, n66473, n66474, n66475,
    n66476, n66477, n66478, n66479, n66480, n66481, n66482, n66483, n66484,
    n66485, n66486, n66487, n66488, n66489, n66490, n66491, n66492, n66493,
    n66494, n66495, n66496, n66497, n66498, n66499, n66500, n66501, n66502,
    n66503, n66504, n66505, n66506, n66507, n66508, n66509, n66510, n66511,
    n66512, n66513, n66514, n66515, n66516, n66517, n66518, n66519, n66520,
    n66521, n66522, n66523, n66524, n66525, n66526, n66527, n66528, n66529,
    n66530, n66531, n66532, n66533, n66534, n66535, n66536, n66537, n66538,
    n66539, n66540, n66541, n66542, n66543, n66544, n66545, n66546, n66547,
    n66548, n66549, n66550, n66551, n66552, n66553, n66554, n66555, n66556,
    n66557, n66558, n66559, n66560, n66561, n66562, n66563, n66564, n66565,
    n66566, n66567, n66568, n66569, n66570, n66571, n66572, n66573, n66574,
    n66575, n66576, n66577, n66578, n66579, n66580, n66581, n66582, n66583,
    n66584, n66585, n66586, n66587, n66588, n66589, n66590, n66591, n66592,
    n66593, n66594, n66595, n66596, n66597, n66598, n66599, n66600, n66601,
    n66602, n66603, n66604, n66605, n66606, n66607, n66608, n66609, n66610,
    n66611, n66612, n66613, n66614, n66615, n66616, n66617, n66618, n66619,
    n66620, n66621, n66622, n66623, n66624, n66625, n66626, n66627, n66628,
    n66629, n66630, n66631, n66632, n66633, n66634, n66635, n66636, n66637,
    n66638, n66639, n66640, n66641, n66642, n66643, n66644, n66645, n66646,
    n66647, n66648, n66649, n66650, n66651, n66652, n66653, n66654, n66655,
    n66656, n66657, n66658, n66659, n66660, n66661, n66662, n66663, n66664,
    n66665, n66666, n66667, n66668, n66669, n66670, n66671, n66672, n66673,
    n66674, n66675, n66676, n66677, n66678, n66679, n66680, n66681, n66682,
    n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690, n66691,
    n66692, n66693, n66694, n66695, n66696, n66697, n66698, n66699, n66700,
    n66701, n66702, n66703, n66704, n66705, n66706, n66707, n66708, n66709,
    n66710, n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718,
    n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726, n66727,
    n66728, n66729, n66730, n66731, n66732, n66733, n66734, n66735, n66736,
    n66737, n66738, n66739, n66740, n66741, n66742, n66743, n66744, n66745,
    n66746, n66747, n66748, n66749, n66750, n66751, n66752, n66753, n66754,
    n66755, n66756, n66757, n66758, n66759, n66760, n66761, n66762, n66763,
    n66764, n66765, n66766, n66767, n66768, n66769, n66770, n66771, n66772,
    n66773, n66774, n66775, n66776, n66777, n66778, n66779, n66780, n66781,
    n66782, n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790,
    n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798, n66799,
    n66800, n66801, n66802, n66803, n66804, n66805, n66806, n66807, n66808,
    n66809, n66810, n66811, n66812, n66813, n66814, n66815, n66816, n66817,
    n66818, n66819, n66820, n66821, n66822, n66823, n66824, n66825, n66826,
    n66827, n66828, n66829, n66830, n66831, n66832, n66833, n66834, n66835,
    n66836, n66837, n66838, n66839, n66840, n66841, n66842, n66843, n66844,
    n66845, n66846, n66847, n66848, n66849, n66850, n66851, n66852, n66853,
    n66854, n66855, n66856, n66857, n66858, n66859, n66860, n66861, n66862,
    n66863, n66864, n66865, n66866, n66867, n66868, n66869, n66870, n66871,
    n66872, n66873, n66874, n66875, n66876, n66877, n66878, n66879, n66880,
    n66881, n66882, n66883, n66884, n66885, n66886, n66887, n66888, n66889,
    n66890, n66891, n66892, n66893, n66894, n66895, n66896, n66897, n66898,
    n66899, n66900, n66901, n66902, n66903, n66904, n66905, n66906, n66907,
    n66908, n66909, n66910, n66911, n66912, n66913, n66914, n66915, n66916,
    n66917, n66918, n66919, n66920, n66921, n66922, n66923, n66924, n66925,
    n66926, n66927, n66928, n66929, n66930, n66931, n66932, n66933, n66934,
    n66935, n66936, n66937, n66938, n66939, n66940, n66941, n66942, n66943,
    n66944, n66945, n66946, n66947, n66948, n66949, n66950, n66951, n66952,
    n66953, n66954, n66955, n66956, n66957, n66958, n66959, n66960, n66961,
    n66962, n66963, n66964, n66965, n66966, n66967, n66968, n66969, n66970,
    n66971, n66972, n66973, n66974, n66975, n66976, n66977, n66978, n66979,
    n66980, n66981, n66982, n66983, n66984, n66985, n66986, n66987, n66988,
    n66989, n66990, n66991, n66992, n66993, n66994, n66995, n66996, n66997,
    n66998, n66999, n67000, n67001, n67002, n67003, n67004, n67005, n67006,
    n67007, n67008, n67009, n67010, n67011, n67012, n67013, n67014, n67015,
    n67016, n67017, n67018, n67019, n67020, n67021, n67022, n67023, n67024,
    n67025, n67026, n67027, n67028, n67029, n67030, n67031, n67032, n67033,
    n67034, n67035, n67036, n67037, n67038, n67039, n67040, n67041, n67042,
    n67043, n67044, n67045, n67046, n67047, n67048, n67049, n67050, n67051,
    n67052, n67053, n67054, n67055, n67056, n67057, n67058, n67059, n67060,
    n67061, n67062, n67063, n67064, n67065, n67066, n67067, n67068, n67069,
    n67070, n67071, n67072, n67073, n67074, n67075, n67076, n67077, n67078,
    n67079, n67080, n67081, n67082, n67083, n67084, n67085, n67086, n67087,
    n67088, n67089, n67090, n67091, n67092, n67093, n67094, n67095, n67096,
    n67097, n67098, n67099, n67100, n67101, n67102, n67103, n67104, n67105,
    n67106, n67107, n67108, n67109, n67110, n67111, n67112, n67113, n67114,
    n67115, n67116, n67117, n67118, n67119, n67120, n67121, n67122, n67123,
    n67124, n67125, n67126, n67127, n67128, n67129, n67130, n67131, n67132,
    n67133, n67134, n67135, n67136, n67137, n67138, n67139, n67140, n67141,
    n67142, n67143, n67144, n67145, n67146, n67147, n67148, n67149, n67150,
    n67151, n67152, n67153, n67154, n67155, n67156, n67157, n67158, n67159,
    n67160, n67161, n67162, n67163, n67164, n67165, n67166, n67167, n67168,
    n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176, n67177,
    n67178, n67179, n67180, n67181, n67182, n67183, n67184, n67185, n67186,
    n67187, n67188, n67189, n67190, n67191, n67192, n67193, n67194, n67195,
    n67196, n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204,
    n67205, n67206, n67207, n67208, n67209, n67210, n67211, n67212, n67213,
    n67214, n67215, n67216, n67217, n67218, n67219, n67220, n67221, n67222,
    n67223, n67224, n67225, n67226, n67227, n67228, n67229, n67230, n67231,
    n67232, n67233, n67234, n67235, n67236, n67237, n67238, n67239, n67240,
    n67241, n67242, n67243, n67244, n67245, n67246, n67247, n67248, n67249,
    n67250, n67251, n67252, n67253, n67254, n67255, n67256, n67257, n67258,
    n67259, n67260, n67261, n67262, n67263, n67264, n67265, n67266, n67267,
    n67268, n67269, n67270, n67271, n67272, n67273, n67274, n67275, n67276,
    n67277, n67278, n67279, n67280, n67281, n67282, n67283, n67284, n67285,
    n67286, n67287, n67288, n67289, n67290, n67291, n67292, n67293, n67294,
    n67295, n67296, n67297, n67298, n67299, n67300, n67301, n67302, n67303,
    n67304, n67305, n67306, n67307, n67308, n67309, n67310, n67311, n67312,
    n67313, n67314, n67315, n67316, n67317, n67318, n67319, n67320, n67321,
    n67322, n67323, n67324, n67325, n67326, n67327, n67328, n67329, n67330,
    n67331, n67332, n67333, n67334, n67335, n67336, n67337, n67338, n67339,
    n67340, n67341, n67342, n67343, n67344, n67345, n67346, n67347, n67348,
    n67349, n67350, n67351, n67352, n67353, n67354, n67355, n67356, n67357,
    n67358, n67359, n67360, n67361, n67362, n67363, n67364, n67365, n67366,
    n67367, n67368, n67369, n67370, n67371, n67372, n67373, n67374, n67375,
    n67376, n67377, n67378, n67379, n67380, n67381, n67382, n67383, n67384,
    n67385, n67386, n67387, n67388, n67389, n67390, n67391, n67392, n67393,
    n67394, n67395, n67396, n67397, n67398, n67399, n67400, n67401, n67402,
    n67403, n67404, n67405, n67406, n67407, n67408, n67409, n67410, n67411,
    n67412, n67413, n67414, n67415, n67416, n67417, n67418, n67419, n67420,
    n67421, n67422, n67423, n67424, n67425, n67426, n67427, n67428, n67429,
    n67430, n67431, n67432, n67433, n67434, n67435, n67436, n67437, n67438,
    n67439, n67440, n67441, n67442, n67443, n67444, n67445, n67446, n67447,
    n67448, n67449, n67450, n67451, n67452, n67453, n67454, n67455, n67456,
    n67457, n67458, n67459, n67460, n67461, n67462, n67463, n67464, n67465,
    n67466, n67467, n67468, n67469, n67470, n67471, n67472, n67473, n67474,
    n67475, n67476, n67477, n67478, n67479, n67480, n67481, n67482, n67483,
    n67484, n67485, n67486, n67487, n67488, n67489, n67490, n67491, n67492,
    n67493, n67494, n67495, n67496, n67497, n67498, n67499, n67500, n67501,
    n67502, n67503, n67504, n67505, n67506, n67507, n67508, n67509, n67510,
    n67511, n67512, n67513, n67514, n67515, n67516, n67517, n67518, n67519,
    n67520, n67521, n67522, n67523, n67524, n67525, n67526, n67527, n67528,
    n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536, n67537,
    n67538, n67539, n67540, n67541, n67542, n67543, n67544, n67545, n67546,
    n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554, n67555,
    n67556, n67557, n67558, n67559, n67560, n67561, n67562, n67563, n67564,
    n67565, n67566, n67567, n67568, n67569, n67570, n67571, n67572, n67573,
    n67574, n67575, n67576, n67577, n67578, n67579, n67580, n67581, n67582,
    n67583, n67584, n67585, n67586, n67587, n67588, n67589, n67590, n67591,
    n67592, n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600,
    n67601, n67602, n67603, n67604, n67605, n67606, n67607, n67608, n67609,
    n67610, n67611, n67612, n67613, n67614, n67615, n67616, n67617, n67618,
    n67619, n67620, n67621, n67622, n67623, n67624, n67625, n67626, n67627,
    n67628, n67629, n67630, n67631, n67632, n67633, n67634, n67635, n67636,
    n67637, n67638, n67639, n67640, n67641, n67642, n67643, n67644, n67645,
    n67646, n67647, n67648, n67649, n67650, n67651, n67652, n67653, n67654,
    n67655, n67656, n67657, n67658, n67659, n67660, n67661, n67662, n67663,
    n67664, n67665, n67666, n67667, n67668, n67669, n67670, n67671, n67672,
    n67673, n67674, n67675, n67676, n67677, n67678, n67679, n67680, n67681,
    n67682, n67683, n67684, n67685, n67686, n67687, n67688, n67689, n67690,
    n67691, n67692, n67693, n67694, n67695, n67696, n67697, n67698, n67699,
    n67700, n67701, n67702, n67703, n67704, n67705, n67706, n67707, n67708,
    n67709, n67710, n67711, n67712, n67713, n67714, n67715, n67716, n67717,
    n67718, n67719, n67720, n67721, n67722, n67723, n67724, n67725, n67726,
    n67727, n67728, n67729, n67730, n67731, n67732, n67733, n67734, n67735,
    n67736, n67737, n67738, n67739, n67740, n67741, n67742, n67743, n67744,
    n67745, n67746, n67747, n67748, n67749, n67750, n67751, n67752, n67753,
    n67754, n67755, n67756, n67757, n67758, n67759, n67760, n67761, n67762,
    n67763, n67764, n67765, n67766, n67767, n67768, n67769, n67770, n67771,
    n67772, n67773, n67774, n67775, n67776, n67777, n67778, n67779, n67780,
    n67781, n67782, n67783, n67784, n67785, n67786, n67787, n67788, n67789,
    n67790, n67791, n67792, n67793, n67794, n67795, n67796, n67797, n67798,
    n67799, n67800, n67801, n67802, n67803, n67804, n67805, n67806, n67807,
    n67808, n67809, n67810, n67811, n67812, n67813, n67814, n67815, n67816,
    n67817, n67818, n67819, n67820, n67821, n67822, n67823, n67824, n67825,
    n67826, n67827, n67828, n67829, n67830, n67831, n67832, n67833, n67834,
    n67835, n67836, n67837, n67838, n67839, n67840, n67841, n67842, n67843,
    n67844, n67845, n67846, n67847, n67848, n67849, n67850, n67851, n67852,
    n67853, n67854, n67855, n67856, n67857, n67858, n67859, n67860, n67861,
    n67862, n67863, n67864, n67865, n67866, n67867, n67868, n67869, n67870,
    n67871, n67872, n67873, n67874, n67875, n67876, n67877, n67878, n67879,
    n67880, n67881, n67882, n67883, n67884, n67885, n67886, n67887, n67888,
    n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896, n67897,
    n67898, n67899, n67900, n67901, n67902, n67903, n67904, n67905, n67906,
    n67907, n67908, n67909, n67910, n67911, n67912, n67913, n67914, n67915,
    n67916, n67917, n67918, n67919, n67920, n67921, n67922, n67923, n67924,
    n67925, n67926, n67927, n67928, n67929, n67930, n67931, n67932, n67933,
    n67934, n67935, n67936, n67937, n67938, n67939, n67940, n67941, n67942,
    n67943, n67944, n67945, n67946, n67947, n67948, n67949, n67950, n67951,
    n67952, n67953, n67954, n67955, n67956, n67957, n67958, n67959, n67960,
    n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968, n67969,
    n67970, n67971, n67972, n67973, n67974, n67975, n67976, n67977, n67978,
    n67979, n67980, n67981, n67982, n67983, n67984, n67985, n67986, n67987,
    n67988, n67989, n67990, n67991, n67992, n67993, n67994, n67995, n67996,
    n67997, n67998, n67999, n68000, n68001, n68002, n68003, n68004, n68005,
    n68006, n68007, n68008, n68009, n68010, n68011, n68012, n68013, n68014,
    n68015, n68016, n68017, n68018, n68019, n68020, n68021, n68022, n68023,
    n68024, n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032,
    n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040, n68041,
    n68042, n68043, n68044, n68045, n68046, n68047, n68048, n68049, n68050,
    n68051, n68052, n68053, n68054, n68055, n68056, n68057, n68058, n68059,
    n68060, n68061, n68062, n68063, n68064, n68065, n68066, n68067, n68068,
    n68069, n68070, n68071, n68072, n68073, n68074, n68075, n68076, n68077,
    n68078, n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086,
    n68087, n68088, n68089, n68090, n68091, n68092, n68093, n68094, n68095,
    n68096, n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104,
    n68105, n68106, n68107, n68108, n68109, n68110, n68111, n68112, n68113,
    n68114, n68115, n68116, n68117, n68118, n68119, n68120, n68121, n68122,
    n68123, n68124, n68125, n68126, n68127, n68128, n68129, n68130, n68131,
    n68132, n68133, n68134, n68135, n68136, n68137, n68138, n68139, n68140,
    n68141, n68142, n68143, n68144, n68145, n68146, n68147, n68148, n68149,
    n68150, n68151, n68152, n68153, n68154, n68155, n68156, n68157, n68158,
    n68159, n68160, n68161, n68162, n68163, n68164, n68165, n68166, n68167,
    n68168, n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176,
    n68177, n68178, n68179, n68180, n68181, n68182, n68183, n68184, n68185,
    n68186, n68187, n68188, n68189, n68190, n68191, n68192, n68193, n68194,
    n68195, n68196, n68197, n68198, n68199, n68200, n68201, n68202, n68203,
    n68204, n68205, n68206, n68207, n68208, n68209, n68210, n68211, n68212,
    n68213, n68214, n68215, n68216, n68217, n68218, n68219, n68220, n68221,
    n68222, n68223, n68224, n68225, n68226, n68227, n68228, n68229, n68230,
    n68231, n68232, n68233, n68234, n68235, n68236, n68237, n68238, n68239,
    n68240, n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248,
    n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256, n68257,
    n68258, n68259, n68260, n68261, n68262, n68263, n68264, n68265, n68266,
    n68267, n68268, n68269, n68270, n68271, n68272, n68273, n68274, n68275,
    n68276, n68277, n68278, n68279, n68280, n68281, n68282, n68283, n68284,
    n68285, n68286, n68287, n68288, n68289, n68290, n68291, n68292, n68293,
    n68294, n68295, n68296, n68297, n68298, n68299, n68300, n68301, n68302,
    n68303, n68304, n68305, n68306, n68307, n68308, n68309, n68310, n68311,
    n68312, n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320,
    n68321, n68322, n68323, n68324, n68325, n68326, n68327, n68328, n68329,
    n68330, n68331, n68332, n68333, n68334, n68335, n68336, n68337, n68338,
    n68339, n68340, n68341, n68342, n68343, n68344, n68345, n68346, n68347,
    n68348, n68349, n68350, n68351, n68352, n68353, n68354, n68355, n68356,
    n68357, n68358, n68359, n68360, n68361, n68362, n68363, n68364, n68365,
    n68366, n68367, n68368, n68369, n68370, n68371, n68372, n68373, n68374,
    n68375, n68376, n68377, n68378, n68379, n68380, n68381, n68382, n68383,
    n68384, n68385, n68386, n68387, n68388, n68389, n68390, n68391, n68392,
    n68393, n68394, n68395, n68396, n68397, n68398, n68399, n68400, n68401,
    n68402, n68403, n68404, n68405, n68406, n68407, n68408, n68409, n68410,
    n68411, n68412, n68413, n68414, n68415, n68416, n68417, n68418, n68419,
    n68420, n68421, n68422, n68423, n68424, n68425, n68426, n68427, n68428,
    n68429, n68430, n68431, n68432, n68433, n68434, n68435, n68436, n68437,
    n68438, n68439, n68440, n68441, n68442, n68443, n68444, n68445, n68446,
    n68447, n68448, n68449, n68450, n68451, n68452, n68453, n68454, n68455,
    n68456, n68457, n68458, n68459, n68460, n68461, n68462, n68463, n68464,
    n68465, n68466, n68467, n68468, n68469, n68470, n68471, n68472, n68473,
    n68474, n68475, n68476, n68477, n68478, n68479, n68480, n68481, n68482,
    n68483, n68484, n68485, n68486, n68487, n68488, n68489, n68490, n68491,
    n68492, n68493, n68494, n68495, n68496, n68497, n68498, n68499, n68500,
    n68501, n68502, n68503, n68504, n68505, n68506, n68507, n68508, n68509,
    n68510, n68511, n68512, n68513, n68514, n68515, n68516, n68517, n68518,
    n68519, n68520, n68521, n68522, n68523, n68524, n68525, n68526, n68527,
    n68528, n68529, n68530, n68531, n68532, n68533, n68534, n68535, n68536,
    n68537, n68538, n68539, n68540, n68541, n68542, n68543, n68544, n68545,
    n68546, n68547, n68548, n68549, n68550, n68551, n68552, n68553, n68554,
    n68555, n68556, n68557, n68558, n68559, n68560, n68561, n68562, n68563,
    n68564, n68565, n68566, n68567, n68568, n68569, n68570, n68571, n68572,
    n68573, n68574, n68575, n68576, n68577, n68578, n68579, n68580, n68581,
    n68582, n68583, n68584, n68585, n68586, n68587, n68588, n68589, n68590,
    n68591, n68592, n68593, n68594, n68595, n68596, n68597, n68598, n68599,
    n68600, n68601, n68602, n68603, n68604, n68605, n68606, n68607, n68608,
    n68609, n68610, n68611, n68612, n68613, n68614, n68615, n68616, n68617,
    n68618, n68619, n68620, n68621, n68622, n68623, n68624, n68625, n68626,
    n68627, n68628, n68629, n68630, n68631, n68632, n68633, n68634, n68635,
    n68636, n68637, n68638, n68639, n68640, n68641, n68642, n68643, n68644,
    n68645, n68646, n68647, n68648, n68649, n68650, n68651, n68652, n68653,
    n68654, n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662,
    n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671,
    n68672, n68673, n68674, n68675, n68676, n68677, n68678, n68679, n68680,
    n68681, n68682, n68683, n68684, n68685, n68686, n68687, n68688, n68689,
    n68690, n68691, n68692, n68693, n68694, n68695, n68696, n68697, n68698,
    n68699, n68700, n68701, n68702, n68703, n68704, n68705, n68706, n68707,
    n68708, n68709, n68710, n68711, n68712, n68713, n68714, n68715, n68716,
    n68717, n68718, n68719, n68720, n68721, n68722, n68723, n68724, n68725,
    n68726, n68727, n68728, n68729, n68730, n68731, n68732, n68733, n68734,
    n68735, n68736, n68737, n68738, n68739, n68740, n68741, n68742, n68743,
    n68744, n68745, n68746, n68747, n68748, n68749, n68750, n68751, n68752,
    n68753, n68754, n68755, n68756, n68757, n68758, n68759, n68760, n68761,
    n68762, n68763, n68764, n68765, n68766, n68767, n68768, n68769, n68770,
    n68771, n68772, n68773, n68774, n68775, n68776, n68777, n68778, n68779,
    n68780, n68781, n68782, n68783, n68784, n68785, n68786, n68787, n68788,
    n68789, n68790, n68791, n68792, n68793, n68794, n68795, n68796, n68797,
    n68798, n68799, n68800, n68801, n68802, n68803, n68804, n68805, n68806,
    n68807, n68808, n68809, n68810, n68811, n68812, n68813, n68814, n68815,
    n68816, n68817, n68818, n68819, n68820, n68821, n68822, n68823, n68824,
    n68825, n68826, n68827, n68828, n68829, n68830, n68831, n68832, n68833,
    n68834, n68835, n68836, n68837, n68838, n68839, n68840, n68841, n68842,
    n68843, n68844, n68845, n68846, n68847, n68848, n68849, n68850, n68851,
    n68852, n68853, n68854, n68855, n68856, n68857, n68858, n68859, n68860,
    n68861, n68862, n68863, n68864, n68865, n68866, n68867, n68868, n68869,
    n68870, n68871, n68872, n68873, n68874, n68875, n68876, n68877, n68878,
    n68879, n68880, n68881, n68882, n68883, n68884, n68885, n68886, n68887,
    n68888, n68889, n68890, n68891, n68892, n68893, n68894, n68895, n68896,
    n68897, n68898, n68899, n68900, n68901, n68902, n68903, n68904, n68905,
    n68906, n68907, n68908, n68909, n68910, n68911, n68912, n68913, n68914,
    n68915, n68916, n68917, n68918, n68919, n68920, n68921, n68922, n68923,
    n68924, n68925, n68926, n68927, n68928, n68929, n68930, n68931, n68932,
    n68933, n68934, n68935, n68936, n68937, n68938, n68939, n68940, n68941,
    n68942, n68943, n68944, n68945, n68946, n68947, n68948, n68949, n68950,
    n68951, n68952, n68953, n68954, n68955, n68956, n68957, n68958, n68959,
    n68960, n68961, n68962, n68963, n68964, n68965, n68966, n68967, n68968,
    n68969, n68970, n68971, n68972, n68973, n68974, n68975, n68976, n68977,
    n68978, n68979, n68980, n68981, n68982, n68983, n68984, n68985, n68986,
    n68987, n68988, n68989, n68990, n68991, n68992, n68993, n68994, n68995,
    n68996, n68997, n68998, n68999, n69000, n69001, n69002, n69003, n69004,
    n69005, n69006, n69007, n69008, n69009, n69010, n69011, n69012, n69013,
    n69014, n69015, n69016, n69017, n69018, n69019, n69020, n69021, n69022,
    n69023, n69024, n69025, n69026, n69027, n69028, n69029, n69030, n69031,
    n69032, n69033, n69034, n69035, n69036, n69037, n69038, n69039, n69040,
    n69041, n69042, n69043, n69044, n69045, n69046, n69047, n69048, n69049,
    n69050, n69051, n69052, n69053, n69054, n69055, n69056, n69057, n69058,
    n69059, n69060, n69061, n69062, n69063, n69064, n69065, n69066, n69067,
    n69068, n69069, n69070, n69071, n69072, n69073, n69074, n69075, n69076,
    n69077, n69078, n69079, n69080, n69081, n69082, n69083, n69084, n69085,
    n69086, n69087, n69088, n69089, n69090, n69091, n69092, n69093, n69094,
    n69095, n69096, n69097, n69098, n69099, n69100, n69101, n69102, n69103,
    n69104, n69105, n69106, n69107, n69108, n69109, n69110, n69111, n69112,
    n69113, n69114, n69115, n69116, n69117, n69118, n69119, n69120, n69121,
    n69122, n69123, n69124, n69125, n69126, n69127, n69128, n69129, n69130,
    n69131, n69132, n69133, n69134, n69135, n69136, n69137, n69138, n69139,
    n69140, n69141, n69142, n69143, n69144, n69145, n69146, n69147, n69148,
    n69149, n69150, n69151, n69152, n69153, n69154, n69155, n69156, n69157,
    n69158, n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69166,
    n69167, n69168, n69169, n69170, n69171, n69172, n69173, n69174, n69175,
    n69176, n69177, n69178, n69179, n69180, n69181, n69182, n69183, n69184,
    n69185, n69186, n69187, n69188, n69189, n69190, n69191, n69192, n69193,
    n69194, n69195, n69196, n69197, n69198, n69199, n69200, n69201, n69202,
    n69203, n69204, n69205, n69206, n69207, n69208, n69209, n69210, n69211,
    n69212, n69213, n69214, n69215, n69216, n69217, n69218, n69219, n69220,
    n69221, n69222, n69223, n69224, n69225, n69226, n69227, n69228, n69229,
    n69230, n69231, n69232, n69233, n69234, n69235, n69236, n69237, n69238,
    n69239, n69240, n69241, n69242, n69243, n69244, n69245, n69246, n69247,
    n69248, n69249, n69250, n69251, n69252, n69253, n69254, n69255, n69256,
    n69257, n69258, n69259, n69260, n69261, n69262, n69263, n69264, n69265,
    n69266, n69267, n69268, n69269, n69270, n69271, n69272, n69273, n69274,
    n69275, n69276, n69277, n69278, n69279, n69280, n69281, n69282, n69283,
    n69284, n69285, n69286, n69287, n69288, n69289, n69290, n69291, n69292,
    n69293, n69294, n69295, n69296, n69297, n69298, n69299, n69300, n69301,
    n69302, n69303, n69304, n69305, n69306, n69307, n69308, n69309, n69310,
    n69311, n69312, n69313, n69314, n69315, n69316, n69317, n69318, n69319,
    n69320, n69321, n69322, n69323, n69324, n69325, n69326, n69327, n69328,
    n69329, n69330, n69331, n69332, n69333, n69334, n69335, n69336, n69337,
    n69338, n69339, n69340, n69341, n69342, n69343, n69344, n69345, n69346,
    n69347, n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355,
    n69356, n69357, n69358, n69359, n69360, n69361, n69362, n69363, n69364,
    n69365, n69366, n69367, n69368, n69369, n69370, n69371, n69372, n69373,
    n69374, n69375, n69376, n69377, n69378, n69379, n69380, n69381, n69382,
    n69383, n69384, n69385, n69386, n69387, n69388, n69389, n69390, n69391,
    n69392, n69393, n69394, n69395, n69396, n69397, n69398, n69399, n69400,
    n69401, n69402, n69403, n69404, n69405, n69406, n69407, n69408, n69409,
    n69410, n69411, n69412, n69413, n69414, n69415, n69416, n69417, n69418,
    n69419, n69420, n69421, n69422, n69423, n69424, n69425, n69426, n69427,
    n69428, n69429, n69430, n69431, n69432, n69433, n69434, n69435, n69436,
    n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444, n69445,
    n69446, n69447, n69448, n69449, n69450, n69451, n69452, n69453, n69454,
    n69455, n69456, n69457, n69458, n69459, n69460, n69461, n69462, n69463,
    n69464, n69465, n69466, n69467, n69468, n69469, n69470, n69471, n69472,
    n69473, n69474, n69475, n69476, n69477, n69478, n69479, n69480, n69481,
    n69482, n69483, n69484, n69485, n69486, n69487, n69488, n69489, n69490,
    n69491, n69492, n69493, n69494, n69495, n69496, n69497, n69498, n69499,
    n69500, n69501, n69502, n69503, n69504, n69505, n69506, n69507, n69508,
    n69509, n69510, n69511, n69512, n69513, n69514, n69515, n69516, n69517,
    n69518, n69519, n69520, n69521, n69522, n69523, n69524, n69525, n69526,
    n69527, n69528, n69529, n69530, n69531, n69532, n69533, n69534, n69535,
    n69536, n69537, n69538, n69539, n69540, n69541, n69542, n69543, n69544,
    n69545, n69546, n69547, n69548, n69549, n69550, n69551, n69552, n69553,
    n69554, n69555, n69556, n69557, n69558, n69559, n69560, n69561, n69562,
    n69563, n69564, n69565, n69566, n69567, n69568, n69569, n69570, n69571,
    n69572, n69573, n69574, n69575, n69576, n69577, n69578, n69579, n69580,
    n69581, n69582, n69583, n69584, n69585, n69586, n69587, n69588, n69589,
    n69590, n69591, n69592, n69593, n69594, n69595, n69596, n69597, n69598,
    n69599, n69600, n69601, n69602, n69603, n69604, n69605, n69606, n69607,
    n69608, n69609, n69610, n69611, n69612, n69613, n69614, n69615, n69616,
    n69617, n69618, n69619, n69620, n69621, n69622, n69623, n69624, n69625,
    n69626, n69627, n69628, n69629, n69630, n69631, n69632, n69633, n69634,
    n69635, n69636, n69637, n69638, n69639, n69640, n69641, n69642, n69643,
    n69644, n69645, n69646, n69647, n69648, n69649, n69650, n69651, n69652,
    n69653, n69654, n69655, n69656, n69657, n69658, n69659, n69660, n69661,
    n69662, n69663, n69664, n69665, n69666, n69667, n69668, n69669, n69670,
    n69671, n69672, n69673, n69674, n69675, n69676, n69677, n69678, n69679,
    n69680, n69681, n69682, n69683, n69684, n69685, n69686, n69687, n69688,
    n69689, n69690, n69691, n69692, n69693, n69694, n69695, n69696, n69697,
    n69698, n69699, n69700, n69701, n69702, n69703, n69704, n69705, n69706,
    n69707, n69708, n69709, n69710, n69711, n69712, n69713, n69714, n69715,
    n69716, n69717, n69718, n69719, n69720, n69721, n69722, n69723, n69724,
    n69725, n69726, n69727, n69728, n69729, n69730, n69731, n69732, n69733,
    n69734, n69735, n69736, n69737, n69738, n69739, n69740, n69741, n69742,
    n69743, n69744, n69745, n69746, n69747, n69748, n69749, n69750, n69751,
    n69752, n69753, n69754, n69755, n69756, n69757, n69758, n69759, n69760,
    n69761, n69762, n69763, n69764, n69765, n69766, n69767, n69768, n69769,
    n69770, n69771, n69772, n69773, n69774, n69775, n69776, n69777, n69778,
    n69779, n69780, n69781, n69782, n69783, n69784, n69785, n69786, n69787,
    n69788, n69789, n69790, n69791, n69792, n69793, n69794, n69795, n69796,
    n69797, n69798, n69799, n69800, n69801, n69802, n69803, n69804, n69805,
    n69806, n69807, n69808, n69809, n69810, n69811, n69812, n69813, n69814,
    n69815, n69816, n69817, n69818, n69819, n69820, n69821, n69822, n69823,
    n69824, n69825, n69826, n69827, n69828, n69829, n69830, n69831, n69832,
    n69833, n69834, n69835, n69836, n69837, n69838, n69839, n69840, n69841,
    n69842, n69843, n69844, n69845, n69846, n69847, n69848, n69849, n69850,
    n69851, n69852, n69853, n69854, n69855, n69856, n69857, n69858, n69859,
    n69860, n69861, n69862, n69863, n69864, n69865, n69866, n69867, n69868,
    n69869, n69870, n69871, n69872, n69873, n69874, n69875, n69876, n69877,
    n69878, n69879, n69880, n69881, n69882, n69883, n69884, n69885, n69886,
    n69887, n69888, n69889, n69890, n69891, n69892, n69893, n69894, n69895,
    n69896, n69897, n69898, n69899, n69900, n69901, n69902, n69903, n69904,
    n69905, n69906, n69907, n69908, n69909, n69910, n69911, n69912, n69913,
    n69914, n69915, n69916, n69917, n69918, n69919, n69920, n69921, n69922,
    n69923, n69924, n69925, n69926, n69927, n69928, n69929, n69930, n69931,
    n69932, n69933, n69934, n69935, n69936, n69937, n69938, n69939, n69940,
    n69941, n69942, n69943, n69944, n69945, n69946, n69947, n69948, n69949,
    n69950, n69951, n69952, n69953, n69954, n69955, n69956, n69957, n69958,
    n69959, n69960, n69961, n69962, n69963, n69964, n69965, n69966, n69967,
    n69968, n69969, n69970, n69971, n69972, n69973, n69974, n69975, n69976,
    n69977, n69978, n69979, n69980, n69981, n69982, n69983, n69984, n69985,
    n69986, n69987, n69988, n69989, n69990, n69991, n69992, n69993, n69994,
    n69995, n69996, n69997, n69998, n69999, n70000, n70001, n70002, n70003,
    n70004, n70005, n70006, n70007, n70008, n70009, n70010, n70011, n70012,
    n70013, n70014, n70015, n70016, n70017, n70018, n70019, n70020, n70021,
    n70022, n70023, n70024, n70025, n70026, n70027, n70028, n70029, n70030,
    n70031, n70032, n70033, n70034, n70035, n70036, n70037, n70038, n70039,
    n70040, n70041, n70042, n70043, n70044, n70045, n70046, n70047, n70048,
    n70049, n70050, n70051, n70052, n70053, n70054, n70055, n70056, n70057,
    n70058, n70059, n70060, n70061, n70062, n70063, n70064, n70065, n70066,
    n70067, n70068, n70069, n70070, n70071, n70072, n70073, n70074, n70075,
    n70076, n70077, n70078, n70079, n70080, n70081, n70082, n70083, n70084,
    n70085, n70086, n70087, n70088, n70089, n70090, n70091, n70092, n70093,
    n70094, n70095, n70096, n70097, n70098, n70099, n70100, n70101, n70102,
    n70103, n70104, n70105, n70106, n70107, n70108, n70109, n70110, n70111,
    n70112, n70113, n70114, n70115, n70116, n70117, n70118, n70119, n70120,
    n70121, n70122, n70123, n70124, n70125, n70126, n70127, n70128, n70129,
    n70130, n70131, n70132, n70133, n70134, n70135, n70136, n70137, n70138,
    n70139, n70140, n70141, n70142, n70143, n70144, n70145, n70146, n70147,
    n70148, n70149, n70150, n70151, n70152, n70153, n70154, n70155, n70156,
    n70157, n70158, n70159, n70160, n70161, n70162, n70163, n70164, n70165,
    n70166, n70167, n70168, n70169, n70170, n70171, n70172, n70173, n70174,
    n70175, n70176, n70177, n70178, n70179, n70180, n70181, n70182, n70183,
    n70184, n70185, n70186, n70187, n70188, n70189, n70190, n70191, n70192,
    n70193, n70194, n70195, n70196, n70197, n70198, n70199, n70200, n70201,
    n70202, n70203, n70204, n70205, n70206, n70207, n70208, n70209, n70210,
    n70211, n70212, n70213, n70214, n70215, n70216, n70217, n70218, n70219,
    n70220, n70221, n70222, n70223, n70224, n70225, n70226, n70227, n70228,
    n70229, n70230, n70231, n70232, n70233, n70234, n70235, n70236, n70237,
    n70238, n70239, n70240, n70241, n70242, n70243, n70244, n70245, n70246,
    n70247, n70248, n70249, n70250, n70251, n70252, n70253, n70254, n70255,
    n70256, n70257, n70258, n70259, n70260, n70261, n70262, n70263, n70264,
    n70265, n70266, n70267, n70268, n70269, n70270, n70271, n70272, n70273,
    n70274, n70275, n70276, n70277, n70278, n70279, n70280, n70281, n70282,
    n70283, n70284, n70285, n70286, n70287, n70288, n70289, n70290, n70291,
    n70292, n70293, n70294, n70295, n70296, n70297, n70298, n70299, n70300,
    n70301, n70302, n70303, n70304, n70305, n70306, n70307, n70308, n70309,
    n70310, n70311, n70312, n70313, n70314, n70315, n70316, n70317, n70318,
    n70319, n70320, n70321, n70322, n70323, n70324, n70325, n70326, n70327,
    n70328, n70329, n70330, n70331, n70332, n70333, n70334, n70335, n70336,
    n70337, n70338, n70339, n70340, n70341, n70342, n70343, n70344, n70345,
    n70346, n70347, n70348, n70349, n70350, n70351, n70352, n70353, n70354,
    n70355, n70356, n70357, n70358, n70359, n70360, n70361, n70362, n70363,
    n70364, n70365, n70366, n70367, n70368, n70369, n70370, n70371, n70372,
    n70373, n70374, n70375, n70376, n70377, n70378, n70379, n70380, n70381,
    n70382, n70383, n70384, n70385, n70386, n70387, n70388, n70389, n70390,
    n70391, n70392, n70393, n70394, n70395, n70396, n70397, n70398, n70399,
    n70400, n70401, n70402, n70403, n70404, n70405, n70406, n70407, n70408,
    n70409, n70410, n70411, n70412, n70413, n70414, n70415, n70416, n70417,
    n70418, n70419, n70420, n70421, n70422, n70423, n70424, n70425, n70426,
    n70427, n70428, n70429, n70430, n70431, n70432, n70433, n70434, n70435,
    n70436, n70437, n70438, n70439, n70440, n70441, n70442, n70443, n70444,
    n70445, n70446, n70447, n70448, n70449, n70450, n70451, n70452, n70453,
    n70454, n70455, n70456, n70457, n70458, n70459, n70460, n70461, n70462,
    n70463, n70464, n70465, n70466, n70467, n70468, n70469, n70470, n70471,
    n70472, n70473, n70474, n70475, n70476, n70477, n70478, n70479, n70480,
    n70481, n70482, n70483, n70484, n70485, n70486, n70487, n70488, n70489,
    n70490, n70491, n70492, n70493, n70494, n70495, n70496, n70497, n70498,
    n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507,
    n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516,
    n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524, n70525,
    n70526, n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534,
    n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542, n70543,
    n70544, n70545, n70546, n70547, n70548, n70549, n70550, n70551, n70552,
    n70553, n70554, n70555, n70556, n70557, n70558, n70559, n70560, n70561,
    n70562, n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570,
    n70571, n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579,
    n70580, n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588,
    n70589, n70590, n70591, n70592, n70593, n70594, n70595, n70596, n70597,
    n70598, n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606,
    n70607, n70608, n70609, n70610, n70611, n70612, n70613, n70614, n70615,
    n70616, n70617, n70618, n70619, n70620, n70621, n70622, n70623, n70624,
    n70625, n70626, n70627, n70628, n70629, n70630, n70631, n70632, n70633,
    n70634, n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642,
    n70643, n70644, n70645, n70646, n70647, n70648, n70649, n70650, n70651,
    n70652, n70653, n70654, n70655, n70656, n70657, n70658, n70659, n70660,
    n70661, n70662, n70663, n70664, n70665, n70666, n70667, n70668, n70669,
    n70670, n70671, n70672, n70673, n70674, n70675, n70676, n70677, n70678,
    n70679, n70680, n70681, n70682, n70683, n70684, n70685, n70686, n70687,
    n70688, n70689, n70690, n70691, n70692, n70693, n70694, n70695, n70696,
    n70697, n70698, n70699, n70700, n70701, n70702, n70703, n70704, n70705,
    n70706, n70707, n70708, n70709, n70710, n70711, n70712, n70713, n70714,
    n70715, n70716, n70717, n70718, n70719, n70720, n70721, n70722, n70723,
    n70724, n70725, n70726, n70727, n70728, n70729, n70730, n70731, n70732,
    n70733, n70734, n70735, n70736, n70737, n70738, n70739, n70740, n70741,
    n70742, n70743, n70744, n70745, n70746, n70747, n70748, n70749, n70750,
    n70751, n70752, n70753, n70754, n70755, n70756, n70757, n70758, n70759,
    n70760, n70761, n70762, n70763, n70764, n70765, n70766, n70767, n70768,
    n70769, n70770, n70771, n70772, n70773, n70774, n70775, n70776, n70777,
    n70778, n70779, n70780, n70781, n70782, n70783, n70784, n70785, n70786,
    n70787, n70788, n70789, n70790, n70791, n70792, n70793, n70794, n70795,
    n70796, n70797, n70798, n70799, n70800, n70801, n70802, n70803, n70804,
    n70805, n70806, n70807, n70808, n70809, n70810, n70811, n70812, n70813,
    n70814, n70815, n70816, n70817, n70818, n70819, n70820, n70821, n70822,
    n70823, n70824, n70825, n70826, n70827, n70828, n70829, n70830, n70831,
    n70832, n70833, n70834, n70835, n70836, n70837, n70838, n70839, n70840,
    n70841, n70842, n70843, n70844, n70845, n70846, n70847, n70848, n70849,
    n70850, n70851, n70852, n70853, n70854, n70855, n70856, n70857, n70858,
    n70859, n70860, n70861, n70862, n70863, n70864, n70865, n70866, n70867,
    n70868, n70869, n70870, n70871, n70872, n70873, n70874, n70875, n70876,
    n70877, n70878, n70879, n70880, n70881, n70882, n70883, n70884, n70885,
    n70886, n70887, n70888, n70889, n70890, n70891, n70892, n70893, n70894,
    n70895, n70896, n70897, n70898, n70899, n70900, n70901, n70902, n70903,
    n70904, n70905, n70906, n70907, n70908, n70909, n70910, n70911, n70912,
    n70913, n70914, n70915, n70916, n70917, n70918, n70919, n70920, n70921,
    n70922, n70923, n70924, n70925, n70926, n70927, n70928, n70929, n70930,
    n70931, n70932, n70933, n70934, n70935, n70936, n70937, n70938, n70939,
    n70940, n70941, n70942, n70943, n70944, n70945, n70946, n70947, n70948,
    n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956, n70957,
    n70958, n70959, n70960, n70961, n70962, n70963, n70964, n70965, n70966,
    n70967, n70968, n70969, n70970, n70971, n70972, n70973, n70974, n70975,
    n70976, n70977, n70978, n70979, n70980, n70981, n70982, n70983, n70984,
    n70985, n70986, n70987, n70988, n70989, n70990, n70991, n70992, n70993,
    n70994, n70995, n70996, n70997, n70998, n70999, n71000, n71001, n71002,
    n71003, n71004, n71005, n71006, n71007, n71008, n71009, n71010, n71011,
    n71012, n71013, n71014, n71015, n71016, n71017, n71018, n71019, n71020,
    n71021, n71022, n71023, n71024, n71025, n71026, n71027, n71028, n71029,
    n71030, n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038,
    n71039, n71040, n71041, n71042, n71043, n71044, n71045, n71046, n71047,
    n71048, n71049, n71050, n71051, n71052, n71053, n71054, n71055, n71056,
    n71057, n71058, n71059, n71060, n71061, n71062, n71063, n71064, n71065,
    n71066, n71067, n71068, n71069, n71070, n71071, n71072, n71073, n71074,
    n71075, n71076, n71077, n71078, n71079, n71080, n71081, n71082, n71083,
    n71084, n71085, n71086, n71087, n71088, n71089, n71090, n71091, n71092,
    n71093, n71094, n71095, n71096, n71097, n71098, n71099, n71100, n71101,
    n71102, n71103, n71104, n71105, n71106, n71107, n71108, n71109, n71110,
    n71111, n71112, n71113, n71114, n71115, n71116, n71117, n71118, n71119,
    n71120, n71121, n71122, n71123, n71124, n71125, n71126, n71127, n71128,
    n71129, n71130, n71131, n71132, n71133, n71134, n71135, n71136, n71137,
    n71138, n71139, n71140, n71141, n71142, n71143, n71144, n71145, n71146,
    n71147, n71148, n71149, n71150, n71151, n71152, n71153, n71154, n71155,
    n71156, n71157, n71158, n71159, n71160, n71161, n71162, n71163, n71164,
    n71165, n71166, n71167, n71168, n71169, n71170, n71171, n71172, n71173,
    n71174, n71175, n71176, n71177, n71178, n71179, n71180, n71181, n71182,
    n71183, n71184, n71185, n71186, n71187, n71188, n71189, n71190, n71191,
    n71192, n71193, n71194, n71195, n71196, n71197, n71198, n71199, n71200,
    n71201, n71202, n71203, n71204, n71205, n71206, n71207, n71208, n71209,
    n71210, n71211, n71212, n71213, n71214, n71215, n71216, n71217, n71218,
    n71219, n71220, n71221, n71222, n71223, n71224, n71225, n71226, n71227,
    n71228, n71229, n71230, n71231, n71232, n71233, n71234, n71235, n71236,
    n71237, n71238, n71239, n71240, n71241, n71242, n71243, n71244, n71245,
    n71246, n71247, n71248, n71249, n71250, n71251, n71252, n71253, n71254,
    n71255, n71256, n71257, n71258, n71259, n71260, n71261, n71262, n71263,
    n71264, n71265, n71266, n71267, n71268, n71269, n71270, n71271, n71272,
    n71273, n71274, n71275, n71276, n71277, n71278, n71279, n71280, n71281,
    n71282, n71283, n71284, n71285, n71286, n71287, n71288, n71289, n71290,
    n71291, n71292, n71293, n71294, n71295, n71296, n71297, n71298, n71299,
    n71300, n71301, n71302, n71303, n71304, n71305, n71306, n71307, n71308,
    n71309, n71310, n71311, n71312, n71313, n71314, n71315, n71316, n71317,
    n71318, n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326,
    n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334, n71335,
    n71336, n71337, n71338, n71339, n71340, n71341, n71342, n71343, n71344,
    n71345, n71346, n71347, n71348, n71349, n71350, n71351, n71352, n71353,
    n71354, n71355, n71356, n71357, n71358, n71359, n71360, n71361, n71362,
    n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370, n71371,
    n71372, n71373, n71374, n71375, n71376, n71377, n71378, n71379, n71380,
    n71381, n71382, n71383, n71384, n71385, n71386, n71387, n71388, n71389,
    n71390, n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398,
    n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406, n71407,
    n71408, n71409, n71410, n71411, n71412, n71413, n71414, n71415, n71416,
    n71417, n71418, n71419, n71420, n71421, n71422, n71423, n71424, n71425,
    n71426, n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434,
    n71435, n71436, n71437, n71438, n71439, n71440, n71441, n71442, n71443,
    n71444, n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452,
    n71453, n71454, n71455, n71456, n71457, n71458, n71459, n71460, n71461,
    n71462, n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470,
    n71471, n71472, n71473, n71474, n71475, n71476, n71477, n71478, n71479,
    n71480, n71481, n71482, n71483, n71484, n71485, n71486, n71487, n71488,
    n71489, n71490, n71491, n71492, n71493, n71494, n71495, n71496, n71497,
    n71498, n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506,
    n71507, n71508, n71509, n71510, n71511, n71512, n71513, n71514, n71515,
    n71516, n71517, n71518, n71519, n71520, n71521, n71522, n71523, n71524,
    n71525, n71526, n71527, n71528, n71529, n71530, n71531, n71532, n71533,
    n71534, n71535, n71536, n71537, n71538, n71539, n71540, n71541, n71542,
    n71543, n71544, n71545, n71546, n71547, n71548, n71549, n71550, n71551,
    n71552, n71553, n71554, n71555, n71556, n71557, n71558, n71559, n71560,
    n71561, n71562, n71563, n71564, n71565, n71566, n71567, n71568, n71569,
    n71570, n71571, n71572, n71573, n71574, n71575, n71576, n71577, n71578,
    n71579, n71580, n71581, n71582, n71583, n71584, n71585, n71586, n71587,
    n71588, n71589, n71590, n71591, n71592, n71593, n71594, n71595, n71596,
    n71597, n71598, n71599, n71600, n71601, n71602, n71603, n71604, n71605,
    n71606, n71607, n71608, n71609, n71610, n71611, n71612, n71613, n71614,
    n71615, n71616, n71617, n71618, n71619, n71620, n71621, n71622, n71623,
    n71624, n71625, n71626, n71627, n71628, n71629, n71630, n71631, n71632,
    n71633, n71634, n71635, n71636, n71637, n71638, n71639, n71640, n71641,
    n71642, n71643, n71644, n71645, n71646, n71647, n71648, n71649, n71650,
    n71651, n71652, n71653, n71654, n71655, n71656, n71657, n71658, n71659,
    n71660, n71661, n71662, n71663, n71664, n71665, n71666, n71667, n71668,
    n71669, n71670, n71671, n71672, n71673, n71674, n71675, n71676, n71677,
    n71678, n71679, n71680, n71681, n71682, n71683, n71684, n71685, n71686,
    n71687, n71688, n71689, n71690, n71691, n71692, n71693, n71694, n71695,
    n71696, n71697, n71698, n71699, n71700, n71701, n71702, n71703, n71704,
    n71705, n71706, n71707, n71708, n71709, n71710, n71711, n71712, n71713,
    n71714, n71715, n71716, n71717, n71718, n71719, n71720, n71721, n71722,
    n71723, n71724, n71725, n71726, n71727, n71728, n71729, n71730, n71731,
    n71732, n71733, n71734, n71735, n71736, n71737, n71738, n71739, n71740,
    n71741, n71742, n71743, n71744, n71745, n71746, n71747, n71748, n71749,
    n71750, n71751, n71752, n71753, n71754, n71755, n71756, n71757, n71758,
    n71759, n71760, n71761, n71762, n71763, n71764, n71765, n71766, n71767,
    n71768, n71769, n71770, n71771, n71772, n71773, n71774, n71775, n71776,
    n71777, n71778, n71779, n71780, n71781, n71782, n71783, n71784, n71785,
    n71786, n71787, n71788, n71789, n71790, n71791, n71792, n71793, n71794,
    n71795, n71796, n71797, n71798, n71799, n71800, n71801, n71802, n71803,
    n71804, n71805, n71806, n71807, n71808, n71809, n71810, n71811, n71812,
    n71813, n71814, n71815, n71816, n71817, n71818, n71819, n71820, n71821,
    n71822, n71823, n71824, n71825, n71826, n71827, n71828, n71829, n71830,
    n71831, n71832, n71833, n71834, n71835, n71836, n71837, n71838, n71839,
    n71840, n71841, n71842, n71843, n71844, n71845, n71846, n71847, n71848,
    n71849, n71850, n71851, n71852, n71853, n71854, n71855, n71856, n71857,
    n71858, n71859, n71860, n71861, n71862, n71863, n71864, n71865, n71866,
    n71867, n71868, n71869, n71870, n71871, n71872, n71873, n71874, n71875,
    n71876, n71877, n71878, n71879, n71880, n71881, n71882, n71883, n71884,
    n71885, n71886, n71887, n71888, n71889, n71890, n71891, n71892, n71893,
    n71894, n71895, n71896, n71897, n71898, n71899, n71900, n71901, n71902,
    n71903, n71904, n71905, n71906, n71907, n71908, n71909, n71910, n71911,
    n71912, n71913, n71914, n71915, n71916, n71917, n71918, n71919, n71920,
    n71921, n71922, n71923, n71924, n71925, n71926, n71927, n71928, n71929,
    n71930, n71931, n71932, n71933, n71934, n71935, n71936, n71937, n71938,
    n71939, n71940, n71941, n71942, n71943, n71944, n71945, n71946, n71947,
    n71948, n71949, n71950, n71951, n71952, n71953, n71954, n71955, n71956,
    n71957, n71958, n71959, n71960, n71961, n71962, n71963, n71964, n71965,
    n71966, n71967, n71968, n71969, n71970, n71971, n71972, n71973, n71974,
    n71975, n71976, n71977, n71978, n71979, n71980, n71981, n71982, n71983,
    n71984, n71985, n71986, n71987, n71988, n71989, n71990, n71991, n71992,
    n71993, n71994, n71995, n71996, n71997, n71998, n71999, n72000, n72001,
    n72002, n72003, n72004, n72005, n72006, n72007, n72008, n72009, n72010,
    n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018, n72019,
    n72020, n72021, n72022, n72023, n72024, n72025, n72026, n72027, n72028,
    n72029, n72030, n72031, n72032, n72033, n72034, n72035, n72036, n72037,
    n72038, n72039, n72040, n72041, n72042, n72043, n72044, n72045, n72046,
    n72047, n72048, n72049, n72050, n72051, n72052, n72053, n72054, n72055,
    n72056, n72057, n72058, n72059, n72060, n72061, n72062, n72063, n72064,
    n72065, n72066, n72067, n72068, n72069, n72070, n72071, n72072, n72073,
    n72074, n72075, n72076, n72077, n72078, n72079, n72080, n72081, n72082,
    n72083, n72084, n72085, n72086, n72087, n72088, n72089, n72090, n72091,
    n72092, n72093, n72094, n72095, n72096, n72097, n72098, n72099, n72100,
    n72101, n72102, n72103, n72104, n72105, n72106, n72107, n72108, n72109,
    n72110, n72111, n72112, n72113, n72114, n72115, n72116, n72117, n72118,
    n72119, n72120, n72121, n72122, n72123, n72124, n72125, n72126, n72127,
    n72128, n72129, n72130, n72131, n72132, n72133, n72134, n72135, n72136,
    n72137, n72138, n72139, n72140, n72141, n72142, n72143, n72144, n72145,
    n72146, n72147, n72148, n72149, n72150, n72151, n72152, n72153, n72154,
    n72155, n72156, n72157, n72158, n72159, n72160, n72161, n72162, n72163,
    n72164, n72165, n72166, n72167, n72168, n72169, n72170, n72171, n72172,
    n72173, n72174, n72175, n72176, n72177, n72178, n72179, n72180, n72181,
    n72182, n72183, n72184, n72185, n72186, n72187, n72188, n72189, n72190,
    n72191, n72192, n72193, n72194, n72195, n72196, n72197, n72198, n72199,
    n72200, n72201, n72202, n72203, n72204, n72205, n72206, n72207, n72208,
    n72209, n72210, n72211, n72212, n72213, n72214, n72215, n72216, n72217,
    n72218, n72219, n72220, n72221, n72222, n72223, n72224, n72225, n72226,
    n72227, n72228, n72229, n72230, n72231, n72232, n72233, n72234, n72235,
    n72236, n72237, n72238, n72239, n72240, n72241, n72242, n72243, n72244,
    n72245, n72246, n72247, n72248, n72249, n72250, n72251, n72252, n72253,
    n72254, n72255, n72256, n72257, n72258, n72259, n72260, n72261, n72262,
    n72263, n72264, n72265, n72266, n72267, n72268, n72269, n72270, n72271,
    n72272, n72273, n72274, n72275, n72276, n72277, n72278, n72279, n72280,
    n72281, n72282, n72283, n72284, n72285, n72286, n72287, n72288, n72289,
    n72290, n72291, n72292, n72293, n72294, n72295, n72296, n72297, n72298,
    n72299, n72300, n72301, n72302, n72303, n72304, n72305, n72306, n72307,
    n72308, n72309, n72310, n72311, n72312, n72313, n72314, n72315, n72316,
    n72317, n72318, n72319, n72320, n72321, n72322, n72323, n72324, n72325,
    n72326, n72327, n72328, n72329, n72330, n72331, n72332, n72333, n72334,
    n72335, n72336, n72337, n72338, n72339, n72340, n72341, n72342, n72343,
    n72344, n72345, n72346, n72347, n72348, n72349, n72350, n72351, n72352,
    n72353, n72354, n72355, n72356, n72357, n72358, n72359, n72360, n72361,
    n72362, n72363, n72364, n72365, n72366, n72367, n72368, n72369, n72370,
    n72371, n72372, n72373, n72374, n72375, n72376, n72377, n72378, n72379,
    n72380, n72381, n72382, n72383, n72384, n72385, n72386, n72387, n72388,
    n72389, n72390, n72391, n72392, n72393, n72394, n72395, n72396, n72397,
    n72398, n72399, n72400, n72401, n72402, n72403, n72404, n72405, n72406,
    n72407, n72408, n72409, n72410, n72411, n72412, n72413, n72414, n72415,
    n72416, n72417, n72418, n72419, n72420, n72421, n72422, n72423, n72424,
    n72425, n72426, n72427, n72428, n72429, n72430, n72431, n72432, n72433,
    n72434, n72435, n72436, n72437, n72438, n72439, n72440, n72441, n72442,
    n72443, n72444, n72445, n72446, n72447, n72448, n72449, n72450, n72451,
    n72452, n72453, n72454, n72455, n72456, n72457, n72458, n72459, n72460,
    n72461, n72462, n72463, n72464, n72465, n72466, n72467, n72468, n72469,
    n72470, n72471, n72472, n72473, n72474, n72475, n72476, n72477, n72478,
    n72479, n72480, n72481, n72482, n72483, n72484, n72485, n72486, n72487,
    n72488, n72489, n72490, n72491, n72492, n72493, n72494, n72495, n72496,
    n72497, n72498, n72499, n72500, n72501, n72502, n72503, n72504, n72505,
    n72506, n72507, n72508, n72509, n72510, n72511, n72512, n72513, n72514,
    n72515, n72516, n72517, n72518, n72519, n72520, n72521, n72522, n72523,
    n72524, n72525, n72526, n72527, n72528, n72529, n72530, n72531, n72532,
    n72533, n72534, n72535, n72536, n72537, n72538, n72539, n72540, n72541,
    n72542, n72543, n72544, n72545, n72546, n72547, n72548, n72549, n72550,
    n72551, n72552, n72553, n72554, n72555, n72556, n72557, n72558, n72559,
    n72560, n72561, n72562, n72563, n72564, n72565, n72566, n72567, n72568,
    n72569, n72570, n72571, n72572, n72573, n72574, n72575, n72576, n72577,
    n72578, n72579, n72580, n72581, n72582, n72583, n72584, n72585, n72586,
    n72587, n72588, n72589, n72590, n72591, n72592, n72593, n72594, n72595,
    n72596, n72597, n72598, n72599, n72600, n72601, n72602, n72603, n72604,
    n72605, n72606, n72607, n72608, n72609, n72610, n72611, n72612, n72613,
    n72614, n72615, n72616, n72617, n72618, n72619, n72620, n72621, n72622,
    n72623, n72624, n72625, n72626, n72627, n72628, n72629, n72630, n72631,
    n72632, n72633, n72634, n72635, n72636, n72637, n72638, n72639, n72640,
    n72641, n72642, n72643, n72644, n72645, n72646, n72647, n72648, n72649,
    n72650, n72651, n72652, n72653, n72654, n72655, n72656, n72657, n72658,
    n72659, n72660, n72661, n72662, n72663, n72664, n72665, n72666, n72667,
    n72668, n72669, n72670, n72671, n72672, n72673, n72674, n72675, n72676,
    n72677, n72678, n72679, n72680, n72681, n72682, n72683, n72684, n72685,
    n72686, n72687, n72688, n72689, n72690, n72691, n72692, n72693, n72694,
    n72695, n72696, n72697, n72698, n72699, n72700, n72701, n72702, n72703,
    n72704, n72705, n72706, n72707, n72708, n72709, n72710, n72711, n72712,
    n72713, n72714, n72715, n72716, n72717, n72718, n72719, n72720, n72721,
    n72722, n72723, n72724, n72725, n72726, n72727, n72728, n72729, n72730,
    n72731, n72732, n72733, n72734, n72735, n72736, n72737, n72738, n72739,
    n72740, n72741, n72742, n72743, n72744, n72745, n72746, n72747, n72748,
    n72749, n72750, n72751, n72752, n72753, n72754, n72755, n72756, n72757,
    n72758, n72759, n72760, n72761, n72762, n72763, n72764, n72765, n72766,
    n72767, n72768, n72769, n72770, n72771, n72772, n72773, n72774, n72775,
    n72776, n72777, n72778, n72779, n72780, n72781, n72782, n72783, n72784,
    n72785, n72786, n72787, n72788, n72789, n72790, n72791, n72792, n72793,
    n72794, n72795, n72796, n72797, n72798, n72799, n72800, n72801, n72802,
    n72803, n72804, n72805, n72806, n72807, n72808, n72809, n72810, n72811,
    n72812, n72813, n72814, n72815, n72816, n72817, n72818, n72819, n72820,
    n72821, n72822, n72823, n72824, n72825, n72826, n72827, n72828, n72829,
    n72830, n72831, n72832, n72833, n72834, n72835, n72836, n72837, n72838,
    n72839, n72840, n72841, n72842, n72843, n72844, n72845, n72846, n72847,
    n72848, n72849, n72850, n72851, n72852, n72853, n72854, n72855, n72856,
    n72857, n72858, n72859, n72860, n72861, n72862, n72863, n72864, n72865,
    n72866, n72867, n72868, n72869, n72870, n72871, n72872, n72873, n72874,
    n72875, n72876, n72877, n72878, n72879, n72880, n72881, n72882, n72883,
    n72884, n72885, n72886, n72887, n72888, n72889, n72890, n72891, n72892,
    n72893, n72894, n72895, n72896, n72897, n72898, n72899, n72900, n72901,
    n72902, n72903, n72904, n72905, n72906, n72907, n72908, n72909, n72910,
    n72911, n72912, n72913, n72914, n72915, n72916, n72917, n72918, n72919,
    n72920, n72921, n72922, n72923, n72924, n72925, n72926, n72927, n72928,
    n72929, n72930, n72931, n72932, n72933, n72934, n72935, n72936, n72937,
    n72938, n72939, n72940, n72941, n72942, n72943, n72944, n72945, n72946,
    n72947, n72948, n72949, n72950, n72951, n72952, n72953, n72954, n72955,
    n72956, n72957, n72958, n72959, n72960, n72961, n72962, n72963, n72964,
    n72965, n72966, n72967, n72968, n72969, n72970, n72971, n72972, n72973,
    n72974, n72975, n72976, n72977, n72978, n72979, n72980, n72981, n72982,
    n72983, n72984, n72985, n72986, n72987, n72988, n72989, n72990, n72991,
    n72992, n72993, n72994, n72995, n72996, n72997, n72998, n72999, n73000,
    n73001, n73002, n73003, n73004, n73005, n73006, n73007, n73008, n73009,
    n73010, n73011, n73012, n73013, n73014, n73015, n73016, n73017, n73018,
    n73019, n73020, n73021, n73022, n73023, n73024, n73025, n73026, n73027,
    n73028, n73029, n73030, n73031, n73032, n73033, n73034, n73035, n73036,
    n73037, n73038, n73039, n73040, n73041, n73042, n73043, n73044, n73045,
    n73046, n73047, n73048, n73049, n73050, n73051, n73052, n73053, n73054,
    n73055, n73056, n73057, n73058, n73059, n73060, n73061, n73062, n73063,
    n73064, n73065, n73066, n73067, n73068, n73069, n73070, n73071, n73072,
    n73073, n73074, n73075, n73076, n73077, n73078, n73079, n73080, n73081,
    n73082, n73083, n73084, n73085, n73086, n73087, n73088, n73089, n73090,
    n73091, n73092, n73093, n73094, n73095, n73096, n73097, n73098, n73099,
    n73100, n73101, n73102, n73103, n73104, n73105, n73106, n73107, n73108,
    n73109, n73110, n73111, n73112, n73113, n73114, n73115, n73116, n73117,
    n73118, n73119, n73120, n73121, n73122, n73123, n73124, n73125, n73126,
    n73127, n73128, n73129, n73130, n73131, n73132, n73133, n73134, n73135,
    n73136, n73137, n73138, n73139, n73140, n73141, n73142, n73143, n73144,
    n73145, n73146, n73147, n73148, n73149, n73150, n73151, n73152, n73153,
    n73154, n73155, n73156, n73157, n73158, n73159, n73160, n73161, n73162,
    n73163, n73164, n73165, n73166, n73167, n73168, n73169, n73170, n73171,
    n73172, n73173, n73174, n73175, n73176, n73177, n73178, n73179, n73180,
    n73181, n73182, n73183, n73184, n73185, n73186, n73187, n73188, n73189,
    n73190, n73191, n73192, n73193, n73194, n73195, n73196, n73197, n73198,
    n73199, n73200, n73201, n73202, n73203, n73204, n73205, n73206, n73207,
    n73208, n73209, n73210, n73211, n73212, n73213, n73214, n73215, n73216,
    n73217, n73218, n73219, n73220, n73221, n73222, n73223, n73224, n73225,
    n73226, n73227, n73228, n73229, n73230, n73231, n73232, n73233, n73234,
    n73235, n73236, n73237, n73238, n73239, n73240, n73241, n73242, n73243,
    n73244, n73245, n73246, n73247, n73248, n73249, n73250, n73251, n73252,
    n73253, n73254, n73255, n73256, n73257, n73258, n73259, n73260, n73261,
    n73262, n73263, n73264, n73265, n73266, n73267, n73268, n73269, n73270,
    n73271, n73272, n73273, n73274, n73275, n73276, n73277, n73278, n73279,
    n73280, n73281, n73282, n73283, n73284, n73285, n73286, n73287, n73288,
    n73289, n73290, n73291, n73292, n73293, n73294, n73295, n73296, n73297,
    n73298, n73299, n73300, n73301, n73302, n73303, n73304, n73305, n73306,
    n73307, n73308, n73309, n73310, n73311, n73312, n73313, n73314, n73315,
    n73316, n73317, n73318, n73319, n73320, n73321, n73322, n73323, n73324,
    n73325, n73326, n73327, n73328, n73329, n73330, n73331, n73332, n73333,
    n73334, n73335, n73336, n73337, n73338, n73339, n73340, n73341, n73342,
    n73343, n73344, n73345, n73346, n73347, n73348, n73349, n73350, n73351,
    n73352, n73353, n73354, n73355, n73356, n73357, n73358, n73359, n73360,
    n73361, n73362, n73363, n73364, n73365, n73366, n73367, n73368, n73369,
    n73370, n73371, n73372, n73373, n73374, n73375, n73376, n73377, n73378,
    n73379, n73380, n73381, n73382, n73383, n73384, n73385, n73386, n73387,
    n73388, n73389, n73390, n73391, n73392, n73393, n73394, n73395, n73396,
    n73397, n73398, n73399, n73400, n73401, n73402, n73403, n73404, n73405,
    n73406, n73407, n73408, n73409, n73410, n73411, n73412, n73413, n73414,
    n73415, n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423,
    n73424, n73425, n73426, n73427, n73428, n73429, n73430, n73431, n73432,
    n73433, n73434, n73435, n73436, n73437, n73438, n73439, n73440, n73441,
    n73442, n73443, n73444, n73445, n73446, n73447, n73448, n73449, n73450,
    n73451, n73452, n73453, n73454, n73455, n73456, n73457, n73458, n73459,
    n73460, n73461, n73462, n73463, n73464, n73465, n73466, n73467, n73468,
    n73469, n73470, n73471, n73472, n73473, n73474, n73475, n73476, n73477,
    n73478, n73479, n73480, n73481, n73482, n73483, n73484, n73485, n73486,
    n73487, n73488, n73489, n73490, n73491, n73492, n73493, n73494, n73495,
    n73496, n73497, n73498, n73499, n73500, n73501, n73502, n73503, n73504,
    n73505, n73506, n73507, n73508, n73509, n73510, n73511, n73512, n73513,
    n73514, n73515, n73516, n73517, n73518, n73519, n73520, n73521, n73522,
    n73523, n73524, n73525, n73526, n73527, n73528, n73529, n73530, n73531,
    n73532, n73533, n73534, n73535, n73536, n73537, n73538, n73539, n73540,
    n73541, n73542, n73543, n73544, n73545, n73546, n73547, n73548, n73549,
    n73550, n73551, n73552, n73553, n73554, n73555, n73556, n73557, n73558,
    n73559, n73560, n73561, n73562, n73563, n73564, n73565, n73566, n73567,
    n73568, n73569, n73570, n73571, n73572, n73573, n73574, n73575, n73576,
    n73577, n73578, n73579, n73580, n73581, n73582, n73583, n73584, n73585,
    n73586, n73587, n73588, n73589, n73590, n73591, n73592, n73593, n73594,
    n73595, n73596, n73597, n73598, n73599, n73600, n73601, n73602, n73603,
    n73604, n73605, n73606, n73607, n73608, n73609, n73610, n73611, n73612,
    n73613, n73614, n73615, n73616, n73617, n73618, n73619, n73620, n73621,
    n73622, n73623, n73624, n73625, n73626, n73627, n73628, n73629, n73630,
    n73631, n73632, n73633, n73634, n73635, n73636, n73637, n73638, n73639,
    n73640, n73641, n73642, n73643, n73644, n73645, n73646, n73647, n73648,
    n73649, n73650, n73651, n73652, n73653, n73654, n73655, n73656, n73657,
    n73658, n73659, n73660, n73661, n73662, n73663, n73664, n73665, n73666,
    n73667, n73668, n73669, n73670, n73671, n73672, n73673, n73674, n73675,
    n73676, n73677, n73678, n73679, n73680, n73681, n73682, n73683, n73684,
    n73685, n73686, n73687, n73688, n73689, n73690, n73691, n73692, n73693,
    n73694, n73695, n73696, n73697, n73698, n73699, n73700, n73701, n73702,
    n73703, n73704, n73705, n73706, n73707, n73708, n73709, n73710, n73711,
    n73712, n73713, n73714, n73715, n73716, n73717, n73718, n73719, n73720,
    n73721, n73722, n73723, n73724, n73725, n73726, n73727, n73728, n73729,
    n73730, n73731, n73732, n73733, n73734, n73735, n73736, n73737, n73738,
    n73739, n73740, n73741, n73742, n73743, n73744, n73745, n73746, n73747,
    n73748, n73749, n73750, n73751, n73752, n73753, n73754, n73755, n73756,
    n73757, n73758, n73759, n73760, n73761, n73762, n73763, n73764, n73765,
    n73766, n73767, n73768, n73769, n73770, n73771, n73772, n73773, n73774,
    n73775, n73776, n73777, n73778, n73779, n73780, n73781, n73782, n73783,
    n73784, n73785, n73786, n73787, n73788, n73789, n73790, n73791, n73792,
    n73793, n73794, n73795, n73796, n73797, n73798, n73799, n73800, n73801,
    n73802, n73803, n73804, n73805, n73806, n73807, n73808, n73809, n73810,
    n73811, n73812, n73813, n73814, n73815, n73816, n73817, n73818, n73819,
    n73820, n73821, n73822, n73823, n73824, n73825, n73826, n73827, n73828,
    n73829, n73830, n73831, n73832, n73833, n73834, n73835, n73836, n73837,
    n73838, n73839, n73840, n73841, n73842, n73843, n73844, n73845, n73846,
    n73847, n73848, n73849, n73850, n73851, n73852, n73853, n73854, n73855,
    n73856, n73857, n73858, n73859, n73860, n73861, n73862, n73863, n73864,
    n73865, n73866, n73867, n73868, n73869, n73870, n73871, n73872, n73873,
    n73874, n73875, n73876, n73877, n73878, n73879, n73880, n73881, n73882,
    n73883, n73884, n73885, n73886, n73887, n73888, n73889, n73890, n73891,
    n73892, n73893, n73894, n73895, n73896, n73897, n73898, n73899, n73900,
    n73901, n73902, n73903, n73904, n73905, n73906, n73907, n73908, n73909,
    n73910, n73911, n73912, n73913, n73914, n73915, n73916, n73917, n73918,
    n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927,
    n73928, n73929, n73930, n73931, n73932, n73933, n73934, n73935, n73936,
    n73937, n73938, n73939, n73940, n73941, n73942, n73943, n73944, n73945,
    n73946, n73947, n73948, n73949, n73950, n73951, n73952, n73953, n73954,
    n73955, n73956, n73957, n73958, n73959, n73960, n73961, n73962, n73963,
    n73964, n73965, n73966, n73967, n73968, n73969, n73970, n73971, n73972,
    n73973, n73974, n73975, n73976, n73977, n73978, n73979, n73980, n73981,
    n73982, n73983, n73984, n73985, n73986, n73987, n73988, n73989, n73990,
    n73991, n73992, n73993, n73994, n73995, n73996, n73997, n73998, n73999,
    n74000, n74001, n74002, n74003, n74004, n74005, n74006, n74007, n74008,
    n74009, n74010, n74011, n74012, n74013, n74014, n74015, n74016, n74017,
    n74018, n74019, n74020, n74021, n74022, n74023, n74024, n74025, n74026,
    n74027, n74028, n74029, n74030, n74031, n74032, n74033, n74034, n74035,
    n74036, n74037, n74038, n74039, n74040, n74041, n74042, n74043, n74044,
    n74045, n74046, n74047, n74048, n74049, n74050, n74051, n74052, n74053,
    n74054, n74055, n74056, n74057, n74058, n74059, n74060, n74061, n74062,
    n74063, n74064, n74065, n74066, n74067, n74068, n74069, n74070, n74071,
    n74072, n74073, n74074, n74075, n74076, n74077, n74078, n74079, n74080,
    n74081, n74082, n74083, n74084, n74085, n74086, n74087, n74088, n74089,
    n74090, n74091, n74092, n74093, n74094, n74095, n74096, n74097, n74098,
    n74099, n74100, n74101, n74102, n74103, n74104, n74105, n74106, n74107,
    n74108, n74109, n74110, n74111, n74112, n74113, n74114, n74115, n74116,
    n74117, n74118, n74119, n74120, n74121, n74122, n74123, n74124, n74125,
    n74126, n74127, n74128, n74129, n74130, n74131, n74132, n74133, n74134,
    n74135, n74136, n74137, n74138, n74139, n74140, n74141, n74142, n74143,
    n74144, n74145, n74146, n74147, n74148, n74149, n74150, n74151, n74152,
    n74153, n74154, n74155, n74156, n74157, n74158, n74159, n74160, n74161,
    n74162, n74163, n74164, n74165, n74166, n74167, n74168, n74169, n74170,
    n74171, n74172, n74173, n74174, n74175, n74176, n74177, n74178, n74179,
    n74180, n74181, n74182, n74183, n74184, n74185, n74186, n74187, n74188,
    n74189, n74190, n74191, n74192, n74193, n74194, n74195, n74196, n74197,
    n74198, n74199, n74200, n74201, n74202, n74203, n74204, n74205, n74206,
    n74207, n74208, n74209, n74210, n74211, n74212, n74213, n74214, n74215,
    n74216, n74217, n74218, n74219, n74220, n74221, n74222, n74223, n74224,
    n74225, n74226, n74227, n74228, n74229, n74230, n74231, n74232, n74233,
    n74234, n74235, n74236, n74237, n74238, n74239, n74240, n74241, n74242,
    n74243, n74244, n74245, n74246, n74247, n74248, n74249, n74250, n74251,
    n74252, n74253, n74254, n74255, n74256, n74257, n74258, n74259, n74260,
    n74261, n74262, n74263, n74264, n74265, n74266, n74267, n74268, n74269,
    n74270, n74271, n74272, n74273, n74274, n74275, n74276, n74277, n74278,
    n74279, n74280, n74281, n74282, n74283, n74284, n74285, n74286, n74287,
    n74288, n74289, n74290, n74291, n74292, n74293, n74294, n74295, n74296,
    n74297, n74298, n74299, n74300, n74301, n74302, n74303, n74304, n74305,
    n74306, n74307, n74308, n74309, n74310, n74311, n74312, n74313, n74314,
    n74315, n74316, n74317, n74318, n74319, n74320, n74321, n74322, n74323,
    n74324, n74325, n74326, n74327, n74328, n74329, n74330, n74331, n74332,
    n74333, n74334, n74335, n74336, n74337, n74338, n74339, n74340, n74341,
    n74342, n74343, n74344, n74345, n74346, n74347, n74348, n74349, n74350,
    n74351, n74352, n74353, n74354, n74355, n74356, n74357, n74358, n74359,
    n74360, n74361, n74362, n74363, n74364, n74365, n74366, n74367, n74368,
    n74369, n74370, n74371, n74372, n74373, n74374, n74375, n74376, n74377,
    n74378, n74379, n74380, n74381, n74382, n74383, n74384, n74385, n74386,
    n74387, n74388, n74389, n74390, n74391, n74392, n74393, n74394, n74395,
    n74396, n74397, n74398, n74399, n74400, n74401, n74402, n74403, n74404,
    n74405, n74406, n74407, n74408, n74409, n74410, n74411, n74412, n74413,
    n74414, n74415, n74416, n74417, n74418, n74419, n74420, n74421, n74422,
    n74423, n74424, n74425, n74426, n74427, n74428, n74429, n74430, n74431,
    n74432, n74433, n74434, n74435, n74436, n74437, n74438, n74439, n74440,
    n74441, n74442, n74443, n74444, n74445, n74446, n74447, n74448, n74449,
    n74450, n74451, n74452, n74453, n74454, n74455, n74456, n74457, n74458,
    n74459, n74460, n74461, n74462, n74463, n74464, n74465, n74466, n74467,
    n74468, n74469, n74470, n74471, n74472, n74473, n74474, n74475, n74476,
    n74477, n74478, n74479, n74480, n74481, n74482, n74483, n74484, n74485,
    n74486, n74487, n74488, n74489, n74490, n74491, n74492, n74493, n74494,
    n74495, n74496, n74497, n74498, n74499, n74500, n74501, n74502, n74503,
    n74504, n74505, n74506, n74507, n74508, n74509, n74510, n74511, n74512,
    n74513, n74514, n74515, n74516, n74517, n74518, n74519, n74520, n74521,
    n74522, n74523, n74524, n74525, n74526, n74527, n74528, n74529, n74530,
    n74531, n74532, n74533, n74534, n74535, n74536, n74537, n74538, n74539,
    n74540, n74541, n74542, n74543, n74544, n74545, n74546, n74547, n74548,
    n74549, n74550, n74551, n74552, n74553, n74554, n74555, n74556, n74557,
    n74558, n74559, n74560, n74561, n74562, n74563, n74564, n74565, n74566,
    n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574, n74575,
    n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583, n74584,
    n74585, n74586, n74587, n74588, n74589, n74590, n74591, n74592, n74593,
    n74594, n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602,
    n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610, n74611,
    n74612, n74613, n74614, n74615, n74616, n74617, n74618, n74619, n74620,
    n74621, n74622, n74623, n74624, n74625, n74626, n74627, n74628, n74629,
    n74630, n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638,
    n74639, n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647,
    n74648, n74649, n74650, n74651, n74652, n74653, n74654, n74655, n74656,
    n74657, n74658, n74659, n74660, n74661, n74662, n74663, n74664, n74665,
    n74666, n74667, n74668, n74669, n74670, n74671, n74672, n74673, n74674,
    n74675, n74676, n74677, n74678, n74679, n74680, n74681, n74682, n74683,
    n74684, n74685, n74686, n74687, n74688, n74689, n74690, n74691, n74692,
    n74693, n74694, n74695, n74696, n74697, n74698, n74699, n74700, n74701,
    n74702, n74703, n74704, n74705, n74706, n74707, n74708, n74709, n74710,
    n74711, n74712, n74713, n74714, n74715, n74716, n74717, n74718, n74719,
    n74720, n74721, n74722, n74723, n74724, n74725, n74726, n74727, n74728,
    n74729, n74730, n74731, n74732, n74733, n74734, n74735, n74736, n74737,
    n74738, n74739, n74740, n74741, n74742, n74743, n74744, n74745, n74746,
    n74747, n74748, n74749, n74750, n74751, n74752, n74753, n74754, n74755,
    n74756, n74757, n74758, n74759, n74760, n74761, n74762, n74763, n74764,
    n74765, n74766, n74767, n74768, n74769, n74770, n74771, n74772, n74773,
    n74774, n74775, n74776, n74777, n74778, n74779, n74780, n74781, n74782,
    n74783, n74784, n74785, n74786, n74787, n74788, n74789, n74790, n74791,
    n74792, n74793, n74794, n74795, n74796, n74797, n74798, n74799, n74800,
    n74801, n74802, n74803, n74804, n74805, n74806, n74807, n74808, n74809,
    n74810, n74811, n74812, n74813, n74814, n74815, n74816, n74817, n74818,
    n74819, n74820, n74821, n74822, n74823, n74824, n74825, n74826, n74827,
    n74828, n74829, n74830, n74831, n74832, n74833, n74834, n74835, n74836,
    n74837, n74838, n74839, n74840, n74841, n74842, n74843, n74844, n74845,
    n74846, n74847, n74848, n74849, n74850, n74851, n74852, n74853, n74854,
    n74855, n74856, n74857, n74858, n74859, n74860, n74861, n74862, n74863,
    n74864, n74865, n74866, n74867, n74868, n74869, n74870, n74871, n74872,
    n74873, n74874, n74875, n74876, n74877, n74878, n74879, n74880, n74881,
    n74882, n74883, n74884, n74885, n74886, n74887, n74888, n74889, n74890,
    n74891, n74892, n74893, n74894, n74895, n74896, n74897, n74898, n74899,
    n74900, n74901, n74902, n74903, n74904, n74905, n74906, n74907, n74908,
    n74909, n74910, n74911, n74912, n74913, n74914, n74915, n74916, n74917,
    n74918, n74919, n74920, n74921, n74922, n74923, n74924, n74925, n74926,
    n74927, n74928, n74929, n74930, n74931, n74932, n74933, n74934, n74935,
    n74936, n74937, n74938, n74939, n74940, n74941, n74942, n74943, n74944,
    n74945, n74946, n74947, n74948, n74949, n74950, n74951, n74952, n74953,
    n74954, n74955, n74956, n74957, n74958, n74959, n74960, n74961, n74962,
    n74963, n74964, n74965, n74966, n74967, n74968, n74969, n74970, n74971,
    n74972, n74973, n74974, n74975, n74976, n74977, n74978, n74979, n74980,
    n74981, n74982, n74983, n74984, n74985, n74986, n74987, n74988, n74989,
    n74990, n74991, n74992, n74993, n74994, n74995, n74996, n74997, n74998,
    n74999, n75000, n75001, n75002, n75003, n75004, n75005, n75006, n75007,
    n75008, n75009, n75010, n75011, n75012, n75013, n75014, n75015, n75016,
    n75017, n75018, n75019, n75020, n75021, n75022, n75023, n75024, n75025,
    n75026, n75027, n75028, n75029, n75030, n75031, n75032, n75033, n75034,
    n75035, n75036, n75037, n75038, n75039, n75040, n75041, n75042, n75043,
    n75044, n75045, n75046, n75047, n75048, n75049, n75050, n75051, n75052,
    n75053, n75054, n75055, n75056, n75057, n75058, n75059, n75060, n75061,
    n75062, n75063, n75064, n75065, n75066, n75067, n75068, n75069, n75070,
    n75071, n75072, n75073, n75074, n75075, n75076, n75077, n75078, n75079,
    n75080, n75081, n75082, n75083, n75084, n75085, n75086, n75087, n75088,
    n75089, n75090, n75091, n75092, n75093, n75094, n75095, n75096, n75097,
    n75098, n75099, n75100, n75101, n75102, n75103, n75104, n75105, n75106,
    n75107, n75108, n75109, n75110, n75111, n75112, n75113, n75114, n75115,
    n75116, n75117, n75118, n75119, n75120, n75121, n75122, n75123, n75124,
    n75125, n75126, n75127, n75128, n75129, n75130, n75131, n75132, n75133,
    n75134, n75135, n75136, n75137, n75138, n75139, n75140, n75141, n75142,
    n75143, n75144, n75145, n75146, n75147, n75148, n75149, n75150, n75151,
    n75152, n75153, n75154, n75155, n75156, n75157, n75158, n75159, n75160,
    n75161, n75162, n75163, n75164, n75165, n75166, n75167, n75168, n75169,
    n75170, n75171, n75172, n75173, n75174, n75175, n75176, n75177, n75178,
    n75179, n75180, n75181, n75182, n75183, n75184, n75185, n75186, n75187,
    n75188, n75189, n75190, n75191, n75192, n75193, n75194, n75195, n75196,
    n75197, n75198, n75199, n75200, n75201, n75202, n75203, n75204, n75205,
    n75206, n75207, n75208, n75209, n75210, n75211, n75212, n75213, n75214,
    n75215, n75216, n75217, n75218, n75219, n75220, n75221, n75222, n75223,
    n75224, n75225, n75226, n75227, n75228, n75229, n75230, n75231, n75232,
    n75233, n75234, n75235, n75236, n75237, n75238, n75239, n75240, n75241,
    n75242, n75243, n75244, n75245, n75246, n75247, n75248, n75249, n75250,
    n75251, n75252, n75253, n75254, n75255, n75256, n75257, n75258, n75259,
    n75260, n75261, n75262, n75263, n75264, n75265, n75266, n75267, n75268,
    n75269, n75270, n75271, n75272, n75273, n75274, n75275, n75276, n75277,
    n75278, n75279, n75280, n75281, n75282, n75283, n75284, n75285, n75286,
    n75287, n75288, n75289, n75290, n75291, n75292, n75293, n75294, n75295,
    n75296, n75297, n75298, n75299, n75300, n75301, n75302, n75303, n75304,
    n75305, n75306, n75307, n75308, n75309, n75310, n75311, n75312, n75313,
    n75314, n75315, n75316, n75317, n75318, n75319, n75320, n75321, n75322,
    n75323, n75324, n75325, n75326, n75327, n75328, n75329, n75330, n75331,
    n75332, n75333, n75334, n75335, n75336, n75337, n75338, n75339, n75340,
    n75341, n75342, n75343, n75344, n75345, n75346, n75347, n75348, n75349,
    n75350, n75351, n75352, n75353, n75354, n75355, n75356, n75357, n75358,
    n75359, n75360, n75361, n75362, n75363, n75364, n75365, n75366, n75367,
    n75368, n75369, n75370, n75371, n75372, n75373, n75374, n75375, n75376,
    n75377, n75378, n75379, n75380, n75381, n75382, n75383, n75384, n75385,
    n75386, n75387, n75388, n75389, n75390, n75391, n75392, n75393, n75394,
    n75395, n75396, n75397, n75398, n75399, n75400, n75401, n75402, n75403,
    n75404, n75405, n75406, n75407, n75408, n75409, n75410, n75411, n75412,
    n75413, n75414, n75415, n75416, n75417, n75418, n75419, n75420, n75421,
    n75422, n75423, n75424, n75425, n75426, n75427, n75428, n75429, n75430,
    n75431, n75432, n75433, n75434, n75435, n75436, n75437, n75438, n75439,
    n75440, n75441, n75442, n75443, n75444, n75445, n75446, n75447, n75448,
    n75449, n75450, n75451, n75452, n75453, n75454, n75455, n75456, n75457,
    n75458, n75459, n75460, n75461, n75462, n75463, n75464, n75465, n75466,
    n75467, n75468, n75469, n75470, n75471, n75472, n75473, n75474, n75475,
    n75476, n75477, n75478, n75479, n75480, n75481, n75482, n75483, n75484,
    n75485, n75486, n75487, n75488, n75489, n75490, n75491, n75492, n75493,
    n75494, n75495, n75496, n75497, n75498, n75499, n75500, n75501, n75502,
    n75503, n75504, n75505, n75506, n75507, n75508, n75509, n75510, n75511,
    n75512, n75513, n75514, n75515, n75516, n75517, n75518, n75519, n75520,
    n75521, n75522, n75523, n75524, n75525, n75526, n75527, n75528, n75529,
    n75530, n75531, n75532, n75533, n75534, n75535, n75536, n75537, n75538,
    n75539, n75540, n75541, n75542, n75543, n75544, n75545, n75546, n75547,
    n75548, n75549, n75550, n75551, n75552, n75553, n75554, n75555, n75556,
    n75557, n75558, n75559, n75560, n75561, n75562, n75563, n75564, n75565,
    n75566, n75567, n75568, n75569, n75570, n75571, n75572, n75573, n75574,
    n75575, n75576, n75577, n75578, n75579, n75580, n75581, n75582, n75583,
    n75584, n75585, n75586, n75587, n75588, n75589, n75590, n75591, n75592,
    n75593, n75594, n75595, n75596, n75597, n75598, n75599, n75600, n75601,
    n75602, n75603, n75604, n75605, n75606, n75607, n75608, n75609, n75610,
    n75611, n75612, n75613, n75614, n75615, n75616, n75617, n75618, n75619,
    n75620, n75621, n75622, n75623, n75624, n75625, n75626, n75627, n75628,
    n75629, n75630, n75631, n75632, n75633, n75634, n75635, n75636, n75637,
    n75638, n75639, n75640, n75641, n75642, n75643, n75644, n75645, n75646,
    n75647, n75648, n75649, n75650, n75651, n75652, n75653, n75654, n75655,
    n75656, n75657, n75658, n75659, n75660, n75661, n75662, n75663, n75664,
    n75665, n75666, n75667, n75668, n75669, n75670, n75671, n75672, n75673,
    n75674, n75675, n75676, n75677, n75678, n75679, n75680, n75681, n75682,
    n75683, n75684, n75685, n75686, n75687, n75688, n75689, n75690, n75691,
    n75692, n75693, n75694, n75695, n75696, n75697, n75698, n75699, n75700,
    n75701, n75702, n75703, n75704, n75705, n75706, n75707, n75708, n75709,
    n75710, n75711, n75712, n75713, n75714, n75715, n75716, n75717, n75718,
    n75719, n75720, n75721, n75722, n75723, n75724, n75725, n75726, n75727,
    n75728, n75729, n75730, n75731, n75732, n75733, n75734, n75735, n75736,
    n75737, n75738, n75739, n75740, n75741, n75742, n75743, n75744, n75745,
    n75746, n75747, n75748, n75749, n75750, n75751, n75752, n75753, n75754,
    n75755, n75756, n75757, n75758, n75759, n75760, n75761, n75762, n75763,
    n75764, n75765, n75766, n75767, n75768, n75769, n75770, n75771, n75772,
    n75773, n75774, n75775, n75776, n75777, n75778, n75779, n75780, n75781,
    n75782, n75783, n75784, n75785, n75786, n75787, n75788, n75789, n75790,
    n75791, n75792, n75793, n75794, n75795, n75796, n75797, n75798, n75799,
    n75800, n75801, n75802, n75803, n75804, n75805, n75806, n75807, n75808,
    n75809, n75810, n75811, n75812, n75813, n75814, n75815, n75816, n75817,
    n75818, n75819, n75820, n75821, n75822, n75823, n75824, n75825, n75826,
    n75827, n75828, n75829, n75830, n75831, n75832, n75833, n75834, n75835,
    n75836, n75837, n75838, n75839, n75840, n75841, n75842, n75843, n75844,
    n75845, n75846, n75847, n75848, n75849, n75850, n75851, n75852, n75853,
    n75854, n75855, n75856, n75857, n75858, n75859, n75860, n75861, n75862,
    n75863, n75864, n75865, n75866, n75867, n75868, n75869, n75870, n75871,
    n75872, n75873, n75874, n75875, n75876, n75877, n75878, n75879, n75880,
    n75881, n75882, n75883, n75884, n75885, n75886, n75887, n75888, n75889,
    n75890, n75891, n75892, n75893, n75894, n75895, n75896, n75897, n75898,
    n75899, n75900, n75901, n75902, n75903, n75904, n75905, n75906, n75907,
    n75908, n75909, n75910, n75911, n75912, n75913, n75914, n75915, n75916,
    n75917, n75918, n75919, n75920, n75921, n75922, n75923, n75924, n75925,
    n75926, n75927, n75928, n75929, n75930, n75931, n75932, n75933, n75934,
    n75935, n75936, n75937, n75938, n75939, n75940, n75941, n75942, n75943,
    n75944, n75945, n75946, n75947, n75948, n75949, n75950, n75951, n75952,
    n75953, n75954, n75955, n75956, n75957, n75958, n75959, n75960, n75961,
    n75962, n75963, n75964, n75965, n75966, n75967, n75968, n75969, n75970,
    n75971, n75972, n75973, n75974, n75975, n75976, n75977, n75978, n75979,
    n75980, n75981, n75982, n75983, n75984, n75985, n75986, n75987, n75988,
    n75989, n75990, n75991, n75992, n75993, n75994, n75995, n75996, n75997,
    n75998, n75999, n76000, n76001, n76002, n76003, n76004, n76005, n76006,
    n76007, n76008, n76009, n76010, n76011, n76012, n76013, n76014, n76015,
    n76016, n76017, n76018, n76019, n76020, n76021, n76022, n76023, n76024,
    n76025, n76026, n76027, n76028, n76029, n76030, n76031, n76032, n76033,
    n76034, n76035, n76036, n76037, n76038, n76039, n76040, n76041, n76042,
    n76043, n76044, n76045, n76046, n76047, n76048, n76049, n76050, n76051,
    n76052, n76053, n76054, n76055, n76056, n76057, n76058, n76059, n76060,
    n76061, n76062, n76063, n76064, n76065, n76066, n76067, n76068, n76069,
    n76070, n76071, n76072, n76073, n76074, n76075, n76076, n76077, n76078,
    n76079, n76080, n76081, n76082, n76083, n76084, n76085, n76086, n76087,
    n76088, n76089, n76090, n76091, n76092, n76093, n76094, n76095, n76096,
    n76097, n76098, n76099, n76100, n76101, n76102, n76103, n76104, n76105,
    n76106, n76107, n76108, n76109, n76110, n76111, n76112, n76113, n76114,
    n76115, n76116, n76117, n76118, n76119, n76120, n76121, n76122, n76123,
    n76124, n76125, n76126, n76127, n76128, n76129, n76130, n76131, n76132,
    n76133, n76134, n76135, n76136, n76137, n76138, n76139, n76140, n76141,
    n76142, n76143, n76144, n76145, n76146, n76147, n76148, n76149, n76150,
    n76151, n76152, n76153, n76154, n76155, n76156, n76157, n76158, n76159,
    n76160, n76161, n76162, n76163, n76164, n76165, n76166, n76167, n76168,
    n76169, n76170, n76171, n76172, n76173, n76174, n76175, n76176, n76177,
    n76178, n76179, n76180, n76181, n76182, n76183, n76184, n76185, n76186,
    n76187, n76188, n76189, n76190, n76191, n76192, n76193, n76194, n76195,
    n76196, n76197, n76198, n76199, n76200, n76201, n76202, n76203, n76204,
    n76205, n76206, n76207, n76208, n76209, n76210, n76211, n76212, n76213,
    n76214, n76215, n76216, n76217, n76218, n76219, n76220, n76221, n76222,
    n76223, n76224, n76225, n76226, n76227, n76228, n76229, n76230, n76231,
    n76232, n76233, n76234, n76235, n76236, n76237, n76238, n76239, n76240,
    n76241, n76242, n76243, n76244, n76245, n76246, n76247, n76248, n76249,
    n76250, n76251, n76252, n76253, n76254, n76255, n76256, n76257, n76258,
    n76259, n76260, n76261, n76262, n76263, n76264, n76265, n76266, n76267,
    n76268, n76269, n76270, n76271, n76272, n76273, n76274, n76275, n76276,
    n76277, n76278, n76279, n76280, n76281, n76282, n76283, n76284, n76285,
    n76286, n76287, n76288, n76289, n76290, n76291, n76292, n76293, n76294,
    n76295, n76296, n76297, n76298, n76299, n76300, n76301, n76302, n76303,
    n76304, n76305, n76306, n76307, n76308, n76309, n76310, n76311, n76312,
    n76313, n76314, n76315, n76316, n76317, n76318, n76319, n76320, n76321,
    n76322, n76323, n76324, n76325, n76326, n76327, n76328, n76329, n76330,
    n76331, n76332, n76333, n76334, n76335, n76336, n76337, n76338, n76339,
    n76340, n76341, n76342, n76343, n76344, n76345, n76346, n76347, n76348,
    n76349, n76350, n76351, n76352, n76353, n76354, n76355, n76356, n76357,
    n76358, n76359, n76360, n76361, n76362, n76363, n76364, n76365, n76366,
    n76367, n76368, n76369, n76370, n76371, n76372, n76373, n76374, n76375,
    n76376, n76377, n76378, n76379, n76380, n76381, n76382, n76383, n76384,
    n76385, n76386, n76387, n76388, n76389, n76390, n76391, n76392, n76393,
    n76394, n76395, n76396, n76397, n76398, n76399, n76400, n76401, n76402,
    n76403, n76404, n76405, n76406, n76407, n76408, n76409, n76410, n76411,
    n76412, n76413, n76414, n76415, n76416, n76417, n76418, n76419, n76420,
    n76421, n76422, n76423, n76424, n76425, n76426, n76427, n76428, n76429,
    n76430, n76431, n76432, n76433, n76434, n76435, n76436, n76437, n76438,
    n76439, n76440, n76441, n76442, n76443, n76444, n76445, n76446, n76447,
    n76448, n76449, n76450, n76451, n76452, n76453, n76454, n76455, n76456,
    n76457, n76458, n76459, n76460, n76461, n76462, n76463, n76464, n76465,
    n76466, n76467, n76468, n76469, n76470, n76471, n76472, n76473, n76474,
    n76475, n76476, n76477, n76478, n76479, n76480, n76481, n76482, n76483,
    n76484, n76485, n76486, n76487, n76488, n76489, n76490, n76491, n76492,
    n76493, n76494, n76495, n76496, n76497, n76498, n76499, n76500, n76501,
    n76502, n76503, n76504, n76505, n76506, n76507, n76508, n76509, n76510,
    n76511, n76512, n76513, n76514, n76515, n76516, n76517, n76518, n76519,
    n76520, n76521, n76522, n76523, n76524, n76525, n76526, n76527, n76528,
    n76529, n76530, n76531, n76532, n76533, n76534, n76535, n76536, n76537,
    n76538, n76539, n76540, n76541, n76542, n76543, n76544, n76545, n76546,
    n76547, n76548, n76549, n76550, n76551, n76552, n76553, n76554, n76555,
    n76556, n76557, n76558, n76559, n76560, n76561, n76562, n76563, n76564,
    n76565, n76566, n76567, n76568, n76569, n76570, n76571, n76572, n76573,
    n76574, n76575, n76576, n76577, n76578, n76579, n76580, n76581, n76582,
    n76583, n76584, n76585, n76586, n76587, n76588, n76589, n76590, n76591,
    n76592, n76593, n76594, n76595, n76596, n76597, n76598, n76599, n76600,
    n76601, n76602, n76603, n76604, n76605, n76606, n76607, n76608, n76609,
    n76610, n76611, n76612, n76613, n76614, n76615, n76616, n76617, n76618,
    n76619, n76620, n76621, n76622, n76623, n76624, n76625, n76626, n76627,
    n76628, n76629, n76630, n76631, n76632, n76633, n76634, n76635, n76636,
    n76637, n76638, n76639, n76640, n76641, n76642, n76643, n76644, n76645,
    n76646, n76647, n76648, n76649, n76650, n76651, n76652, n76653, n76654,
    n76655, n76656, n76657, n76658, n76659, n76660, n76661, n76662, n76663,
    n76664, n76665, n76666, n76667, n76668, n76669, n76670, n76671, n76672,
    n76673, n76674, n76675, n76676, n76677, n76678, n76679, n76680, n76681,
    n76682, n76683, n76684, n76685, n76686, n76687, n76688, n76689, n76690,
    n76691, n76692, n76693, n76694, n76695, n76696, n76697, n76698, n76699,
    n76700, n76701, n76702, n76703, n76704, n76705, n76706, n76707, n76708,
    n76709, n76710, n76711, n76712, n76713, n76714, n76715, n76716, n76717,
    n76718, n76719, n76720, n76721, n76722, n76723, n76724, n76725, n76726,
    n76727, n76728, n76729, n76730, n76731, n76732, n76733, n76734, n76735,
    n76736, n76737, n76738, n76739, n76740, n76741, n76742, n76743, n76744,
    n76745, n76746, n76747, n76748, n76749, n76750, n76751, n76752, n76753,
    n76754, n76755, n76756, n76757, n76758, n76759, n76760, n76761, n76762,
    n76763, n76764, n76765, n76766, n76767, n76768, n76769, n76770, n76771,
    n76772, n76773, n76774, n76775, n76776, n76777, n76778, n76779, n76780,
    n76781, n76782, n76783, n76784, n76785, n76786, n76787, n76788, n76789,
    n76790, n76791, n76792, n76793, n76794, n76795, n76796, n76797, n76798,
    n76799, n76800, n76801, n76802, n76803, n76804, n76805, n76806, n76807,
    n76808, n76809, n76810, n76811, n76812, n76813, n76814, n76815, n76816,
    n76817, n76818, n76819, n76820, n76821, n76822, n76823, n76824, n76825,
    n76826, n76827, n76828, n76829, n76830, n76831, n76832, n76833, n76834,
    n76835, n76836, n76837, n76838, n76839, n76840, n76841, n76842, n76843,
    n76844, n76845, n76846, n76847, n76848, n76849, n76850, n76851, n76852,
    n76853, n76854, n76855, n76856, n76857, n76858, n76859, n76860, n76861,
    n76862, n76863, n76864, n76865, n76866, n76867, n76868, n76869, n76870,
    n76871, n76872, n76873, n76874, n76875, n76876, n76877, n76878, n76879,
    n76880, n76881, n76882, n76883, n76884, n76885, n76886, n76887, n76888,
    n76889, n76890, n76891, n76892, n76893, n76894, n76895, n76896, n76897,
    n76898, n76899, n76900, n76901, n76902, n76903, n76904, n76905, n76906,
    n76907, n76908, n76909, n76910, n76911, n76912, n76913, n76914, n76915,
    n76916, n76917, n76918, n76919, n76920, n76921, n76922, n76923, n76924,
    n76925, n76926, n76927, n76928, n76929, n76930, n76931, n76932, n76933,
    n76934, n76935, n76936, n76937, n76938, n76939, n76940, n76941, n76942,
    n76943, n76944, n76945, n76946, n76947, n76948, n76949, n76950, n76951,
    n76952, n76953, n76954, n76955, n76956, n76957, n76958, n76959, n76960,
    n76961, n76962, n76963, n76964, n76965, n76966, n76967, n76968, n76969,
    n76970, n76971, n76972, n76973, n76974, n76975, n76976, n76977, n76978,
    n76979, n76980, n76981, n76982, n76983, n76984, n76985, n76986, n76987,
    n76988, n76989, n76990, n76991, n76992, n76993, n76994, n76995, n76996,
    n76997, n76998, n76999, n77000, n77001, n77002, n77003, n77004, n77005,
    n77006, n77007, n77008, n77009, n77010, n77011, n77012, n77013, n77014,
    n77015, n77016, n77017, n77018, n77019, n77020, n77021, n77022, n77023,
    n77024, n77025, n77026, n77027, n77028, n77029, n77030, n77031, n77032,
    n77033, n77034, n77035, n77036, n77037, n77038, n77039, n77040, n77041,
    n77042, n77043, n77044, n77045, n77046, n77047, n77048, n77049, n77050,
    n77051, n77052, n77053, n77054, n77055, n77056, n77057, n77058, n77059,
    n77060, n77061, n77062, n77063, n77064, n77065, n77066, n77067, n77068,
    n77069, n77070, n77071, n77072, n77073, n77074, n77075, n77076, n77077,
    n77078, n77079, n77080, n77081, n77082, n77083, n77084, n77085, n77086,
    n77087, n77088, n77089, n77090, n77091, n77092, n77093, n77094, n77095,
    n77096, n77097, n77098, n77099, n77100, n77101, n77102, n77103, n77104,
    n77105, n77106, n77107, n77108, n77109, n77110, n77111, n77112, n77113,
    n77114, n77115, n77116, n77117, n77118, n77119, n77120, n77121, n77122,
    n77123, n77124, n77125, n77126, n77127, n77128, n77129, n77130, n77131,
    n77132, n77133, n77134, n77135, n77136, n77137, n77138, n77139, n77140,
    n77141, n77142, n77143, n77144, n77145, n77146, n77147, n77148, n77149,
    n77150, n77151, n77152, n77153, n77154, n77155, n77156, n77157, n77158,
    n77159, n77160, n77161, n77162, n77163, n77164, n77165, n77166, n77167,
    n77168, n77169, n77170, n77171, n77172, n77173, n77174, n77175, n77176,
    n77177, n77178, n77179, n77180, n77181, n77182, n77183, n77184, n77185,
    n77186, n77187, n77188, n77189, n77190, n77191, n77192, n77193, n77194,
    n77195, n77196, n77197, n77198, n77199, n77200, n77201, n77202, n77203,
    n77204, n77205, n77206, n77207, n77208, n77209, n77210, n77211, n77212,
    n77213, n77214, n77215, n77216, n77217, n77218, n77219, n77220, n77221,
    n77222, n77223, n77224, n77225, n77226, n77227, n77228, n77229, n77230,
    n77231, n77232, n77233, n77234, n77235, n77236, n77237, n77238, n77239,
    n77240, n77241, n77242, n77243, n77244, n77245, n77246, n77247, n77248,
    n77249, n77250, n77251, n77252, n77253, n77254, n77255, n77256, n77257,
    n77258, n77259, n77260, n77261, n77262, n77263, n77264, n77265, n77266,
    n77267, n77268, n77269, n77270, n77271, n77272, n77273, n77274, n77275,
    n77276, n77277, n77278, n77279, n77280, n77281, n77282, n77283, n77284,
    n77285, n77286, n77287, n77288, n77289, n77290, n77291, n77292, n77293,
    n77294, n77295, n77296, n77297, n77298, n77299, n77300, n77301, n77302,
    n77303, n77304, n77305, n77306, n77307, n77308, n77309, n77310, n77311,
    n77312, n77313, n77314, n77315, n77316, n77317, n77318, n77319, n77320,
    n77321, n77322, n77323, n77324, n77325, n77326, n77327, n77328, n77329,
    n77330, n77331, n77332, n77333, n77334, n77335, n77336, n77337, n77338,
    n77339, n77340, n77341, n77342, n77343, n77344, n77345, n77346, n77347,
    n77348, n77349, n77350, n77351, n77352, n77353, n77354, n77355, n77356,
    n77357, n77358, n77359, n77360, n77361, n77362, n77363, n77364, n77365,
    n77366, n77367, n77368, n77369, n77370, n77371, n77372, n77373, n77374,
    n77375, n77376, n77377, n77378, n77379, n77380, n77381, n77382, n77383,
    n77384, n77385, n77386, n77387, n77388, n77389, n77390, n77391, n77392,
    n77393, n77394, n77395, n77396, n77397, n77398, n77399, n77400, n77401,
    n77402, n77403, n77404, n77405, n77406, n77407, n77408, n77409, n77410,
    n77411, n77412, n77413, n77414, n77415, n77416, n77417, n77418, n77419,
    n77420, n77421, n77422, n77423, n77424, n77425, n77426, n77427, n77428,
    n77429, n77430, n77431, n77432, n77433, n77434, n77435, n77436, n77437,
    n77438, n77439, n77440, n77441, n77442, n77443, n77444, n77445, n77446,
    n77447, n77448, n77449, n77450, n77451, n77452, n77453, n77454, n77455,
    n77456, n77457, n77458, n77459, n77460, n77461, n77462, n77463, n77464,
    n77465, n77466, n77467, n77468, n77469, n77470, n77471, n77472, n77473,
    n77474, n77475, n77476, n77477, n77478, n77479, n77480, n77481, n77482,
    n77483, n77484, n77485, n77486, n77487, n77488, n77489, n77490, n77491,
    n77492, n77493, n77494, n77495, n77496, n77497, n77498, n77499, n77500,
    n77501, n77502, n77503, n77504, n77505, n77506, n77507, n77508, n77509,
    n77510, n77511, n77512, n77513, n77514, n77515, n77516, n77517, n77518,
    n77519, n77520, n77521, n77522, n77523, n77524, n77525, n77526, n77527,
    n77528, n77529, n77530, n77531, n77532, n77533, n77534, n77535, n77536,
    n77537, n77538, n77539, n77540, n77541, n77542, n77543, n77544, n77545,
    n77546, n77547, n77548, n77549, n77550, n77551, n77552, n77553, n77554,
    n77555, n77556, n77557, n77558, n77559, n77560, n77561, n77562, n77563,
    n77564, n77565, n77566, n77567, n77568, n77569, n77570, n77571, n77572,
    n77573, n77574, n77575, n77576, n77577, n77578, n77579, n77580, n77581,
    n77582, n77583, n77584, n77585, n77586, n77587, n77588, n77589, n77590,
    n77591, n77592, n77593, n77594, n77595, n77596, n77597, n77598, n77599,
    n77600, n77601, n77602, n77603, n77604, n77605, n77606, n77607, n77608,
    n77609, n77610, n77611, n77612, n77613, n77614, n77615, n77616, n77617,
    n77618, n77619, n77620, n77621, n77622, n77623, n77624, n77625, n77626,
    n77627, n77628, n77629, n77630, n77631, n77632, n77633, n77634, n77635,
    n77636, n77637, n77638, n77639, n77640, n77641, n77642, n77643, n77644,
    n77645, n77646, n77647, n77648, n77649, n77650, n77651, n77652, n77653,
    n77654, n77655, n77656, n77657, n77658, n77659, n77660, n77661, n77662,
    n77663, n77664, n77665, n77666, n77667, n77668, n77669, n77670, n77671,
    n77672, n77673, n77674, n77675, n77676, n77677, n77678, n77679, n77680,
    n77681, n77682, n77683, n77684, n77685, n77686, n77687, n77688, n77689,
    n77690, n77691, n77692, n77693, n77694, n77695, n77696, n77697, n77698,
    n77699, n77700, n77701, n77702, n77703, n77704, n77705, n77706, n77707,
    n77708, n77709, n77710, n77711, n77712, n77713, n77714, n77715, n77716,
    n77717, n77718, n77719, n77720, n77721, n77722, n77723, n77724, n77725,
    n77726, n77727, n77728, n77729, n77730, n77731, n77732, n77733, n77734,
    n77735, n77736, n77737, n77738, n77739, n77740, n77741, n77742, n77743,
    n77744, n77745, n77746, n77747, n77748, n77749, n77750, n77751, n77752,
    n77753, n77754, n77755, n77756, n77757, n77758, n77759, n77760, n77761,
    n77762, n77763, n77764, n77765, n77766, n77767, n77768, n77769, n77770,
    n77771, n77772, n77773, n77774, n77775, n77776, n77777, n77778, n77779,
    n77780, n77781, n77782, n77783, n77784, n77785, n77786, n77787, n77788,
    n77789, n77790, n77791, n77792, n77793, n77794, n77795, n77796, n77797,
    n77798, n77799, n77800, n77801, n77802, n77803, n77804, n77805, n77806,
    n77807, n77808, n77809, n77810, n77811, n77812, n77813, n77814, n77815,
    n77816, n77817, n77818, n77819, n77820, n77821, n77822, n77823, n77824,
    n77825, n77826, n77827, n77828, n77829, n77830, n77831, n77832, n77833,
    n77834, n77835, n77836, n77837, n77838, n77839, n77840, n77841, n77842,
    n77843, n77844, n77845, n77846, n77847, n77848, n77849, n77850, n77851,
    n77852, n77853, n77854, n77855, n77856, n77857, n77858, n77859, n77860,
    n77861, n77862, n77863, n77864, n77865, n77866, n77867, n77868, n77869,
    n77870, n77871, n77872, n77873, n77874, n77875, n77876, n77877, n77878,
    n77879, n77880, n77881, n77882, n77883, n77884, n77885, n77886, n77887,
    n77888, n77889, n77890, n77891, n77892, n77893, n77894, n77895, n77896,
    n77897, n77898, n77899, n77900, n77901, n77902, n77903, n77904, n77905,
    n77906, n77907, n77908, n77909, n77910, n77911, n77912, n77913, n77914,
    n77915, n77916, n77917, n77918, n77919, n77920, n77921, n77922, n77923,
    n77924, n77925, n77926, n77927, n77928, n77929, n77930, n77931, n77932,
    n77933, n77934, n77935, n77936, n77937, n77938, n77939, n77940, n77941,
    n77942, n77943, n77944, n77945, n77946, n77947, n77948, n77949, n77950,
    n77951, n77952, n77953, n77954, n77955, n77956, n77957, n77958, n77959,
    n77960, n77961, n77962, n77963, n77964, n77965, n77966, n77967, n77968,
    n77969, n77970, n77971, n77972, n77973, n77974, n77975, n77976, n77977,
    n77978, n77979, n77980, n77981, n77982, n77983, n77984, n77985, n77986,
    n77987, n77988, n77989, n77990, n77991, n77992, n77993;
  assign n32 = 1'b1;
  assign n33 = pi29 ? n32 : ~n32;
  assign n34 = pi28 ? n32 : n33;
  assign n35 = pi27 ? n32 : n34;
  assign n36 = pi26 ? n32 : n35;
  assign n37 = pi25 ? n32 : n36;
  assign n38 = pi24 ? n32 : n37;
  assign n39 = pi23 ? n32 : n38;
  assign n40 = pi22 ? n32 : n39;
  assign n41 = pi21 ? n40 : n37;
  assign n42 = pi20 ? n41 : n37;
  assign n43 = pi19 ? n42 : n37;
  assign n44 = pi18 ? n32 : n43;
  assign n45 = pi17 ? n32 : n44;
  assign n46 = pi24 ? n37 : n32;
  assign n47 = pi23 ? n46 : n32;
  assign n48 = pi22 ? n37 : n47;
  assign n49 = pi21 ? n37 : n48;
  assign n50 = pi20 ? n37 : n49;
  assign n51 = pi19 ? n37 : n50;
  assign n52 = pi18 ? n51 : n32;
  assign n53 = pi17 ? n37 : n52;
  assign n54 = pi16 ? n45 : n53;
  assign n55 = pi23 ? n38 : n37;
  assign n56 = pi22 ? n32 : n55;
  assign n57 = pi21 ? n56 : n37;
  assign n58 = pi20 ? n57 : n37;
  assign n59 = pi19 ? n58 : n37;
  assign n60 = pi18 ? n32 : n59;
  assign n61 = pi17 ? n32 : n60;
  assign n62 = pi16 ? n61 : n53;
  assign n63 = pi15 ? n54 : n62;
  assign n64 = pi23 ? n32 : n37;
  assign n65 = pi22 ? n64 : n37;
  assign n66 = pi21 ? n65 : n37;
  assign n67 = pi20 ? n66 : n37;
  assign n68 = pi19 ? n67 : n37;
  assign n69 = pi18 ? n32 : n68;
  assign n70 = pi17 ? n32 : n69;
  assign n71 = pi16 ? n70 : n53;
  assign n72 = pi18 ? n32 : n37;
  assign n73 = pi17 ? n32 : n72;
  assign n74 = pi16 ? n73 : n53;
  assign n75 = pi15 ? n71 : n74;
  assign n76 = pi14 ? n63 : n75;
  assign n77 = pi13 ? n32 : n76;
  assign n78 = pi22 ? n32 : n64;
  assign n79 = pi21 ? n32 : n78;
  assign n80 = pi20 ? n32 : n79;
  assign n81 = pi19 ? n32 : n80;
  assign n82 = pi18 ? n81 : n37;
  assign n83 = pi17 ? n32 : n82;
  assign n84 = pi23 ? n37 : n32;
  assign n85 = pi22 ? n37 : n84;
  assign n86 = pi21 ? n37 : n85;
  assign n87 = pi20 ? n37 : n86;
  assign n88 = pi19 ? n37 : n87;
  assign n89 = pi18 ? n88 : n32;
  assign n90 = pi17 ? n37 : n89;
  assign n91 = pi16 ? n83 : n90;
  assign n92 = pi22 ? n32 : n37;
  assign n93 = pi21 ? n32 : n92;
  assign n94 = pi20 ? n32 : n93;
  assign n95 = pi19 ? n32 : n94;
  assign n96 = pi28 ? n32 : ~n33;
  assign n97 = pi27 ? n32 : n96;
  assign n98 = pi26 ? n32 : n97;
  assign n99 = pi25 ? n32 : n98;
  assign n100 = pi18 ? n95 : n99;
  assign n101 = pi17 ? n32 : n100;
  assign n102 = pi24 ? n99 : n32;
  assign n103 = pi23 ? n102 : n32;
  assign n104 = pi22 ? n99 : n103;
  assign n105 = pi21 ? n99 : n104;
  assign n106 = pi20 ? n99 : n105;
  assign n107 = pi19 ? n99 : n106;
  assign n108 = pi18 ? n107 : n32;
  assign n109 = pi17 ? n99 : n108;
  assign n110 = pi16 ? n101 : n109;
  assign n111 = pi15 ? n91 : n110;
  assign n112 = pi23 ? n37 : n99;
  assign n113 = pi22 ? n32 : n112;
  assign n114 = pi21 ? n32 : n113;
  assign n115 = pi20 ? n32 : n114;
  assign n116 = pi19 ? n32 : n115;
  assign n117 = pi18 ? n116 : n99;
  assign n118 = pi17 ? n32 : n117;
  assign n119 = pi23 ? n99 : n32;
  assign n120 = pi22 ? n99 : n119;
  assign n121 = pi21 ? n99 : n120;
  assign n122 = pi20 ? n99 : n121;
  assign n123 = pi19 ? n99 : n122;
  assign n124 = pi18 ? n123 : n32;
  assign n125 = pi17 ? n99 : n124;
  assign n126 = pi16 ? n118 : n125;
  assign n127 = pi22 ? n64 : n99;
  assign n128 = pi21 ? n32 : n127;
  assign n129 = pi20 ? n32 : n128;
  assign n130 = pi19 ? n32 : n129;
  assign n131 = pi18 ? n130 : n99;
  assign n132 = pi17 ? n32 : n131;
  assign n133 = pi16 ? n132 : n125;
  assign n134 = pi15 ? n126 : n133;
  assign n135 = pi14 ? n111 : n134;
  assign n136 = pi28 ? n33 : n32;
  assign n137 = pi27 ? n32 : n136;
  assign n138 = pi26 ? n32 : n137;
  assign n139 = pi25 ? n32 : n138;
  assign n140 = pi23 ? n139 : n32;
  assign n141 = pi22 ? n99 : n140;
  assign n142 = pi21 ? n99 : n141;
  assign n143 = pi20 ? n99 : n142;
  assign n144 = pi19 ? n99 : n143;
  assign n145 = pi18 ? n144 : n32;
  assign n146 = pi17 ? n99 : n145;
  assign n147 = pi16 ? n132 : n146;
  assign n148 = pi23 ? n32 : n99;
  assign n149 = pi22 ? n148 : n99;
  assign n150 = pi21 ? n32 : n149;
  assign n151 = pi20 ? n32 : n150;
  assign n152 = pi19 ? n32 : n151;
  assign n153 = pi18 ? n152 : n99;
  assign n154 = pi17 ? n32 : n153;
  assign n155 = pi27 ? n96 : n32;
  assign n156 = pi26 ? n32 : n155;
  assign n157 = pi25 ? n32 : n156;
  assign n158 = pi23 ? n99 : n157;
  assign n159 = pi22 ? n99 : n158;
  assign n160 = pi21 ? n159 : n99;
  assign n161 = pi20 ? n99 : n160;
  assign n162 = pi19 ? n161 : n99;
  assign n163 = pi18 ? n99 : n162;
  assign n164 = pi23 ? n157 : n99;
  assign n165 = pi22 ? n99 : n164;
  assign n166 = pi21 ? n99 : n165;
  assign n167 = pi20 ? n99 : n166;
  assign n168 = pi22 ? n158 : n99;
  assign n169 = pi21 ? n168 : n99;
  assign n170 = pi24 ? n99 : n157;
  assign n171 = pi23 ? n170 : n32;
  assign n172 = pi22 ? n99 : n171;
  assign n173 = pi21 ? n99 : n172;
  assign n174 = pi20 ? n169 : n173;
  assign n175 = pi19 ? n167 : n174;
  assign n176 = pi18 ? n175 : n32;
  assign n177 = pi17 ? n163 : n176;
  assign n178 = pi16 ? n154 : n177;
  assign n179 = pi15 ? n147 : n178;
  assign n180 = pi22 ? n55 : n37;
  assign n181 = pi22 ? n37 : n99;
  assign n182 = pi21 ? n180 : n181;
  assign n183 = pi20 ? n32 : n182;
  assign n184 = pi19 ? n32 : n183;
  assign n185 = pi18 ? n184 : n99;
  assign n186 = pi17 ? n32 : n185;
  assign n187 = pi16 ? n186 : n177;
  assign n188 = pi20 ? n99 : n173;
  assign n189 = pi19 ? n99 : n188;
  assign n190 = pi18 ? n189 : n32;
  assign n191 = pi17 ? n99 : n190;
  assign n192 = pi16 ? n186 : n191;
  assign n193 = pi15 ? n187 : n192;
  assign n194 = pi14 ? n179 : n193;
  assign n195 = pi13 ? n135 : n194;
  assign n196 = pi12 ? n77 : n195;
  assign n197 = pi21 ? n180 : n99;
  assign n198 = pi20 ? n32 : n197;
  assign n199 = pi19 ? n32 : n198;
  assign n200 = pi18 ? n199 : n99;
  assign n201 = pi17 ? n32 : n200;
  assign n202 = pi27 ? n136 : n32;
  assign n203 = pi26 ? n32 : n202;
  assign n204 = pi25 ? n32 : n203;
  assign n205 = pi24 ? n99 : n204;
  assign n206 = pi23 ? n205 : n32;
  assign n207 = pi22 ? n99 : n206;
  assign n208 = pi21 ? n99 : n207;
  assign n209 = pi20 ? n99 : n208;
  assign n210 = pi19 ? n99 : n209;
  assign n211 = pi18 ? n210 : n32;
  assign n212 = pi17 ? n99 : n211;
  assign n213 = pi16 ? n201 : n212;
  assign n214 = pi22 ? n37 : n158;
  assign n215 = pi21 ? n180 : n214;
  assign n216 = pi20 ? n32 : n215;
  assign n217 = pi19 ? n32 : n216;
  assign n218 = pi22 ? n99 : n37;
  assign n219 = pi21 ? n218 : n99;
  assign n220 = pi21 ? n99 : n181;
  assign n221 = pi21 ? n99 : n218;
  assign n222 = pi20 ? n220 : n221;
  assign n223 = pi19 ? n219 : n222;
  assign n224 = pi18 ? n217 : n223;
  assign n225 = pi17 ? n32 : n224;
  assign n226 = pi21 ? n181 : n99;
  assign n227 = pi20 ? n99 : n226;
  assign n228 = pi19 ? n227 : n99;
  assign n229 = pi18 ? n228 : n99;
  assign n230 = pi28 ? n33 : ~n32;
  assign n231 = pi27 ? n230 : ~n32;
  assign n232 = pi26 ? n32 : ~n231;
  assign n233 = pi25 ? n32 : n232;
  assign n234 = pi24 ? n99 : n233;
  assign n235 = pi23 ? n234 : n32;
  assign n236 = pi22 ? n99 : n235;
  assign n237 = pi21 ? n99 : n236;
  assign n238 = pi20 ? n99 : n237;
  assign n239 = pi19 ? n99 : n238;
  assign n240 = pi18 ? n239 : n32;
  assign n241 = pi17 ? n229 : n240;
  assign n242 = pi16 ? n225 : n241;
  assign n243 = pi15 ? n213 : n242;
  assign n244 = pi22 ? n37 : n157;
  assign n245 = pi21 ? n180 : n244;
  assign n246 = pi20 ? n32 : n245;
  assign n247 = pi19 ? n32 : n246;
  assign n248 = pi22 ? n139 : n157;
  assign n249 = pi21 ? n248 : n157;
  assign n250 = pi20 ? n249 : n157;
  assign n251 = pi19 ? n250 : n157;
  assign n252 = pi18 ? n247 : n251;
  assign n253 = pi17 ? n32 : n252;
  assign n254 = pi20 ? n157 : n249;
  assign n255 = pi19 ? n157 : n254;
  assign n256 = pi19 ? n157 : n250;
  assign n257 = pi18 ? n255 : n256;
  assign n258 = pi22 ? n157 : n139;
  assign n259 = pi21 ? n157 : n258;
  assign n260 = pi24 ? n139 : n32;
  assign n261 = pi23 ? n260 : n32;
  assign n262 = pi22 ? n157 : n261;
  assign n263 = pi21 ? n157 : n262;
  assign n264 = pi20 ? n259 : n263;
  assign n265 = pi19 ? n254 : n264;
  assign n266 = pi18 ? n265 : n32;
  assign n267 = pi17 ? n257 : n266;
  assign n268 = pi16 ? n253 : n267;
  assign n269 = pi21 ? n248 : n244;
  assign n270 = pi21 ? n157 : n244;
  assign n271 = pi20 ? n269 : n270;
  assign n272 = pi22 ? n157 : n37;
  assign n273 = pi21 ? n157 : n272;
  assign n274 = pi20 ? n273 : n157;
  assign n275 = pi19 ? n271 : n274;
  assign n276 = pi18 ? n247 : n275;
  assign n277 = pi17 ? n32 : n276;
  assign n278 = pi21 ? n244 : n157;
  assign n279 = pi21 ? n272 : n157;
  assign n280 = pi20 ? n278 : n279;
  assign n281 = pi19 ? n280 : n254;
  assign n282 = pi21 ? n258 : n157;
  assign n283 = pi20 ? n269 : n279;
  assign n284 = pi19 ? n282 : n283;
  assign n285 = pi18 ? n281 : n284;
  assign n286 = pi20 ? n279 : n249;
  assign n287 = pi21 ? n248 : n258;
  assign n288 = pi20 ? n287 : n263;
  assign n289 = pi19 ? n286 : n288;
  assign n290 = pi18 ? n289 : n32;
  assign n291 = pi17 ? n285 : n290;
  assign n292 = pi16 ? n277 : n291;
  assign n293 = pi15 ? n268 : n292;
  assign n294 = pi14 ? n243 : n293;
  assign n295 = pi23 ? n37 : n139;
  assign n296 = pi22 ? n55 : n295;
  assign n297 = pi22 ? n37 : n139;
  assign n298 = pi21 ? n296 : n297;
  assign n299 = pi20 ? n32 : n298;
  assign n300 = pi19 ? n32 : n299;
  assign n301 = pi18 ? n300 : n139;
  assign n302 = pi17 ? n32 : n301;
  assign n303 = pi22 ? n139 : n261;
  assign n304 = pi21 ? n139 : n303;
  assign n305 = pi20 ? n139 : n304;
  assign n306 = pi19 ? n139 : n305;
  assign n307 = pi18 ? n306 : n32;
  assign n308 = pi17 ? n139 : n307;
  assign n309 = pi16 ? n302 : n308;
  assign n310 = pi21 ? n296 : n139;
  assign n311 = pi20 ? n32 : n310;
  assign n312 = pi19 ? n32 : n311;
  assign n313 = pi18 ? n312 : n139;
  assign n314 = pi17 ? n32 : n313;
  assign n315 = pi26 ? n97 : n32;
  assign n316 = pi25 ? n32 : n315;
  assign n317 = pi23 ? n316 : n32;
  assign n318 = pi22 ? n139 : n317;
  assign n319 = pi21 ? n139 : n318;
  assign n320 = pi20 ? n139 : n319;
  assign n321 = pi19 ? n139 : n320;
  assign n322 = pi18 ? n321 : n32;
  assign n323 = pi17 ? n139 : n322;
  assign n324 = pi16 ? n314 : n323;
  assign n325 = pi15 ? n309 : n324;
  assign n326 = pi22 ? n55 : n139;
  assign n327 = pi21 ? n326 : n139;
  assign n328 = pi20 ? n32 : n327;
  assign n329 = pi19 ? n32 : n328;
  assign n330 = pi18 ? n329 : n139;
  assign n331 = pi17 ? n32 : n330;
  assign n332 = pi16 ? n331 : n323;
  assign n333 = pi27 ? n32 : ~n230;
  assign n334 = pi26 ? n32 : n333;
  assign n335 = pi25 ? n32 : n334;
  assign n336 = pi22 ? n335 : n317;
  assign n337 = pi21 ? n139 : n336;
  assign n338 = pi20 ? n139 : n337;
  assign n339 = pi19 ? n139 : n338;
  assign n340 = pi18 ? n339 : n32;
  assign n341 = pi17 ? n139 : n340;
  assign n342 = pi16 ? n331 : n341;
  assign n343 = pi15 ? n332 : n342;
  assign n344 = pi14 ? n325 : n343;
  assign n345 = pi13 ? n294 : n344;
  assign n346 = pi22 ? n139 : n316;
  assign n347 = pi21 ? n139 : n346;
  assign n348 = pi23 ? n316 : n139;
  assign n349 = pi22 ? n139 : n348;
  assign n350 = pi21 ? n349 : n139;
  assign n351 = pi20 ? n347 : n350;
  assign n352 = pi19 ? n351 : n139;
  assign n353 = pi18 ? n139 : n352;
  assign n354 = pi22 ? n348 : n316;
  assign n355 = pi21 ? n139 : n354;
  assign n356 = pi22 ? n316 : n139;
  assign n357 = pi21 ? n349 : n356;
  assign n358 = pi20 ? n355 : n357;
  assign n359 = pi22 ? n348 : n139;
  assign n360 = pi21 ? n359 : n139;
  assign n361 = pi27 ? n34 : n32;
  assign n362 = pi26 ? n32 : n361;
  assign n363 = pi25 ? n32 : n362;
  assign n364 = pi23 ? n139 : n363;
  assign n365 = pi22 ? n364 : n317;
  assign n366 = pi21 ? n139 : n365;
  assign n367 = pi20 ? n360 : n366;
  assign n368 = pi19 ? n358 : n367;
  assign n369 = pi18 ? n368 : n32;
  assign n370 = pi17 ? n353 : n369;
  assign n371 = pi16 ? n331 : n370;
  assign n372 = pi21 ? n180 : n37;
  assign n373 = pi20 ? n32 : n372;
  assign n374 = pi19 ? n32 : n373;
  assign n375 = pi22 ? n295 : n37;
  assign n376 = pi21 ? n37 : n375;
  assign n377 = pi20 ? n376 : n37;
  assign n378 = pi19 ? n377 : n37;
  assign n379 = pi18 ? n374 : n378;
  assign n380 = pi17 ? n32 : n379;
  assign n381 = pi22 ? n37 : n316;
  assign n382 = pi21 ? n37 : n381;
  assign n383 = pi23 ? n37 : n316;
  assign n384 = pi22 ? n383 : n37;
  assign n385 = pi21 ? n384 : n37;
  assign n386 = pi20 ? n382 : n385;
  assign n387 = pi19 ? n386 : n37;
  assign n388 = pi18 ? n37 : n387;
  assign n389 = pi21 ? n37 : n316;
  assign n390 = pi23 ? n316 : n37;
  assign n391 = pi22 ? n37 : n390;
  assign n392 = pi22 ? n316 : n383;
  assign n393 = pi21 ? n391 : n392;
  assign n394 = pi20 ? n389 : n393;
  assign n395 = pi24 ? n316 : n32;
  assign n396 = pi23 ? n316 : n395;
  assign n397 = pi22 ? n316 : n396;
  assign n398 = pi21 ? n37 : n397;
  assign n399 = pi20 ? n37 : n398;
  assign n400 = pi19 ? n394 : n399;
  assign n401 = pi18 ? n400 : n32;
  assign n402 = pi17 ? n388 : n401;
  assign n403 = pi16 ? n380 : n402;
  assign n404 = pi15 ? n371 : n403;
  assign n405 = pi21 ? n180 : n391;
  assign n406 = pi20 ? n32 : n405;
  assign n407 = pi19 ? n32 : n406;
  assign n408 = pi21 ? n37 : n391;
  assign n409 = pi20 ? n408 : n37;
  assign n410 = pi19 ? n409 : n37;
  assign n411 = pi18 ? n407 : n410;
  assign n412 = pi17 ? n32 : n411;
  assign n413 = pi21 ? n37 : n390;
  assign n414 = pi20 ? n413 : n408;
  assign n415 = pi19 ? n37 : n414;
  assign n416 = pi21 ? n384 : n381;
  assign n417 = pi22 ? n390 : n37;
  assign n418 = pi21 ? n384 : n417;
  assign n419 = pi20 ? n416 : n418;
  assign n420 = pi21 ? n392 : n37;
  assign n421 = pi20 ? n37 : n420;
  assign n422 = pi19 ? n419 : n421;
  assign n423 = pi18 ? n415 : n422;
  assign n424 = pi22 ? n390 : n316;
  assign n425 = pi21 ? n392 : n424;
  assign n426 = pi21 ? n384 : n392;
  assign n427 = pi20 ? n425 : n426;
  assign n428 = pi22 ? n37 : n383;
  assign n429 = pi21 ? n391 : n428;
  assign n430 = pi23 ? n204 : n395;
  assign n431 = pi22 ? n316 : n430;
  assign n432 = pi21 ? n391 : n431;
  assign n433 = pi20 ? n429 : n432;
  assign n434 = pi19 ? n427 : n433;
  assign n435 = pi18 ? n434 : n32;
  assign n436 = pi17 ? n423 : n435;
  assign n437 = pi16 ? n412 : n436;
  assign n438 = pi18 ? n374 : n37;
  assign n439 = pi17 ? n32 : n438;
  assign n440 = pi21 ? n428 : n381;
  assign n441 = pi20 ? n440 : n426;
  assign n442 = pi19 ? n441 : n399;
  assign n443 = pi18 ? n442 : n32;
  assign n444 = pi17 ? n388 : n443;
  assign n445 = pi16 ? n439 : n444;
  assign n446 = pi15 ? n437 : n445;
  assign n447 = pi14 ? n404 : n446;
  assign n448 = pi23 ? n335 : n204;
  assign n449 = pi22 ? n55 : n448;
  assign n450 = pi23 ? n204 : n335;
  assign n451 = pi22 ? n37 : n450;
  assign n452 = pi21 ? n449 : n451;
  assign n453 = pi20 ? n32 : n452;
  assign n454 = pi19 ? n32 : n453;
  assign n455 = pi23 ? n204 : n37;
  assign n456 = pi23 ? n37 : n204;
  assign n457 = pi22 ? n455 : n456;
  assign n458 = pi22 ? n448 : n450;
  assign n459 = pi21 ? n457 : n458;
  assign n460 = pi22 ? n448 : n37;
  assign n461 = pi21 ? n457 : n460;
  assign n462 = pi20 ? n459 : n461;
  assign n463 = pi22 ? n450 : n455;
  assign n464 = pi22 ? n456 : n448;
  assign n465 = pi21 ? n463 : n464;
  assign n466 = pi21 ? n451 : n457;
  assign n467 = pi20 ? n465 : n466;
  assign n468 = pi19 ? n462 : n467;
  assign n469 = pi18 ? n454 : n468;
  assign n470 = pi17 ? n32 : n469;
  assign n471 = pi21 ? n460 : n463;
  assign n472 = pi21 ? n464 : n451;
  assign n473 = pi20 ? n471 : n472;
  assign n474 = pi22 ? n204 : n448;
  assign n475 = pi21 ? n474 : n451;
  assign n476 = pi22 ? n335 : n450;
  assign n477 = pi21 ? n457 : n476;
  assign n478 = pi20 ? n475 : n477;
  assign n479 = pi19 ? n473 : n478;
  assign n480 = pi22 ? n316 : n448;
  assign n481 = pi21 ? n480 : n451;
  assign n482 = pi20 ? n477 : n481;
  assign n483 = pi19 ? n482 : n459;
  assign n484 = pi18 ? n479 : n483;
  assign n485 = pi22 ? n456 : n335;
  assign n486 = pi22 ? n450 : n316;
  assign n487 = pi21 ? n485 : n486;
  assign n488 = pi20 ? n477 : n487;
  assign n489 = pi22 ? n450 : n456;
  assign n490 = pi21 ? n460 : n489;
  assign n491 = pi22 ? n204 : n396;
  assign n492 = pi21 ? n460 : n491;
  assign n493 = pi20 ? n490 : n492;
  assign n494 = pi19 ? n488 : n493;
  assign n495 = pi18 ? n494 : n32;
  assign n496 = pi17 ? n484 : n495;
  assign n497 = pi16 ? n470 : n496;
  assign n498 = pi22 ? n55 : n456;
  assign n499 = pi22 ? n456 : n37;
  assign n500 = pi21 ? n498 : n499;
  assign n501 = pi20 ? n32 : n500;
  assign n502 = pi19 ? n32 : n501;
  assign n503 = pi21 ? n455 : n460;
  assign n504 = pi21 ? n455 : n456;
  assign n505 = pi20 ? n503 : n504;
  assign n506 = pi22 ? n37 : n455;
  assign n507 = pi21 ? n506 : n457;
  assign n508 = pi21 ? n499 : n455;
  assign n509 = pi20 ? n507 : n508;
  assign n510 = pi19 ? n505 : n509;
  assign n511 = pi18 ? n502 : n510;
  assign n512 = pi17 ? n32 : n511;
  assign n513 = pi21 ? n456 : n506;
  assign n514 = pi21 ? n457 : n499;
  assign n515 = pi20 ? n513 : n514;
  assign n516 = pi22 ? n455 : n204;
  assign n517 = pi21 ? n516 : n499;
  assign n518 = pi20 ? n514 : n517;
  assign n519 = pi19 ? n515 : n518;
  assign n520 = pi22 ? n456 : n455;
  assign n521 = pi21 ? n516 : n520;
  assign n522 = pi22 ? n204 : n456;
  assign n523 = pi21 ? n522 : n499;
  assign n524 = pi20 ? n521 : n523;
  assign n525 = pi21 ? n455 : n499;
  assign n526 = pi19 ? n524 : n525;
  assign n527 = pi18 ? n519 : n526;
  assign n528 = pi21 ? n522 : n516;
  assign n529 = pi20 ? n521 : n528;
  assign n530 = pi21 ? n456 : n516;
  assign n531 = pi24 ? n204 : n32;
  assign n532 = pi23 ? n531 : n32;
  assign n533 = pi22 ? n450 : n532;
  assign n534 = pi21 ? n456 : n533;
  assign n535 = pi20 ? n530 : n534;
  assign n536 = pi19 ? n529 : n535;
  assign n537 = pi18 ? n536 : n32;
  assign n538 = pi17 ? n527 : n537;
  assign n539 = pi16 ? n512 : n538;
  assign n540 = pi15 ? n497 : n539;
  assign n541 = pi20 ? n525 : n504;
  assign n542 = pi19 ? n541 : n509;
  assign n543 = pi18 ? n502 : n542;
  assign n544 = pi17 ? n32 : n543;
  assign n545 = pi20 ? n517 : n514;
  assign n546 = pi19 ? n545 : n525;
  assign n547 = pi18 ? n519 : n546;
  assign n548 = pi21 ? n522 : n506;
  assign n549 = pi20 ? n517 : n548;
  assign n550 = pi20 ? n513 : n534;
  assign n551 = pi19 ? n549 : n550;
  assign n552 = pi18 ? n551 : n32;
  assign n553 = pi17 ? n547 : n552;
  assign n554 = pi16 ? n544 : n553;
  assign n555 = pi22 ? n55 : n335;
  assign n556 = pi21 ? n555 : n37;
  assign n557 = pi20 ? n32 : n556;
  assign n558 = pi19 ? n32 : n557;
  assign n559 = pi23 ? n37 : n233;
  assign n560 = pi22 ? n559 : n37;
  assign n561 = pi21 ? n37 : n560;
  assign n562 = pi20 ? n561 : n37;
  assign n563 = pi19 ? n562 : n37;
  assign n564 = pi18 ? n558 : n563;
  assign n565 = pi17 ? n32 : n564;
  assign n566 = pi23 ? n335 : n37;
  assign n567 = pi22 ? n566 : n335;
  assign n568 = pi21 ? n567 : n37;
  assign n569 = pi22 ? n37 : n335;
  assign n570 = pi22 ? n335 : n37;
  assign n571 = pi21 ? n569 : n570;
  assign n572 = pi20 ? n568 : n571;
  assign n573 = pi19 ? n37 : n572;
  assign n574 = pi22 ? n566 : n37;
  assign n575 = pi21 ? n574 : n37;
  assign n576 = pi20 ? n571 : n575;
  assign n577 = pi21 ? n37 : n335;
  assign n578 = pi19 ? n576 : n577;
  assign n579 = pi18 ? n573 : n578;
  assign n580 = pi22 ? n37 : n566;
  assign n581 = pi21 ? n335 : n580;
  assign n582 = pi20 ? n571 : n581;
  assign n583 = pi23 ? n37 : n335;
  assign n584 = pi22 ? n37 : n583;
  assign n585 = pi21 ? n584 : n580;
  assign n586 = pi24 ? n335 : n32;
  assign n587 = pi23 ? n586 : n32;
  assign n588 = pi22 ? n335 : n587;
  assign n589 = pi21 ? n584 : n588;
  assign n590 = pi20 ? n585 : n589;
  assign n591 = pi19 ? n582 : n590;
  assign n592 = pi18 ? n591 : n32;
  assign n593 = pi17 ? n579 : n592;
  assign n594 = pi16 ? n565 : n593;
  assign n595 = pi15 ? n554 : n594;
  assign n596 = pi14 ? n540 : n595;
  assign n597 = pi13 ? n447 : n596;
  assign n598 = pi12 ? n345 : n597;
  assign n599 = pi11 ? n196 : n598;
  assign n600 = pi21 ? n555 : n335;
  assign n601 = pi20 ? n32 : n600;
  assign n602 = pi19 ? n32 : n601;
  assign n603 = pi21 ? n569 : n335;
  assign n604 = pi21 ? n570 : n335;
  assign n605 = pi21 ? n335 : n569;
  assign n606 = pi20 ? n604 : n605;
  assign n607 = pi19 ? n603 : n606;
  assign n608 = pi18 ? n602 : n607;
  assign n609 = pi17 ? n32 : n608;
  assign n610 = pi21 ? n335 : n570;
  assign n611 = pi20 ? n610 : n335;
  assign n612 = pi20 ? n335 : n603;
  assign n613 = pi19 ? n611 : n612;
  assign n614 = pi20 ? n571 : n335;
  assign n615 = pi19 ? n614 : n603;
  assign n616 = pi18 ? n613 : n615;
  assign n617 = pi20 ? n571 : n605;
  assign n618 = pi21 ? n335 : n588;
  assign n619 = pi20 ? n605 : n618;
  assign n620 = pi19 ? n617 : n619;
  assign n621 = pi18 ? n620 : n32;
  assign n622 = pi17 ? n616 : n621;
  assign n623 = pi16 ? n609 : n622;
  assign n624 = pi24 ? n233 : n32;
  assign n625 = pi23 ? n624 : n32;
  assign n626 = pi22 ? n335 : n625;
  assign n627 = pi21 ? n335 : n626;
  assign n628 = pi20 ? n605 : n627;
  assign n629 = pi19 ? n617 : n628;
  assign n630 = pi18 ? n629 : n32;
  assign n631 = pi17 ? n616 : n630;
  assign n632 = pi16 ? n609 : n631;
  assign n633 = pi15 ? n623 : n632;
  assign n634 = pi20 ? n571 : n37;
  assign n635 = pi19 ? n634 : n37;
  assign n636 = pi18 ? n558 : n635;
  assign n637 = pi17 ? n32 : n636;
  assign n638 = pi21 ? n569 : n37;
  assign n639 = pi21 ? n37 : n570;
  assign n640 = pi20 ? n638 : n639;
  assign n641 = pi19 ? n37 : n640;
  assign n642 = pi21 ? n570 : n37;
  assign n643 = pi20 ? n639 : n642;
  assign n644 = pi20 ? n37 : n642;
  assign n645 = pi19 ? n643 : n644;
  assign n646 = pi18 ? n641 : n645;
  assign n647 = pi21 ? n335 : n37;
  assign n648 = pi20 ? n647 : n605;
  assign n649 = pi21 ? n37 : n569;
  assign n650 = pi22 ? n233 : n625;
  assign n651 = pi21 ? n37 : n650;
  assign n652 = pi20 ? n649 : n651;
  assign n653 = pi19 ? n648 : n652;
  assign n654 = pi18 ? n653 : n32;
  assign n655 = pi17 ? n646 : n654;
  assign n656 = pi16 ? n637 : n655;
  assign n657 = pi20 ? n37 : n651;
  assign n658 = pi19 ? n37 : n657;
  assign n659 = pi18 ? n658 : n32;
  assign n660 = pi17 ? n37 : n659;
  assign n661 = pi16 ? n439 : n660;
  assign n662 = pi15 ? n656 : n661;
  assign n663 = pi14 ? n633 : n662;
  assign n664 = pi23 ? n233 : n32;
  assign n665 = pi22 ? n233 : n664;
  assign n666 = pi21 ? n37 : n665;
  assign n667 = pi20 ? n37 : n666;
  assign n668 = pi19 ? n37 : n667;
  assign n669 = pi18 ? n668 : n32;
  assign n670 = pi17 ? n37 : n669;
  assign n671 = pi16 ? n439 : n670;
  assign n672 = pi15 ? n661 : n671;
  assign n673 = pi23 ? n363 : n233;
  assign n674 = pi22 ? n673 : n625;
  assign n675 = pi21 ? n37 : n674;
  assign n676 = pi20 ? n37 : n675;
  assign n677 = pi19 ? n37 : n676;
  assign n678 = pi18 ? n677 : n32;
  assign n679 = pi17 ? n37 : n678;
  assign n680 = pi16 ? n439 : n679;
  assign n681 = pi15 ? n661 : n680;
  assign n682 = pi14 ? n672 : n681;
  assign n683 = pi13 ? n663 : n682;
  assign n684 = pi26 ? n35 : n32;
  assign n685 = pi25 ? n32 : n684;
  assign n686 = pi23 ? n363 : n685;
  assign n687 = pi24 ? n685 : n32;
  assign n688 = pi23 ? n687 : n32;
  assign n689 = pi22 ? n686 : n688;
  assign n690 = pi21 ? n37 : n689;
  assign n691 = pi20 ? n37 : n690;
  assign n692 = pi19 ? n37 : n691;
  assign n693 = pi18 ? n692 : n32;
  assign n694 = pi17 ? n37 : n693;
  assign n695 = pi16 ? n439 : n694;
  assign n696 = pi22 ? n685 : n688;
  assign n697 = pi21 ? n37 : n696;
  assign n698 = pi20 ? n37 : n697;
  assign n699 = pi19 ? n37 : n698;
  assign n700 = pi18 ? n699 : n32;
  assign n701 = pi17 ? n37 : n700;
  assign n702 = pi16 ? n439 : n701;
  assign n703 = pi15 ? n695 : n702;
  assign n704 = pi14 ? n680 : n703;
  assign n705 = pi23 ? n363 : n316;
  assign n706 = pi23 ? n395 : n32;
  assign n707 = pi22 ? n705 : n706;
  assign n708 = pi21 ? n37 : n707;
  assign n709 = pi20 ? n37 : n708;
  assign n710 = pi19 ? n37 : n709;
  assign n711 = pi18 ? n710 : n32;
  assign n712 = pi17 ? n37 : n711;
  assign n713 = pi16 ? n439 : n712;
  assign n714 = pi24 ? n32 : n99;
  assign n715 = pi23 ? n714 : n99;
  assign n716 = pi22 ? n715 : n99;
  assign n717 = pi21 ? n716 : n99;
  assign n718 = pi20 ? n32 : n717;
  assign n719 = pi19 ? n32 : n718;
  assign n720 = pi18 ? n719 : n99;
  assign n721 = pi17 ? n32 : n720;
  assign n722 = pi22 ? n99 : n363;
  assign n723 = pi21 ? n722 : n707;
  assign n724 = pi20 ? n99 : n723;
  assign n725 = pi19 ? n227 : n724;
  assign n726 = pi18 ? n725 : n32;
  assign n727 = pi17 ? n99 : n726;
  assign n728 = pi16 ? n721 : n727;
  assign n729 = pi15 ? n713 : n728;
  assign n730 = pi23 ? n685 : n531;
  assign n731 = pi22 ? n730 : n32;
  assign n732 = pi21 ? n99 : n731;
  assign n733 = pi20 ? n99 : n732;
  assign n734 = pi19 ? n99 : n733;
  assign n735 = pi18 ? n734 : n32;
  assign n736 = pi17 ? n99 : n735;
  assign n737 = pi16 ? n721 : n736;
  assign n738 = pi23 ? n38 : n99;
  assign n739 = pi22 ? n738 : n99;
  assign n740 = pi21 ? n739 : n99;
  assign n741 = pi20 ? n32 : n740;
  assign n742 = pi19 ? n32 : n741;
  assign n743 = pi18 ? n742 : n99;
  assign n744 = pi17 ? n32 : n743;
  assign n745 = pi23 ? n99 : n139;
  assign n746 = pi22 ? n99 : n745;
  assign n747 = pi23 ? n157 : n624;
  assign n748 = pi22 ? n747 : n32;
  assign n749 = pi21 ? n746 : n748;
  assign n750 = pi20 ? n99 : n749;
  assign n751 = pi19 ? n99 : n750;
  assign n752 = pi18 ? n751 : n32;
  assign n753 = pi17 ? n99 : n752;
  assign n754 = pi16 ? n744 : n753;
  assign n755 = pi15 ? n737 : n754;
  assign n756 = pi14 ? n729 : n755;
  assign n757 = pi13 ? n704 : n756;
  assign n758 = pi12 ? n683 : n757;
  assign n759 = pi23 ? n685 : n687;
  assign n760 = pi22 ? n759 : n32;
  assign n761 = pi21 ? n746 : n760;
  assign n762 = pi20 ? n99 : n761;
  assign n763 = pi19 ? n99 : n762;
  assign n764 = pi18 ? n763 : n32;
  assign n765 = pi17 ? n99 : n764;
  assign n766 = pi16 ? n744 : n765;
  assign n767 = pi22 ? n99 : n685;
  assign n768 = pi21 ? n767 : n760;
  assign n769 = pi20 ? n99 : n768;
  assign n770 = pi19 ? n99 : n769;
  assign n771 = pi18 ? n770 : n32;
  assign n772 = pi17 ? n99 : n771;
  assign n773 = pi16 ? n721 : n772;
  assign n774 = pi15 ? n766 : n773;
  assign n775 = pi22 ? n157 : n99;
  assign n776 = pi21 ? n99 : n775;
  assign n777 = pi22 ? n99 : n157;
  assign n778 = pi24 ? n157 : n685;
  assign n779 = pi23 ? n778 : n687;
  assign n780 = pi22 ? n779 : n32;
  assign n781 = pi21 ? n777 : n780;
  assign n782 = pi20 ? n776 : n781;
  assign n783 = pi19 ? n99 : n782;
  assign n784 = pi18 ? n783 : n32;
  assign n785 = pi17 ? n99 : n784;
  assign n786 = pi16 ? n744 : n785;
  assign n787 = pi21 ? n777 : n157;
  assign n788 = pi21 ? n157 : n780;
  assign n789 = pi20 ? n787 : n788;
  assign n790 = pi19 ? n99 : n789;
  assign n791 = pi18 ? n790 : n32;
  assign n792 = pi17 ? n99 : n791;
  assign n793 = pi16 ? n744 : n792;
  assign n794 = pi15 ? n786 : n793;
  assign n795 = pi14 ? n774 : n794;
  assign n796 = pi22 ? n55 : n99;
  assign n797 = pi21 ? n796 : n99;
  assign n798 = pi20 ? n32 : n797;
  assign n799 = pi19 ? n32 : n798;
  assign n800 = pi18 ? n799 : n99;
  assign n801 = pi17 ? n32 : n800;
  assign n802 = pi21 ? n775 : n99;
  assign n803 = pi20 ? n776 : n802;
  assign n804 = pi19 ? n99 : n803;
  assign n805 = pi18 ? n804 : n99;
  assign n806 = pi20 ? n776 : n788;
  assign n807 = pi19 ? n99 : n806;
  assign n808 = pi18 ? n807 : n32;
  assign n809 = pi17 ? n805 : n808;
  assign n810 = pi16 ? n801 : n809;
  assign n811 = pi22 ? n55 : n745;
  assign n812 = pi23 ? n139 : n99;
  assign n813 = pi22 ? n112 : n812;
  assign n814 = pi21 ? n811 : n813;
  assign n815 = pi20 ? n32 : n814;
  assign n816 = pi19 ? n32 : n815;
  assign n817 = pi22 ? n139 : n158;
  assign n818 = pi21 ? n817 : n258;
  assign n819 = pi22 ? n745 : n157;
  assign n820 = pi22 ? n139 : n37;
  assign n821 = pi21 ? n819 : n820;
  assign n822 = pi20 ? n818 : n821;
  assign n823 = pi22 ? n745 : n812;
  assign n824 = pi21 ? n823 : n248;
  assign n825 = pi22 ? n139 : n745;
  assign n826 = pi21 ? n813 : n825;
  assign n827 = pi20 ? n824 : n826;
  assign n828 = pi19 ? n822 : n827;
  assign n829 = pi18 ? n816 : n828;
  assign n830 = pi17 ? n32 : n829;
  assign n831 = pi22 ? n745 : n112;
  assign n832 = pi21 ? n258 : n831;
  assign n833 = pi20 ? n832 : n287;
  assign n834 = pi19 ? n833 : n157;
  assign n835 = pi22 ? n164 : n139;
  assign n836 = pi21 ? n157 : n835;
  assign n837 = pi22 ? n745 : n99;
  assign n838 = pi21 ? n837 : n157;
  assign n839 = pi20 ? n836 : n838;
  assign n840 = pi19 ? n157 : n839;
  assign n841 = pi18 ? n834 : n840;
  assign n842 = pi24 ? n157 : n316;
  assign n843 = pi23 ? n842 : n395;
  assign n844 = pi22 ? n843 : n32;
  assign n845 = pi21 ? n157 : n844;
  assign n846 = pi20 ? n157 : n845;
  assign n847 = pi19 ? n157 : n846;
  assign n848 = pi18 ? n847 : n32;
  assign n849 = pi17 ? n841 : n848;
  assign n850 = pi16 ? n830 : n849;
  assign n851 = pi15 ? n810 : n850;
  assign n852 = pi23 ? n157 : n139;
  assign n853 = pi22 ? n852 : n139;
  assign n854 = pi21 ? n326 : n853;
  assign n855 = pi20 ? n32 : n854;
  assign n856 = pi19 ? n32 : n855;
  assign n857 = pi22 ? n852 : n157;
  assign n858 = pi22 ? n139 : n852;
  assign n859 = pi21 ? n857 : n858;
  assign n860 = pi20 ? n287 : n859;
  assign n861 = pi23 ? n139 : n157;
  assign n862 = pi22 ? n139 : n861;
  assign n863 = pi21 ? n862 : n858;
  assign n864 = pi21 ? n139 : n858;
  assign n865 = pi20 ? n863 : n864;
  assign n866 = pi19 ? n860 : n865;
  assign n867 = pi18 ? n856 : n866;
  assign n868 = pi17 ? n32 : n867;
  assign n869 = pi21 ? n258 : n858;
  assign n870 = pi21 ? n258 : n857;
  assign n871 = pi20 ? n869 : n870;
  assign n872 = pi19 ? n871 : n250;
  assign n873 = pi21 ? n157 : n248;
  assign n874 = pi20 ? n873 : n157;
  assign n875 = pi21 ? n248 : n139;
  assign n876 = pi21 ? n139 : n258;
  assign n877 = pi20 ? n875 : n876;
  assign n878 = pi19 ? n874 : n877;
  assign n879 = pi18 ? n872 : n878;
  assign n880 = pi21 ? n157 : n139;
  assign n881 = pi20 ? n873 : n880;
  assign n882 = pi22 ? n396 : n32;
  assign n883 = pi21 ? n157 : n882;
  assign n884 = pi20 ? n287 : n883;
  assign n885 = pi19 ? n881 : n884;
  assign n886 = pi18 ? n885 : n32;
  assign n887 = pi17 ? n879 : n886;
  assign n888 = pi16 ? n868 : n887;
  assign n889 = pi23 ? n157 : n37;
  assign n890 = pi22 ? n139 : n889;
  assign n891 = pi21 ? n857 : n890;
  assign n892 = pi20 ? n287 : n891;
  assign n893 = pi23 ? n37 : n157;
  assign n894 = pi22 ? n139 : n893;
  assign n895 = pi21 ? n894 : n858;
  assign n896 = pi20 ? n895 : n864;
  assign n897 = pi19 ? n892 : n896;
  assign n898 = pi18 ? n856 : n897;
  assign n899 = pi17 ? n32 : n898;
  assign n900 = pi21 ? n857 : n882;
  assign n901 = pi20 ? n875 : n900;
  assign n902 = pi19 ? n881 : n901;
  assign n903 = pi18 ? n902 : n32;
  assign n904 = pi17 ? n879 : n903;
  assign n905 = pi16 ? n899 : n904;
  assign n906 = pi15 ? n888 : n905;
  assign n907 = pi14 ? n851 : n906;
  assign n908 = pi13 ? n795 : n907;
  assign n909 = pi23 ? n38 : n139;
  assign n910 = pi22 ? n909 : n139;
  assign n911 = pi21 ? n910 : n139;
  assign n912 = pi20 ? n32 : n911;
  assign n913 = pi19 ? n32 : n912;
  assign n914 = pi18 ? n913 : n139;
  assign n915 = pi17 ? n32 : n914;
  assign n916 = pi22 ? n139 : n204;
  assign n917 = pi19 ? n139 : n916;
  assign n918 = pi23 ? n204 : n139;
  assign n919 = pi22 ? n139 : n918;
  assign n920 = pi21 ? n919 : n139;
  assign n921 = pi22 ? n204 : n139;
  assign n922 = pi21 ? n921 : n139;
  assign n923 = pi20 ? n920 : n922;
  assign n924 = pi19 ? n923 : n139;
  assign n925 = pi18 ? n917 : n924;
  assign n926 = pi20 ? n139 : n922;
  assign n927 = pi21 ? n916 : n139;
  assign n928 = pi22 ? n317 : n32;
  assign n929 = pi21 ? n346 : n928;
  assign n930 = pi20 ? n927 : n929;
  assign n931 = pi19 ? n926 : n930;
  assign n932 = pi18 ? n931 : n32;
  assign n933 = pi17 ? n925 : n932;
  assign n934 = pi16 ? n915 : n933;
  assign n935 = pi22 ? n909 : n37;
  assign n936 = pi21 ? n935 : n297;
  assign n937 = pi20 ? n32 : n936;
  assign n938 = pi19 ? n32 : n937;
  assign n939 = pi21 ? n139 : n297;
  assign n940 = pi20 ? n139 : n939;
  assign n941 = pi21 ? n139 : n37;
  assign n942 = pi21 ? n297 : n139;
  assign n943 = pi20 ? n941 : n942;
  assign n944 = pi19 ? n940 : n943;
  assign n945 = pi18 ? n938 : n944;
  assign n946 = pi17 ? n32 : n945;
  assign n947 = pi21 ? n820 : n139;
  assign n948 = pi20 ? n297 : n947;
  assign n949 = pi19 ? n948 : n139;
  assign n950 = pi19 ? n139 : n943;
  assign n951 = pi18 ? n949 : n950;
  assign n952 = pi22 ? n37 : n348;
  assign n953 = pi21 ? n139 : n952;
  assign n954 = pi21 ? n916 : n928;
  assign n955 = pi20 ? n953 : n954;
  assign n956 = pi19 ? n139 : n955;
  assign n957 = pi18 ? n956 : n32;
  assign n958 = pi17 ? n951 : n957;
  assign n959 = pi16 ? n946 : n958;
  assign n960 = pi15 ? n934 : n959;
  assign n961 = pi24 ? n32 : n139;
  assign n962 = pi23 ? n961 : n139;
  assign n963 = pi22 ? n962 : n139;
  assign n964 = pi21 ? n963 : n139;
  assign n965 = pi20 ? n32 : n964;
  assign n966 = pi19 ? n32 : n965;
  assign n967 = pi19 ? n940 : n139;
  assign n968 = pi18 ? n966 : n967;
  assign n969 = pi17 ? n32 : n968;
  assign n970 = pi20 ? n139 : n929;
  assign n971 = pi19 ? n139 : n970;
  assign n972 = pi18 ? n971 : n32;
  assign n973 = pi17 ? n139 : n972;
  assign n974 = pi16 ? n969 : n973;
  assign n975 = pi21 ? n139 : n316;
  assign n976 = pi21 ? n346 : n139;
  assign n977 = pi20 ? n975 : n976;
  assign n978 = pi19 ? n139 : n977;
  assign n979 = pi18 ? n978 : n139;
  assign n980 = pi21 ? n316 : n928;
  assign n981 = pi20 ? n139 : n980;
  assign n982 = pi19 ? n139 : n981;
  assign n983 = pi18 ? n982 : n32;
  assign n984 = pi17 ? n979 : n983;
  assign n985 = pi16 ? n969 : n984;
  assign n986 = pi15 ? n974 : n985;
  assign n987 = pi14 ? n960 : n986;
  assign n988 = pi21 ? n180 : n139;
  assign n989 = pi20 ? n32 : n988;
  assign n990 = pi19 ? n32 : n989;
  assign n991 = pi20 ? n942 : n939;
  assign n992 = pi21 ? n139 : n820;
  assign n993 = pi20 ? n941 : n992;
  assign n994 = pi19 ? n991 : n993;
  assign n995 = pi18 ? n990 : n994;
  assign n996 = pi17 ? n32 : n995;
  assign n997 = pi21 ? n297 : n820;
  assign n998 = pi20 ? n997 : n139;
  assign n999 = pi20 ? n975 : n316;
  assign n1000 = pi19 ? n998 : n999;
  assign n1001 = pi21 ? n346 : n356;
  assign n1002 = pi20 ? n356 : n1001;
  assign n1003 = pi21 ? n297 : n37;
  assign n1004 = pi20 ? n1003 : n947;
  assign n1005 = pi19 ? n1002 : n1004;
  assign n1006 = pi18 ? n1000 : n1005;
  assign n1007 = pi20 ? n942 : n1001;
  assign n1008 = pi21 ? n139 : n356;
  assign n1009 = pi22 ? n706 : n32;
  assign n1010 = pi21 ? n316 : n1009;
  assign n1011 = pi20 ? n1008 : n1010;
  assign n1012 = pi19 ? n1007 : n1011;
  assign n1013 = pi18 ? n1012 : n32;
  assign n1014 = pi17 ? n1006 : n1013;
  assign n1015 = pi16 ? n996 : n1014;
  assign n1016 = pi21 ? n139 : n204;
  assign n1017 = pi20 ? n139 : n1016;
  assign n1018 = pi22 ? n316 : n204;
  assign n1019 = pi21 ? n1018 : n316;
  assign n1020 = pi20 ? n1019 : n356;
  assign n1021 = pi19 ? n1017 : n1020;
  assign n1022 = pi21 ? n316 : n139;
  assign n1023 = pi20 ? n1022 : n976;
  assign n1024 = pi19 ? n1023 : n139;
  assign n1025 = pi18 ? n1021 : n1024;
  assign n1026 = pi21 ? n139 : n916;
  assign n1027 = pi22 ? n204 : n316;
  assign n1028 = pi21 ? n1027 : n1018;
  assign n1029 = pi20 ? n1026 : n1028;
  assign n1030 = pi21 ? n1027 : n1009;
  assign n1031 = pi20 ? n976 : n1030;
  assign n1032 = pi19 ? n1029 : n1031;
  assign n1033 = pi18 ? n1032 : n32;
  assign n1034 = pi17 ? n1025 : n1033;
  assign n1035 = pi16 ? n331 : n1034;
  assign n1036 = pi15 ? n1015 : n1035;
  assign n1037 = pi22 ? n55 : n204;
  assign n1038 = pi23 ? n139 : n204;
  assign n1039 = pi22 ? n1038 : n204;
  assign n1040 = pi21 ? n1037 : n1039;
  assign n1041 = pi20 ? n32 : n1040;
  assign n1042 = pi19 ? n32 : n1041;
  assign n1043 = pi23 ? n139 : n37;
  assign n1044 = pi22 ? n204 : n1043;
  assign n1045 = pi21 ? n1044 : n204;
  assign n1046 = pi22 ? n204 : n37;
  assign n1047 = pi21 ? n1046 : n375;
  assign n1048 = pi20 ? n1045 : n1047;
  assign n1049 = pi22 ? n1043 : n204;
  assign n1050 = pi21 ? n1049 : n204;
  assign n1051 = pi20 ? n1046 : n1050;
  assign n1052 = pi19 ? n1048 : n1051;
  assign n1053 = pi18 ? n1042 : n1052;
  assign n1054 = pi17 ? n32 : n1053;
  assign n1055 = pi21 ? n375 : n204;
  assign n1056 = pi22 ? n37 : n204;
  assign n1057 = pi21 ? n1056 : n204;
  assign n1058 = pi20 ? n1055 : n1057;
  assign n1059 = pi21 ? n204 : n1018;
  assign n1060 = pi21 ? n1018 : n204;
  assign n1061 = pi20 ? n1059 : n1060;
  assign n1062 = pi19 ? n1058 : n1061;
  assign n1063 = pi21 ? n204 : n1046;
  assign n1064 = pi20 ? n204 : n1063;
  assign n1065 = pi20 ? n1046 : n1056;
  assign n1066 = pi19 ? n1064 : n1065;
  assign n1067 = pi18 ? n1062 : n1066;
  assign n1068 = pi21 ? n1027 : n204;
  assign n1069 = pi20 ? n204 : n1068;
  assign n1070 = pi23 ? n233 : n316;
  assign n1071 = pi22 ? n204 : n1070;
  assign n1072 = pi21 ? n1071 : n32;
  assign n1073 = pi20 ? n1068 : n1072;
  assign n1074 = pi19 ? n1069 : n1073;
  assign n1075 = pi18 ? n1074 : n32;
  assign n1076 = pi17 ? n1067 : n1075;
  assign n1077 = pi16 ? n1054 : n1076;
  assign n1078 = pi22 ? n715 : n335;
  assign n1079 = pi22 ? n335 : n204;
  assign n1080 = pi21 ? n1078 : n1079;
  assign n1081 = pi20 ? n32 : n1080;
  assign n1082 = pi19 ? n32 : n1081;
  assign n1083 = pi22 ? n204 : n335;
  assign n1084 = pi21 ? n1083 : n335;
  assign n1085 = pi20 ? n1084 : n335;
  assign n1086 = pi19 ? n1085 : n335;
  assign n1087 = pi18 ? n1082 : n1086;
  assign n1088 = pi17 ? n32 : n1087;
  assign n1089 = pi21 ? n335 : n204;
  assign n1090 = pi20 ? n335 : n1089;
  assign n1091 = pi22 ? n316 : n335;
  assign n1092 = pi21 ? n1091 : n1083;
  assign n1093 = pi20 ? n1059 : n1092;
  assign n1094 = pi19 ? n1090 : n1093;
  assign n1095 = pi21 ? n1079 : n335;
  assign n1096 = pi20 ? n204 : n1095;
  assign n1097 = pi19 ? n1096 : n335;
  assign n1098 = pi18 ? n1094 : n1097;
  assign n1099 = pi21 ? n1083 : n204;
  assign n1100 = pi20 ? n1099 : n204;
  assign n1101 = pi21 ? n1027 : n32;
  assign n1102 = pi20 ? n204 : n1101;
  assign n1103 = pi19 ? n1100 : n1102;
  assign n1104 = pi18 ? n1103 : n32;
  assign n1105 = pi17 ? n1098 : n1104;
  assign n1106 = pi16 ? n1088 : n1105;
  assign n1107 = pi15 ? n1077 : n1106;
  assign n1108 = pi14 ? n1036 : n1107;
  assign n1109 = pi13 ? n987 : n1108;
  assign n1110 = pi12 ? n908 : n1109;
  assign n1111 = pi11 ? n758 : n1110;
  assign n1112 = pi10 ? n599 : n1111;
  assign n1113 = pi09 ? n32 : n1112;
  assign n1114 = pi21 ? n78 : n37;
  assign n1115 = pi20 ? n1114 : n37;
  assign n1116 = pi19 ? n1115 : n37;
  assign n1117 = pi18 ? n32 : n1116;
  assign n1118 = pi17 ? n32 : n1117;
  assign n1119 = pi16 ? n1118 : n90;
  assign n1120 = pi15 ? n32 : n1119;
  assign n1121 = pi14 ? n32 : n1120;
  assign n1122 = pi16 ? n61 : n90;
  assign n1123 = pi16 ? n70 : n90;
  assign n1124 = pi15 ? n1122 : n1123;
  assign n1125 = pi16 ? n73 : n90;
  assign n1126 = pi15 ? n1125 : n91;
  assign n1127 = pi14 ? n1124 : n1126;
  assign n1128 = pi13 ? n1121 : n1127;
  assign n1129 = pi18 ? n95 : n37;
  assign n1130 = pi17 ? n32 : n1129;
  assign n1131 = pi16 ? n1130 : n90;
  assign n1132 = pi22 ? n99 : n84;
  assign n1133 = pi21 ? n99 : n1132;
  assign n1134 = pi20 ? n99 : n1133;
  assign n1135 = pi19 ? n99 : n1134;
  assign n1136 = pi18 ? n1135 : n32;
  assign n1137 = pi17 ? n99 : n1136;
  assign n1138 = pi16 ? n118 : n1137;
  assign n1139 = pi15 ? n1131 : n1138;
  assign n1140 = pi16 ? n154 : n125;
  assign n1141 = pi15 ? n133 : n1140;
  assign n1142 = pi14 ? n1139 : n1141;
  assign n1143 = pi22 ? n112 : n99;
  assign n1144 = pi21 ? n180 : n1143;
  assign n1145 = pi20 ? n32 : n1144;
  assign n1146 = pi19 ? n32 : n1145;
  assign n1147 = pi18 ? n1146 : n99;
  assign n1148 = pi17 ? n32 : n1147;
  assign n1149 = pi24 ? n157 : n32;
  assign n1150 = pi23 ? n335 : n1149;
  assign n1151 = pi22 ? n99 : n1150;
  assign n1152 = pi21 ? n99 : n1151;
  assign n1153 = pi20 ? n169 : n1152;
  assign n1154 = pi19 ? n167 : n1153;
  assign n1155 = pi18 ? n1154 : n32;
  assign n1156 = pi17 ? n163 : n1155;
  assign n1157 = pi16 ? n1148 : n1156;
  assign n1158 = pi15 ? n147 : n1157;
  assign n1159 = pi23 ? n363 : n1149;
  assign n1160 = pi22 ? n99 : n1159;
  assign n1161 = pi21 ? n99 : n1160;
  assign n1162 = pi20 ? n169 : n1161;
  assign n1163 = pi19 ? n167 : n1162;
  assign n1164 = pi18 ? n1163 : n32;
  assign n1165 = pi17 ? n163 : n1164;
  assign n1166 = pi16 ? n186 : n1165;
  assign n1167 = pi23 ? n99 : n1149;
  assign n1168 = pi22 ? n99 : n1167;
  assign n1169 = pi21 ? n99 : n1168;
  assign n1170 = pi20 ? n99 : n1169;
  assign n1171 = pi19 ? n99 : n1170;
  assign n1172 = pi18 ? n1171 : n32;
  assign n1173 = pi17 ? n99 : n1172;
  assign n1174 = pi16 ? n186 : n1173;
  assign n1175 = pi15 ? n1166 : n1174;
  assign n1176 = pi14 ? n1158 : n1175;
  assign n1177 = pi13 ? n1142 : n1176;
  assign n1178 = pi12 ? n1128 : n1177;
  assign n1179 = pi22 ? n715 : n112;
  assign n1180 = pi21 ? n1179 : n99;
  assign n1181 = pi20 ? n32 : n1180;
  assign n1182 = pi19 ? n32 : n1181;
  assign n1183 = pi18 ? n1182 : n99;
  assign n1184 = pi17 ? n32 : n1183;
  assign n1185 = pi23 ? n99 : n531;
  assign n1186 = pi22 ? n99 : n1185;
  assign n1187 = pi21 ? n99 : n1186;
  assign n1188 = pi20 ? n99 : n1187;
  assign n1189 = pi19 ? n99 : n1188;
  assign n1190 = pi18 ? n1189 : n32;
  assign n1191 = pi17 ? n99 : n1190;
  assign n1192 = pi16 ? n1184 : n1191;
  assign n1193 = pi17 ? n229 : n1172;
  assign n1194 = pi16 ? n225 : n1193;
  assign n1195 = pi15 ? n1192 : n1194;
  assign n1196 = pi23 ? n139 : n1149;
  assign n1197 = pi22 ? n157 : n1196;
  assign n1198 = pi21 ? n157 : n1197;
  assign n1199 = pi20 ? n259 : n1198;
  assign n1200 = pi19 ? n254 : n1199;
  assign n1201 = pi18 ? n1200 : n32;
  assign n1202 = pi17 ? n257 : n1201;
  assign n1203 = pi16 ? n253 : n1202;
  assign n1204 = pi20 ? n287 : n1198;
  assign n1205 = pi19 ? n286 : n1204;
  assign n1206 = pi18 ? n1205 : n32;
  assign n1207 = pi17 ? n285 : n1206;
  assign n1208 = pi16 ? n277 : n1207;
  assign n1209 = pi15 ? n1203 : n1208;
  assign n1210 = pi14 ? n1195 : n1209;
  assign n1211 = pi22 ? n1043 : n139;
  assign n1212 = pi21 ? n296 : n1211;
  assign n1213 = pi20 ? n32 : n1212;
  assign n1214 = pi19 ? n32 : n1213;
  assign n1215 = pi18 ? n1214 : n139;
  assign n1216 = pi17 ? n32 : n1215;
  assign n1217 = pi23 ? n139 : n531;
  assign n1218 = pi22 ? n139 : n1217;
  assign n1219 = pi21 ? n139 : n1218;
  assign n1220 = pi20 ? n139 : n1219;
  assign n1221 = pi19 ? n139 : n1220;
  assign n1222 = pi18 ? n1221 : n32;
  assign n1223 = pi17 ? n139 : n1222;
  assign n1224 = pi16 ? n1216 : n1223;
  assign n1225 = pi16 ? n314 : n1223;
  assign n1226 = pi15 ? n1224 : n1225;
  assign n1227 = pi16 ? n331 : n1223;
  assign n1228 = pi23 ? n316 : n531;
  assign n1229 = pi22 ? n335 : n1228;
  assign n1230 = pi21 ? n139 : n1229;
  assign n1231 = pi20 ? n139 : n1230;
  assign n1232 = pi19 ? n139 : n1231;
  assign n1233 = pi18 ? n1232 : n32;
  assign n1234 = pi17 ? n139 : n1233;
  assign n1235 = pi16 ? n331 : n1234;
  assign n1236 = pi15 ? n1227 : n1235;
  assign n1237 = pi14 ? n1226 : n1236;
  assign n1238 = pi13 ? n1210 : n1237;
  assign n1239 = pi22 ? n364 : n396;
  assign n1240 = pi21 ? n139 : n1239;
  assign n1241 = pi20 ? n360 : n1240;
  assign n1242 = pi19 ? n358 : n1241;
  assign n1243 = pi18 ? n1242 : n32;
  assign n1244 = pi17 ? n353 : n1243;
  assign n1245 = pi16 ? n331 : n1244;
  assign n1246 = pi22 ? n316 : n1228;
  assign n1247 = pi21 ? n37 : n1246;
  assign n1248 = pi20 ? n37 : n1247;
  assign n1249 = pi19 ? n394 : n1248;
  assign n1250 = pi18 ? n1249 : n32;
  assign n1251 = pi17 ? n388 : n1250;
  assign n1252 = pi16 ? n380 : n1251;
  assign n1253 = pi15 ? n1245 : n1252;
  assign n1254 = pi24 ? n37 : n316;
  assign n1255 = pi23 ? n1254 : n531;
  assign n1256 = pi22 ? n316 : n1255;
  assign n1257 = pi21 ? n391 : n1256;
  assign n1258 = pi20 ? n429 : n1257;
  assign n1259 = pi19 ? n427 : n1258;
  assign n1260 = pi18 ? n1259 : n32;
  assign n1261 = pi17 ? n423 : n1260;
  assign n1262 = pi16 ? n412 : n1261;
  assign n1263 = pi23 ? n316 : n624;
  assign n1264 = pi22 ? n316 : n1263;
  assign n1265 = pi21 ? n37 : n1264;
  assign n1266 = pi20 ? n37 : n1265;
  assign n1267 = pi19 ? n441 : n1266;
  assign n1268 = pi18 ? n1267 : n32;
  assign n1269 = pi17 ? n388 : n1268;
  assign n1270 = pi16 ? n439 : n1269;
  assign n1271 = pi15 ? n1262 : n1270;
  assign n1272 = pi14 ? n1253 : n1271;
  assign n1273 = pi22 ? n566 : n450;
  assign n1274 = pi21 ? n449 : n1273;
  assign n1275 = pi20 ? n32 : n1274;
  assign n1276 = pi19 ? n32 : n1275;
  assign n1277 = pi21 ? n489 : n458;
  assign n1278 = pi22 ? n448 : n566;
  assign n1279 = pi21 ? n489 : n1278;
  assign n1280 = pi20 ? n1277 : n1279;
  assign n1281 = pi21 ? n450 : n464;
  assign n1282 = pi21 ? n1273 : n489;
  assign n1283 = pi20 ? n1281 : n1282;
  assign n1284 = pi19 ? n1280 : n1283;
  assign n1285 = pi18 ? n1276 : n1284;
  assign n1286 = pi17 ? n32 : n1285;
  assign n1287 = pi21 ? n1278 : n450;
  assign n1288 = pi21 ? n464 : n1273;
  assign n1289 = pi20 ? n1287 : n1288;
  assign n1290 = pi21 ? n474 : n1273;
  assign n1291 = pi21 ? n489 : n476;
  assign n1292 = pi20 ? n1290 : n1291;
  assign n1293 = pi19 ? n1289 : n1292;
  assign n1294 = pi21 ? n480 : n1273;
  assign n1295 = pi20 ? n1291 : n1294;
  assign n1296 = pi19 ? n1295 : n1277;
  assign n1297 = pi18 ? n1293 : n1296;
  assign n1298 = pi20 ? n1291 : n487;
  assign n1299 = pi21 ? n1278 : n489;
  assign n1300 = pi21 ? n1278 : n486;
  assign n1301 = pi20 ? n1299 : n1300;
  assign n1302 = pi19 ? n1298 : n1301;
  assign n1303 = pi18 ? n1302 : n32;
  assign n1304 = pi17 ? n1297 : n1303;
  assign n1305 = pi16 ? n1286 : n1304;
  assign n1306 = pi21 ? n498 : n37;
  assign n1307 = pi20 ? n32 : n1306;
  assign n1308 = pi19 ? n32 : n1307;
  assign n1309 = pi22 ? n455 : n37;
  assign n1310 = pi21 ? n1309 : n460;
  assign n1311 = pi21 ? n1309 : n499;
  assign n1312 = pi20 ? n1310 : n1311;
  assign n1313 = pi22 ? n37 : n456;
  assign n1314 = pi21 ? n506 : n1313;
  assign n1315 = pi21 ? n37 : n1309;
  assign n1316 = pi20 ? n1314 : n1315;
  assign n1317 = pi19 ? n1312 : n1316;
  assign n1318 = pi18 ? n1308 : n1317;
  assign n1319 = pi17 ? n32 : n1318;
  assign n1320 = pi21 ? n499 : n506;
  assign n1321 = pi21 ? n1313 : n37;
  assign n1322 = pi20 ? n1320 : n1321;
  assign n1323 = pi21 ? n457 : n37;
  assign n1324 = pi20 ? n1323 : n514;
  assign n1325 = pi19 ? n1322 : n1324;
  assign n1326 = pi21 ? n457 : n520;
  assign n1327 = pi21 ? n522 : n37;
  assign n1328 = pi20 ? n1326 : n1327;
  assign n1329 = pi19 ? n1328 : n1311;
  assign n1330 = pi18 ? n1325 : n1329;
  assign n1331 = pi20 ? n1326 : n528;
  assign n1332 = pi21 ? n499 : n516;
  assign n1333 = pi23 ? n335 : n395;
  assign n1334 = pi22 ? n450 : n1333;
  assign n1335 = pi21 ? n499 : n1334;
  assign n1336 = pi20 ? n1332 : n1335;
  assign n1337 = pi19 ? n1331 : n1336;
  assign n1338 = pi18 ? n1337 : n32;
  assign n1339 = pi17 ? n1330 : n1338;
  assign n1340 = pi16 ? n1319 : n1339;
  assign n1341 = pi15 ? n1305 : n1340;
  assign n1342 = pi24 ? n37 : n335;
  assign n1343 = pi23 ? n204 : n1342;
  assign n1344 = pi23 ? n335 : n32;
  assign n1345 = pi22 ? n1343 : n1344;
  assign n1346 = pi21 ? n456 : n1345;
  assign n1347 = pi20 ? n513 : n1346;
  assign n1348 = pi19 ? n549 : n1347;
  assign n1349 = pi18 ? n1348 : n32;
  assign n1350 = pi17 ? n547 : n1349;
  assign n1351 = pi16 ? n544 : n1350;
  assign n1352 = pi22 ? n335 : n1344;
  assign n1353 = pi21 ? n584 : n1352;
  assign n1354 = pi20 ? n585 : n1353;
  assign n1355 = pi19 ? n582 : n1354;
  assign n1356 = pi18 ? n1355 : n32;
  assign n1357 = pi17 ? n579 : n1356;
  assign n1358 = pi16 ? n565 : n1357;
  assign n1359 = pi15 ? n1351 : n1358;
  assign n1360 = pi14 ? n1341 : n1359;
  assign n1361 = pi13 ? n1272 : n1360;
  assign n1362 = pi12 ? n1238 : n1361;
  assign n1363 = pi11 ? n1178 : n1362;
  assign n1364 = pi21 ? n335 : n1352;
  assign n1365 = pi20 ? n605 : n1364;
  assign n1366 = pi19 ? n617 : n1365;
  assign n1367 = pi18 ? n1366 : n32;
  assign n1368 = pi17 ? n616 : n1367;
  assign n1369 = pi16 ? n609 : n1368;
  assign n1370 = pi23 ? n363 : n32;
  assign n1371 = pi22 ? n233 : n1370;
  assign n1372 = pi21 ? n37 : n1371;
  assign n1373 = pi20 ? n649 : n1372;
  assign n1374 = pi19 ? n648 : n1373;
  assign n1375 = pi18 ? n1374 : n32;
  assign n1376 = pi17 ? n646 : n1375;
  assign n1377 = pi16 ? n637 : n1376;
  assign n1378 = pi23 ? n157 : n32;
  assign n1379 = pi22 ? n233 : n1378;
  assign n1380 = pi21 ? n37 : n1379;
  assign n1381 = pi20 ? n37 : n1380;
  assign n1382 = pi19 ? n37 : n1381;
  assign n1383 = pi18 ? n1382 : n32;
  assign n1384 = pi17 ? n37 : n1383;
  assign n1385 = pi16 ? n439 : n1384;
  assign n1386 = pi15 ? n1377 : n1385;
  assign n1387 = pi14 ? n1369 : n1386;
  assign n1388 = pi23 ? n233 : n624;
  assign n1389 = pi22 ? n233 : n1388;
  assign n1390 = pi21 ? n37 : n1389;
  assign n1391 = pi20 ? n37 : n1390;
  assign n1392 = pi19 ? n37 : n1391;
  assign n1393 = pi18 ? n1392 : n32;
  assign n1394 = pi17 ? n37 : n1393;
  assign n1395 = pi16 ? n439 : n1394;
  assign n1396 = pi15 ? n671 : n1395;
  assign n1397 = pi22 ? n673 : n664;
  assign n1398 = pi21 ? n37 : n1397;
  assign n1399 = pi20 ? n37 : n1398;
  assign n1400 = pi19 ? n37 : n1399;
  assign n1401 = pi18 ? n1400 : n32;
  assign n1402 = pi17 ? n37 : n1401;
  assign n1403 = pi16 ? n439 : n1402;
  assign n1404 = pi15 ? n671 : n1403;
  assign n1405 = pi14 ? n1396 : n1404;
  assign n1406 = pi13 ? n1387 : n1405;
  assign n1407 = pi23 ? n685 : n32;
  assign n1408 = pi22 ? n363 : n1407;
  assign n1409 = pi21 ? n37 : n1408;
  assign n1410 = pi20 ? n37 : n1409;
  assign n1411 = pi19 ? n37 : n1410;
  assign n1412 = pi18 ? n1411 : n32;
  assign n1413 = pi17 ? n37 : n1412;
  assign n1414 = pi16 ? n439 : n1413;
  assign n1415 = pi15 ? n1403 : n1414;
  assign n1416 = pi22 ? n686 : n1407;
  assign n1417 = pi21 ? n37 : n1416;
  assign n1418 = pi20 ? n37 : n1417;
  assign n1419 = pi19 ? n37 : n1418;
  assign n1420 = pi18 ? n1419 : n32;
  assign n1421 = pi17 ? n37 : n1420;
  assign n1422 = pi16 ? n439 : n1421;
  assign n1423 = pi22 ? n685 : n1407;
  assign n1424 = pi21 ? n37 : n1423;
  assign n1425 = pi20 ? n37 : n1424;
  assign n1426 = pi19 ? n37 : n1425;
  assign n1427 = pi18 ? n1426 : n32;
  assign n1428 = pi17 ? n37 : n1427;
  assign n1429 = pi16 ? n439 : n1428;
  assign n1430 = pi15 ? n1422 : n1429;
  assign n1431 = pi14 ? n1415 : n1430;
  assign n1432 = pi24 ? n37 : n363;
  assign n1433 = pi23 ? n1432 : n316;
  assign n1434 = pi22 ? n1433 : n317;
  assign n1435 = pi21 ? n37 : n1434;
  assign n1436 = pi20 ? n37 : n1435;
  assign n1437 = pi19 ? n37 : n1436;
  assign n1438 = pi18 ? n1437 : n32;
  assign n1439 = pi17 ? n37 : n1438;
  assign n1440 = pi16 ? n439 : n1439;
  assign n1441 = pi22 ? n705 : n317;
  assign n1442 = pi21 ? n722 : n1441;
  assign n1443 = pi20 ? n99 : n1442;
  assign n1444 = pi19 ? n227 : n1443;
  assign n1445 = pi18 ? n1444 : n32;
  assign n1446 = pi17 ? n99 : n1445;
  assign n1447 = pi16 ? n721 : n1446;
  assign n1448 = pi15 ? n1440 : n1447;
  assign n1449 = pi23 ? n685 : n204;
  assign n1450 = pi22 ? n1449 : n688;
  assign n1451 = pi21 ? n99 : n1450;
  assign n1452 = pi20 ? n99 : n1451;
  assign n1453 = pi19 ? n99 : n1452;
  assign n1454 = pi18 ? n1453 : n32;
  assign n1455 = pi17 ? n99 : n1454;
  assign n1456 = pi16 ? n721 : n1455;
  assign n1457 = pi23 ? n157 : n233;
  assign n1458 = pi22 ? n1457 : n688;
  assign n1459 = pi21 ? n99 : n1458;
  assign n1460 = pi20 ? n99 : n1459;
  assign n1461 = pi19 ? n99 : n1460;
  assign n1462 = pi18 ? n1461 : n32;
  assign n1463 = pi17 ? n99 : n1462;
  assign n1464 = pi16 ? n744 : n1463;
  assign n1465 = pi15 ? n1456 : n1464;
  assign n1466 = pi14 ? n1448 : n1465;
  assign n1467 = pi13 ? n1431 : n1466;
  assign n1468 = pi12 ? n1406 : n1467;
  assign n1469 = pi21 ? n99 : n696;
  assign n1470 = pi20 ? n99 : n1469;
  assign n1471 = pi19 ? n99 : n1470;
  assign n1472 = pi18 ? n1471 : n32;
  assign n1473 = pi17 ? n99 : n1472;
  assign n1474 = pi16 ? n744 : n1473;
  assign n1475 = pi23 ? n685 : n316;
  assign n1476 = pi22 ? n1475 : n706;
  assign n1477 = pi21 ? n767 : n1476;
  assign n1478 = pi20 ? n99 : n1477;
  assign n1479 = pi19 ? n99 : n1478;
  assign n1480 = pi18 ? n1479 : n32;
  assign n1481 = pi17 ? n99 : n1480;
  assign n1482 = pi16 ? n744 : n1481;
  assign n1483 = pi15 ? n1474 : n1482;
  assign n1484 = pi23 ? n157 : n316;
  assign n1485 = pi22 ? n1484 : n32;
  assign n1486 = pi21 ? n777 : n1485;
  assign n1487 = pi20 ? n776 : n1486;
  assign n1488 = pi19 ? n99 : n1487;
  assign n1489 = pi18 ? n1488 : n32;
  assign n1490 = pi17 ? n99 : n1489;
  assign n1491 = pi16 ? n744 : n1490;
  assign n1492 = pi21 ? n99 : n168;
  assign n1493 = pi20 ? n1492 : n99;
  assign n1494 = pi19 ? n99 : n1493;
  assign n1495 = pi18 ? n1494 : n99;
  assign n1496 = pi21 ? n157 : n748;
  assign n1497 = pi20 ? n787 : n1496;
  assign n1498 = pi19 ? n99 : n1497;
  assign n1499 = pi18 ? n1498 : n32;
  assign n1500 = pi17 ? n1495 : n1499;
  assign n1501 = pi16 ? n721 : n1500;
  assign n1502 = pi15 ? n1491 : n1501;
  assign n1503 = pi14 ? n1483 : n1502;
  assign n1504 = pi23 ? n714 : n37;
  assign n1505 = pi22 ? n1504 : n99;
  assign n1506 = pi21 ? n1505 : n99;
  assign n1507 = pi20 ? n32 : n1506;
  assign n1508 = pi19 ? n32 : n1507;
  assign n1509 = pi18 ? n1508 : n99;
  assign n1510 = pi17 ? n32 : n1509;
  assign n1511 = pi23 ? n157 : n687;
  assign n1512 = pi22 ? n1511 : n32;
  assign n1513 = pi21 ? n157 : n1512;
  assign n1514 = pi20 ? n776 : n1513;
  assign n1515 = pi19 ? n99 : n1514;
  assign n1516 = pi18 ? n1515 : n32;
  assign n1517 = pi17 ? n805 : n1516;
  assign n1518 = pi16 ? n1510 : n1517;
  assign n1519 = pi23 ? n961 : n37;
  assign n1520 = pi22 ? n1519 : n745;
  assign n1521 = pi22 ? n112 : n1043;
  assign n1522 = pi21 ? n1520 : n1521;
  assign n1523 = pi20 ? n32 : n1522;
  assign n1524 = pi19 ? n32 : n1523;
  assign n1525 = pi21 ? n894 : n258;
  assign n1526 = pi22 ? n295 : n157;
  assign n1527 = pi21 ? n1526 : n820;
  assign n1528 = pi20 ? n1525 : n1527;
  assign n1529 = pi22 ? n295 : n1043;
  assign n1530 = pi21 ? n1529 : n248;
  assign n1531 = pi22 ? n139 : n295;
  assign n1532 = pi21 ? n1521 : n1531;
  assign n1533 = pi20 ? n1530 : n1532;
  assign n1534 = pi19 ? n1528 : n1533;
  assign n1535 = pi18 ? n1524 : n1534;
  assign n1536 = pi17 ? n32 : n1535;
  assign n1537 = pi22 ? n889 : n139;
  assign n1538 = pi21 ? n157 : n1537;
  assign n1539 = pi21 ? n831 : n157;
  assign n1540 = pi20 ? n1538 : n1539;
  assign n1541 = pi19 ? n157 : n1540;
  assign n1542 = pi18 ? n834 : n1541;
  assign n1543 = pi20 ? n157 : n1513;
  assign n1544 = pi19 ? n157 : n1543;
  assign n1545 = pi18 ? n1544 : n32;
  assign n1546 = pi17 ? n1542 : n1545;
  assign n1547 = pi16 ? n1536 : n1546;
  assign n1548 = pi15 ? n1518 : n1547;
  assign n1549 = pi22 ? n1519 : n139;
  assign n1550 = pi21 ? n1549 : n853;
  assign n1551 = pi20 ? n32 : n1550;
  assign n1552 = pi19 ? n32 : n1551;
  assign n1553 = pi18 ? n1552 : n866;
  assign n1554 = pi17 ? n32 : n1553;
  assign n1555 = pi16 ? n1554 : n887;
  assign n1556 = pi15 ? n1555 : n905;
  assign n1557 = pi14 ? n1548 : n1556;
  assign n1558 = pi13 ? n1503 : n1557;
  assign n1559 = pi18 ? n913 : n967;
  assign n1560 = pi17 ? n32 : n1559;
  assign n1561 = pi16 ? n1560 : n973;
  assign n1562 = pi15 ? n1561 : n985;
  assign n1563 = pi14 ? n960 : n1562;
  assign n1564 = pi22 ? n1519 : n37;
  assign n1565 = pi21 ? n1564 : n139;
  assign n1566 = pi20 ? n32 : n1565;
  assign n1567 = pi19 ? n32 : n1566;
  assign n1568 = pi18 ? n1567 : n994;
  assign n1569 = pi17 ? n32 : n1568;
  assign n1570 = pi16 ? n1569 : n1014;
  assign n1571 = pi21 ? n1549 : n139;
  assign n1572 = pi20 ? n32 : n1571;
  assign n1573 = pi19 ? n32 : n1572;
  assign n1574 = pi18 ? n1573 : n139;
  assign n1575 = pi17 ? n32 : n1574;
  assign n1576 = pi16 ? n1575 : n1034;
  assign n1577 = pi15 ? n1570 : n1576;
  assign n1578 = pi22 ? n456 : n204;
  assign n1579 = pi21 ? n1037 : n1578;
  assign n1580 = pi20 ? n32 : n1579;
  assign n1581 = pi19 ? n32 : n1580;
  assign n1582 = pi21 ? n1046 : n204;
  assign n1583 = pi21 ? n1046 : n37;
  assign n1584 = pi20 ? n1582 : n1583;
  assign n1585 = pi20 ? n1046 : n1057;
  assign n1586 = pi19 ? n1584 : n1585;
  assign n1587 = pi18 ? n1581 : n1586;
  assign n1588 = pi17 ? n32 : n1587;
  assign n1589 = pi16 ? n1588 : n1076;
  assign n1590 = pi24 ? n32 : n335;
  assign n1591 = pi23 ? n1590 : n99;
  assign n1592 = pi22 ? n1591 : n335;
  assign n1593 = pi21 ? n1592 : n1079;
  assign n1594 = pi20 ? n32 : n1593;
  assign n1595 = pi19 ? n32 : n1594;
  assign n1596 = pi18 ? n1595 : n1086;
  assign n1597 = pi17 ? n32 : n1596;
  assign n1598 = pi24 ? n204 : n685;
  assign n1599 = pi23 ? n1598 : n316;
  assign n1600 = pi22 ? n204 : n1599;
  assign n1601 = pi21 ? n1600 : n32;
  assign n1602 = pi20 ? n204 : n1601;
  assign n1603 = pi19 ? n1100 : n1602;
  assign n1604 = pi18 ? n1603 : n32;
  assign n1605 = pi17 ? n1098 : n1604;
  assign n1606 = pi16 ? n1597 : n1605;
  assign n1607 = pi15 ? n1589 : n1606;
  assign n1608 = pi14 ? n1577 : n1607;
  assign n1609 = pi13 ? n1563 : n1608;
  assign n1610 = pi12 ? n1558 : n1609;
  assign n1611 = pi11 ? n1468 : n1610;
  assign n1612 = pi10 ? n1363 : n1611;
  assign n1613 = pi09 ? n32 : n1612;
  assign n1614 = pi08 ? n1113 : n1613;
  assign n1615 = pi07 ? n32 : n1614;
  assign n1616 = pi06 ? n32 : n1615;
  assign n1617 = pi23 ? n37 : n46;
  assign n1618 = pi22 ? n37 : n1617;
  assign n1619 = pi21 ? n37 : n1618;
  assign n1620 = pi20 ? n37 : n1619;
  assign n1621 = pi19 ? n37 : n1620;
  assign n1622 = pi18 ? n1621 : n32;
  assign n1623 = pi17 ? n37 : n1622;
  assign n1624 = pi16 ? n1118 : n1623;
  assign n1625 = pi15 ? n32 : n1624;
  assign n1626 = pi14 ? n32 : n1625;
  assign n1627 = pi16 ? n61 : n1623;
  assign n1628 = pi16 ? n70 : n1623;
  assign n1629 = pi15 ? n1627 : n1628;
  assign n1630 = pi16 ? n73 : n1623;
  assign n1631 = pi18 ? n37 : n32;
  assign n1632 = pi17 ? n37 : n1631;
  assign n1633 = pi16 ? n83 : n1632;
  assign n1634 = pi15 ? n1630 : n1633;
  assign n1635 = pi14 ? n1629 : n1634;
  assign n1636 = pi13 ? n1626 : n1635;
  assign n1637 = pi16 ? n1130 : n1632;
  assign n1638 = pi22 ? n64 : n112;
  assign n1639 = pi21 ? n32 : n1638;
  assign n1640 = pi20 ? n32 : n1639;
  assign n1641 = pi19 ? n32 : n1640;
  assign n1642 = pi18 ? n1641 : n99;
  assign n1643 = pi17 ? n32 : n1642;
  assign n1644 = pi18 ? n99 : n32;
  assign n1645 = pi17 ? n99 : n1644;
  assign n1646 = pi16 ? n1643 : n1645;
  assign n1647 = pi15 ? n1637 : n1646;
  assign n1648 = pi16 ? n132 : n1645;
  assign n1649 = pi14 ? n1647 : n1648;
  assign n1650 = pi21 ? n99 : n746;
  assign n1651 = pi20 ? n169 : n1650;
  assign n1652 = pi19 ? n167 : n1651;
  assign n1653 = pi18 ? n1652 : n32;
  assign n1654 = pi17 ? n163 : n1653;
  assign n1655 = pi16 ? n1148 : n1654;
  assign n1656 = pi23 ? n99 : n335;
  assign n1657 = pi22 ? n99 : n1656;
  assign n1658 = pi21 ? n99 : n1657;
  assign n1659 = pi20 ? n169 : n1658;
  assign n1660 = pi19 ? n167 : n1659;
  assign n1661 = pi18 ? n1660 : n32;
  assign n1662 = pi17 ? n163 : n1661;
  assign n1663 = pi16 ? n744 : n1662;
  assign n1664 = pi15 ? n1655 : n1663;
  assign n1665 = pi21 ? n99 : n159;
  assign n1666 = pi20 ? n99 : n1665;
  assign n1667 = pi19 ? n99 : n1666;
  assign n1668 = pi18 ? n1667 : n32;
  assign n1669 = pi17 ? n99 : n1668;
  assign n1670 = pi16 ? n801 : n1669;
  assign n1671 = pi22 ? n738 : n37;
  assign n1672 = pi21 ? n1671 : n99;
  assign n1673 = pi20 ? n32 : n1672;
  assign n1674 = pi19 ? n32 : n1673;
  assign n1675 = pi18 ? n1674 : n99;
  assign n1676 = pi17 ? n32 : n1675;
  assign n1677 = pi16 ? n1676 : n1669;
  assign n1678 = pi15 ? n1670 : n1677;
  assign n1679 = pi14 ? n1664 : n1678;
  assign n1680 = pi13 ? n1649 : n1679;
  assign n1681 = pi12 ? n1636 : n1680;
  assign n1682 = pi23 ? n99 : n205;
  assign n1683 = pi22 ? n99 : n1682;
  assign n1684 = pi21 ? n99 : n1683;
  assign n1685 = pi20 ? n99 : n1684;
  assign n1686 = pi19 ? n99 : n1685;
  assign n1687 = pi18 ? n1686 : n32;
  assign n1688 = pi17 ? n99 : n1687;
  assign n1689 = pi16 ? n744 : n1688;
  assign n1690 = pi21 ? n180 : n297;
  assign n1691 = pi20 ? n32 : n1690;
  assign n1692 = pi19 ? n32 : n1691;
  assign n1693 = pi21 ? n375 : n1211;
  assign n1694 = pi21 ? n375 : n1043;
  assign n1695 = pi20 ? n1693 : n1694;
  assign n1696 = pi22 ? n37 : n1043;
  assign n1697 = pi21 ? n295 : n1696;
  assign n1698 = pi22 ? n1043 : n295;
  assign n1699 = pi21 ? n1698 : n375;
  assign n1700 = pi20 ? n1697 : n1699;
  assign n1701 = pi19 ? n1695 : n1700;
  assign n1702 = pi18 ? n1692 : n1701;
  assign n1703 = pi17 ? n32 : n1702;
  assign n1704 = pi21 ? n1043 : n295;
  assign n1705 = pi21 ? n1696 : n1698;
  assign n1706 = pi20 ? n1704 : n1705;
  assign n1707 = pi21 ? n1529 : n1211;
  assign n1708 = pi21 ? n295 : n139;
  assign n1709 = pi20 ? n1707 : n1708;
  assign n1710 = pi19 ? n1706 : n1709;
  assign n1711 = pi22 ? n139 : n1043;
  assign n1712 = pi21 ? n1711 : n1211;
  assign n1713 = pi20 ? n1708 : n1712;
  assign n1714 = pi21 ? n295 : n1211;
  assign n1715 = pi21 ? n1531 : n1211;
  assign n1716 = pi20 ? n1714 : n1715;
  assign n1717 = pi19 ? n1713 : n1716;
  assign n1718 = pi18 ? n1710 : n1717;
  assign n1719 = pi21 ? n1531 : n139;
  assign n1720 = pi20 ? n1719 : n139;
  assign n1721 = pi22 ? n295 : n139;
  assign n1722 = pi21 ? n1043 : n1721;
  assign n1723 = pi23 ? n139 : n234;
  assign n1724 = pi22 ? n295 : n1723;
  assign n1725 = pi21 ? n1043 : n1724;
  assign n1726 = pi20 ? n1722 : n1725;
  assign n1727 = pi19 ? n1720 : n1726;
  assign n1728 = pi18 ? n1727 : n32;
  assign n1729 = pi17 ? n1718 : n1728;
  assign n1730 = pi16 ? n1703 : n1729;
  assign n1731 = pi15 ? n1689 : n1730;
  assign n1732 = pi21 ? n180 : n1211;
  assign n1733 = pi20 ? n32 : n1732;
  assign n1734 = pi19 ? n32 : n1733;
  assign n1735 = pi21 ? n295 : n1043;
  assign n1736 = pi20 ? n1714 : n1735;
  assign n1737 = pi21 ? n1531 : n1529;
  assign n1738 = pi21 ? n1211 : n295;
  assign n1739 = pi20 ? n1737 : n1738;
  assign n1740 = pi19 ? n1736 : n1739;
  assign n1741 = pi18 ? n1734 : n1740;
  assign n1742 = pi17 ? n32 : n1741;
  assign n1743 = pi21 ? n1043 : n1531;
  assign n1744 = pi20 ? n1743 : n1707;
  assign n1745 = pi19 ? n1744 : n1709;
  assign n1746 = pi18 ? n1745 : n1717;
  assign n1747 = pi21 ? n1043 : n139;
  assign n1748 = pi24 ? n139 : n685;
  assign n1749 = pi23 ? n37 : n1748;
  assign n1750 = pi22 ? n139 : n1749;
  assign n1751 = pi21 ? n1043 : n1750;
  assign n1752 = pi20 ? n1747 : n1751;
  assign n1753 = pi19 ? n1720 : n1752;
  assign n1754 = pi18 ? n1753 : n32;
  assign n1755 = pi17 ? n1746 : n1754;
  assign n1756 = pi16 ? n1742 : n1755;
  assign n1757 = pi21 ? n820 : n1211;
  assign n1758 = pi20 ? n1708 : n1757;
  assign n1759 = pi19 ? n1758 : n1716;
  assign n1760 = pi18 ? n1745 : n1759;
  assign n1761 = pi21 ? n1696 : n139;
  assign n1762 = pi23 ? n37 : n260;
  assign n1763 = pi22 ? n139 : n1762;
  assign n1764 = pi21 ? n1043 : n1763;
  assign n1765 = pi20 ? n1761 : n1764;
  assign n1766 = pi19 ? n1720 : n1765;
  assign n1767 = pi18 ? n1766 : n32;
  assign n1768 = pi17 ? n1760 : n1767;
  assign n1769 = pi16 ? n1742 : n1768;
  assign n1770 = pi15 ? n1756 : n1769;
  assign n1771 = pi14 ? n1731 : n1770;
  assign n1772 = pi18 ? n990 : n139;
  assign n1773 = pi17 ? n32 : n1772;
  assign n1774 = pi22 ? n139 : n390;
  assign n1775 = pi21 ? n139 : n1774;
  assign n1776 = pi20 ? n139 : n1775;
  assign n1777 = pi22 ? n139 : n383;
  assign n1778 = pi21 ? n139 : n1777;
  assign n1779 = pi20 ? n139 : n1778;
  assign n1780 = pi19 ? n1776 : n1779;
  assign n1781 = pi18 ? n1780 : n32;
  assign n1782 = pi17 ? n139 : n1781;
  assign n1783 = pi16 ? n1773 : n1782;
  assign n1784 = pi23 ? n139 : n316;
  assign n1785 = pi22 ? n139 : n1784;
  assign n1786 = pi21 ? n139 : n1785;
  assign n1787 = pi20 ? n139 : n1786;
  assign n1788 = pi19 ? n139 : n1787;
  assign n1789 = pi18 ? n1788 : n32;
  assign n1790 = pi17 ? n139 : n1789;
  assign n1791 = pi16 ? n331 : n1790;
  assign n1792 = pi15 ? n1783 : n1791;
  assign n1793 = pi22 ? n139 : n1038;
  assign n1794 = pi21 ? n139 : n1793;
  assign n1795 = pi20 ? n139 : n1794;
  assign n1796 = pi19 ? n139 : n1795;
  assign n1797 = pi18 ? n1796 : n32;
  assign n1798 = pi17 ? n139 : n1797;
  assign n1799 = pi16 ? n331 : n1798;
  assign n1800 = pi20 ? n992 : n139;
  assign n1801 = pi19 ? n1800 : n139;
  assign n1802 = pi18 ? n329 : n1801;
  assign n1803 = pi17 ? n32 : n1802;
  assign n1804 = pi20 ? n947 : n939;
  assign n1805 = pi19 ? n139 : n1804;
  assign n1806 = pi20 ? n939 : n139;
  assign n1807 = pi19 ? n1806 : n992;
  assign n1808 = pi18 ? n1805 : n1807;
  assign n1809 = pi20 ? n139 : n942;
  assign n1810 = pi22 ? n139 : n456;
  assign n1811 = pi21 ? n139 : n1810;
  assign n1812 = pi20 ? n992 : n1811;
  assign n1813 = pi19 ? n1809 : n1812;
  assign n1814 = pi18 ? n1813 : n32;
  assign n1815 = pi17 ? n1808 : n1814;
  assign n1816 = pi16 ? n1803 : n1815;
  assign n1817 = pi15 ? n1799 : n1816;
  assign n1818 = pi14 ? n1792 : n1817;
  assign n1819 = pi13 ? n1771 : n1818;
  assign n1820 = pi20 ? n139 : n347;
  assign n1821 = pi19 ? n139 : n1820;
  assign n1822 = pi21 ? n1009 : n32;
  assign n1823 = pi20 ? n1822 : n32;
  assign n1824 = pi19 ? n1823 : n32;
  assign n1825 = pi18 ? n1821 : n1824;
  assign n1826 = pi17 ? n139 : n1825;
  assign n1827 = pi16 ? n331 : n1826;
  assign n1828 = pi22 ? n1043 : n455;
  assign n1829 = pi21 ? n296 : n1828;
  assign n1830 = pi20 ? n32 : n1829;
  assign n1831 = pi19 ? n32 : n1830;
  assign n1832 = pi22 ? n918 : n456;
  assign n1833 = pi21 ? n1832 : n520;
  assign n1834 = pi22 ? n456 : n1043;
  assign n1835 = pi21 ? n1832 : n1834;
  assign n1836 = pi20 ? n1833 : n1835;
  assign n1837 = pi22 ? n455 : n918;
  assign n1838 = pi21 ? n1837 : n456;
  assign n1839 = pi21 ? n1828 : n1832;
  assign n1840 = pi20 ? n1838 : n1839;
  assign n1841 = pi19 ? n1836 : n1840;
  assign n1842 = pi18 ? n1831 : n1841;
  assign n1843 = pi17 ? n32 : n1842;
  assign n1844 = pi21 ? n1834 : n1837;
  assign n1845 = pi21 ? n456 : n1828;
  assign n1846 = pi20 ? n1844 : n1845;
  assign n1847 = pi22 ? n918 : n295;
  assign n1848 = pi21 ? n1847 : n1828;
  assign n1849 = pi21 ? n1832 : n1696;
  assign n1850 = pi20 ? n1848 : n1849;
  assign n1851 = pi19 ? n1846 : n1850;
  assign n1852 = pi21 ? n1810 : n1828;
  assign n1853 = pi20 ? n1849 : n1852;
  assign n1854 = pi21 ? n1810 : n1834;
  assign n1855 = pi20 ? n1835 : n1854;
  assign n1856 = pi19 ? n1853 : n1855;
  assign n1857 = pi18 ? n1851 : n1856;
  assign n1858 = pi21 ? n1810 : n506;
  assign n1859 = pi20 ? n1858 : n1757;
  assign n1860 = pi22 ? n455 : n139;
  assign n1861 = pi21 ? n1834 : n1860;
  assign n1862 = pi21 ? n1834 : n522;
  assign n1863 = pi20 ? n1861 : n1862;
  assign n1864 = pi19 ? n1859 : n1863;
  assign n1865 = pi18 ? n1864 : n1824;
  assign n1866 = pi17 ? n1857 : n1865;
  assign n1867 = pi16 ? n1843 : n1866;
  assign n1868 = pi15 ? n1827 : n1867;
  assign n1869 = pi22 ? n55 : n583;
  assign n1870 = pi21 ? n1869 : n506;
  assign n1871 = pi20 ? n32 : n1870;
  assign n1872 = pi19 ? n32 : n1871;
  assign n1873 = pi20 ? n1326 : n514;
  assign n1874 = pi20 ? n504 : n507;
  assign n1875 = pi19 ? n1873 : n1874;
  assign n1876 = pi18 ? n1872 : n1875;
  assign n1877 = pi17 ? n32 : n1876;
  assign n1878 = pi20 ? n508 : n513;
  assign n1879 = pi22 ? n450 : n583;
  assign n1880 = pi21 ? n1879 : n506;
  assign n1881 = pi21 ? n457 : n580;
  assign n1882 = pi20 ? n1880 : n1881;
  assign n1883 = pi19 ? n1878 : n1882;
  assign n1884 = pi22 ? n335 : n456;
  assign n1885 = pi21 ? n1884 : n506;
  assign n1886 = pi20 ? n1881 : n1885;
  assign n1887 = pi22 ? n566 : n456;
  assign n1888 = pi21 ? n1887 : n499;
  assign n1889 = pi20 ? n514 : n1888;
  assign n1890 = pi19 ? n1886 : n1889;
  assign n1891 = pi18 ? n1883 : n1890;
  assign n1892 = pi21 ? n1887 : n506;
  assign n1893 = pi21 ? n570 : n567;
  assign n1894 = pi20 ? n1892 : n1893;
  assign n1895 = pi22 ? n455 : n335;
  assign n1896 = pi21 ? n499 : n1895;
  assign n1897 = pi21 ? n499 : n457;
  assign n1898 = pi20 ? n1896 : n1897;
  assign n1899 = pi19 ? n1894 : n1898;
  assign n1900 = pi18 ? n1899 : n1824;
  assign n1901 = pi17 ? n1891 : n1900;
  assign n1902 = pi16 ? n1877 : n1901;
  assign n1903 = pi21 ? n180 : n1046;
  assign n1904 = pi20 ? n32 : n1903;
  assign n1905 = pi19 ? n32 : n1904;
  assign n1906 = pi21 ? n1056 : n1046;
  assign n1907 = pi20 ? n1906 : n37;
  assign n1908 = pi19 ? n1907 : n37;
  assign n1909 = pi18 ? n1905 : n1908;
  assign n1910 = pi17 ? n32 : n1909;
  assign n1911 = pi21 ? n37 : n1046;
  assign n1912 = pi21 ? n37 : n1056;
  assign n1913 = pi20 ? n1911 : n1912;
  assign n1914 = pi19 ? n37 : n1913;
  assign n1915 = pi20 ? n1912 : n1583;
  assign n1916 = pi20 ? n37 : n1583;
  assign n1917 = pi19 ? n1915 : n1916;
  assign n1918 = pi18 ? n1914 : n1917;
  assign n1919 = pi20 ? n204 : n1582;
  assign n1920 = pi22 ? n37 : n559;
  assign n1921 = pi21 ? n37 : n1920;
  assign n1922 = pi20 ? n1912 : n1921;
  assign n1923 = pi19 ? n1919 : n1922;
  assign n1924 = pi18 ? n1923 : n1824;
  assign n1925 = pi17 ? n1918 : n1924;
  assign n1926 = pi16 ? n1910 : n1925;
  assign n1927 = pi15 ? n1902 : n1926;
  assign n1928 = pi14 ? n1868 : n1927;
  assign n1929 = pi22 ? n450 : n335;
  assign n1930 = pi21 ? n555 : n1929;
  assign n1931 = pi20 ? n32 : n1930;
  assign n1932 = pi19 ? n32 : n1931;
  assign n1933 = pi18 ? n1932 : n335;
  assign n1934 = pi17 ? n32 : n1933;
  assign n1935 = pi21 ? n567 : n1929;
  assign n1936 = pi22 ? n583 : n204;
  assign n1937 = pi21 ? n335 : n1936;
  assign n1938 = pi20 ? n1935 : n1937;
  assign n1939 = pi19 ? n335 : n1938;
  assign n1940 = pi22 ? n448 : n335;
  assign n1941 = pi21 ? n1940 : n335;
  assign n1942 = pi20 ? n1937 : n1941;
  assign n1943 = pi22 ? n335 : n583;
  assign n1944 = pi21 ? n335 : n1943;
  assign n1945 = pi21 ? n485 : n1943;
  assign n1946 = pi20 ? n1944 : n1945;
  assign n1947 = pi19 ? n1942 : n1946;
  assign n1948 = pi18 ? n1939 : n1947;
  assign n1949 = pi22 ? n450 : n204;
  assign n1950 = pi21 ? n485 : n1949;
  assign n1951 = pi22 ? n448 : n583;
  assign n1952 = pi21 ? n1951 : n474;
  assign n1953 = pi20 ? n1950 : n1952;
  assign n1954 = pi21 ? n335 : n474;
  assign n1955 = pi23 ? n335 : n1598;
  assign n1956 = pi22 ? n204 : n1955;
  assign n1957 = pi21 ? n335 : n1956;
  assign n1958 = pi20 ? n1954 : n1957;
  assign n1959 = pi19 ? n1953 : n1958;
  assign n1960 = pi18 ? n1959 : n32;
  assign n1961 = pi17 ? n1948 : n1960;
  assign n1962 = pi16 ? n1934 : n1961;
  assign n1963 = pi21 ? n449 : n583;
  assign n1964 = pi20 ? n32 : n1963;
  assign n1965 = pi19 ? n32 : n1964;
  assign n1966 = pi22 ? n204 : n566;
  assign n1967 = pi21 ? n1966 : n1943;
  assign n1968 = pi21 ? n1936 : n567;
  assign n1969 = pi21 ? n583 : n1966;
  assign n1970 = pi20 ? n1968 : n1969;
  assign n1971 = pi19 ? n1967 : n1970;
  assign n1972 = pi18 ? n1965 : n1971;
  assign n1973 = pi17 ? n32 : n1972;
  assign n1974 = pi21 ? n1943 : n1936;
  assign n1975 = pi21 ? n567 : n583;
  assign n1976 = pi20 ? n1974 : n1975;
  assign n1977 = pi21 ? n474 : n583;
  assign n1978 = pi22 ? n583 : n450;
  assign n1979 = pi21 ? n474 : n1978;
  assign n1980 = pi20 ? n1977 : n1979;
  assign n1981 = pi19 ? n1976 : n1980;
  assign n1982 = pi21 ? n474 : n1936;
  assign n1983 = pi21 ? n1940 : n583;
  assign n1984 = pi20 ? n1982 : n1983;
  assign n1985 = pi21 ? n1966 : n476;
  assign n1986 = pi19 ? n1984 : n1985;
  assign n1987 = pi18 ? n1981 : n1986;
  assign n1988 = pi21 ? n1940 : n474;
  assign n1989 = pi20 ? n1982 : n1988;
  assign n1990 = pi21 ? n1943 : n474;
  assign n1991 = pi24 ? n335 : n316;
  assign n1992 = pi23 ? n335 : n1991;
  assign n1993 = pi22 ? n204 : n1992;
  assign n1994 = pi21 ? n1943 : n1993;
  assign n1995 = pi20 ? n1990 : n1994;
  assign n1996 = pi19 ? n1989 : n1995;
  assign n1997 = pi18 ? n1996 : n32;
  assign n1998 = pi17 ? n1987 : n1997;
  assign n1999 = pi16 ? n1973 : n1998;
  assign n2000 = pi15 ? n1962 : n1999;
  assign n2001 = pi21 ? n555 : n583;
  assign n2002 = pi20 ? n32 : n2001;
  assign n2003 = pi19 ? n32 : n2002;
  assign n2004 = pi21 ? n580 : n335;
  assign n2005 = pi21 ? n580 : n1943;
  assign n2006 = pi20 ? n2004 : n2005;
  assign n2007 = pi22 ? n583 : n37;
  assign n2008 = pi21 ? n2007 : n567;
  assign n2009 = pi21 ? n583 : n580;
  assign n2010 = pi20 ? n2008 : n2009;
  assign n2011 = pi19 ? n2006 : n2010;
  assign n2012 = pi18 ? n2003 : n2011;
  assign n2013 = pi17 ? n32 : n2012;
  assign n2014 = pi21 ? n1943 : n2007;
  assign n2015 = pi20 ? n2014 : n1975;
  assign n2016 = pi21 ? n569 : n583;
  assign n2017 = pi20 ? n2016 : n2005;
  assign n2018 = pi19 ? n2015 : n2017;
  assign n2019 = pi21 ? n580 : n570;
  assign n2020 = pi20 ? n2019 : n1975;
  assign n2021 = pi19 ? n2020 : n2005;
  assign n2022 = pi18 ? n2018 : n2021;
  assign n2023 = pi21 ? n567 : n580;
  assign n2024 = pi20 ? n571 : n2023;
  assign n2025 = pi21 ? n1943 : n580;
  assign n2026 = pi23 ? n335 : n586;
  assign n2027 = pi22 ? n37 : n2026;
  assign n2028 = pi21 ? n1943 : n2027;
  assign n2029 = pi20 ? n2025 : n2028;
  assign n2030 = pi19 ? n2024 : n2029;
  assign n2031 = pi18 ? n2030 : n32;
  assign n2032 = pi17 ? n2022 : n2031;
  assign n2033 = pi16 ? n2013 : n2032;
  assign n2034 = pi18 ? n602 : n335;
  assign n2035 = pi17 ? n32 : n2034;
  assign n2036 = pi22 ? n335 : n2026;
  assign n2037 = pi21 ? n335 : n2036;
  assign n2038 = pi20 ? n335 : n2037;
  assign n2039 = pi19 ? n335 : n2038;
  assign n2040 = pi18 ? n2039 : n32;
  assign n2041 = pi17 ? n335 : n2040;
  assign n2042 = pi16 ? n2035 : n2041;
  assign n2043 = pi15 ? n2033 : n2042;
  assign n2044 = pi14 ? n2000 : n2043;
  assign n2045 = pi13 ? n1928 : n2044;
  assign n2046 = pi12 ? n1819 : n2045;
  assign n2047 = pi11 ? n1681 : n2046;
  assign n2048 = pi22 ? n233 : n37;
  assign n2049 = pi21 ? n37 : n2048;
  assign n2050 = pi20 ? n2049 : n37;
  assign n2051 = pi19 ? n2050 : n37;
  assign n2052 = pi18 ? n558 : n2051;
  assign n2053 = pi17 ? n32 : n2052;
  assign n2054 = pi20 ? n647 : n603;
  assign n2055 = pi19 ? n37 : n2054;
  assign n2056 = pi20 ? n571 : n647;
  assign n2057 = pi19 ? n2056 : n577;
  assign n2058 = pi18 ? n2055 : n2057;
  assign n2059 = pi20 ? n610 : n605;
  assign n2060 = pi23 ? n335 : n233;
  assign n2061 = pi22 ? n335 : n2060;
  assign n2062 = pi21 ? n335 : n2061;
  assign n2063 = pi20 ? n605 : n2062;
  assign n2064 = pi19 ? n2059 : n2063;
  assign n2065 = pi18 ? n2064 : n32;
  assign n2066 = pi17 ? n2058 : n2065;
  assign n2067 = pi16 ? n2053 : n2066;
  assign n2068 = pi20 ? n647 : n577;
  assign n2069 = pi19 ? n37 : n2068;
  assign n2070 = pi20 ? n577 : n647;
  assign n2071 = pi19 ? n2070 : n577;
  assign n2072 = pi18 ? n2069 : n2071;
  assign n2073 = pi20 ? n647 : n335;
  assign n2074 = pi22 ? n37 : n2060;
  assign n2075 = pi21 ? n335 : n2074;
  assign n2076 = pi20 ? n335 : n2075;
  assign n2077 = pi19 ? n2073 : n2076;
  assign n2078 = pi18 ? n2077 : n32;
  assign n2079 = pi17 ? n2072 : n2078;
  assign n2080 = pi16 ? n439 : n2079;
  assign n2081 = pi15 ? n2067 : n2080;
  assign n2082 = pi19 ? n643 : n577;
  assign n2083 = pi18 ? n641 : n2082;
  assign n2084 = pi22 ? n37 : n673;
  assign n2085 = pi21 ? n37 : n2084;
  assign n2086 = pi20 ? n577 : n2085;
  assign n2087 = pi19 ? n2073 : n2086;
  assign n2088 = pi18 ? n2087 : n32;
  assign n2089 = pi17 ? n2083 : n2088;
  assign n2090 = pi16 ? n439 : n2089;
  assign n2091 = pi22 ? n37 : n233;
  assign n2092 = pi21 ? n2091 : n37;
  assign n2093 = pi20 ? n2092 : n37;
  assign n2094 = pi21 ? n37 : n2091;
  assign n2095 = pi20 ? n37 : n2094;
  assign n2096 = pi19 ? n2093 : n2095;
  assign n2097 = pi18 ? n2096 : n32;
  assign n2098 = pi17 ? n37 : n2097;
  assign n2099 = pi16 ? n439 : n2098;
  assign n2100 = pi15 ? n2090 : n2099;
  assign n2101 = pi14 ? n2081 : n2100;
  assign n2102 = pi19 ? n37 : n2095;
  assign n2103 = pi18 ? n2102 : n32;
  assign n2104 = pi17 ? n37 : n2103;
  assign n2105 = pi16 ? n439 : n2104;
  assign n2106 = pi22 ? n37 : n685;
  assign n2107 = pi21 ? n37 : n2106;
  assign n2108 = pi20 ? n37 : n2107;
  assign n2109 = pi19 ? n37 : n2108;
  assign n2110 = pi18 ? n2109 : n32;
  assign n2111 = pi17 ? n37 : n2110;
  assign n2112 = pi16 ? n439 : n2111;
  assign n2113 = pi20 ? n37 : n1921;
  assign n2114 = pi19 ? n37 : n2113;
  assign n2115 = pi18 ? n37 : n2114;
  assign n2116 = pi23 ? n233 : n37;
  assign n2117 = pi22 ? n2116 : n559;
  assign n2118 = pi21 ? n2117 : n37;
  assign n2119 = pi20 ? n37 : n2118;
  assign n2120 = pi24 ? n233 : n316;
  assign n2121 = pi23 ? n233 : n2120;
  assign n2122 = pi22 ? n363 : n2121;
  assign n2123 = pi21 ? n37 : n2122;
  assign n2124 = pi20 ? n37 : n2123;
  assign n2125 = pi19 ? n2119 : n2124;
  assign n2126 = pi18 ? n2125 : n32;
  assign n2127 = pi17 ? n2115 : n2126;
  assign n2128 = pi16 ? n439 : n2127;
  assign n2129 = pi15 ? n2112 : n2128;
  assign n2130 = pi14 ? n2105 : n2129;
  assign n2131 = pi13 ? n2101 : n2130;
  assign n2132 = pi22 ? n363 : n1388;
  assign n2133 = pi21 ? n37 : n2132;
  assign n2134 = pi20 ? n37 : n2133;
  assign n2135 = pi19 ? n37 : n2134;
  assign n2136 = pi18 ? n2135 : n32;
  assign n2137 = pi17 ? n37 : n2136;
  assign n2138 = pi16 ? n439 : n2137;
  assign n2139 = pi22 ? n363 : n759;
  assign n2140 = pi21 ? n37 : n2139;
  assign n2141 = pi20 ? n37 : n2140;
  assign n2142 = pi19 ? n37 : n2141;
  assign n2143 = pi18 ? n2142 : n32;
  assign n2144 = pi17 ? n37 : n2143;
  assign n2145 = pi16 ? n439 : n2144;
  assign n2146 = pi15 ? n2138 : n2145;
  assign n2147 = pi22 ? n685 : n759;
  assign n2148 = pi21 ? n37 : n2147;
  assign n2149 = pi20 ? n37 : n2148;
  assign n2150 = pi19 ? n37 : n2149;
  assign n2151 = pi18 ? n2150 : n32;
  assign n2152 = pi17 ? n37 : n2151;
  assign n2153 = pi16 ? n439 : n2152;
  assign n2154 = pi15 ? n2145 : n2153;
  assign n2155 = pi14 ? n2146 : n2154;
  assign n2156 = pi22 ? n112 : n37;
  assign n2157 = pi21 ? n796 : n2156;
  assign n2158 = pi20 ? n32 : n2157;
  assign n2159 = pi19 ? n32 : n2158;
  assign n2160 = pi23 ? n99 : n37;
  assign n2161 = pi22 ? n2160 : n99;
  assign n2162 = pi22 ? n112 : n2160;
  assign n2163 = pi21 ? n2161 : n2162;
  assign n2164 = pi22 ? n99 : n112;
  assign n2165 = pi21 ? n2164 : n2161;
  assign n2166 = pi20 ? n2163 : n2165;
  assign n2167 = pi21 ? n2162 : n2161;
  assign n2168 = pi22 ? n2160 : n112;
  assign n2169 = pi21 ? n2162 : n2168;
  assign n2170 = pi20 ? n2167 : n2169;
  assign n2171 = pi19 ? n2166 : n2170;
  assign n2172 = pi18 ? n2159 : n2171;
  assign n2173 = pi17 ? n32 : n2172;
  assign n2174 = pi21 ? n2162 : n2164;
  assign n2175 = pi22 ? n37 : n2160;
  assign n2176 = pi21 ? n2175 : n218;
  assign n2177 = pi20 ? n2174 : n2176;
  assign n2178 = pi21 ? n2161 : n181;
  assign n2179 = pi20 ? n2178 : n2161;
  assign n2180 = pi19 ? n2177 : n2179;
  assign n2181 = pi21 ? n181 : n1143;
  assign n2182 = pi21 ? n2162 : n218;
  assign n2183 = pi20 ? n2181 : n2182;
  assign n2184 = pi21 ? n2161 : n2175;
  assign n2185 = pi21 ? n2164 : n2175;
  assign n2186 = pi20 ? n2184 : n2185;
  assign n2187 = pi19 ? n2183 : n2186;
  assign n2188 = pi18 ? n2180 : n2187;
  assign n2189 = pi21 ? n2162 : n99;
  assign n2190 = pi20 ? n2165 : n2189;
  assign n2191 = pi21 ? n99 : n1143;
  assign n2192 = pi23 ? n685 : n395;
  assign n2193 = pi22 ? n363 : n2192;
  assign n2194 = pi21 ? n99 : n2193;
  assign n2195 = pi20 ? n2191 : n2194;
  assign n2196 = pi19 ? n2190 : n2195;
  assign n2197 = pi18 ? n2196 : n32;
  assign n2198 = pi17 ? n2188 : n2197;
  assign n2199 = pi16 ? n2173 : n2198;
  assign n2200 = pi22 ? n685 : n2192;
  assign n2201 = pi21 ? n99 : n2200;
  assign n2202 = pi20 ? n99 : n2201;
  assign n2203 = pi19 ? n99 : n2202;
  assign n2204 = pi18 ? n2203 : n32;
  assign n2205 = pi17 ? n99 : n2204;
  assign n2206 = pi16 ? n744 : n2205;
  assign n2207 = pi15 ? n2199 : n2206;
  assign n2208 = pi21 ? n99 : n1423;
  assign n2209 = pi20 ? n99 : n2208;
  assign n2210 = pi19 ? n99 : n2209;
  assign n2211 = pi18 ? n2210 : n32;
  assign n2212 = pi17 ? n99 : n2211;
  assign n2213 = pi16 ? n744 : n2212;
  assign n2214 = pi21 ? n685 : n1423;
  assign n2215 = pi20 ? n99 : n2214;
  assign n2216 = pi19 ? n99 : n2215;
  assign n2217 = pi18 ? n2216 : n32;
  assign n2218 = pi17 ? n99 : n2217;
  assign n2219 = pi16 ? n744 : n2218;
  assign n2220 = pi15 ? n2213 : n2219;
  assign n2221 = pi14 ? n2207 : n2220;
  assign n2222 = pi13 ? n2155 : n2221;
  assign n2223 = pi12 ? n2131 : n2222;
  assign n2224 = pi21 ? n767 : n1423;
  assign n2225 = pi20 ? n99 : n2224;
  assign n2226 = pi19 ? n99 : n2225;
  assign n2227 = pi18 ? n2226 : n32;
  assign n2228 = pi17 ? n99 : n2227;
  assign n2229 = pi16 ? n721 : n2228;
  assign n2230 = pi22 ? n685 : n317;
  assign n2231 = pi21 ? n99 : n2230;
  assign n2232 = pi20 ? n99 : n2231;
  assign n2233 = pi19 ? n99 : n2232;
  assign n2234 = pi18 ? n2233 : n32;
  assign n2235 = pi17 ? n99 : n2234;
  assign n2236 = pi16 ? n801 : n2235;
  assign n2237 = pi15 ? n2229 : n2236;
  assign n2238 = pi21 ? n99 : n777;
  assign n2239 = pi20 ? n2238 : n802;
  assign n2240 = pi19 ? n99 : n2239;
  assign n2241 = pi18 ? n2240 : n99;
  assign n2242 = pi20 ? n99 : n2238;
  assign n2243 = pi21 ? n99 : n157;
  assign n2244 = pi23 ? n157 : n685;
  assign n2245 = pi22 ? n2244 : n706;
  assign n2246 = pi21 ? n99 : n2245;
  assign n2247 = pi20 ? n2243 : n2246;
  assign n2248 = pi19 ? n2242 : n2247;
  assign n2249 = pi18 ? n2248 : n32;
  assign n2250 = pi17 ? n2241 : n2249;
  assign n2251 = pi16 ? n801 : n2250;
  assign n2252 = pi20 ? n2238 : n99;
  assign n2253 = pi19 ? n99 : n2252;
  assign n2254 = pi18 ? n2253 : n99;
  assign n2255 = pi20 ? n99 : n776;
  assign n2256 = pi22 ? n2244 : n32;
  assign n2257 = pi21 ? n777 : n2256;
  assign n2258 = pi20 ? n787 : n2257;
  assign n2259 = pi19 ? n2255 : n2258;
  assign n2260 = pi18 ? n2259 : n32;
  assign n2261 = pi17 ? n2254 : n2260;
  assign n2262 = pi16 ? n744 : n2261;
  assign n2263 = pi15 ? n2251 : n2262;
  assign n2264 = pi14 ? n2237 : n2263;
  assign n2265 = pi20 ? n2243 : n99;
  assign n2266 = pi19 ? n99 : n2265;
  assign n2267 = pi18 ? n2266 : n99;
  assign n2268 = pi20 ? n157 : n1486;
  assign n2269 = pi19 ? n2255 : n2268;
  assign n2270 = pi18 ? n2269 : n32;
  assign n2271 = pi17 ? n2267 : n2270;
  assign n2272 = pi16 ? n721 : n2271;
  assign n2273 = pi20 ? n876 : n139;
  assign n2274 = pi19 ? n2273 : n139;
  assign n2275 = pi18 ? n913 : n2274;
  assign n2276 = pi17 ? n32 : n2275;
  assign n2277 = pi19 ? n139 : n157;
  assign n2278 = pi20 ? n259 : n157;
  assign n2279 = pi19 ? n2278 : n139;
  assign n2280 = pi18 ? n2277 : n2279;
  assign n2281 = pi21 ? n139 : n248;
  assign n2282 = pi20 ? n2281 : n157;
  assign n2283 = pi21 ? n157 : n1485;
  assign n2284 = pi20 ? n157 : n2283;
  assign n2285 = pi19 ? n2282 : n2284;
  assign n2286 = pi18 ? n2285 : n32;
  assign n2287 = pi17 ? n2280 : n2286;
  assign n2288 = pi16 ? n2276 : n2287;
  assign n2289 = pi15 ? n2272 : n2288;
  assign n2290 = pi18 ? n966 : n139;
  assign n2291 = pi17 ? n32 : n2290;
  assign n2292 = pi21 ? n258 : n139;
  assign n2293 = pi20 ? n157 : n2292;
  assign n2294 = pi19 ? n139 : n2293;
  assign n2295 = pi20 ? n2292 : n139;
  assign n2296 = pi19 ? n2295 : n139;
  assign n2297 = pi18 ? n2294 : n2296;
  assign n2298 = pi20 ? n139 : n249;
  assign n2299 = pi23 ? n204 : n316;
  assign n2300 = pi22 ? n2299 : n32;
  assign n2301 = pi21 ? n346 : n2300;
  assign n2302 = pi20 ? n157 : n2301;
  assign n2303 = pi19 ? n2298 : n2302;
  assign n2304 = pi18 ? n2303 : n32;
  assign n2305 = pi17 ? n2297 : n2304;
  assign n2306 = pi16 ? n2291 : n2305;
  assign n2307 = pi20 ? n139 : n992;
  assign n2308 = pi19 ? n2307 : n139;
  assign n2309 = pi18 ? n966 : n2308;
  assign n2310 = pi17 ? n32 : n2309;
  assign n2311 = pi20 ? n204 : n922;
  assign n2312 = pi19 ? n139 : n2311;
  assign n2313 = pi20 ? n922 : n139;
  assign n2314 = pi19 ? n2313 : n139;
  assign n2315 = pi18 ? n2312 : n2314;
  assign n2316 = pi21 ? n916 : n204;
  assign n2317 = pi20 ? n139 : n2316;
  assign n2318 = pi21 ? n204 : n139;
  assign n2319 = pi22 ? n1784 : n316;
  assign n2320 = pi22 ? n316 : n32;
  assign n2321 = pi21 ? n2319 : n2320;
  assign n2322 = pi20 ? n2318 : n2321;
  assign n2323 = pi19 ? n2317 : n2322;
  assign n2324 = pi18 ? n2323 : n32;
  assign n2325 = pi17 ? n2315 : n2324;
  assign n2326 = pi16 ? n2310 : n2325;
  assign n2327 = pi15 ? n2306 : n2326;
  assign n2328 = pi14 ? n2289 : n2327;
  assign n2329 = pi13 ? n2264 : n2328;
  assign n2330 = pi21 ? n316 : n882;
  assign n2331 = pi20 ? n139 : n2330;
  assign n2332 = pi19 ? n1017 : n2331;
  assign n2333 = pi18 ? n2332 : n32;
  assign n2334 = pi17 ? n139 : n2333;
  assign n2335 = pi16 ? n915 : n2334;
  assign n2336 = pi19 ? n992 : n139;
  assign n2337 = pi18 ? n913 : n2336;
  assign n2338 = pi17 ? n32 : n2337;
  assign n2339 = pi20 ? n975 : n2330;
  assign n2340 = pi19 ? n139 : n2339;
  assign n2341 = pi18 ? n2340 : n32;
  assign n2342 = pi17 ? n139 : n2341;
  assign n2343 = pi16 ? n2338 : n2342;
  assign n2344 = pi15 ? n2335 : n2343;
  assign n2345 = pi20 ? n1786 : n139;
  assign n2346 = pi19 ? n139 : n2345;
  assign n2347 = pi18 ? n2346 : n139;
  assign n2348 = pi17 ? n2347 : n2341;
  assign n2349 = pi16 ? n915 : n2348;
  assign n2350 = pi19 ? n1806 : n139;
  assign n2351 = pi18 ? n2346 : n2350;
  assign n2352 = pi20 ? n139 : n975;
  assign n2353 = pi21 ? n346 : n316;
  assign n2354 = pi21 ? n346 : n882;
  assign n2355 = pi20 ? n2353 : n2354;
  assign n2356 = pi19 ? n2352 : n2355;
  assign n2357 = pi18 ? n2356 : n32;
  assign n2358 = pi17 ? n2351 : n2357;
  assign n2359 = pi16 ? n915 : n2358;
  assign n2360 = pi15 ? n2349 : n2359;
  assign n2361 = pi14 ? n2344 : n2360;
  assign n2362 = pi21 ? n935 : n139;
  assign n2363 = pi20 ? n32 : n2362;
  assign n2364 = pi19 ? n32 : n2363;
  assign n2365 = pi21 ? n139 : n1531;
  assign n2366 = pi20 ? n2365 : n939;
  assign n2367 = pi19 ? n2366 : n942;
  assign n2368 = pi18 ? n2364 : n2367;
  assign n2369 = pi17 ? n32 : n2368;
  assign n2370 = pi21 ? n1777 : n346;
  assign n2371 = pi21 ? n1777 : n139;
  assign n2372 = pi20 ? n2370 : n2371;
  assign n2373 = pi19 ? n139 : n2372;
  assign n2374 = pi20 ? n297 : n139;
  assign n2375 = pi20 ? n297 : n820;
  assign n2376 = pi19 ? n2374 : n2375;
  assign n2377 = pi18 ? n2373 : n2376;
  assign n2378 = pi20 ? n1022 : n929;
  assign n2379 = pi19 ? n2352 : n2378;
  assign n2380 = pi18 ? n2379 : n32;
  assign n2381 = pi17 ? n2377 : n2380;
  assign n2382 = pi16 ? n2369 : n2381;
  assign n2383 = pi21 ? n1027 : n316;
  assign n2384 = pi20 ? n1026 : n2383;
  assign n2385 = pi19 ? n2384 : n2378;
  assign n2386 = pi18 ? n2385 : n32;
  assign n2387 = pi17 ? n139 : n2386;
  assign n2388 = pi16 ? n2291 : n2387;
  assign n2389 = pi15 ? n2382 : n2388;
  assign n2390 = pi23 ? n38 : n204;
  assign n2391 = pi22 ? n2390 : n204;
  assign n2392 = pi21 ? n2391 : n204;
  assign n2393 = pi20 ? n32 : n2392;
  assign n2394 = pi19 ? n32 : n2393;
  assign n2395 = pi22 ? n204 : n455;
  assign n2396 = pi21 ? n204 : n2395;
  assign n2397 = pi20 ? n204 : n2396;
  assign n2398 = pi19 ? n2397 : n204;
  assign n2399 = pi18 ? n2394 : n2398;
  assign n2400 = pi17 ? n32 : n2399;
  assign n2401 = pi23 ? n316 : n204;
  assign n2402 = pi22 ? n204 : n2401;
  assign n2403 = pi20 ? n2402 : n204;
  assign n2404 = pi19 ? n204 : n2403;
  assign n2405 = pi21 ? n204 : n1083;
  assign n2406 = pi20 ? n2405 : n204;
  assign n2407 = pi19 ? n2406 : n204;
  assign n2408 = pi18 ? n2404 : n2407;
  assign n2409 = pi22 ? n2401 : n316;
  assign n2410 = pi21 ? n1027 : n2409;
  assign n2411 = pi20 ? n204 : n2410;
  assign n2412 = pi22 ? n2299 : n316;
  assign n2413 = pi21 ? n2412 : n204;
  assign n2414 = pi20 ? n2413 : n1030;
  assign n2415 = pi19 ? n2411 : n2414;
  assign n2416 = pi18 ? n2415 : n32;
  assign n2417 = pi17 ? n2408 : n2416;
  assign n2418 = pi16 ? n2400 : n2417;
  assign n2419 = pi23 ? n1590 : n335;
  assign n2420 = pi22 ? n2419 : n335;
  assign n2421 = pi21 ? n2420 : n335;
  assign n2422 = pi20 ? n32 : n2421;
  assign n2423 = pi19 ? n32 : n2422;
  assign n2424 = pi18 ? n2423 : n335;
  assign n2425 = pi17 ? n32 : n2424;
  assign n2426 = pi21 ? n476 : n1079;
  assign n2427 = pi22 ? n2401 : n204;
  assign n2428 = pi21 ? n204 : n2427;
  assign n2429 = pi20 ? n2426 : n2428;
  assign n2430 = pi20 ? n204 : n1030;
  assign n2431 = pi19 ? n2429 : n2430;
  assign n2432 = pi18 ? n2431 : n32;
  assign n2433 = pi17 ? n335 : n2432;
  assign n2434 = pi16 ? n2425 : n2433;
  assign n2435 = pi15 ? n2418 : n2434;
  assign n2436 = pi14 ? n2389 : n2435;
  assign n2437 = pi13 ? n2361 : n2436;
  assign n2438 = pi12 ? n2329 : n2437;
  assign n2439 = pi11 ? n2223 : n2438;
  assign n2440 = pi10 ? n2047 : n2439;
  assign n2441 = pi09 ? n32 : n2440;
  assign n2442 = pi16 ? n61 : n1632;
  assign n2443 = pi21 ? n92 : n37;
  assign n2444 = pi20 ? n2443 : n37;
  assign n2445 = pi19 ? n2444 : n37;
  assign n2446 = pi18 ? n32 : n2445;
  assign n2447 = pi17 ? n32 : n2446;
  assign n2448 = pi16 ? n2447 : n1632;
  assign n2449 = pi15 ? n2442 : n2448;
  assign n2450 = pi14 ? n32 : n2449;
  assign n2451 = pi16 ? n70 : n1632;
  assign n2452 = pi16 ? n73 : n1632;
  assign n2453 = pi15 ? n2451 : n2452;
  assign n2454 = pi15 ? n1633 : n1637;
  assign n2455 = pi14 ? n2453 : n2454;
  assign n2456 = pi13 ? n2450 : n2455;
  assign n2457 = pi21 ? n32 : n65;
  assign n2458 = pi20 ? n32 : n2457;
  assign n2459 = pi19 ? n32 : n2458;
  assign n2460 = pi18 ? n2459 : n37;
  assign n2461 = pi17 ? n32 : n2460;
  assign n2462 = pi16 ? n2461 : n1632;
  assign n2463 = pi15 ? n2462 : n1648;
  assign n2464 = pi16 ? n154 : n1645;
  assign n2465 = pi16 ? n186 : n1645;
  assign n2466 = pi15 ? n2464 : n2465;
  assign n2467 = pi14 ? n2463 : n2466;
  assign n2468 = pi23 ? n1149 : n32;
  assign n2469 = pi22 ? n2468 : n32;
  assign n2470 = pi21 ? n2469 : n32;
  assign n2471 = pi20 ? n2470 : n32;
  assign n2472 = pi19 ? n2471 : n32;
  assign n2473 = pi18 ? n1652 : n2472;
  assign n2474 = pi17 ? n163 : n2473;
  assign n2475 = pi16 ? n1148 : n2474;
  assign n2476 = pi18 ? n1660 : n2472;
  assign n2477 = pi17 ? n163 : n2476;
  assign n2478 = pi16 ? n721 : n2477;
  assign n2479 = pi15 ? n2475 : n2478;
  assign n2480 = pi18 ? n1667 : n2472;
  assign n2481 = pi17 ? n99 : n2480;
  assign n2482 = pi16 ? n801 : n2481;
  assign n2483 = pi22 ? n715 : n37;
  assign n2484 = pi21 ? n2483 : n99;
  assign n2485 = pi20 ? n32 : n2484;
  assign n2486 = pi19 ? n32 : n2485;
  assign n2487 = pi18 ? n2486 : n99;
  assign n2488 = pi17 ? n32 : n2487;
  assign n2489 = pi18 ? n99 : n2472;
  assign n2490 = pi17 ? n99 : n2489;
  assign n2491 = pi16 ? n2488 : n2490;
  assign n2492 = pi15 ? n2482 : n2491;
  assign n2493 = pi14 ? n2479 : n2492;
  assign n2494 = pi13 ? n2467 : n2493;
  assign n2495 = pi12 ? n2456 : n2494;
  assign n2496 = pi16 ? n721 : n2490;
  assign n2497 = pi22 ? n1519 : n295;
  assign n2498 = pi21 ? n2497 : n139;
  assign n2499 = pi20 ? n32 : n2498;
  assign n2500 = pi19 ? n32 : n2499;
  assign n2501 = pi18 ? n2500 : n139;
  assign n2502 = pi17 ? n32 : n2501;
  assign n2503 = pi18 ? n139 : n2472;
  assign n2504 = pi17 ? n139 : n2503;
  assign n2505 = pi16 ? n2502 : n2504;
  assign n2506 = pi15 ? n2496 : n2505;
  assign n2507 = pi21 ? n2497 : n1211;
  assign n2508 = pi20 ? n32 : n2507;
  assign n2509 = pi19 ? n32 : n2508;
  assign n2510 = pi21 ? n1531 : n1711;
  assign n2511 = pi20 ? n1719 : n2510;
  assign n2512 = pi21 ? n139 : n1721;
  assign n2513 = pi21 ? n1211 : n1531;
  assign n2514 = pi20 ? n2512 : n2513;
  assign n2515 = pi19 ? n2511 : n2514;
  assign n2516 = pi18 ? n2509 : n2515;
  assign n2517 = pi17 ? n32 : n2516;
  assign n2518 = pi21 ? n1711 : n139;
  assign n2519 = pi21 ? n1721 : n1211;
  assign n2520 = pi20 ? n2518 : n2519;
  assign n2521 = pi21 ? n139 : n1211;
  assign n2522 = pi20 ? n2521 : n1719;
  assign n2523 = pi19 ? n2520 : n2522;
  assign n2524 = pi20 ? n1719 : n2521;
  assign n2525 = pi19 ? n2524 : n1719;
  assign n2526 = pi18 ? n2523 : n2525;
  assign n2527 = pi21 ? n1711 : n1531;
  assign n2528 = pi20 ? n2518 : n2527;
  assign n2529 = pi19 ? n1720 : n2528;
  assign n2530 = pi23 ? n842 : n32;
  assign n2531 = pi22 ? n2530 : n32;
  assign n2532 = pi21 ? n2531 : n32;
  assign n2533 = pi20 ? n2532 : n32;
  assign n2534 = pi19 ? n2533 : n32;
  assign n2535 = pi18 ? n2529 : n2534;
  assign n2536 = pi17 ? n2526 : n2535;
  assign n2537 = pi16 ? n2517 : n2536;
  assign n2538 = pi18 ? n1214 : n2515;
  assign n2539 = pi17 ? n32 : n2538;
  assign n2540 = pi20 ? n1719 : n1715;
  assign n2541 = pi19 ? n2540 : n1719;
  assign n2542 = pi18 ? n2523 : n2541;
  assign n2543 = pi21 ? n1529 : n139;
  assign n2544 = pi20 ? n2543 : n2527;
  assign n2545 = pi19 ? n1720 : n2544;
  assign n2546 = pi18 ? n2545 : n2534;
  assign n2547 = pi17 ? n2542 : n2546;
  assign n2548 = pi16 ? n2539 : n2547;
  assign n2549 = pi15 ? n2537 : n2548;
  assign n2550 = pi14 ? n2506 : n2549;
  assign n2551 = pi20 ? n139 : n2365;
  assign n2552 = pi19 ? n1776 : n2551;
  assign n2553 = pi22 ? n532 : n32;
  assign n2554 = pi21 ? n2553 : n32;
  assign n2555 = pi20 ? n2554 : n32;
  assign n2556 = pi19 ? n2555 : n32;
  assign n2557 = pi18 ? n2552 : n2556;
  assign n2558 = pi17 ? n139 : n2557;
  assign n2559 = pi16 ? n1773 : n2558;
  assign n2560 = pi18 ? n139 : n2556;
  assign n2561 = pi17 ? n139 : n2560;
  assign n2562 = pi16 ? n331 : n2561;
  assign n2563 = pi15 ? n2559 : n2562;
  assign n2564 = pi23 ? n204 : n32;
  assign n2565 = pi22 ? n2564 : n32;
  assign n2566 = pi21 ? n2565 : n32;
  assign n2567 = pi20 ? n2566 : n32;
  assign n2568 = pi19 ? n2567 : n32;
  assign n2569 = pi18 ? n1796 : n2568;
  assign n2570 = pi17 ? n139 : n2569;
  assign n2571 = pi16 ? n331 : n2570;
  assign n2572 = pi18 ? n1813 : n2568;
  assign n2573 = pi17 ? n1808 : n2572;
  assign n2574 = pi16 ? n1803 : n2573;
  assign n2575 = pi15 ? n2571 : n2574;
  assign n2576 = pi14 ? n2563 : n2575;
  assign n2577 = pi13 ? n2550 : n2576;
  assign n2578 = pi22 ? n664 : n32;
  assign n2579 = pi21 ? n2578 : n32;
  assign n2580 = pi20 ? n2579 : n32;
  assign n2581 = pi19 ? n2580 : n32;
  assign n2582 = pi18 ? n1821 : n2581;
  assign n2583 = pi17 ? n139 : n2582;
  assign n2584 = pi16 ? n331 : n2583;
  assign n2585 = pi22 ? n295 : n456;
  assign n2586 = pi21 ? n2585 : n506;
  assign n2587 = pi21 ? n2585 : n1696;
  assign n2588 = pi20 ? n2586 : n2587;
  assign n2589 = pi22 ? n455 : n295;
  assign n2590 = pi21 ? n2589 : n499;
  assign n2591 = pi21 ? n1828 : n2585;
  assign n2592 = pi20 ? n2590 : n2591;
  assign n2593 = pi19 ? n2588 : n2592;
  assign n2594 = pi18 ? n1831 : n2593;
  assign n2595 = pi17 ? n32 : n2594;
  assign n2596 = pi21 ? n1696 : n2589;
  assign n2597 = pi21 ? n499 : n1828;
  assign n2598 = pi20 ? n2596 : n2597;
  assign n2599 = pi21 ? n295 : n1828;
  assign n2600 = pi20 ? n2599 : n2587;
  assign n2601 = pi19 ? n2598 : n2600;
  assign n2602 = pi21 ? n820 : n1828;
  assign n2603 = pi20 ? n2587 : n2602;
  assign n2604 = pi21 ? n1810 : n1696;
  assign n2605 = pi20 ? n2587 : n2604;
  assign n2606 = pi19 ? n2603 : n2605;
  assign n2607 = pi18 ? n2601 : n2606;
  assign n2608 = pi21 ? n1696 : n1860;
  assign n2609 = pi21 ? n1696 : n522;
  assign n2610 = pi20 ? n2608 : n2609;
  assign n2611 = pi19 ? n1859 : n2610;
  assign n2612 = pi18 ? n2611 : n2581;
  assign n2613 = pi17 ? n2607 : n2612;
  assign n2614 = pi16 ? n2595 : n2613;
  assign n2615 = pi15 ? n2584 : n2614;
  assign n2616 = pi21 ? n1313 : n506;
  assign n2617 = pi20 ? n2616 : n1321;
  assign n2618 = pi20 ? n1311 : n1314;
  assign n2619 = pi19 ? n2617 : n2618;
  assign n2620 = pi18 ? n1872 : n2619;
  assign n2621 = pi17 ? n32 : n2620;
  assign n2622 = pi20 ? n1315 : n1320;
  assign n2623 = pi21 ? n584 : n506;
  assign n2624 = pi21 ? n1313 : n580;
  assign n2625 = pi20 ? n2623 : n2624;
  assign n2626 = pi19 ? n2622 : n2625;
  assign n2627 = pi21 ? n570 : n506;
  assign n2628 = pi20 ? n2624 : n2627;
  assign n2629 = pi21 ? n1887 : n37;
  assign n2630 = pi20 ? n1321 : n2629;
  assign n2631 = pi19 ? n2628 : n2630;
  assign n2632 = pi18 ? n2626 : n2631;
  assign n2633 = pi21 ? n37 : n1895;
  assign n2634 = pi21 ? n37 : n457;
  assign n2635 = pi20 ? n2633 : n2634;
  assign n2636 = pi19 ? n1894 : n2635;
  assign n2637 = pi22 ? n1407 : n32;
  assign n2638 = pi21 ? n2637 : n32;
  assign n2639 = pi20 ? n2638 : n32;
  assign n2640 = pi19 ? n2639 : n32;
  assign n2641 = pi18 ? n2636 : n2640;
  assign n2642 = pi17 ? n2632 : n2641;
  assign n2643 = pi16 ? n2621 : n2642;
  assign n2644 = pi21 ? n37 : n1313;
  assign n2645 = pi20 ? n1912 : n2644;
  assign n2646 = pi19 ? n1919 : n2645;
  assign n2647 = pi18 ? n2646 : n2640;
  assign n2648 = pi17 ? n1918 : n2647;
  assign n2649 = pi16 ? n1910 : n2648;
  assign n2650 = pi15 ? n2643 : n2649;
  assign n2651 = pi14 ? n2615 : n2650;
  assign n2652 = pi19 ? n1953 : n1954;
  assign n2653 = pi21 ? n928 : n32;
  assign n2654 = pi20 ? n2653 : n32;
  assign n2655 = pi19 ? n2654 : n32;
  assign n2656 = pi18 ? n2652 : n2655;
  assign n2657 = pi17 ? n1948 : n2656;
  assign n2658 = pi16 ? n1934 : n2657;
  assign n2659 = pi19 ? n1989 : n1990;
  assign n2660 = pi18 ? n2659 : n2655;
  assign n2661 = pi17 ? n1987 : n2660;
  assign n2662 = pi16 ? n1973 : n2661;
  assign n2663 = pi15 ? n2658 : n2662;
  assign n2664 = pi21 ? n1943 : n2074;
  assign n2665 = pi20 ? n2025 : n2664;
  assign n2666 = pi19 ? n2024 : n2665;
  assign n2667 = pi18 ? n2666 : n32;
  assign n2668 = pi17 ? n2022 : n2667;
  assign n2669 = pi16 ? n2013 : n2668;
  assign n2670 = pi18 ? n335 : n32;
  assign n2671 = pi17 ? n335 : n2670;
  assign n2672 = pi16 ? n2035 : n2671;
  assign n2673 = pi15 ? n2669 : n2672;
  assign n2674 = pi14 ? n2663 : n2673;
  assign n2675 = pi13 ? n2651 : n2674;
  assign n2676 = pi12 ? n2577 : n2675;
  assign n2677 = pi11 ? n2495 : n2676;
  assign n2678 = pi22 ? n625 : n32;
  assign n2679 = pi21 ? n2678 : n32;
  assign n2680 = pi20 ? n2679 : n32;
  assign n2681 = pi19 ? n2680 : n32;
  assign n2682 = pi18 ? n2064 : n2681;
  assign n2683 = pi17 ? n2058 : n2682;
  assign n2684 = pi16 ? n2053 : n2683;
  assign n2685 = pi18 ? n2077 : n2681;
  assign n2686 = pi17 ? n2072 : n2685;
  assign n2687 = pi16 ? n439 : n2686;
  assign n2688 = pi15 ? n2684 : n2687;
  assign n2689 = pi18 ? n2087 : n2681;
  assign n2690 = pi17 ? n2083 : n2689;
  assign n2691 = pi16 ? n439 : n2690;
  assign n2692 = pi18 ? n2096 : n2681;
  assign n2693 = pi17 ? n37 : n2692;
  assign n2694 = pi16 ? n439 : n2693;
  assign n2695 = pi15 ? n2691 : n2694;
  assign n2696 = pi14 ? n2688 : n2695;
  assign n2697 = pi18 ? n2102 : n2681;
  assign n2698 = pi17 ? n37 : n2697;
  assign n2699 = pi16 ? n439 : n2698;
  assign n2700 = pi22 ? n688 : n32;
  assign n2701 = pi21 ? n2700 : n32;
  assign n2702 = pi20 ? n2701 : n32;
  assign n2703 = pi19 ? n2702 : n32;
  assign n2704 = pi18 ? n2109 : n2703;
  assign n2705 = pi17 ? n37 : n2704;
  assign n2706 = pi16 ? n439 : n2705;
  assign n2707 = pi22 ? n363 : n233;
  assign n2708 = pi21 ? n37 : n2707;
  assign n2709 = pi20 ? n37 : n2708;
  assign n2710 = pi19 ? n2119 : n2709;
  assign n2711 = pi18 ? n2710 : n1824;
  assign n2712 = pi17 ? n2115 : n2711;
  assign n2713 = pi16 ? n439 : n2712;
  assign n2714 = pi15 ? n2706 : n2713;
  assign n2715 = pi14 ? n2699 : n2714;
  assign n2716 = pi13 ? n2696 : n2715;
  assign n2717 = pi19 ? n37 : n2709;
  assign n2718 = pi18 ? n2717 : n32;
  assign n2719 = pi17 ? n37 : n2718;
  assign n2720 = pi16 ? n439 : n2719;
  assign n2721 = pi22 ? n363 : n685;
  assign n2722 = pi21 ? n37 : n2721;
  assign n2723 = pi20 ? n37 : n2722;
  assign n2724 = pi19 ? n37 : n2723;
  assign n2725 = pi18 ? n2724 : n32;
  assign n2726 = pi17 ? n37 : n2725;
  assign n2727 = pi16 ? n439 : n2726;
  assign n2728 = pi15 ? n2720 : n2727;
  assign n2729 = pi21 ? n37 : n685;
  assign n2730 = pi20 ? n37 : n2729;
  assign n2731 = pi19 ? n37 : n2730;
  assign n2732 = pi18 ? n2731 : n32;
  assign n2733 = pi17 ? n37 : n2732;
  assign n2734 = pi16 ? n439 : n2733;
  assign n2735 = pi15 ? n2727 : n2734;
  assign n2736 = pi14 ? n2728 : n2735;
  assign n2737 = pi21 ? n716 : n2162;
  assign n2738 = pi20 ? n32 : n2737;
  assign n2739 = pi19 ? n32 : n2738;
  assign n2740 = pi21 ? n99 : n2162;
  assign n2741 = pi20 ? n2740 : n2165;
  assign n2742 = pi20 ? n2167 : n2174;
  assign n2743 = pi19 ? n2741 : n2742;
  assign n2744 = pi18 ? n2739 : n2743;
  assign n2745 = pi17 ? n32 : n2744;
  assign n2746 = pi22 ? n99 : n2160;
  assign n2747 = pi21 ? n2161 : n2746;
  assign n2748 = pi20 ? n2174 : n2747;
  assign n2749 = pi21 ? n99 : n2161;
  assign n2750 = pi20 ? n2749 : n2161;
  assign n2751 = pi19 ? n2748 : n2750;
  assign n2752 = pi21 ? n2161 : n1143;
  assign n2753 = pi21 ? n2162 : n2746;
  assign n2754 = pi20 ? n2752 : n2753;
  assign n2755 = pi21 ? n2164 : n2160;
  assign n2756 = pi20 ? n2749 : n2755;
  assign n2757 = pi19 ? n2754 : n2756;
  assign n2758 = pi18 ? n2751 : n2757;
  assign n2759 = pi22 ? n363 : n1475;
  assign n2760 = pi21 ? n99 : n2759;
  assign n2761 = pi20 ? n2191 : n2760;
  assign n2762 = pi19 ? n2190 : n2761;
  assign n2763 = pi18 ? n2762 : n32;
  assign n2764 = pi17 ? n2758 : n2763;
  assign n2765 = pi16 ? n2745 : n2764;
  assign n2766 = pi24 ? n685 : n316;
  assign n2767 = pi23 ? n685 : n2766;
  assign n2768 = pi22 ? n685 : n2767;
  assign n2769 = pi21 ? n99 : n2768;
  assign n2770 = pi20 ? n99 : n2769;
  assign n2771 = pi19 ? n99 : n2770;
  assign n2772 = pi18 ? n2771 : n32;
  assign n2773 = pi17 ? n99 : n2772;
  assign n2774 = pi16 ? n721 : n2773;
  assign n2775 = pi15 ? n2765 : n2774;
  assign n2776 = pi21 ? n99 : n2147;
  assign n2777 = pi20 ? n99 : n2776;
  assign n2778 = pi19 ? n99 : n2777;
  assign n2779 = pi18 ? n2778 : n32;
  assign n2780 = pi17 ? n99 : n2779;
  assign n2781 = pi16 ? n744 : n2780;
  assign n2782 = pi21 ? n685 : n2200;
  assign n2783 = pi20 ? n99 : n2782;
  assign n2784 = pi19 ? n99 : n2783;
  assign n2785 = pi18 ? n2784 : n32;
  assign n2786 = pi17 ? n99 : n2785;
  assign n2787 = pi16 ? n744 : n2786;
  assign n2788 = pi15 ? n2781 : n2787;
  assign n2789 = pi14 ? n2775 : n2788;
  assign n2790 = pi13 ? n2736 : n2789;
  assign n2791 = pi12 ? n2716 : n2790;
  assign n2792 = pi21 ? n767 : n2200;
  assign n2793 = pi20 ? n99 : n2792;
  assign n2794 = pi19 ? n99 : n2793;
  assign n2795 = pi18 ? n2794 : n32;
  assign n2796 = pi17 ? n99 : n2795;
  assign n2797 = pi16 ? n721 : n2796;
  assign n2798 = pi16 ? n1510 : n2235;
  assign n2799 = pi15 ? n2797 : n2798;
  assign n2800 = pi14 ? n2799 : n2263;
  assign n2801 = pi16 ? n744 : n2271;
  assign n2802 = pi15 ? n2801 : n2288;
  assign n2803 = pi21 ? n346 : n1485;
  assign n2804 = pi20 ? n157 : n2803;
  assign n2805 = pi19 ? n2298 : n2804;
  assign n2806 = pi18 ? n2805 : n32;
  assign n2807 = pi17 ? n2297 : n2806;
  assign n2808 = pi16 ? n915 : n2807;
  assign n2809 = pi18 ? n913 : n2308;
  assign n2810 = pi17 ? n32 : n2809;
  assign n2811 = pi16 ? n2810 : n2325;
  assign n2812 = pi15 ? n2808 : n2811;
  assign n2813 = pi14 ? n2802 : n2812;
  assign n2814 = pi13 ? n2800 : n2813;
  assign n2815 = pi22 ? n1263 : n32;
  assign n2816 = pi21 ? n316 : n2815;
  assign n2817 = pi20 ? n139 : n2816;
  assign n2818 = pi19 ? n1017 : n2817;
  assign n2819 = pi18 ? n2818 : n32;
  assign n2820 = pi17 ? n139 : n2819;
  assign n2821 = pi16 ? n2291 : n2820;
  assign n2822 = pi18 ? n966 : n2336;
  assign n2823 = pi17 ? n32 : n2822;
  assign n2824 = pi20 ? n975 : n2816;
  assign n2825 = pi19 ? n1787 : n2824;
  assign n2826 = pi18 ? n2825 : n32;
  assign n2827 = pi17 ? n139 : n2826;
  assign n2828 = pi16 ? n2823 : n2827;
  assign n2829 = pi15 ? n2821 : n2828;
  assign n2830 = pi21 ? n139 : n1711;
  assign n2831 = pi20 ? n2830 : n139;
  assign n2832 = pi19 ? n139 : n2831;
  assign n2833 = pi18 ? n2832 : n139;
  assign n2834 = pi23 ? n316 : n687;
  assign n2835 = pi22 ? n2834 : n32;
  assign n2836 = pi21 ? n316 : n2835;
  assign n2837 = pi20 ? n975 : n2836;
  assign n2838 = pi19 ? n139 : n2837;
  assign n2839 = pi18 ? n2838 : n32;
  assign n2840 = pi17 ? n2833 : n2839;
  assign n2841 = pi16 ? n2291 : n2840;
  assign n2842 = pi18 ? n2832 : n2350;
  assign n2843 = pi21 ? n346 : n2835;
  assign n2844 = pi20 ? n2353 : n2843;
  assign n2845 = pi19 ? n2352 : n2844;
  assign n2846 = pi18 ? n2845 : n32;
  assign n2847 = pi17 ? n2842 : n2846;
  assign n2848 = pi16 ? n2291 : n2847;
  assign n2849 = pi15 ? n2841 : n2848;
  assign n2850 = pi14 ? n2829 : n2849;
  assign n2851 = pi20 ? n820 : n1719;
  assign n2852 = pi19 ? n139 : n2851;
  assign n2853 = pi18 ? n2852 : n2376;
  assign n2854 = pi17 ? n2853 : n2380;
  assign n2855 = pi16 ? n2369 : n2854;
  assign n2856 = pi22 ? n909 : n918;
  assign n2857 = pi21 ? n2856 : n139;
  assign n2858 = pi20 ? n32 : n2857;
  assign n2859 = pi19 ? n32 : n2858;
  assign n2860 = pi18 ? n2859 : n139;
  assign n2861 = pi17 ? n32 : n2860;
  assign n2862 = pi20 ? n139 : n921;
  assign n2863 = pi22 ? n918 : n139;
  assign n2864 = pi22 ? n918 : n1038;
  assign n2865 = pi21 ? n2863 : n2864;
  assign n2866 = pi21 ? n2863 : n919;
  assign n2867 = pi20 ? n2865 : n2866;
  assign n2868 = pi19 ? n2862 : n2867;
  assign n2869 = pi22 ? n1038 : n139;
  assign n2870 = pi21 ? n919 : n2869;
  assign n2871 = pi20 ? n2870 : n1794;
  assign n2872 = pi21 ? n139 : n2869;
  assign n2873 = pi20 ? n2872 : n1794;
  assign n2874 = pi19 ? n2871 : n2873;
  assign n2875 = pi18 ? n2868 : n2874;
  assign n2876 = pi22 ? n918 : n204;
  assign n2877 = pi21 ? n2864 : n2876;
  assign n2878 = pi20 ? n2877 : n2383;
  assign n2879 = pi19 ? n2878 : n2378;
  assign n2880 = pi18 ? n2879 : n32;
  assign n2881 = pi17 ? n2875 : n2880;
  assign n2882 = pi16 ? n2861 : n2881;
  assign n2883 = pi15 ? n2855 : n2882;
  assign n2884 = pi21 ? n522 : n204;
  assign n2885 = pi20 ? n2884 : n204;
  assign n2886 = pi19 ? n204 : n2885;
  assign n2887 = pi18 ? n2886 : n2407;
  assign n2888 = pi20 ? n204 : n1027;
  assign n2889 = pi21 ? n1027 : n2700;
  assign n2890 = pi20 ? n2413 : n2889;
  assign n2891 = pi19 ? n2888 : n2890;
  assign n2892 = pi18 ? n2891 : n32;
  assign n2893 = pi17 ? n2887 : n2892;
  assign n2894 = pi16 ? n2400 : n2893;
  assign n2895 = pi23 ? n714 : n204;
  assign n2896 = pi22 ? n2895 : n450;
  assign n2897 = pi21 ? n2896 : n448;
  assign n2898 = pi20 ? n32 : n2897;
  assign n2899 = pi19 ? n32 : n2898;
  assign n2900 = pi21 ? n1949 : n1940;
  assign n2901 = pi21 ? n1079 : n458;
  assign n2902 = pi20 ? n2900 : n2901;
  assign n2903 = pi22 ? n450 : n448;
  assign n2904 = pi21 ? n2903 : n458;
  assign n2905 = pi21 ? n474 : n476;
  assign n2906 = pi20 ? n2904 : n2905;
  assign n2907 = pi19 ? n2902 : n2906;
  assign n2908 = pi18 ? n2899 : n2907;
  assign n2909 = pi17 ? n32 : n2908;
  assign n2910 = pi21 ? n1940 : n2903;
  assign n2911 = pi20 ? n2910 : n474;
  assign n2912 = pi21 ? n2903 : n1949;
  assign n2913 = pi21 ? n1949 : n458;
  assign n2914 = pi20 ? n2912 : n2913;
  assign n2915 = pi19 ? n2911 : n2914;
  assign n2916 = pi21 ? n458 : n1083;
  assign n2917 = pi21 ? n2903 : n1079;
  assign n2918 = pi20 ? n2916 : n2917;
  assign n2919 = pi18 ? n2915 : n2918;
  assign n2920 = pi20 ? n1949 : n204;
  assign n2921 = pi19 ? n2920 : n2430;
  assign n2922 = pi18 ? n2921 : n32;
  assign n2923 = pi17 ? n2919 : n2922;
  assign n2924 = pi16 ? n2909 : n2923;
  assign n2925 = pi15 ? n2894 : n2924;
  assign n2926 = pi14 ? n2883 : n2925;
  assign n2927 = pi13 ? n2850 : n2926;
  assign n2928 = pi12 ? n2814 : n2927;
  assign n2929 = pi11 ? n2791 : n2928;
  assign n2930 = pi10 ? n2677 : n2929;
  assign n2931 = pi09 ? n32 : n2930;
  assign n2932 = pi08 ? n2441 : n2931;
  assign n2933 = pi22 ? n47 : n32;
  assign n2934 = pi21 ? n2933 : n32;
  assign n2935 = pi20 ? n2934 : n32;
  assign n2936 = pi19 ? n2935 : n32;
  assign n2937 = pi18 ? n37 : n2936;
  assign n2938 = pi17 ? n37 : n2937;
  assign n2939 = pi16 ? n61 : n2938;
  assign n2940 = pi16 ? n2447 : n2938;
  assign n2941 = pi15 ? n2939 : n2940;
  assign n2942 = pi14 ? n32 : n2941;
  assign n2943 = pi16 ? n70 : n2938;
  assign n2944 = pi16 ? n73 : n2938;
  assign n2945 = pi15 ? n2943 : n2944;
  assign n2946 = pi22 ? n84 : n32;
  assign n2947 = pi21 ? n2946 : n32;
  assign n2948 = pi20 ? n2947 : n32;
  assign n2949 = pi19 ? n2948 : n32;
  assign n2950 = pi18 ? n37 : n2949;
  assign n2951 = pi17 ? n37 : n2950;
  assign n2952 = pi16 ? n83 : n2951;
  assign n2953 = pi16 ? n1130 : n2951;
  assign n2954 = pi15 ? n2952 : n2953;
  assign n2955 = pi14 ? n2945 : n2954;
  assign n2956 = pi13 ? n2942 : n2955;
  assign n2957 = pi22 ? n37 : n112;
  assign n2958 = pi21 ? n2957 : n2175;
  assign n2959 = pi21 ? n2168 : n2175;
  assign n2960 = pi20 ? n2958 : n2959;
  assign n2961 = pi21 ? n2161 : n2156;
  assign n2962 = pi21 ? n2160 : n2164;
  assign n2963 = pi20 ? n2961 : n2962;
  assign n2964 = pi19 ? n2960 : n2963;
  assign n2965 = pi18 ? n2459 : n2964;
  assign n2966 = pi17 ? n32 : n2965;
  assign n2967 = pi21 ? n2175 : n2161;
  assign n2968 = pi21 ? n2156 : n2160;
  assign n2969 = pi20 ? n2967 : n2968;
  assign n2970 = pi21 ? n2957 : n37;
  assign n2971 = pi20 ? n2185 : n2970;
  assign n2972 = pi19 ? n2969 : n2971;
  assign n2973 = pi21 ? n181 : n37;
  assign n2974 = pi21 ? n37 : n2175;
  assign n2975 = pi20 ? n2973 : n2974;
  assign n2976 = pi21 ? n2161 : n37;
  assign n2977 = pi20 ? n2970 : n2976;
  assign n2978 = pi19 ? n2975 : n2977;
  assign n2979 = pi18 ? n2972 : n2978;
  assign n2980 = pi20 ? n2976 : n37;
  assign n2981 = pi22 ? n2160 : n37;
  assign n2982 = pi21 ? n37 : n2981;
  assign n2983 = pi21 ? n37 : n2161;
  assign n2984 = pi20 ? n2982 : n2983;
  assign n2985 = pi19 ? n2980 : n2984;
  assign n2986 = pi18 ? n2985 : n2949;
  assign n2987 = pi17 ? n2979 : n2986;
  assign n2988 = pi16 ? n2966 : n2987;
  assign n2989 = pi22 ? n119 : n32;
  assign n2990 = pi21 ? n2989 : n32;
  assign n2991 = pi20 ? n2990 : n32;
  assign n2992 = pi19 ? n2991 : n32;
  assign n2993 = pi18 ? n99 : n2992;
  assign n2994 = pi17 ? n99 : n2993;
  assign n2995 = pi16 ? n132 : n2994;
  assign n2996 = pi15 ? n2988 : n2995;
  assign n2997 = pi16 ? n1148 : n2994;
  assign n2998 = pi22 ? n164 : n99;
  assign n2999 = pi21 ? n2998 : n99;
  assign n3000 = pi20 ? n1492 : n2999;
  assign n3001 = pi19 ? n99 : n3000;
  assign n3002 = pi22 ? n164 : n157;
  assign n3003 = pi21 ? n3002 : n99;
  assign n3004 = pi21 ? n3002 : n168;
  assign n3005 = pi20 ? n3003 : n3004;
  assign n3006 = pi21 ? n777 : n168;
  assign n3007 = pi20 ? n99 : n3006;
  assign n3008 = pi19 ? n3005 : n3007;
  assign n3009 = pi18 ? n3001 : n3008;
  assign n3010 = pi22 ? n158 : n164;
  assign n3011 = pi21 ? n3002 : n3010;
  assign n3012 = pi20 ? n3006 : n3011;
  assign n3013 = pi22 ? n157 : n158;
  assign n3014 = pi21 ? n3013 : n99;
  assign n3015 = pi19 ? n3012 : n3014;
  assign n3016 = pi18 ? n3015 : n2992;
  assign n3017 = pi17 ? n3009 : n3016;
  assign n3018 = pi16 ? n186 : n3017;
  assign n3019 = pi15 ? n2997 : n3018;
  assign n3020 = pi14 ? n2996 : n3019;
  assign n3021 = pi16 ? n744 : n2994;
  assign n3022 = pi22 ? n140 : n32;
  assign n3023 = pi21 ? n3022 : n32;
  assign n3024 = pi20 ? n3023 : n32;
  assign n3025 = pi19 ? n3024 : n32;
  assign n3026 = pi18 ? n99 : n3025;
  assign n3027 = pi17 ? n99 : n3026;
  assign n3028 = pi16 ? n744 : n3027;
  assign n3029 = pi21 ? n180 : n218;
  assign n3030 = pi20 ? n32 : n3029;
  assign n3031 = pi19 ? n32 : n3030;
  assign n3032 = pi21 ? n2156 : n181;
  assign n3033 = pi21 ? n218 : n2156;
  assign n3034 = pi20 ? n2970 : n3033;
  assign n3035 = pi19 ? n3032 : n3034;
  assign n3036 = pi18 ? n3031 : n3035;
  assign n3037 = pi17 ? n32 : n3036;
  assign n3038 = pi21 ? n181 : n2957;
  assign n3039 = pi21 ? n37 : n218;
  assign n3040 = pi20 ? n3038 : n3039;
  assign n3041 = pi21 ? n2156 : n218;
  assign n3042 = pi21 ? n2156 : n99;
  assign n3043 = pi20 ? n3041 : n3042;
  assign n3044 = pi19 ? n3040 : n3043;
  assign n3045 = pi20 ? n3042 : n218;
  assign n3046 = pi21 ? n218 : n181;
  assign n3047 = pi20 ? n3032 : n3046;
  assign n3048 = pi19 ? n3045 : n3047;
  assign n3049 = pi18 ? n3044 : n3048;
  assign n3050 = pi20 ? n219 : n99;
  assign n3051 = pi20 ? n181 : n2973;
  assign n3052 = pi19 ? n3050 : n3051;
  assign n3053 = pi18 ? n3052 : n3025;
  assign n3054 = pi17 ? n3049 : n3053;
  assign n3055 = pi16 ? n3037 : n3054;
  assign n3056 = pi15 ? n3028 : n3055;
  assign n3057 = pi14 ? n3021 : n3056;
  assign n3058 = pi13 ? n3020 : n3057;
  assign n3059 = pi12 ? n2956 : n3058;
  assign n3060 = pi22 ? n55 : n112;
  assign n3061 = pi21 ? n3060 : n99;
  assign n3062 = pi20 ? n32 : n3061;
  assign n3063 = pi19 ? n32 : n3062;
  assign n3064 = pi18 ? n3063 : n99;
  assign n3065 = pi17 ? n32 : n3064;
  assign n3066 = pi22 ? n1344 : n32;
  assign n3067 = pi21 ? n3066 : n32;
  assign n3068 = pi20 ? n3067 : n32;
  assign n3069 = pi19 ? n3068 : n32;
  assign n3070 = pi18 ? n99 : n3069;
  assign n3071 = pi17 ? n99 : n3070;
  assign n3072 = pi16 ? n3065 : n3071;
  assign n3073 = pi22 ? n37 : n295;
  assign n3074 = pi21 ? n3073 : n297;
  assign n3075 = pi21 ? n3073 : n37;
  assign n3076 = pi20 ? n3074 : n3075;
  assign n3077 = pi21 ? n820 : n375;
  assign n3078 = pi21 ? n297 : n3073;
  assign n3079 = pi20 ? n3077 : n3078;
  assign n3080 = pi19 ? n3076 : n3079;
  assign n3081 = pi18 ? n1692 : n3080;
  assign n3082 = pi17 ? n32 : n3081;
  assign n3083 = pi21 ? n37 : n820;
  assign n3084 = pi21 ? n375 : n297;
  assign n3085 = pi20 ? n3083 : n3084;
  assign n3086 = pi21 ? n37 : n297;
  assign n3087 = pi21 ? n3073 : n139;
  assign n3088 = pi20 ? n3086 : n3087;
  assign n3089 = pi19 ? n3085 : n3088;
  assign n3090 = pi21 ? n820 : n297;
  assign n3091 = pi20 ? n3087 : n3090;
  assign n3092 = pi21 ? n1531 : n297;
  assign n3093 = pi20 ? n3074 : n3092;
  assign n3094 = pi19 ? n3091 : n3093;
  assign n3095 = pi18 ? n3089 : n3094;
  assign n3096 = pi21 ? n37 : n139;
  assign n3097 = pi20 ? n3096 : n3083;
  assign n3098 = pi19 ? n1720 : n3097;
  assign n3099 = pi18 ? n3098 : n3069;
  assign n3100 = pi17 ? n3095 : n3099;
  assign n3101 = pi16 ? n3082 : n3100;
  assign n3102 = pi15 ? n3072 : n3101;
  assign n3103 = pi20 ? n3086 : n37;
  assign n3104 = pi21 ? n820 : n37;
  assign n3105 = pi20 ? n3104 : n1003;
  assign n3106 = pi19 ? n3103 : n3105;
  assign n3107 = pi18 ? n1692 : n3106;
  assign n3108 = pi17 ? n32 : n3107;
  assign n3109 = pi20 ? n3083 : n3086;
  assign n3110 = pi20 ? n3086 : n3096;
  assign n3111 = pi19 ? n3109 : n3110;
  assign n3112 = pi21 ? n390 : n297;
  assign n3113 = pi20 ? n3096 : n3112;
  assign n3114 = pi20 ? n3086 : n3090;
  assign n3115 = pi19 ? n3113 : n3114;
  assign n3116 = pi18 ? n3111 : n3115;
  assign n3117 = pi21 ? n820 : n356;
  assign n3118 = pi22 ? n383 : n390;
  assign n3119 = pi21 ? n424 : n3118;
  assign n3120 = pi20 ? n3117 : n3119;
  assign n3121 = pi21 ? n417 : n139;
  assign n3122 = pi20 ? n3121 : n3083;
  assign n3123 = pi19 ? n3120 : n3122;
  assign n3124 = pi23 ? n363 : n395;
  assign n3125 = pi22 ? n3124 : n32;
  assign n3126 = pi21 ? n3125 : n32;
  assign n3127 = pi20 ? n3126 : n32;
  assign n3128 = pi19 ? n3127 : n32;
  assign n3129 = pi18 ? n3123 : n3128;
  assign n3130 = pi17 ? n3116 : n3129;
  assign n3131 = pi16 ? n3108 : n3130;
  assign n3132 = pi18 ? n1567 : n139;
  assign n3133 = pi17 ? n32 : n3132;
  assign n3134 = pi24 ? n139 : n363;
  assign n3135 = pi23 ? n3134 : n32;
  assign n3136 = pi22 ? n3135 : n32;
  assign n3137 = pi21 ? n3136 : n32;
  assign n3138 = pi20 ? n3137 : n32;
  assign n3139 = pi19 ? n3138 : n32;
  assign n3140 = pi18 ? n139 : n3139;
  assign n3141 = pi17 ? n139 : n3140;
  assign n3142 = pi16 ? n3133 : n3141;
  assign n3143 = pi15 ? n3131 : n3142;
  assign n3144 = pi14 ? n3102 : n3143;
  assign n3145 = pi24 ? n139 : n157;
  assign n3146 = pi23 ? n3145 : n32;
  assign n3147 = pi22 ? n3146 : n32;
  assign n3148 = pi21 ? n3147 : n32;
  assign n3149 = pi20 ? n3148 : n32;
  assign n3150 = pi19 ? n3149 : n32;
  assign n3151 = pi18 ? n139 : n3150;
  assign n3152 = pi17 ? n139 : n3151;
  assign n3153 = pi16 ? n1773 : n3152;
  assign n3154 = pi16 ? n331 : n3152;
  assign n3155 = pi15 ? n3153 : n3154;
  assign n3156 = pi22 ? n1217 : n32;
  assign n3157 = pi21 ? n3156 : n32;
  assign n3158 = pi20 ? n3157 : n32;
  assign n3159 = pi19 ? n3158 : n32;
  assign n3160 = pi18 ? n139 : n3159;
  assign n3161 = pi17 ? n139 : n3160;
  assign n3162 = pi16 ? n331 : n3161;
  assign n3163 = pi19 ? n2345 : n139;
  assign n3164 = pi18 ? n329 : n3163;
  assign n3165 = pi17 ? n32 : n3164;
  assign n3166 = pi20 ? n350 : n1008;
  assign n3167 = pi19 ? n139 : n3166;
  assign n3168 = pi20 ? n1008 : n139;
  assign n3169 = pi19 ? n3168 : n1786;
  assign n3170 = pi18 ? n3167 : n3169;
  assign n3171 = pi20 ? n1008 : n360;
  assign n3172 = pi21 ? n139 : n349;
  assign n3173 = pi19 ? n3171 : n3172;
  assign n3174 = pi23 ? n204 : n531;
  assign n3175 = pi22 ? n3174 : n32;
  assign n3176 = pi21 ? n3175 : n32;
  assign n3177 = pi20 ? n3176 : n32;
  assign n3178 = pi19 ? n3177 : n32;
  assign n3179 = pi18 ? n3173 : n3178;
  assign n3180 = pi17 ? n3170 : n3179;
  assign n3181 = pi16 ? n3165 : n3180;
  assign n3182 = pi15 ? n3162 : n3181;
  assign n3183 = pi14 ? n3155 : n3182;
  assign n3184 = pi13 ? n3144 : n3183;
  assign n3185 = pi21 ? n296 : n1027;
  assign n3186 = pi20 ? n32 : n3185;
  assign n3187 = pi19 ? n32 : n3186;
  assign n3188 = pi22 ? n316 : n918;
  assign n3189 = pi22 ? n918 : n316;
  assign n3190 = pi21 ? n3188 : n3189;
  assign n3191 = pi22 ? n1038 : n1784;
  assign n3192 = pi21 ? n3191 : n918;
  assign n3193 = pi22 ? n316 : n1038;
  assign n3194 = pi22 ? n1784 : n918;
  assign n3195 = pi21 ? n3193 : n3194;
  assign n3196 = pi20 ? n3192 : n3195;
  assign n3197 = pi19 ? n3190 : n3196;
  assign n3198 = pi18 ? n3187 : n3197;
  assign n3199 = pi17 ? n32 : n3198;
  assign n3200 = pi21 ? n3189 : n3191;
  assign n3201 = pi21 ? n918 : n3193;
  assign n3202 = pi20 ? n3200 : n3201;
  assign n3203 = pi21 ? n2319 : n1027;
  assign n3204 = pi20 ? n3203 : n316;
  assign n3205 = pi19 ? n3202 : n3204;
  assign n3206 = pi18 ? n3205 : n316;
  assign n3207 = pi22 ? n1038 : n316;
  assign n3208 = pi21 ? n316 : n3207;
  assign n3209 = pi19 ? n316 : n3208;
  assign n3210 = pi21 ? n2320 : n32;
  assign n3211 = pi20 ? n3210 : n32;
  assign n3212 = pi19 ? n3211 : n32;
  assign n3213 = pi18 ? n3209 : n3212;
  assign n3214 = pi17 ? n3206 : n3213;
  assign n3215 = pi16 ? n3199 : n3214;
  assign n3216 = pi21 ? n296 : n346;
  assign n3217 = pi20 ? n32 : n3216;
  assign n3218 = pi19 ? n32 : n3217;
  assign n3219 = pi22 ? n295 : n383;
  assign n3220 = pi22 ? n295 : n316;
  assign n3221 = pi21 ? n3219 : n3220;
  assign n3222 = pi21 ? n3219 : n297;
  assign n3223 = pi20 ? n3221 : n3222;
  assign n3224 = pi22 ? n316 : n295;
  assign n3225 = pi21 ? n3224 : n384;
  assign n3226 = pi21 ? n346 : n3219;
  assign n3227 = pi20 ? n3225 : n3226;
  assign n3228 = pi19 ? n3223 : n3227;
  assign n3229 = pi18 ? n3218 : n3228;
  assign n3230 = pi17 ? n32 : n3229;
  assign n3231 = pi21 ? n297 : n3224;
  assign n3232 = pi21 ? n384 : n346;
  assign n3233 = pi20 ? n3231 : n3232;
  assign n3234 = pi21 ? n295 : n346;
  assign n3235 = pi21 ? n3219 : n1211;
  assign n3236 = pi20 ? n3234 : n3235;
  assign n3237 = pi19 ? n3233 : n3236;
  assign n3238 = pi21 ? n375 : n346;
  assign n3239 = pi20 ? n3235 : n3238;
  assign n3240 = pi21 ? n3219 : n1696;
  assign n3241 = pi21 ? n1777 : n1696;
  assign n3242 = pi20 ? n3240 : n3241;
  assign n3243 = pi19 ? n3239 : n3242;
  assign n3244 = pi18 ? n3237 : n3243;
  assign n3245 = pi21 ? n1529 : n1531;
  assign n3246 = pi20 ? n2370 : n3245;
  assign n3247 = pi19 ? n3246 : n3231;
  assign n3248 = pi18 ? n3247 : n3212;
  assign n3249 = pi17 ? n3244 : n3248;
  assign n3250 = pi16 ? n3230 : n3249;
  assign n3251 = pi15 ? n3215 : n3250;
  assign n3252 = pi21 ? n180 : n381;
  assign n3253 = pi20 ? n32 : n3252;
  assign n3254 = pi19 ? n32 : n3253;
  assign n3255 = pi21 ? n428 : n316;
  assign n3256 = pi21 ? n428 : n37;
  assign n3257 = pi20 ? n3255 : n3256;
  assign n3258 = pi22 ? n316 : n37;
  assign n3259 = pi21 ? n3258 : n384;
  assign n3260 = pi21 ? n381 : n428;
  assign n3261 = pi20 ? n3259 : n3260;
  assign n3262 = pi19 ? n3257 : n3261;
  assign n3263 = pi18 ? n3254 : n3262;
  assign n3264 = pi17 ? n32 : n3263;
  assign n3265 = pi21 ? n37 : n3258;
  assign n3266 = pi20 ? n3265 : n416;
  assign n3267 = pi20 ? n416 : n440;
  assign n3268 = pi19 ? n3266 : n3267;
  assign n3269 = pi20 ? n440 : n416;
  assign n3270 = pi21 ? n428 : n391;
  assign n3271 = pi21 ? n392 : n391;
  assign n3272 = pi20 ? n3270 : n3271;
  assign n3273 = pi19 ? n3269 : n3272;
  assign n3274 = pi18 ? n3268 : n3273;
  assign n3275 = pi21 ? n392 : n381;
  assign n3276 = pi20 ? n3275 : n426;
  assign n3277 = pi21 ? n37 : n392;
  assign n3278 = pi19 ? n3276 : n3277;
  assign n3279 = pi18 ? n3278 : n3212;
  assign n3280 = pi17 ? n3274 : n3279;
  assign n3281 = pi16 ? n3264 : n3280;
  assign n3282 = pi21 ? n1869 : n37;
  assign n3283 = pi20 ? n32 : n3282;
  assign n3284 = pi19 ? n32 : n3283;
  assign n3285 = pi20 ? n639 : n37;
  assign n3286 = pi19 ? n3285 : n37;
  assign n3287 = pi18 ? n3284 : n3286;
  assign n3288 = pi17 ? n32 : n3287;
  assign n3289 = pi21 ? n584 : n37;
  assign n3290 = pi20 ? n3289 : n649;
  assign n3291 = pi19 ? n37 : n3290;
  assign n3292 = pi21 ? n2007 : n37;
  assign n3293 = pi20 ? n649 : n3292;
  assign n3294 = pi19 ? n3293 : n644;
  assign n3295 = pi18 ? n3291 : n3294;
  assign n3296 = pi22 ? n204 : n583;
  assign n3297 = pi21 ? n2007 : n3296;
  assign n3298 = pi20 ? n1089 : n3297;
  assign n3299 = pi21 ? n37 : n584;
  assign n3300 = pi19 ? n3298 : n3299;
  assign n3301 = pi23 ? n204 : n624;
  assign n3302 = pi22 ? n3301 : n32;
  assign n3303 = pi21 ? n3302 : n32;
  assign n3304 = pi20 ? n3303 : n32;
  assign n3305 = pi19 ? n3304 : n32;
  assign n3306 = pi18 ? n3300 : n3305;
  assign n3307 = pi17 ? n3295 : n3306;
  assign n3308 = pi16 ? n3288 : n3307;
  assign n3309 = pi15 ? n3281 : n3308;
  assign n3310 = pi14 ? n3251 : n3309;
  assign n3311 = pi21 ? n335 : n1079;
  assign n3312 = pi20 ? n3311 : n335;
  assign n3313 = pi19 ? n3312 : n610;
  assign n3314 = pi18 ? n335 : n3313;
  assign n3315 = pi21 ? n335 : n1083;
  assign n3316 = pi20 ? n3311 : n3315;
  assign n3317 = pi19 ? n3316 : n3315;
  assign n3318 = pi23 ? n204 : n687;
  assign n3319 = pi22 ? n3318 : n32;
  assign n3320 = pi21 ? n3319 : n32;
  assign n3321 = pi20 ? n3320 : n32;
  assign n3322 = pi19 ? n3321 : n32;
  assign n3323 = pi18 ? n3317 : n3322;
  assign n3324 = pi17 ? n3314 : n3323;
  assign n3325 = pi16 ? n2035 : n3324;
  assign n3326 = pi20 ? n649 : n37;
  assign n3327 = pi19 ? n639 : n3326;
  assign n3328 = pi18 ? n374 : n3327;
  assign n3329 = pi17 ? n32 : n3328;
  assign n3330 = pi20 ? n642 : n638;
  assign n3331 = pi19 ? n3330 : n37;
  assign n3332 = pi20 ? n37 : n638;
  assign n3333 = pi19 ? n3332 : n639;
  assign n3334 = pi18 ? n3331 : n3333;
  assign n3335 = pi21 ? n570 : n569;
  assign n3336 = pi20 ? n642 : n3335;
  assign n3337 = pi19 ? n37 : n3336;
  assign n3338 = pi23 ? n233 : n395;
  assign n3339 = pi22 ? n3338 : n32;
  assign n3340 = pi21 ? n3339 : n32;
  assign n3341 = pi20 ? n3340 : n32;
  assign n3342 = pi19 ? n3341 : n32;
  assign n3343 = pi18 ? n3337 : n3342;
  assign n3344 = pi17 ? n3334 : n3343;
  assign n3345 = pi16 ? n3329 : n3344;
  assign n3346 = pi15 ? n3325 : n3345;
  assign n3347 = pi21 ? n180 : n335;
  assign n3348 = pi20 ? n32 : n3347;
  assign n3349 = pi19 ? n32 : n3348;
  assign n3350 = pi18 ? n3349 : n335;
  assign n3351 = pi17 ? n32 : n3350;
  assign n3352 = pi19 ? n611 : n335;
  assign n3353 = pi18 ? n335 : n3352;
  assign n3354 = pi19 ? n2059 : n605;
  assign n3355 = pi18 ? n3354 : n2581;
  assign n3356 = pi17 ? n3353 : n3355;
  assign n3357 = pi16 ? n3351 : n3356;
  assign n3358 = pi19 ? n37 : n3326;
  assign n3359 = pi18 ? n374 : n3358;
  assign n3360 = pi17 ? n32 : n3359;
  assign n3361 = pi19 ? n3330 : n3332;
  assign n3362 = pi19 ? n638 : n639;
  assign n3363 = pi18 ? n3361 : n3362;
  assign n3364 = pi20 ? n638 : n642;
  assign n3365 = pi19 ? n3364 : n3336;
  assign n3366 = pi18 ? n3365 : n2640;
  assign n3367 = pi17 ? n3363 : n3366;
  assign n3368 = pi16 ? n3360 : n3367;
  assign n3369 = pi15 ? n3357 : n3368;
  assign n3370 = pi14 ? n3346 : n3369;
  assign n3371 = pi13 ? n3310 : n3370;
  assign n3372 = pi12 ? n3184 : n3371;
  assign n3373 = pi11 ? n3059 : n3372;
  assign n3374 = pi20 ? n638 : n577;
  assign n3375 = pi19 ? n37 : n3374;
  assign n3376 = pi20 ? n639 : n647;
  assign n3377 = pi19 ? n3376 : n639;
  assign n3378 = pi18 ? n3375 : n3377;
  assign n3379 = pi20 ? n610 : n569;
  assign n3380 = pi19 ? n3379 : n605;
  assign n3381 = pi18 ? n3380 : n2640;
  assign n3382 = pi17 ? n3378 : n3381;
  assign n3383 = pi16 ? n439 : n3382;
  assign n3384 = pi20 ? n335 : n605;
  assign n3385 = pi19 ? n2073 : n3384;
  assign n3386 = pi18 ? n3385 : n2655;
  assign n3387 = pi17 ? n2072 : n3386;
  assign n3388 = pi16 ? n439 : n3387;
  assign n3389 = pi15 ? n3383 : n3388;
  assign n3390 = pi19 ? n37 : n577;
  assign n3391 = pi18 ? n37 : n3390;
  assign n3392 = pi22 ? n37 : n363;
  assign n3393 = pi21 ? n37 : n3392;
  assign n3394 = pi20 ? n577 : n3393;
  assign n3395 = pi19 ? n2073 : n3394;
  assign n3396 = pi23 ? n2120 : n32;
  assign n3397 = pi22 ? n3396 : n32;
  assign n3398 = pi21 ? n3397 : n32;
  assign n3399 = pi20 ? n3398 : n32;
  assign n3400 = pi19 ? n3399 : n32;
  assign n3401 = pi18 ? n3395 : n3400;
  assign n3402 = pi17 ? n3391 : n3401;
  assign n3403 = pi16 ? n439 : n3402;
  assign n3404 = pi22 ? n2116 : n37;
  assign n3405 = pi21 ? n3404 : n37;
  assign n3406 = pi20 ? n37 : n3405;
  assign n3407 = pi19 ? n37 : n3406;
  assign n3408 = pi18 ? n37 : n3407;
  assign n3409 = pi22 ? n2116 : n233;
  assign n3410 = pi21 ? n3409 : n37;
  assign n3411 = pi22 ? n233 : n559;
  assign n3412 = pi21 ? n3411 : n2091;
  assign n3413 = pi20 ? n3410 : n3412;
  assign n3414 = pi19 ? n3413 : n2094;
  assign n3415 = pi18 ? n3414 : n2681;
  assign n3416 = pi17 ? n3408 : n3415;
  assign n3417 = pi16 ? n439 : n3416;
  assign n3418 = pi15 ? n3403 : n3417;
  assign n3419 = pi14 ? n3389 : n3418;
  assign n3420 = pi20 ? n2094 : n2091;
  assign n3421 = pi19 ? n37 : n3420;
  assign n3422 = pi18 ? n3421 : n2703;
  assign n3423 = pi17 ? n37 : n3422;
  assign n3424 = pi16 ? n439 : n3423;
  assign n3425 = pi18 ? n2102 : n1824;
  assign n3426 = pi17 ? n37 : n3425;
  assign n3427 = pi16 ? n439 : n3426;
  assign n3428 = pi15 ? n3424 : n3427;
  assign n3429 = pi14 ? n2699 : n3428;
  assign n3430 = pi13 ? n3419 : n3429;
  assign n3431 = pi18 ? n2109 : n1824;
  assign n3432 = pi17 ? n37 : n3431;
  assign n3433 = pi16 ? n439 : n3432;
  assign n3434 = pi15 ? n2112 : n3433;
  assign n3435 = pi14 ? n3434 : n2735;
  assign n3436 = pi22 ? n363 : n316;
  assign n3437 = pi21 ? n722 : n3436;
  assign n3438 = pi20 ? n99 : n3437;
  assign n3439 = pi19 ? n99 : n3438;
  assign n3440 = pi18 ? n3439 : n32;
  assign n3441 = pi17 ? n99 : n3440;
  assign n3442 = pi16 ? n721 : n3441;
  assign n3443 = pi23 ? n99 : n685;
  assign n3444 = pi22 ? n99 : n3443;
  assign n3445 = pi22 ? n685 : n316;
  assign n3446 = pi21 ? n3444 : n3445;
  assign n3447 = pi20 ? n99 : n3446;
  assign n3448 = pi19 ? n99 : n3447;
  assign n3449 = pi18 ? n3448 : n32;
  assign n3450 = pi17 ? n99 : n3449;
  assign n3451 = pi16 ? n721 : n3450;
  assign n3452 = pi15 ? n3442 : n3451;
  assign n3453 = pi22 ? n3443 : n759;
  assign n3454 = pi21 ? n99 : n3453;
  assign n3455 = pi20 ? n99 : n3454;
  assign n3456 = pi19 ? n99 : n3455;
  assign n3457 = pi18 ? n3456 : n32;
  assign n3458 = pi17 ? n99 : n3457;
  assign n3459 = pi16 ? n801 : n3458;
  assign n3460 = pi22 ? n158 : n759;
  assign n3461 = pi21 ? n99 : n3460;
  assign n3462 = pi20 ? n99 : n3461;
  assign n3463 = pi19 ? n99 : n3462;
  assign n3464 = pi18 ? n3463 : n32;
  assign n3465 = pi17 ? n99 : n3464;
  assign n3466 = pi16 ? n801 : n3465;
  assign n3467 = pi15 ? n3459 : n3466;
  assign n3468 = pi14 ? n3452 : n3467;
  assign n3469 = pi13 ? n3435 : n3468;
  assign n3470 = pi12 ? n3430 : n3469;
  assign n3471 = pi16 ? n744 : n3458;
  assign n3472 = pi23 ? n139 : n685;
  assign n3473 = pi22 ? n3472 : n396;
  assign n3474 = pi21 ? n99 : n3473;
  assign n3475 = pi20 ? n99 : n3474;
  assign n3476 = pi19 ? n99 : n3475;
  assign n3477 = pi18 ? n3476 : n32;
  assign n3478 = pi17 ? n99 : n3477;
  assign n3479 = pi16 ? n721 : n3478;
  assign n3480 = pi15 ? n3471 : n3479;
  assign n3481 = pi20 ? n99 : n2999;
  assign n3482 = pi19 ? n99 : n3481;
  assign n3483 = pi18 ? n3482 : n99;
  assign n3484 = pi21 ? n159 : n157;
  assign n3485 = pi21 ? n2998 : n2230;
  assign n3486 = pi20 ? n3484 : n3485;
  assign n3487 = pi19 ? n99 : n3486;
  assign n3488 = pi18 ? n3487 : n32;
  assign n3489 = pi17 ? n3483 : n3488;
  assign n3490 = pi16 ? n721 : n3489;
  assign n3491 = pi24 ? n99 : n139;
  assign n3492 = pi23 ? n99 : n3491;
  assign n3493 = pi22 ? n99 : n3492;
  assign n3494 = pi22 ? n316 : n688;
  assign n3495 = pi21 ? n3493 : n3494;
  assign n3496 = pi20 ? n787 : n3495;
  assign n3497 = pi19 ? n99 : n3496;
  assign n3498 = pi18 ? n3497 : n32;
  assign n3499 = pi17 ? n99 : n3498;
  assign n3500 = pi16 ? n721 : n3499;
  assign n3501 = pi15 ? n3490 : n3500;
  assign n3502 = pi14 ? n3480 : n3501;
  assign n3503 = pi21 ? n796 : n2162;
  assign n3504 = pi20 ? n32 : n3503;
  assign n3505 = pi19 ? n32 : n3504;
  assign n3506 = pi21 ? n1143 : n2161;
  assign n3507 = pi20 ? n2165 : n3506;
  assign n3508 = pi21 ? n112 : n2161;
  assign n3509 = pi20 ? n3508 : n2189;
  assign n3510 = pi19 ? n3507 : n3509;
  assign n3511 = pi18 ? n3505 : n3510;
  assign n3512 = pi17 ? n32 : n3511;
  assign n3513 = pi20 ? n2174 : n2746;
  assign n3514 = pi20 ? n2164 : n2165;
  assign n3515 = pi19 ? n3513 : n3514;
  assign n3516 = pi21 ? n1143 : n2162;
  assign n3517 = pi20 ? n3516 : n2165;
  assign n3518 = pi19 ? n3517 : n2166;
  assign n3519 = pi18 ? n3515 : n3518;
  assign n3520 = pi22 ? n812 : n157;
  assign n3521 = pi21 ? n746 : n3520;
  assign n3522 = pi20 ? n2164 : n3521;
  assign n3523 = pi22 ? n316 : n706;
  assign n3524 = pi21 ? n819 : n3523;
  assign n3525 = pi20 ? n157 : n3524;
  assign n3526 = pi19 ? n3522 : n3525;
  assign n3527 = pi18 ? n3526 : n32;
  assign n3528 = pi17 ? n3519 : n3527;
  assign n3529 = pi16 ? n3512 : n3528;
  assign n3530 = pi21 ? n326 : n1711;
  assign n3531 = pi20 ? n32 : n3530;
  assign n3532 = pi19 ? n32 : n3531;
  assign n3533 = pi20 ? n139 : n1719;
  assign n3534 = pi20 ? n1715 : n2521;
  assign n3535 = pi19 ? n3533 : n3534;
  assign n3536 = pi18 ? n3532 : n3535;
  assign n3537 = pi17 ? n32 : n3536;
  assign n3538 = pi20 ? n3245 : n2518;
  assign n3539 = pi19 ? n3538 : n139;
  assign n3540 = pi20 ? n139 : n1715;
  assign n3541 = pi18 ? n3539 : n3540;
  assign n3542 = pi20 ? n1719 : n249;
  assign n3543 = pi21 ? n157 : n2245;
  assign n3544 = pi20 ? n157 : n3543;
  assign n3545 = pi19 ? n3542 : n3544;
  assign n3546 = pi18 ? n3545 : n32;
  assign n3547 = pi17 ? n3541 : n3546;
  assign n3548 = pi16 ? n3537 : n3547;
  assign n3549 = pi15 ? n3529 : n3548;
  assign n3550 = pi20 ? n1719 : n1712;
  assign n3551 = pi19 ? n2522 : n3550;
  assign n3552 = pi18 ? n913 : n3551;
  assign n3553 = pi17 ? n32 : n3552;
  assign n3554 = pi20 ? n139 : n2518;
  assign n3555 = pi20 ? n2365 : n1715;
  assign n3556 = pi19 ? n3554 : n3555;
  assign n3557 = pi21 ? n139 : n1529;
  assign n3558 = pi20 ? n3557 : n139;
  assign n3559 = pi19 ? n3558 : n2831;
  assign n3560 = pi18 ? n3556 : n3559;
  assign n3561 = pi20 ? n1531 : n249;
  assign n3562 = pi22 ? n157 : n316;
  assign n3563 = pi21 ? n3562 : n3523;
  assign n3564 = pi20 ? n157 : n3563;
  assign n3565 = pi19 ? n3561 : n3564;
  assign n3566 = pi18 ? n3565 : n32;
  assign n3567 = pi17 ? n3560 : n3566;
  assign n3568 = pi16 ? n3553 : n3567;
  assign n3569 = pi21 ? n910 : n1531;
  assign n3570 = pi20 ? n32 : n3569;
  assign n3571 = pi19 ? n32 : n3570;
  assign n3572 = pi21 ? n139 : n1696;
  assign n3573 = pi20 ? n3572 : n2510;
  assign n3574 = pi20 ? n1719 : n1757;
  assign n3575 = pi19 ? n3573 : n3574;
  assign n3576 = pi18 ? n3571 : n3575;
  assign n3577 = pi17 ? n32 : n3576;
  assign n3578 = pi20 ? n139 : n947;
  assign n3579 = pi21 ? n1698 : n297;
  assign n3580 = pi20 ? n2365 : n3579;
  assign n3581 = pi19 ? n3578 : n3580;
  assign n3582 = pi20 ? n1711 : n139;
  assign n3583 = pi19 ? n3558 : n3582;
  assign n3584 = pi18 ? n3581 : n3583;
  assign n3585 = pi20 ? n1531 : n2316;
  assign n3586 = pi21 ? n346 : n3523;
  assign n3587 = pi20 ? n2318 : n3586;
  assign n3588 = pi19 ? n3585 : n3587;
  assign n3589 = pi18 ? n3588 : n32;
  assign n3590 = pi17 ? n3584 : n3589;
  assign n3591 = pi16 ? n3577 : n3590;
  assign n3592 = pi15 ? n3568 : n3591;
  assign n3593 = pi14 ? n3549 : n3592;
  assign n3594 = pi13 ? n3502 : n3593;
  assign n3595 = pi21 ? n326 : n820;
  assign n3596 = pi20 ? n32 : n3595;
  assign n3597 = pi19 ? n32 : n3596;
  assign n3598 = pi21 ? n3073 : n1711;
  assign n3599 = pi20 ? n3572 : n3598;
  assign n3600 = pi20 ? n947 : n3090;
  assign n3601 = pi19 ? n3599 : n3600;
  assign n3602 = pi18 ? n3597 : n3601;
  assign n3603 = pi17 ? n32 : n3602;
  assign n3604 = pi20 ? n1757 : n947;
  assign n3605 = pi21 ? n1211 : n1698;
  assign n3606 = pi21 ? n1698 : n1696;
  assign n3607 = pi20 ? n3605 : n3606;
  assign n3608 = pi19 ? n3604 : n3607;
  assign n3609 = pi21 ? n1711 : n375;
  assign n3610 = pi21 ? n1211 : n297;
  assign n3611 = pi20 ? n3609 : n3610;
  assign n3612 = pi21 ? n1711 : n820;
  assign n3613 = pi20 ? n3612 : n3610;
  assign n3614 = pi19 ? n3611 : n3613;
  assign n3615 = pi18 ? n3608 : n3614;
  assign n3616 = pi22 ? n2401 : n139;
  assign n3617 = pi22 ? n1784 : n139;
  assign n3618 = pi21 ? n3616 : n3617;
  assign n3619 = pi21 ? n316 : n2320;
  assign n3620 = pi20 ? n3618 : n3619;
  assign n3621 = pi19 ? n3585 : n3620;
  assign n3622 = pi18 ? n3621 : n32;
  assign n3623 = pi17 ? n3615 : n3622;
  assign n3624 = pi16 ? n3603 : n3623;
  assign n3625 = pi21 ? n1721 : n139;
  assign n3626 = pi20 ? n139 : n3625;
  assign n3627 = pi19 ? n3626 : n139;
  assign n3628 = pi18 ? n329 : n3627;
  assign n3629 = pi17 ? n32 : n3628;
  assign n3630 = pi20 ? n316 : n3619;
  assign n3631 = pi19 ? n139 : n3630;
  assign n3632 = pi18 ? n3631 : n32;
  assign n3633 = pi17 ? n139 : n3632;
  assign n3634 = pi16 ? n3629 : n3633;
  assign n3635 = pi15 ? n3624 : n3634;
  assign n3636 = pi20 ? n975 : n3619;
  assign n3637 = pi19 ? n139 : n3636;
  assign n3638 = pi18 ? n3637 : n32;
  assign n3639 = pi17 ? n139 : n3638;
  assign n3640 = pi16 ? n915 : n3639;
  assign n3641 = pi21 ? n296 : n820;
  assign n3642 = pi20 ? n32 : n3641;
  assign n3643 = pi19 ? n32 : n3642;
  assign n3644 = pi20 ? n2519 : n3625;
  assign n3645 = pi21 ? n375 : n139;
  assign n3646 = pi20 ? n3645 : n3612;
  assign n3647 = pi19 ? n3644 : n3646;
  assign n3648 = pi18 ? n3643 : n3647;
  assign n3649 = pi17 ? n32 : n3648;
  assign n3650 = pi20 ? n3572 : n139;
  assign n3651 = pi21 ? n139 : n295;
  assign n3652 = pi20 ? n3651 : n2521;
  assign n3653 = pi19 ? n3650 : n3652;
  assign n3654 = pi21 ? n1531 : n1721;
  assign n3655 = pi20 ? n3654 : n3612;
  assign n3656 = pi21 ? n1211 : n1721;
  assign n3657 = pi20 ? n3656 : n3612;
  assign n3658 = pi19 ? n3655 : n3657;
  assign n3659 = pi18 ? n3653 : n3658;
  assign n3660 = pi21 ? n346 : n2320;
  assign n3661 = pi20 ? n2353 : n3660;
  assign n3662 = pi19 ? n2352 : n3661;
  assign n3663 = pi18 ? n3662 : n32;
  assign n3664 = pi17 ? n3659 : n3663;
  assign n3665 = pi16 ? n3649 : n3664;
  assign n3666 = pi15 ? n3640 : n3665;
  assign n3667 = pi14 ? n3635 : n3666;
  assign n3668 = pi22 ? n1043 : n37;
  assign n3669 = pi21 ? n1721 : n3668;
  assign n3670 = pi20 ? n3669 : n942;
  assign n3671 = pi21 ? n1696 : n820;
  assign n3672 = pi20 ? n3096 : n3671;
  assign n3673 = pi19 ? n3670 : n3672;
  assign n3674 = pi18 ? n3643 : n3673;
  assign n3675 = pi17 ? n32 : n3674;
  assign n3676 = pi21 ? n1711 : n1529;
  assign n3677 = pi20 ? n3572 : n3676;
  assign n3678 = pi21 ? n1529 : n375;
  assign n3679 = pi20 ? n3678 : n1757;
  assign n3680 = pi19 ? n3677 : n3679;
  assign n3681 = pi20 ? n3579 : n3612;
  assign n3682 = pi20 ? n3610 : n3612;
  assign n3683 = pi19 ? n3681 : n3682;
  assign n3684 = pi18 ? n3680 : n3683;
  assign n3685 = pi20 ? n1022 : n3660;
  assign n3686 = pi19 ? n2352 : n3685;
  assign n3687 = pi18 ? n3686 : n32;
  assign n3688 = pi17 ? n3684 : n3687;
  assign n3689 = pi16 ? n3675 : n3688;
  assign n3690 = pi24 ? n32 : n316;
  assign n3691 = pi23 ? n3690 : n37;
  assign n3692 = pi22 ? n3691 : n316;
  assign n3693 = pi22 ? n335 : n316;
  assign n3694 = pi21 ? n3692 : n3693;
  assign n3695 = pi20 ? n32 : n3694;
  assign n3696 = pi19 ? n32 : n3695;
  assign n3697 = pi21 ? n3258 : n316;
  assign n3698 = pi22 ? n335 : n383;
  assign n3699 = pi21 ? n3258 : n3698;
  assign n3700 = pi20 ? n3697 : n3699;
  assign n3701 = pi21 ? n316 : n569;
  assign n3702 = pi21 ? n381 : n316;
  assign n3703 = pi20 ? n3701 : n3702;
  assign n3704 = pi19 ? n3700 : n3703;
  assign n3705 = pi18 ? n3696 : n3704;
  assign n3706 = pi17 ? n32 : n3705;
  assign n3707 = pi21 ? n3693 : n316;
  assign n3708 = pi20 ? n3707 : n316;
  assign n3709 = pi19 ? n3708 : n316;
  assign n3710 = pi18 ? n3709 : n316;
  assign n3711 = pi22 ? n348 : n37;
  assign n3712 = pi21 ? n316 : n3711;
  assign n3713 = pi20 ? n3712 : n2330;
  assign n3714 = pi19 ? n316 : n3713;
  assign n3715 = pi18 ? n3714 : n32;
  assign n3716 = pi17 ? n3710 : n3715;
  assign n3717 = pi16 ? n3706 : n3716;
  assign n3718 = pi15 ? n3689 : n3717;
  assign n3719 = pi24 ? n32 : n204;
  assign n3720 = pi23 ? n3719 : n99;
  assign n3721 = pi22 ? n3720 : n204;
  assign n3722 = pi21 ? n3721 : n1027;
  assign n3723 = pi20 ? n32 : n3722;
  assign n3724 = pi19 ? n32 : n3723;
  assign n3725 = pi18 ? n3724 : n204;
  assign n3726 = pi17 ? n32 : n3725;
  assign n3727 = pi20 ? n204 : n2383;
  assign n3728 = pi21 ? n316 : n1018;
  assign n3729 = pi20 ? n316 : n3728;
  assign n3730 = pi19 ? n3727 : n3729;
  assign n3731 = pi21 ? n316 : n204;
  assign n3732 = pi20 ? n2383 : n3731;
  assign n3733 = pi20 ? n1028 : n3731;
  assign n3734 = pi19 ? n3732 : n3733;
  assign n3735 = pi18 ? n3730 : n3734;
  assign n3736 = pi20 ? n2383 : n316;
  assign n3737 = pi21 ? n1027 : n928;
  assign n3738 = pi20 ? n3731 : n3737;
  assign n3739 = pi19 ? n3736 : n3738;
  assign n3740 = pi18 ? n3739 : n32;
  assign n3741 = pi17 ? n3735 : n3740;
  assign n3742 = pi16 ? n3726 : n3741;
  assign n3743 = pi21 ? n3721 : n1079;
  assign n3744 = pi20 ? n32 : n3743;
  assign n3745 = pi19 ? n32 : n3744;
  assign n3746 = pi22 ? n335 : n99;
  assign n3747 = pi21 ? n3746 : n204;
  assign n3748 = pi20 ? n1099 : n3747;
  assign n3749 = pi21 ? n1079 : n204;
  assign n3750 = pi19 ? n3748 : n3749;
  assign n3751 = pi18 ? n3745 : n3750;
  assign n3752 = pi17 ? n32 : n3751;
  assign n3753 = pi21 ? n1079 : n1083;
  assign n3754 = pi20 ? n3753 : n1083;
  assign n3755 = pi20 ? n1083 : n1099;
  assign n3756 = pi19 ? n3754 : n3755;
  assign n3757 = pi20 ? n1079 : n1099;
  assign n3758 = pi18 ? n3756 : n3757;
  assign n3759 = pi22 ? n99 : n204;
  assign n3760 = pi21 ? n204 : n3759;
  assign n3761 = pi20 ? n3749 : n3760;
  assign n3762 = pi23 ? n204 : n685;
  assign n3763 = pi22 ? n204 : n3762;
  assign n3764 = pi21 ? n3763 : n2700;
  assign n3765 = pi20 ? n204 : n3764;
  assign n3766 = pi19 ? n3761 : n3765;
  assign n3767 = pi18 ? n3766 : n32;
  assign n3768 = pi17 ? n3758 : n3767;
  assign n3769 = pi16 ? n3752 : n3768;
  assign n3770 = pi15 ? n3742 : n3769;
  assign n3771 = pi14 ? n3718 : n3770;
  assign n3772 = pi13 ? n3667 : n3771;
  assign n3773 = pi12 ? n3594 : n3772;
  assign n3774 = pi11 ? n3470 : n3773;
  assign n3775 = pi10 ? n3373 : n3774;
  assign n3776 = pi09 ? n32 : n3775;
  assign n3777 = pi16 ? n2447 : n2951;
  assign n3778 = pi15 ? n32 : n3777;
  assign n3779 = pi22 ? n39 : n37;
  assign n3780 = pi21 ? n3779 : n37;
  assign n3781 = pi20 ? n3780 : n37;
  assign n3782 = pi19 ? n3781 : n37;
  assign n3783 = pi18 ? n32 : n3782;
  assign n3784 = pi17 ? n32 : n3783;
  assign n3785 = pi16 ? n3784 : n2951;
  assign n3786 = pi16 ? n70 : n2951;
  assign n3787 = pi15 ? n3785 : n3786;
  assign n3788 = pi14 ? n3778 : n3787;
  assign n3789 = pi16 ? n73 : n2951;
  assign n3790 = pi15 ? n3789 : n2952;
  assign n3791 = pi22 ? n1617 : n32;
  assign n3792 = pi21 ? n3791 : n32;
  assign n3793 = pi20 ? n3792 : n32;
  assign n3794 = pi19 ? n3793 : n32;
  assign n3795 = pi18 ? n37 : n3794;
  assign n3796 = pi17 ? n37 : n3795;
  assign n3797 = pi16 ? n2461 : n3796;
  assign n3798 = pi15 ? n2953 : n3797;
  assign n3799 = pi14 ? n3790 : n3798;
  assign n3800 = pi13 ? n3788 : n3799;
  assign n3801 = pi22 ? n64 : n2160;
  assign n3802 = pi21 ? n32 : n3801;
  assign n3803 = pi20 ? n32 : n3802;
  assign n3804 = pi19 ? n32 : n3803;
  assign n3805 = pi21 ? n112 : n2160;
  assign n3806 = pi20 ? n3805 : n2755;
  assign n3807 = pi21 ? n2161 : n2164;
  assign n3808 = pi20 ? n2740 : n3807;
  assign n3809 = pi19 ? n3806 : n3808;
  assign n3810 = pi18 ? n3804 : n3809;
  assign n3811 = pi17 ? n32 : n3810;
  assign n3812 = pi21 ? n2160 : n99;
  assign n3813 = pi20 ? n3812 : n2167;
  assign n3814 = pi21 ? n112 : n2175;
  assign n3815 = pi20 ? n2755 : n3814;
  assign n3816 = pi19 ? n3813 : n3815;
  assign n3817 = pi21 ? n1143 : n2175;
  assign n3818 = pi20 ? n3817 : n2968;
  assign n3819 = pi20 ? n3814 : n2184;
  assign n3820 = pi19 ? n3818 : n3819;
  assign n3821 = pi18 ? n3816 : n3820;
  assign n3822 = pi21 ? n2156 : n2168;
  assign n3823 = pi20 ? n2184 : n3822;
  assign n3824 = pi21 ? n2175 : n2164;
  assign n3825 = pi21 ? n2175 : n99;
  assign n3826 = pi20 ? n3824 : n3825;
  assign n3827 = pi19 ? n3823 : n3826;
  assign n3828 = pi18 ? n3827 : n2949;
  assign n3829 = pi17 ? n3821 : n3828;
  assign n3830 = pi16 ? n3811 : n3829;
  assign n3831 = pi23 ? n99 : n102;
  assign n3832 = pi22 ? n3831 : n32;
  assign n3833 = pi21 ? n3832 : n32;
  assign n3834 = pi20 ? n3833 : n32;
  assign n3835 = pi19 ? n3834 : n32;
  assign n3836 = pi18 ? n99 : n3835;
  assign n3837 = pi17 ? n99 : n3836;
  assign n3838 = pi16 ? n1148 : n3837;
  assign n3839 = pi15 ? n3830 : n3838;
  assign n3840 = pi23 ? n99 : n46;
  assign n3841 = pi22 ? n3840 : n32;
  assign n3842 = pi21 ? n3841 : n32;
  assign n3843 = pi20 ? n3842 : n32;
  assign n3844 = pi19 ? n3843 : n32;
  assign n3845 = pi18 ? n99 : n3844;
  assign n3846 = pi17 ? n99 : n3845;
  assign n3847 = pi16 ? n721 : n3846;
  assign n3848 = pi22 ? n1167 : n32;
  assign n3849 = pi21 ? n3848 : n32;
  assign n3850 = pi20 ? n3849 : n32;
  assign n3851 = pi19 ? n3850 : n32;
  assign n3852 = pi18 ? n3015 : n3851;
  assign n3853 = pi17 ? n3009 : n3852;
  assign n3854 = pi16 ? n186 : n3853;
  assign n3855 = pi15 ? n3847 : n3854;
  assign n3856 = pi14 ? n3839 : n3855;
  assign n3857 = pi16 ? n721 : n3837;
  assign n3858 = pi23 ? n139 : n102;
  assign n3859 = pi22 ? n3858 : n32;
  assign n3860 = pi21 ? n3859 : n32;
  assign n3861 = pi20 ? n3860 : n32;
  assign n3862 = pi19 ? n3861 : n32;
  assign n3863 = pi18 ? n99 : n3862;
  assign n3864 = pi17 ? n99 : n3863;
  assign n3865 = pi16 ? n721 : n3864;
  assign n3866 = pi21 ? n180 : n2746;
  assign n3867 = pi20 ? n32 : n3866;
  assign n3868 = pi19 ? n32 : n3867;
  assign n3869 = pi21 ? n112 : n181;
  assign n3870 = pi21 ? n2168 : n2156;
  assign n3871 = pi21 ? n2746 : n112;
  assign n3872 = pi20 ? n3870 : n3871;
  assign n3873 = pi19 ? n3869 : n3872;
  assign n3874 = pi18 ? n3868 : n3873;
  assign n3875 = pi17 ? n32 : n3874;
  assign n3876 = pi21 ? n181 : n2168;
  assign n3877 = pi21 ? n2156 : n2746;
  assign n3878 = pi20 ? n3876 : n3877;
  assign n3879 = pi21 ? n112 : n99;
  assign n3880 = pi20 ? n3877 : n3879;
  assign n3881 = pi19 ? n3878 : n3880;
  assign n3882 = pi21 ? n218 : n2746;
  assign n3883 = pi20 ? n3879 : n3882;
  assign n3884 = pi21 ? n2164 : n181;
  assign n3885 = pi20 ? n3869 : n3884;
  assign n3886 = pi19 ? n3883 : n3885;
  assign n3887 = pi18 ? n3881 : n3886;
  assign n3888 = pi21 ? n2164 : n99;
  assign n3889 = pi20 ? n3888 : n99;
  assign n3890 = pi21 ? n181 : n2161;
  assign n3891 = pi21 ? n181 : n2981;
  assign n3892 = pi20 ? n3890 : n3891;
  assign n3893 = pi19 ? n3889 : n3892;
  assign n3894 = pi22 ? n861 : n32;
  assign n3895 = pi21 ? n3894 : n32;
  assign n3896 = pi20 ? n3895 : n32;
  assign n3897 = pi19 ? n3896 : n32;
  assign n3898 = pi18 ? n3893 : n3897;
  assign n3899 = pi17 ? n3887 : n3898;
  assign n3900 = pi16 ? n3875 : n3899;
  assign n3901 = pi15 ? n3865 : n3900;
  assign n3902 = pi14 ? n3857 : n3901;
  assign n3903 = pi13 ? n3856 : n3902;
  assign n3904 = pi12 ? n3800 : n3903;
  assign n3905 = pi23 ? n335 : n102;
  assign n3906 = pi22 ? n3905 : n32;
  assign n3907 = pi21 ? n3906 : n32;
  assign n3908 = pi20 ? n3907 : n32;
  assign n3909 = pi19 ? n3908 : n32;
  assign n3910 = pi18 ? n99 : n3909;
  assign n3911 = pi17 ? n99 : n3910;
  assign n3912 = pi16 ? n3065 : n3911;
  assign n3913 = pi21 ? n1698 : n1721;
  assign n3914 = pi20 ? n3913 : n1699;
  assign n3915 = pi21 ? n1711 : n295;
  assign n3916 = pi21 ? n297 : n1698;
  assign n3917 = pi20 ? n3915 : n3916;
  assign n3918 = pi19 ? n3914 : n3917;
  assign n3919 = pi18 ? n1692 : n3918;
  assign n3920 = pi17 ? n32 : n3919;
  assign n3921 = pi21 ? n375 : n1711;
  assign n3922 = pi21 ? n295 : n297;
  assign n3923 = pi20 ? n3921 : n3922;
  assign n3924 = pi21 ? n3668 : n297;
  assign n3925 = pi21 ? n1698 : n139;
  assign n3926 = pi20 ? n3924 : n3925;
  assign n3927 = pi19 ? n3923 : n3926;
  assign n3928 = pi20 ? n3925 : n3092;
  assign n3929 = pi20 ? n3913 : n3654;
  assign n3930 = pi19 ? n3928 : n3929;
  assign n3931 = pi18 ? n3927 : n3930;
  assign n3932 = pi21 ? n375 : n820;
  assign n3933 = pi20 ? n3645 : n3932;
  assign n3934 = pi19 ? n1720 : n3933;
  assign n3935 = pi23 ? n335 : n157;
  assign n3936 = pi22 ? n3935 : n32;
  assign n3937 = pi21 ? n3936 : n32;
  assign n3938 = pi20 ? n3937 : n32;
  assign n3939 = pi19 ? n3938 : n32;
  assign n3940 = pi18 ? n3934 : n3939;
  assign n3941 = pi17 ? n3931 : n3940;
  assign n3942 = pi16 ? n3920 : n3941;
  assign n3943 = pi15 ? n3912 : n3942;
  assign n3944 = pi23 ? n363 : n157;
  assign n3945 = pi22 ? n3944 : n32;
  assign n3946 = pi21 ? n3945 : n32;
  assign n3947 = pi20 ? n3946 : n32;
  assign n3948 = pi19 ? n3947 : n32;
  assign n3949 = pi18 ? n3123 : n3948;
  assign n3950 = pi17 ? n3116 : n3949;
  assign n3951 = pi16 ? n3108 : n3950;
  assign n3952 = pi22 ? n456 : n32;
  assign n3953 = pi21 ? n3952 : n32;
  assign n3954 = pi20 ? n3953 : n32;
  assign n3955 = pi19 ? n3954 : n32;
  assign n3956 = pi18 ? n139 : n3955;
  assign n3957 = pi17 ? n139 : n3956;
  assign n3958 = pi16 ? n1773 : n3957;
  assign n3959 = pi15 ? n3951 : n3958;
  assign n3960 = pi14 ? n3943 : n3959;
  assign n3961 = pi23 ? n99 : n204;
  assign n3962 = pi22 ? n3961 : n32;
  assign n3963 = pi21 ? n3962 : n32;
  assign n3964 = pi20 ? n3963 : n32;
  assign n3965 = pi19 ? n3964 : n32;
  assign n3966 = pi18 ? n139 : n3965;
  assign n3967 = pi17 ? n139 : n3966;
  assign n3968 = pi16 ? n331 : n3967;
  assign n3969 = pi15 ? n3958 : n3968;
  assign n3970 = pi22 ? n1038 : n32;
  assign n3971 = pi21 ? n3970 : n32;
  assign n3972 = pi20 ? n3971 : n32;
  assign n3973 = pi19 ? n3972 : n32;
  assign n3974 = pi18 ? n139 : n3973;
  assign n3975 = pi17 ? n139 : n3974;
  assign n3976 = pi16 ? n331 : n3975;
  assign n3977 = pi21 ? n2300 : n32;
  assign n3978 = pi20 ? n3977 : n32;
  assign n3979 = pi19 ? n3978 : n32;
  assign n3980 = pi18 ? n3173 : n3979;
  assign n3981 = pi17 ? n3170 : n3980;
  assign n3982 = pi16 ? n3165 : n3981;
  assign n3983 = pi15 ? n3976 : n3982;
  assign n3984 = pi14 ? n3969 : n3983;
  assign n3985 = pi13 ? n3960 : n3984;
  assign n3986 = pi22 ? n55 : n383;
  assign n3987 = pi21 ? n3986 : n1027;
  assign n3988 = pi20 ? n32 : n3987;
  assign n3989 = pi19 ? n32 : n3988;
  assign n3990 = pi22 ? n316 : n2299;
  assign n3991 = pi21 ? n3990 : n2412;
  assign n3992 = pi21 ? n2409 : n2299;
  assign n3993 = pi22 ? n316 : n2401;
  assign n3994 = pi21 ? n3993 : n3990;
  assign n3995 = pi20 ? n3992 : n3994;
  assign n3996 = pi19 ? n3991 : n3995;
  assign n3997 = pi18 ? n3989 : n3996;
  assign n3998 = pi17 ? n32 : n3997;
  assign n3999 = pi21 ? n2412 : n2409;
  assign n4000 = pi21 ? n2299 : n3993;
  assign n4001 = pi20 ? n3999 : n4000;
  assign n4002 = pi21 ? n316 : n1027;
  assign n4003 = pi20 ? n4002 : n316;
  assign n4004 = pi19 ? n4001 : n4003;
  assign n4005 = pi18 ? n4004 : n316;
  assign n4006 = pi21 ? n316 : n2409;
  assign n4007 = pi19 ? n316 : n4006;
  assign n4008 = pi21 ? n3523 : n32;
  assign n4009 = pi20 ? n4008 : n32;
  assign n4010 = pi19 ? n4009 : n32;
  assign n4011 = pi18 ? n4007 : n4010;
  assign n4012 = pi17 ? n4005 : n4011;
  assign n4013 = pi16 ? n3998 : n4012;
  assign n4014 = pi22 ? n348 : n383;
  assign n4015 = pi22 ? n383 : n316;
  assign n4016 = pi21 ? n4014 : n4015;
  assign n4017 = pi22 ? n383 : n139;
  assign n4018 = pi21 ? n4014 : n4017;
  assign n4019 = pi20 ? n4016 : n4018;
  assign n4020 = pi22 ? n316 : n348;
  assign n4021 = pi21 ? n4020 : n383;
  assign n4022 = pi21 ? n346 : n4014;
  assign n4023 = pi20 ? n4021 : n4022;
  assign n4024 = pi19 ? n4019 : n4023;
  assign n4025 = pi18 ? n3218 : n4024;
  assign n4026 = pi17 ? n32 : n4025;
  assign n4027 = pi21 ? n4017 : n4020;
  assign n4028 = pi21 ? n383 : n346;
  assign n4029 = pi20 ? n4027 : n4028;
  assign n4030 = pi22 ? n348 : n295;
  assign n4031 = pi21 ? n4030 : n346;
  assign n4032 = pi21 ? n4014 : n1211;
  assign n4033 = pi20 ? n4031 : n4032;
  assign n4034 = pi19 ? n4029 : n4033;
  assign n4035 = pi21 ? n3219 : n346;
  assign n4036 = pi20 ? n4032 : n4035;
  assign n4037 = pi22 ? n383 : n1043;
  assign n4038 = pi21 ? n4014 : n4037;
  assign n4039 = pi21 ? n1777 : n4037;
  assign n4040 = pi20 ? n4038 : n4039;
  assign n4041 = pi19 ? n4036 : n4040;
  assign n4042 = pi18 ? n4034 : n4041;
  assign n4043 = pi21 ? n4017 : n3224;
  assign n4044 = pi19 ? n3246 : n4043;
  assign n4045 = pi18 ? n4044 : n4010;
  assign n4046 = pi17 ? n4042 : n4045;
  assign n4047 = pi16 ? n4026 : n4046;
  assign n4048 = pi15 ? n4013 : n4047;
  assign n4049 = pi21 ? n3986 : n381;
  assign n4050 = pi20 ? n32 : n4049;
  assign n4051 = pi19 ? n32 : n4050;
  assign n4052 = pi22 ? n390 : n383;
  assign n4053 = pi21 ? n4052 : n316;
  assign n4054 = pi21 ? n4052 : n384;
  assign n4055 = pi20 ? n4053 : n4054;
  assign n4056 = pi22 ? n316 : n390;
  assign n4057 = pi21 ? n4056 : n383;
  assign n4058 = pi21 ? n381 : n4052;
  assign n4059 = pi20 ? n4057 : n4058;
  assign n4060 = pi19 ? n4055 : n4059;
  assign n4061 = pi18 ? n4051 : n4060;
  assign n4062 = pi17 ? n32 : n4061;
  assign n4063 = pi21 ? n384 : n4056;
  assign n4064 = pi21 ? n383 : n381;
  assign n4065 = pi20 ? n4063 : n4064;
  assign n4066 = pi21 ? n4052 : n381;
  assign n4067 = pi20 ? n3275 : n4066;
  assign n4068 = pi19 ? n4065 : n4067;
  assign n4069 = pi20 ? n4066 : n4064;
  assign n4070 = pi21 ? n4052 : n3118;
  assign n4071 = pi21 ? n392 : n3118;
  assign n4072 = pi20 ? n4070 : n4071;
  assign n4073 = pi19 ? n4069 : n4072;
  assign n4074 = pi18 ? n4068 : n4073;
  assign n4075 = pi19 ? n3276 : n426;
  assign n4076 = pi18 ? n4075 : n4010;
  assign n4077 = pi17 ? n4074 : n4076;
  assign n4078 = pi16 ? n4062 : n4077;
  assign n4079 = pi23 ? n204 : n233;
  assign n4080 = pi22 ? n4079 : n32;
  assign n4081 = pi21 ? n4080 : n32;
  assign n4082 = pi20 ? n4081 : n32;
  assign n4083 = pi19 ? n4082 : n32;
  assign n4084 = pi18 ? n3300 : n4083;
  assign n4085 = pi17 ? n3295 : n4084;
  assign n4086 = pi16 ? n3288 : n4085;
  assign n4087 = pi15 ? n4078 : n4086;
  assign n4088 = pi14 ? n4048 : n4087;
  assign n4089 = pi21 ? n335 : n1940;
  assign n4090 = pi20 ? n4089 : n335;
  assign n4091 = pi19 ? n4090 : n335;
  assign n4092 = pi18 ? n602 : n4091;
  assign n4093 = pi17 ? n32 : n4092;
  assign n4094 = pi22 ? n3762 : n32;
  assign n4095 = pi21 ? n4094 : n32;
  assign n4096 = pi20 ? n4095 : n32;
  assign n4097 = pi19 ? n4096 : n32;
  assign n4098 = pi18 ? n3317 : n4097;
  assign n4099 = pi17 ? n3314 : n4098;
  assign n4100 = pi16 ? n4093 : n4099;
  assign n4101 = pi22 ? n1070 : n32;
  assign n4102 = pi21 ? n4101 : n32;
  assign n4103 = pi20 ? n4102 : n32;
  assign n4104 = pi19 ? n4103 : n32;
  assign n4105 = pi18 ? n3337 : n4104;
  assign n4106 = pi17 ? n3334 : n4105;
  assign n4107 = pi16 ? n3329 : n4106;
  assign n4108 = pi15 ? n4100 : n4107;
  assign n4109 = pi22 ? n1388 : n32;
  assign n4110 = pi21 ? n4109 : n32;
  assign n4111 = pi20 ? n4110 : n32;
  assign n4112 = pi19 ? n4111 : n32;
  assign n4113 = pi18 ? n3354 : n4112;
  assign n4114 = pi17 ? n3353 : n4113;
  assign n4115 = pi16 ? n3351 : n4114;
  assign n4116 = pi21 ? n760 : n32;
  assign n4117 = pi20 ? n4116 : n32;
  assign n4118 = pi19 ? n4117 : n32;
  assign n4119 = pi18 ? n3365 : n4118;
  assign n4120 = pi17 ? n3363 : n4119;
  assign n4121 = pi16 ? n3360 : n4120;
  assign n4122 = pi15 ? n4115 : n4121;
  assign n4123 = pi14 ? n4108 : n4122;
  assign n4124 = pi13 ? n4088 : n4123;
  assign n4125 = pi12 ? n3985 : n4124;
  assign n4126 = pi11 ? n3904 : n4125;
  assign n4127 = pi18 ? n3380 : n4118;
  assign n4128 = pi17 ? n3378 : n4127;
  assign n4129 = pi16 ? n439 : n4128;
  assign n4130 = pi18 ? n3385 : n3342;
  assign n4131 = pi17 ? n2072 : n4130;
  assign n4132 = pi16 ? n439 : n4131;
  assign n4133 = pi15 ? n4129 : n4132;
  assign n4134 = pi18 ? n3395 : n3342;
  assign n4135 = pi17 ? n3391 : n4134;
  assign n4136 = pi16 ? n439 : n4135;
  assign n4137 = pi18 ? n3414 : n2581;
  assign n4138 = pi17 ? n3408 : n4137;
  assign n4139 = pi16 ? n439 : n4138;
  assign n4140 = pi15 ? n4136 : n4139;
  assign n4141 = pi14 ? n4133 : n4140;
  assign n4142 = pi18 ? n2102 : n2581;
  assign n4143 = pi17 ? n37 : n4142;
  assign n4144 = pi16 ? n439 : n4143;
  assign n4145 = pi24 ? n233 : n685;
  assign n4146 = pi23 ? n4145 : n32;
  assign n4147 = pi22 ? n4146 : n32;
  assign n4148 = pi21 ? n4147 : n32;
  assign n4149 = pi20 ? n4148 : n32;
  assign n4150 = pi19 ? n4149 : n32;
  assign n4151 = pi18 ? n3421 : n4150;
  assign n4152 = pi17 ? n37 : n4151;
  assign n4153 = pi16 ? n439 : n4152;
  assign n4154 = pi18 ? n2102 : n3400;
  assign n4155 = pi17 ? n37 : n4154;
  assign n4156 = pi16 ? n439 : n4155;
  assign n4157 = pi15 ? n4153 : n4156;
  assign n4158 = pi14 ? n4144 : n4157;
  assign n4159 = pi13 ? n4141 : n4158;
  assign n4160 = pi18 ? n2724 : n2703;
  assign n4161 = pi17 ? n37 : n4160;
  assign n4162 = pi16 ? n439 : n4161;
  assign n4163 = pi18 ? n2731 : n2703;
  assign n4164 = pi17 ? n37 : n4163;
  assign n4165 = pi16 ? n439 : n4164;
  assign n4166 = pi15 ? n4162 : n4165;
  assign n4167 = pi14 ? n2706 : n4166;
  assign n4168 = pi18 ? n3439 : n1824;
  assign n4169 = pi17 ? n99 : n4168;
  assign n4170 = pi16 ? n744 : n4169;
  assign n4171 = pi18 ? n3448 : n1824;
  assign n4172 = pi17 ? n99 : n4171;
  assign n4173 = pi16 ? n721 : n4172;
  assign n4174 = pi15 ? n4170 : n4173;
  assign n4175 = pi22 ? n3443 : n685;
  assign n4176 = pi21 ? n99 : n4175;
  assign n4177 = pi20 ? n99 : n4176;
  assign n4178 = pi19 ? n99 : n4177;
  assign n4179 = pi18 ? n4178 : n32;
  assign n4180 = pi17 ? n99 : n4179;
  assign n4181 = pi16 ? n1510 : n4180;
  assign n4182 = pi22 ? n158 : n1475;
  assign n4183 = pi21 ? n99 : n4182;
  assign n4184 = pi20 ? n99 : n4183;
  assign n4185 = pi19 ? n99 : n4184;
  assign n4186 = pi18 ? n4185 : n32;
  assign n4187 = pi17 ? n99 : n4186;
  assign n4188 = pi16 ? n801 : n4187;
  assign n4189 = pi15 ? n4181 : n4188;
  assign n4190 = pi14 ? n4174 : n4189;
  assign n4191 = pi13 ? n4167 : n4190;
  assign n4192 = pi12 ? n4159 : n4191;
  assign n4193 = pi22 ? n3443 : n1475;
  assign n4194 = pi21 ? n99 : n4193;
  assign n4195 = pi20 ? n99 : n4194;
  assign n4196 = pi19 ? n99 : n4195;
  assign n4197 = pi18 ? n4196 : n32;
  assign n4198 = pi17 ? n99 : n4197;
  assign n4199 = pi16 ? n721 : n4198;
  assign n4200 = pi16 ? n744 : n3478;
  assign n4201 = pi15 ? n4199 : n4200;
  assign n4202 = pi21 ? n1143 : n99;
  assign n4203 = pi20 ? n99 : n4202;
  assign n4204 = pi19 ? n99 : n4203;
  assign n4205 = pi18 ? n4204 : n99;
  assign n4206 = pi17 ? n4205 : n3488;
  assign n4207 = pi16 ? n744 : n4206;
  assign n4208 = pi22 ? n316 : n625;
  assign n4209 = pi21 ? n99 : n4208;
  assign n4210 = pi20 ? n787 : n4209;
  assign n4211 = pi19 ? n99 : n4210;
  assign n4212 = pi18 ? n4211 : n32;
  assign n4213 = pi17 ? n99 : n4212;
  assign n4214 = pi16 ? n744 : n4213;
  assign n4215 = pi15 ? n4207 : n4214;
  assign n4216 = pi14 ? n4201 : n4215;
  assign n4217 = pi22 ? n909 : n99;
  assign n4218 = pi21 ? n4217 : n825;
  assign n4219 = pi20 ? n32 : n4218;
  assign n4220 = pi19 ? n32 : n4219;
  assign n4221 = pi22 ? n99 : n812;
  assign n4222 = pi21 ? n4221 : n837;
  assign n4223 = pi22 ? n812 : n99;
  assign n4224 = pi21 ? n4223 : n837;
  assign n4225 = pi20 ? n4222 : n4224;
  assign n4226 = pi22 ? n812 : n295;
  assign n4227 = pi21 ? n4226 : n837;
  assign n4228 = pi22 ? n812 : n745;
  assign n4229 = pi21 ? n4228 : n4221;
  assign n4230 = pi20 ? n4227 : n4229;
  assign n4231 = pi19 ? n4225 : n4230;
  assign n4232 = pi18 ? n4220 : n4231;
  assign n4233 = pi17 ? n32 : n4232;
  assign n4234 = pi22 ? n812 : n139;
  assign n4235 = pi21 ? n825 : n4234;
  assign n4236 = pi22 ? n745 : n139;
  assign n4237 = pi22 ? n99 : n139;
  assign n4238 = pi21 ? n4236 : n4237;
  assign n4239 = pi20 ? n4235 : n4238;
  assign n4240 = pi21 ? n4237 : n823;
  assign n4241 = pi21 ? n823 : n837;
  assign n4242 = pi20 ? n4240 : n4241;
  assign n4243 = pi19 ? n4239 : n4242;
  assign n4244 = pi21 ? n825 : n4228;
  assign n4245 = pi21 ? n4234 : n823;
  assign n4246 = pi20 ? n4244 : n4245;
  assign n4247 = pi22 ? n139 : n99;
  assign n4248 = pi21 ? n4247 : n4228;
  assign n4249 = pi20 ? n4248 : n4245;
  assign n4250 = pi19 ? n4246 : n4249;
  assign n4251 = pi18 ? n4243 : n4250;
  assign n4252 = pi22 ? n139 : n812;
  assign n4253 = pi21 ? n4252 : n823;
  assign n4254 = pi21 ? n4236 : n3520;
  assign n4255 = pi20 ? n4253 : n4254;
  assign n4256 = pi21 ? n819 : n3494;
  assign n4257 = pi20 ? n157 : n4256;
  assign n4258 = pi19 ? n4255 : n4257;
  assign n4259 = pi18 ? n4258 : n32;
  assign n4260 = pi17 ? n4251 : n4259;
  assign n4261 = pi16 ? n4233 : n4260;
  assign n4262 = pi24 ? n32 : n157;
  assign n4263 = pi23 ? n4262 : n157;
  assign n4264 = pi22 ? n4263 : n861;
  assign n4265 = pi21 ? n4264 : n248;
  assign n4266 = pi20 ? n32 : n4265;
  assign n4267 = pi19 ? n32 : n4266;
  assign n4268 = pi22 ? n861 : n139;
  assign n4269 = pi22 ? n852 : n861;
  assign n4270 = pi21 ? n4268 : n4269;
  assign n4271 = pi21 ? n858 : n862;
  assign n4272 = pi20 ? n4270 : n4271;
  assign n4273 = pi21 ? n858 : n861;
  assign n4274 = pi21 ? n858 : n4268;
  assign n4275 = pi20 ? n4273 : n4274;
  assign n4276 = pi19 ? n4272 : n4275;
  assign n4277 = pi18 ? n4267 : n4276;
  assign n4278 = pi17 ? n32 : n4277;
  assign n4279 = pi22 ? n861 : n852;
  assign n4280 = pi21 ? n857 : n4279;
  assign n4281 = pi22 ? n157 : n861;
  assign n4282 = pi21 ? n4281 : n258;
  assign n4283 = pi20 ? n4280 : n4282;
  assign n4284 = pi21 ? n258 : n4281;
  assign n4285 = pi20 ? n4284 : n4269;
  assign n4286 = pi19 ? n4283 : n4285;
  assign n4287 = pi21 ? n248 : n4279;
  assign n4288 = pi21 ? n4279 : n4281;
  assign n4289 = pi20 ? n4287 : n4288;
  assign n4290 = pi20 ? n859 : n4288;
  assign n4291 = pi19 ? n4289 : n4290;
  assign n4292 = pi18 ? n4286 : n4291;
  assign n4293 = pi21 ? n857 : n4269;
  assign n4294 = pi21 ? n857 : n157;
  assign n4295 = pi20 ? n4293 : n4294;
  assign n4296 = pi22 ? n2244 : n688;
  assign n4297 = pi21 ? n157 : n4296;
  assign n4298 = pi20 ? n157 : n4297;
  assign n4299 = pi19 ? n4295 : n4298;
  assign n4300 = pi18 ? n4299 : n32;
  assign n4301 = pi17 ? n4292 : n4300;
  assign n4302 = pi16 ? n4278 : n4301;
  assign n4303 = pi15 ? n4261 : n4302;
  assign n4304 = pi23 ? n4262 : n139;
  assign n4305 = pi22 ? n4304 : n139;
  assign n4306 = pi21 ? n4305 : n858;
  assign n4307 = pi20 ? n32 : n4306;
  assign n4308 = pi19 ? n32 : n4307;
  assign n4309 = pi22 ? n889 : n861;
  assign n4310 = pi21 ? n139 : n4309;
  assign n4311 = pi20 ? n4310 : n4271;
  assign n4312 = pi21 ? n858 : n139;
  assign n4313 = pi21 ? n890 : n4268;
  assign n4314 = pi20 ? n4312 : n4313;
  assign n4315 = pi19 ? n4311 : n4314;
  assign n4316 = pi18 ? n4308 : n4315;
  assign n4317 = pi17 ? n32 : n4316;
  assign n4318 = pi21 ? n4269 : n258;
  assign n4319 = pi20 ? n4274 : n4318;
  assign n4320 = pi22 ? n852 : n893;
  assign n4321 = pi21 ? n258 : n4320;
  assign n4322 = pi21 ? n4320 : n4309;
  assign n4323 = pi20 ? n4321 : n4322;
  assign n4324 = pi19 ? n4319 : n4323;
  assign n4325 = pi22 ? n893 : n889;
  assign n4326 = pi21 ? n858 : n4325;
  assign n4327 = pi20 ? n4326 : n4270;
  assign n4328 = pi21 ? n248 : n890;
  assign n4329 = pi20 ? n4328 : n4270;
  assign n4330 = pi19 ? n4327 : n4329;
  assign n4331 = pi18 ? n4324 : n4330;
  assign n4332 = pi21 ? n248 : n4320;
  assign n4333 = pi20 ? n4332 : n4294;
  assign n4334 = pi19 ? n4333 : n3564;
  assign n4335 = pi18 ? n4334 : n32;
  assign n4336 = pi17 ? n4331 : n4335;
  assign n4337 = pi16 ? n4317 : n4336;
  assign n4338 = pi23 ? n3719 : n139;
  assign n4339 = pi22 ? n4338 : n139;
  assign n4340 = pi21 ? n4339 : n919;
  assign n4341 = pi20 ? n32 : n4340;
  assign n4342 = pi19 ? n32 : n4341;
  assign n4343 = pi22 ? n455 : n1038;
  assign n4344 = pi21 ? n139 : n4343;
  assign n4345 = pi21 ? n919 : n1793;
  assign n4346 = pi20 ? n4344 : n4345;
  assign n4347 = pi22 ? n139 : n455;
  assign n4348 = pi21 ? n4347 : n2869;
  assign n4349 = pi20 ? n920 : n4348;
  assign n4350 = pi19 ? n4346 : n4349;
  assign n4351 = pi18 ? n4342 : n4350;
  assign n4352 = pi17 ? n32 : n4351;
  assign n4353 = pi21 ? n1832 : n921;
  assign n4354 = pi20 ? n2870 : n4353;
  assign n4355 = pi21 ? n921 : n1832;
  assign n4356 = pi21 ? n457 : n4343;
  assign n4357 = pi20 ? n4355 : n4356;
  assign n4358 = pi19 ? n4354 : n4357;
  assign n4359 = pi21 ? n919 : n520;
  assign n4360 = pi21 ? n2869 : n2864;
  assign n4361 = pi20 ? n4359 : n4360;
  assign n4362 = pi21 ? n916 : n4347;
  assign n4363 = pi20 ? n4362 : n4360;
  assign n4364 = pi19 ? n4361 : n4363;
  assign n4365 = pi18 ? n4358 : n4364;
  assign n4366 = pi21 ? n916 : n1810;
  assign n4367 = pi20 ? n4366 : n2316;
  assign n4368 = pi19 ? n4367 : n3587;
  assign n4369 = pi18 ? n4368 : n32;
  assign n4370 = pi17 ? n4365 : n4369;
  assign n4371 = pi16 ? n4352 : n4370;
  assign n4372 = pi15 ? n4337 : n4371;
  assign n4373 = pi14 ? n4303 : n4372;
  assign n4374 = pi13 ? n4216 : n4373;
  assign n4375 = pi23 ? n3719 : n37;
  assign n4376 = pi22 ? n4375 : n139;
  assign n4377 = pi21 ? n4376 : n4347;
  assign n4378 = pi20 ? n32 : n4377;
  assign n4379 = pi19 ? n32 : n4378;
  assign n4380 = pi21 ? n3073 : n1793;
  assign n4381 = pi20 ? n4344 : n4380;
  assign n4382 = pi21 ? n4347 : n139;
  assign n4383 = pi22 ? n456 : n139;
  assign n4384 = pi21 ? n4347 : n4383;
  assign n4385 = pi20 ? n4382 : n4384;
  assign n4386 = pi19 ? n4381 : n4385;
  assign n4387 = pi18 ? n4379 : n4386;
  assign n4388 = pi17 ? n32 : n4387;
  assign n4389 = pi20 ? n4348 : n4353;
  assign n4390 = pi21 ? n921 : n457;
  assign n4391 = pi20 ? n4390 : n4356;
  assign n4392 = pi19 ? n4389 : n4391;
  assign n4393 = pi21 ? n4347 : n520;
  assign n4394 = pi21 ? n2869 : n4343;
  assign n4395 = pi20 ? n4393 : n4394;
  assign n4396 = pi20 ? n4362 : n4394;
  assign n4397 = pi19 ? n4395 : n4396;
  assign n4398 = pi18 ? n4392 : n4397;
  assign n4399 = pi19 ? n4367 : n3620;
  assign n4400 = pi18 ? n4399 : n32;
  assign n4401 = pi17 ? n4398 : n4400;
  assign n4402 = pi16 ? n4388 : n4401;
  assign n4403 = pi18 ? n1573 : n3627;
  assign n4404 = pi17 ? n32 : n4403;
  assign n4405 = pi16 ? n4404 : n3633;
  assign n4406 = pi15 ? n4402 : n4405;
  assign n4407 = pi22 ? n55 : n348;
  assign n4408 = pi21 ? n4407 : n1777;
  assign n4409 = pi20 ? n32 : n4408;
  assign n4410 = pi19 ? n32 : n4409;
  assign n4411 = pi21 ? n359 : n3617;
  assign n4412 = pi20 ? n4411 : n360;
  assign n4413 = pi21 ? n4014 : n139;
  assign n4414 = pi21 ? n1785 : n1774;
  assign n4415 = pi20 ? n4413 : n4414;
  assign n4416 = pi19 ? n4412 : n4415;
  assign n4417 = pi18 ? n4410 : n4416;
  assign n4418 = pi17 ? n32 : n4417;
  assign n4419 = pi22 ? n390 : n1784;
  assign n4420 = pi21 ? n139 : n4419;
  assign n4421 = pi22 ? n1784 : n348;
  assign n4422 = pi21 ? n349 : n4421;
  assign n4423 = pi20 ? n4420 : n4422;
  assign n4424 = pi22 ? n383 : n348;
  assign n4425 = pi21 ? n4421 : n4424;
  assign n4426 = pi21 ? n3617 : n356;
  assign n4427 = pi20 ? n4425 : n4426;
  assign n4428 = pi19 ? n4423 : n4427;
  assign n4429 = pi22 ? n348 : n1784;
  assign n4430 = pi21 ? n4014 : n4429;
  assign n4431 = pi21 ? n346 : n1774;
  assign n4432 = pi20 ? n4430 : n4431;
  assign n4433 = pi21 ? n3617 : n4429;
  assign n4434 = pi20 ? n4433 : n4431;
  assign n4435 = pi19 ? n4432 : n4434;
  assign n4436 = pi18 ? n4428 : n4435;
  assign n4437 = pi21 ? n356 : n316;
  assign n4438 = pi20 ? n4426 : n4437;
  assign n4439 = pi19 ? n4438 : n3661;
  assign n4440 = pi18 ? n4439 : n32;
  assign n4441 = pi17 ? n4436 : n4440;
  assign n4442 = pi16 ? n4418 : n4441;
  assign n4443 = pi15 ? n3640 : n4442;
  assign n4444 = pi14 ? n4406 : n4443;
  assign n4445 = pi22 ? n1784 : n37;
  assign n4446 = pi21 ? n359 : n4445;
  assign n4447 = pi22 ? n390 : n139;
  assign n4448 = pi21 ? n4447 : n139;
  assign n4449 = pi20 ? n4446 : n4448;
  assign n4450 = pi21 ? n4052 : n139;
  assign n4451 = pi22 ? n37 : n1784;
  assign n4452 = pi21 ? n4451 : n1774;
  assign n4453 = pi20 ? n4450 : n4452;
  assign n4454 = pi19 ? n4449 : n4453;
  assign n4455 = pi18 ? n4410 : n4454;
  assign n4456 = pi17 ? n32 : n4455;
  assign n4457 = pi21 ? n1774 : n3118;
  assign n4458 = pi20 ? n4420 : n4457;
  assign n4459 = pi21 ? n4445 : n356;
  assign n4460 = pi20 ? n3118 : n4459;
  assign n4461 = pi19 ? n4458 : n4460;
  assign n4462 = pi21 ? n4052 : n4419;
  assign n4463 = pi20 ? n4462 : n4431;
  assign n4464 = pi21 ? n3617 : n4419;
  assign n4465 = pi20 ? n4464 : n4431;
  assign n4466 = pi19 ? n4463 : n4465;
  assign n4467 = pi18 ? n4461 : n4466;
  assign n4468 = pi19 ? n4438 : n3685;
  assign n4469 = pi18 ? n4468 : n32;
  assign n4470 = pi17 ? n4467 : n4469;
  assign n4471 = pi16 ? n4456 : n4470;
  assign n4472 = pi22 ? n55 : n316;
  assign n4473 = pi21 ? n4472 : n3693;
  assign n4474 = pi20 ? n32 : n4473;
  assign n4475 = pi19 ? n32 : n4474;
  assign n4476 = pi18 ? n4475 : n3704;
  assign n4477 = pi17 ? n32 : n4476;
  assign n4478 = pi21 ? n316 : n417;
  assign n4479 = pi20 ? n4478 : n2330;
  assign n4480 = pi19 ? n316 : n4479;
  assign n4481 = pi18 ? n4480 : n32;
  assign n4482 = pi17 ? n3710 : n4481;
  assign n4483 = pi16 ? n4477 : n4482;
  assign n4484 = pi15 ? n4471 : n4483;
  assign n4485 = pi22 ? n715 : n204;
  assign n4486 = pi21 ? n4485 : n1027;
  assign n4487 = pi20 ? n32 : n4486;
  assign n4488 = pi19 ? n32 : n4487;
  assign n4489 = pi18 ? n4488 : n204;
  assign n4490 = pi17 ? n32 : n4489;
  assign n4491 = pi16 ? n4490 : n3741;
  assign n4492 = pi21 ? n4485 : n1079;
  assign n4493 = pi20 ? n32 : n4492;
  assign n4494 = pi19 ? n32 : n4493;
  assign n4495 = pi18 ? n4494 : n3750;
  assign n4496 = pi17 ? n32 : n4495;
  assign n4497 = pi21 ? n3763 : n928;
  assign n4498 = pi20 ? n204 : n4497;
  assign n4499 = pi19 ? n3761 : n4498;
  assign n4500 = pi18 ? n4499 : n32;
  assign n4501 = pi17 ? n3758 : n4500;
  assign n4502 = pi16 ? n4496 : n4501;
  assign n4503 = pi15 ? n4491 : n4502;
  assign n4504 = pi14 ? n4484 : n4503;
  assign n4505 = pi13 ? n4444 : n4504;
  assign n4506 = pi12 ? n4374 : n4505;
  assign n4507 = pi11 ? n4192 : n4506;
  assign n4508 = pi10 ? n4126 : n4507;
  assign n4509 = pi09 ? n32 : n4508;
  assign n4510 = pi08 ? n3776 : n4509;
  assign n4511 = pi07 ? n2932 : n4510;
  assign n4512 = pi16 ? n2447 : n3796;
  assign n4513 = pi15 ? n32 : n4512;
  assign n4514 = pi16 ? n3784 : n3796;
  assign n4515 = pi16 ? n70 : n3796;
  assign n4516 = pi15 ? n4514 : n4515;
  assign n4517 = pi14 ? n4513 : n4516;
  assign n4518 = pi16 ? n73 : n3796;
  assign n4519 = pi22 ? n37 : n32;
  assign n4520 = pi21 ? n4519 : n32;
  assign n4521 = pi20 ? n4520 : n32;
  assign n4522 = pi19 ? n4521 : n32;
  assign n4523 = pi18 ? n37 : n4522;
  assign n4524 = pi17 ? n37 : n4523;
  assign n4525 = pi16 ? n83 : n4524;
  assign n4526 = pi15 ? n4518 : n4525;
  assign n4527 = pi16 ? n1130 : n4524;
  assign n4528 = pi21 ? n48 : n32;
  assign n4529 = pi20 ? n4528 : n32;
  assign n4530 = pi19 ? n4529 : n32;
  assign n4531 = pi18 ? n37 : n4530;
  assign n4532 = pi17 ? n37 : n4531;
  assign n4533 = pi16 ? n2461 : n4532;
  assign n4534 = pi15 ? n4527 : n4533;
  assign n4535 = pi14 ? n4526 : n4534;
  assign n4536 = pi13 ? n4517 : n4535;
  assign n4537 = pi23 ? n99 : n363;
  assign n4538 = pi22 ? n4537 : n99;
  assign n4539 = pi21 ? n4538 : n99;
  assign n4540 = pi19 ? n4539 : n99;
  assign n4541 = pi18 ? n184 : n4540;
  assign n4542 = pi17 ? n32 : n4541;
  assign n4543 = pi23 ? n363 : n99;
  assign n4544 = pi21 ? n4538 : n4543;
  assign n4545 = pi20 ? n99 : n4544;
  assign n4546 = pi19 ? n99 : n4545;
  assign n4547 = pi21 ? n99 : n4543;
  assign n4548 = pi22 ? n99 : n4537;
  assign n4549 = pi21 ? n99 : n4548;
  assign n4550 = pi20 ? n4547 : n4549;
  assign n4551 = pi22 ? n99 : n4543;
  assign n4552 = pi21 ? n4538 : n4551;
  assign n4553 = pi20 ? n4544 : n4552;
  assign n4554 = pi19 ? n4550 : n4553;
  assign n4555 = pi18 ? n4546 : n4554;
  assign n4556 = pi20 ? n4552 : n4539;
  assign n4557 = pi20 ? n4549 : n99;
  assign n4558 = pi19 ? n4556 : n4557;
  assign n4559 = pi22 ? n99 : n32;
  assign n4560 = pi21 ? n4559 : n32;
  assign n4561 = pi20 ? n4560 : n32;
  assign n4562 = pi19 ? n4561 : n32;
  assign n4563 = pi18 ? n4558 : n4562;
  assign n4564 = pi17 ? n4555 : n4563;
  assign n4565 = pi16 ? n4542 : n4564;
  assign n4566 = pi21 ? n104 : n32;
  assign n4567 = pi20 ? n4566 : n32;
  assign n4568 = pi19 ? n4567 : n32;
  assign n4569 = pi18 ? n99 : n4568;
  assign n4570 = pi17 ? n99 : n4569;
  assign n4571 = pi16 ? n1148 : n4570;
  assign n4572 = pi15 ? n4565 : n4571;
  assign n4573 = pi16 ? n744 : n4570;
  assign n4574 = pi14 ? n4572 : n4573;
  assign n4575 = pi22 ? n99 : n261;
  assign n4576 = pi21 ? n4575 : n32;
  assign n4577 = pi20 ? n4576 : n32;
  assign n4578 = pi19 ? n4577 : n32;
  assign n4579 = pi18 ? n99 : n4578;
  assign n4580 = pi17 ? n99 : n4579;
  assign n4581 = pi16 ? n801 : n4580;
  assign n4582 = pi19 ? n99 : n3050;
  assign n4583 = pi20 ? n99 : n219;
  assign n4584 = pi19 ? n4583 : n99;
  assign n4585 = pi18 ? n4582 : n4584;
  assign n4586 = pi19 ? n4583 : n226;
  assign n4587 = pi22 ? n99 : n587;
  assign n4588 = pi21 ? n4587 : n32;
  assign n4589 = pi20 ? n4588 : n32;
  assign n4590 = pi19 ? n4589 : n32;
  assign n4591 = pi18 ? n4586 : n4590;
  assign n4592 = pi17 ? n4585 : n4591;
  assign n4593 = pi16 ? n801 : n4592;
  assign n4594 = pi15 ? n4581 : n4593;
  assign n4595 = pi18 ? n99 : n4562;
  assign n4596 = pi17 ? n99 : n4595;
  assign n4597 = pi16 ? n721 : n4596;
  assign n4598 = pi19 ? n99 : n167;
  assign n4599 = pi20 ? n166 : n99;
  assign n4600 = pi19 ? n4599 : n4203;
  assign n4601 = pi18 ? n4598 : n4600;
  assign n4602 = pi21 ? n1143 : n165;
  assign n4603 = pi20 ? n4602 : n169;
  assign n4604 = pi20 ? n1665 : n99;
  assign n4605 = pi19 ? n4603 : n4604;
  assign n4606 = pi18 ? n4605 : n4562;
  assign n4607 = pi17 ? n4601 : n4606;
  assign n4608 = pi16 ? n2488 : n4607;
  assign n4609 = pi15 ? n4597 : n4608;
  assign n4610 = pi14 ? n4594 : n4609;
  assign n4611 = pi13 ? n4574 : n4610;
  assign n4612 = pi12 ? n4536 : n4611;
  assign n4613 = pi21 ? n1179 : n2164;
  assign n4614 = pi20 ? n32 : n4613;
  assign n4615 = pi19 ? n32 : n4614;
  assign n4616 = pi21 ? n2746 : n2164;
  assign n4617 = pi21 ? n2746 : n99;
  assign n4618 = pi20 ? n4616 : n4617;
  assign n4619 = pi21 ? n2164 : n2746;
  assign n4620 = pi20 ? n3506 : n4619;
  assign n4621 = pi19 ? n4618 : n4620;
  assign n4622 = pi18 ? n4615 : n4621;
  assign n4623 = pi17 ? n32 : n4622;
  assign n4624 = pi20 ? n2191 : n3807;
  assign n4625 = pi21 ? n99 : n2164;
  assign n4626 = pi20 ? n4625 : n4617;
  assign n4627 = pi19 ? n4624 : n4626;
  assign n4628 = pi20 ? n4617 : n4625;
  assign n4629 = pi20 ? n4617 : n2189;
  assign n4630 = pi19 ? n4628 : n4629;
  assign n4631 = pi18 ? n4627 : n4630;
  assign n4632 = pi20 ? n2174 : n99;
  assign n4633 = pi19 ? n4632 : n2191;
  assign n4634 = pi18 ? n4633 : n4562;
  assign n4635 = pi17 ? n4631 : n4634;
  assign n4636 = pi16 ? n4623 : n4635;
  assign n4637 = pi22 ? n962 : n37;
  assign n4638 = pi22 ? n157 : n852;
  assign n4639 = pi21 ? n4637 : n4638;
  assign n4640 = pi20 ? n32 : n4639;
  assign n4641 = pi19 ? n32 : n4640;
  assign n4642 = pi22 ? n893 : n861;
  assign n4643 = pi21 ? n4642 : n248;
  assign n4644 = pi21 ? n4320 : n4268;
  assign n4645 = pi21 ? n4638 : n4642;
  assign n4646 = pi20 ? n4644 : n4645;
  assign n4647 = pi19 ? n4643 : n4646;
  assign n4648 = pi18 ? n4641 : n4647;
  assign n4649 = pi17 ? n32 : n4648;
  assign n4650 = pi21 ? n4268 : n4638;
  assign n4651 = pi20 ? n4332 : n4650;
  assign n4652 = pi22 ? n893 : n139;
  assign n4653 = pi21 ? n4652 : n4638;
  assign n4654 = pi21 ? n4642 : n157;
  assign n4655 = pi20 ? n4653 : n4654;
  assign n4656 = pi19 ? n4651 : n4655;
  assign n4657 = pi21 ? n139 : n4638;
  assign n4658 = pi20 ? n4654 : n4657;
  assign n4659 = pi21 ? n4281 : n248;
  assign n4660 = pi20 ? n4643 : n4659;
  assign n4661 = pi19 ? n4658 : n4660;
  assign n4662 = pi18 ? n4656 : n4661;
  assign n4663 = pi21 ? n4281 : n157;
  assign n4664 = pi20 ? n4663 : n258;
  assign n4665 = pi21 ? n248 : n857;
  assign n4666 = pi21 ? n248 : n853;
  assign n4667 = pi20 ? n4665 : n4666;
  assign n4668 = pi19 ? n4664 : n4667;
  assign n4669 = pi22 ? n139 : n2468;
  assign n4670 = pi21 ? n4669 : n32;
  assign n4671 = pi20 ? n4670 : n32;
  assign n4672 = pi19 ? n4671 : n32;
  assign n4673 = pi18 ? n4668 : n4672;
  assign n4674 = pi17 ? n4662 : n4673;
  assign n4675 = pi16 ? n4649 : n4674;
  assign n4676 = pi15 ? n4636 : n4675;
  assign n4677 = pi22 ? n204 : n852;
  assign n4678 = pi21 ? n1564 : n4677;
  assign n4679 = pi20 ? n32 : n4678;
  assign n4680 = pi19 ? n32 : n4679;
  assign n4681 = pi21 ? n4642 : n916;
  assign n4682 = pi21 ? n4677 : n4642;
  assign n4683 = pi20 ? n4644 : n4682;
  assign n4684 = pi19 ? n4681 : n4683;
  assign n4685 = pi18 ? n4680 : n4684;
  assign n4686 = pi17 ? n32 : n4685;
  assign n4687 = pi21 ? n916 : n4320;
  assign n4688 = pi21 ? n4268 : n4677;
  assign n4689 = pi20 ? n4687 : n4688;
  assign n4690 = pi21 ? n4652 : n4677;
  assign n4691 = pi21 ? n4642 : n139;
  assign n4692 = pi20 ? n4690 : n4691;
  assign n4693 = pi19 ? n4689 : n4692;
  assign n4694 = pi21 ? n139 : n4677;
  assign n4695 = pi20 ? n4691 : n4694;
  assign n4696 = pi21 ? n862 : n916;
  assign n4697 = pi20 ? n4681 : n4696;
  assign n4698 = pi19 ? n4695 : n4697;
  assign n4699 = pi18 ? n4693 : n4698;
  assign n4700 = pi20 ? n4696 : n139;
  assign n4701 = pi21 ? n916 : n853;
  assign n4702 = pi19 ? n4700 : n4701;
  assign n4703 = pi18 ? n4702 : n4672;
  assign n4704 = pi17 ? n4699 : n4703;
  assign n4705 = pi16 ? n4686 : n4704;
  assign n4706 = pi21 ? n180 : n919;
  assign n4707 = pi20 ? n32 : n4706;
  assign n4708 = pi19 ? n32 : n4707;
  assign n4709 = pi22 ? n456 : n1038;
  assign n4710 = pi21 ? n4709 : n916;
  assign n4711 = pi21 ? n1832 : n2869;
  assign n4712 = pi22 ? n204 : n918;
  assign n4713 = pi21 ? n4712 : n4709;
  assign n4714 = pi20 ? n4711 : n4713;
  assign n4715 = pi19 ? n4710 : n4714;
  assign n4716 = pi18 ? n4708 : n4715;
  assign n4717 = pi17 ? n32 : n4716;
  assign n4718 = pi21 ? n916 : n1832;
  assign n4719 = pi21 ? n2869 : n4712;
  assign n4720 = pi20 ? n4718 : n4719;
  assign n4721 = pi21 ? n1834 : n139;
  assign n4722 = pi21 ? n4709 : n139;
  assign n4723 = pi20 ? n4721 : n4722;
  assign n4724 = pi19 ? n4720 : n4723;
  assign n4725 = pi22 ? n295 : n1038;
  assign n4726 = pi21 ? n4725 : n139;
  assign n4727 = pi21 ? n1711 : n919;
  assign n4728 = pi20 ? n4726 : n4727;
  assign n4729 = pi21 ? n1721 : n916;
  assign n4730 = pi20 ? n4710 : n4729;
  assign n4731 = pi19 ? n4728 : n4730;
  assign n4732 = pi18 ? n4724 : n4731;
  assign n4733 = pi20 ? n3625 : n139;
  assign n4734 = pi21 ? n1211 : n2863;
  assign n4735 = pi19 ? n4733 : n4734;
  assign n4736 = pi22 ? n139 : n532;
  assign n4737 = pi21 ? n4736 : n32;
  assign n4738 = pi20 ? n4737 : n32;
  assign n4739 = pi19 ? n4738 : n32;
  assign n4740 = pi18 ? n4735 : n4739;
  assign n4741 = pi17 ? n4732 : n4740;
  assign n4742 = pi16 ? n4717 : n4741;
  assign n4743 = pi15 ? n4705 : n4742;
  assign n4744 = pi14 ? n4676 : n4743;
  assign n4745 = pi18 ? n139 : n4739;
  assign n4746 = pi17 ? n139 : n4745;
  assign n4747 = pi16 ? n314 : n4746;
  assign n4748 = pi22 ? n204 : n532;
  assign n4749 = pi21 ? n4748 : n32;
  assign n4750 = pi20 ? n4749 : n32;
  assign n4751 = pi19 ? n4750 : n32;
  assign n4752 = pi18 ? n139 : n4751;
  assign n4753 = pi17 ? n139 : n4752;
  assign n4754 = pi16 ? n1773 : n4753;
  assign n4755 = pi15 ? n4747 : n4754;
  assign n4756 = pi22 ? n335 : n532;
  assign n4757 = pi21 ? n4756 : n32;
  assign n4758 = pi20 ? n4757 : n32;
  assign n4759 = pi19 ? n4758 : n32;
  assign n4760 = pi18 ? n139 : n4759;
  assign n4761 = pi17 ? n139 : n4760;
  assign n4762 = pi16 ? n1773 : n4761;
  assign n4763 = pi21 ? n180 : n346;
  assign n4764 = pi20 ? n32 : n4763;
  assign n4765 = pi19 ? n32 : n4764;
  assign n4766 = pi21 ? n356 : n346;
  assign n4767 = pi21 ? n1785 : n139;
  assign n4768 = pi21 ? n356 : n3617;
  assign n4769 = pi20 ? n4767 : n4768;
  assign n4770 = pi19 ? n4766 : n4769;
  assign n4771 = pi18 ? n4765 : n4770;
  assign n4772 = pi17 ? n32 : n4771;
  assign n4773 = pi21 ? n346 : n1785;
  assign n4774 = pi20 ? n4773 : n1008;
  assign n4775 = pi21 ? n3617 : n346;
  assign n4776 = pi20 ? n4775 : n316;
  assign n4777 = pi19 ? n4774 : n4776;
  assign n4778 = pi21 ? n2319 : n316;
  assign n4779 = pi20 ? n4778 : n4437;
  assign n4780 = pi22 ? n316 : n1784;
  assign n4781 = pi21 ? n4780 : n316;
  assign n4782 = pi20 ? n316 : n4781;
  assign n4783 = pi19 ? n4779 : n4782;
  assign n4784 = pi18 ? n4777 : n4783;
  assign n4785 = pi20 ? n4781 : n316;
  assign n4786 = pi20 ? n346 : n4773;
  assign n4787 = pi19 ? n4785 : n4786;
  assign n4788 = pi22 ? n316 : n532;
  assign n4789 = pi21 ? n4788 : n32;
  assign n4790 = pi20 ? n4789 : n32;
  assign n4791 = pi19 ? n4790 : n32;
  assign n4792 = pi18 ? n4787 : n4791;
  assign n4793 = pi17 ? n4784 : n4792;
  assign n4794 = pi16 ? n4772 : n4793;
  assign n4795 = pi15 ? n4762 : n4794;
  assign n4796 = pi14 ? n4755 : n4795;
  assign n4797 = pi13 ? n4744 : n4796;
  assign n4798 = pi20 ? n440 : n3256;
  assign n4799 = pi19 ? n4798 : n3261;
  assign n4800 = pi18 ? n3254 : n4799;
  assign n4801 = pi17 ? n32 : n4800;
  assign n4802 = pi20 ? n382 : n3255;
  assign n4803 = pi19 ? n3266 : n4802;
  assign n4804 = pi21 ? n3258 : n381;
  assign n4805 = pi20 ? n3255 : n4804;
  assign n4806 = pi20 ? n440 : n3275;
  assign n4807 = pi19 ? n4805 : n4806;
  assign n4808 = pi18 ? n4803 : n4807;
  assign n4809 = pi21 ? n392 : n316;
  assign n4810 = pi20 ? n4809 : n316;
  assign n4811 = pi20 ? n389 : n3265;
  assign n4812 = pi19 ? n4810 : n4811;
  assign n4813 = pi18 ? n4812 : n4791;
  assign n4814 = pi17 ? n4808 : n4813;
  assign n4815 = pi16 ? n4801 : n4814;
  assign n4816 = pi20 ? n382 : n37;
  assign n4817 = pi19 ? n4816 : n37;
  assign n4818 = pi18 ? n37 : n4817;
  assign n4819 = pi20 ? n382 : n3265;
  assign n4820 = pi19 ? n4819 : n3265;
  assign n4821 = pi18 ? n4820 : n4791;
  assign n4822 = pi17 ? n4818 : n4821;
  assign n4823 = pi16 ? n439 : n4822;
  assign n4824 = pi15 ? n4815 : n4823;
  assign n4825 = pi21 ? n180 : n392;
  assign n4826 = pi20 ? n32 : n4825;
  assign n4827 = pi19 ? n32 : n4826;
  assign n4828 = pi21 ? n384 : n4052;
  assign n4829 = pi21 ? n384 : n390;
  assign n4830 = pi20 ? n4828 : n4829;
  assign n4831 = pi21 ? n383 : n391;
  assign n4832 = pi20 ? n4831 : n4054;
  assign n4833 = pi19 ? n4830 : n4832;
  assign n4834 = pi18 ? n4827 : n4833;
  assign n4835 = pi17 ? n32 : n4834;
  assign n4836 = pi21 ? n390 : n383;
  assign n4837 = pi21 ? n391 : n4052;
  assign n4838 = pi20 ? n4836 : n4837;
  assign n4839 = pi21 ? n384 : n424;
  assign n4840 = pi20 ? n426 : n4839;
  assign n4841 = pi19 ? n4838 : n4840;
  assign n4842 = pi21 ? n3118 : n4052;
  assign n4843 = pi20 ? n4839 : n4842;
  assign n4844 = pi19 ? n4843 : n4829;
  assign n4845 = pi18 ? n4841 : n4844;
  assign n4846 = pi21 ? n3118 : n392;
  assign n4847 = pi20 ? n426 : n4846;
  assign n4848 = pi19 ? n4847 : n4836;
  assign n4849 = pi18 ? n4848 : n4791;
  assign n4850 = pi17 ? n4845 : n4849;
  assign n4851 = pi16 ? n4835 : n4850;
  assign n4852 = pi21 ? n650 : n32;
  assign n4853 = pi20 ? n4852 : n32;
  assign n4854 = pi19 ? n4853 : n32;
  assign n4855 = pi18 ? n37 : n4854;
  assign n4856 = pi17 ? n37 : n4855;
  assign n4857 = pi16 ? n439 : n4856;
  assign n4858 = pi15 ? n4851 : n4857;
  assign n4859 = pi14 ? n4824 : n4858;
  assign n4860 = pi21 ? n180 : n457;
  assign n4861 = pi20 ? n32 : n4860;
  assign n4862 = pi19 ? n32 : n4861;
  assign n4863 = pi20 ? n1897 : n508;
  assign n4864 = pi21 ? n204 : n1056;
  assign n4865 = pi20 ? n4864 : n1063;
  assign n4866 = pi19 ? n4863 : n4865;
  assign n4867 = pi18 ? n4862 : n4866;
  assign n4868 = pi17 ? n32 : n4867;
  assign n4869 = pi20 ? n204 : n1057;
  assign n4870 = pi21 ? n1083 : n516;
  assign n4871 = pi20 ? n1582 : n4870;
  assign n4872 = pi19 ? n4869 : n4871;
  assign n4873 = pi20 ? n4870 : n204;
  assign n4874 = pi21 ? n485 : n204;
  assign n4875 = pi20 ? n1099 : n4874;
  assign n4876 = pi19 ? n4873 : n4875;
  assign n4877 = pi18 ? n4872 : n4876;
  assign n4878 = pi21 ? n1578 : n204;
  assign n4879 = pi20 ? n4874 : n4878;
  assign n4880 = pi21 ? n204 : n522;
  assign n4881 = pi19 ? n4879 : n4880;
  assign n4882 = pi24 ? n204 : n233;
  assign n4883 = pi23 ? n204 : n4882;
  assign n4884 = pi22 ? n4883 : n688;
  assign n4885 = pi21 ? n4884 : n32;
  assign n4886 = pi20 ? n4885 : n32;
  assign n4887 = pi19 ? n4886 : n32;
  assign n4888 = pi18 ? n4881 : n4887;
  assign n4889 = pi17 ? n4877 : n4888;
  assign n4890 = pi16 ? n4868 : n4889;
  assign n4891 = pi22 ? n37 : n2116;
  assign n4892 = pi21 ? n559 : n4891;
  assign n4893 = pi22 ? n559 : n335;
  assign n4894 = pi21 ? n2117 : n4893;
  assign n4895 = pi20 ? n4892 : n4894;
  assign n4896 = pi19 ? n37 : n4895;
  assign n4897 = pi18 ? n374 : n4896;
  assign n4898 = pi17 ? n32 : n4897;
  assign n4899 = pi23 ? n233 : n335;
  assign n4900 = pi22 ? n233 : n2060;
  assign n4901 = pi21 ? n4899 : n4900;
  assign n4902 = pi22 ? n335 : n4899;
  assign n4903 = pi22 ? n4899 : n233;
  assign n4904 = pi21 ? n4902 : n4903;
  assign n4905 = pi20 ? n4901 : n4904;
  assign n4906 = pi22 ? n2060 : n37;
  assign n4907 = pi21 ? n4906 : n4903;
  assign n4908 = pi22 ? n2060 : n335;
  assign n4909 = pi21 ? n4908 : n3409;
  assign n4910 = pi20 ? n4907 : n4909;
  assign n4911 = pi19 ? n4905 : n4910;
  assign n4912 = pi22 ? n233 : n4899;
  assign n4913 = pi21 ? n4912 : n4903;
  assign n4914 = pi20 ? n4909 : n4913;
  assign n4915 = pi21 ? n4908 : n4903;
  assign n4916 = pi21 ? n4893 : n4903;
  assign n4917 = pi20 ? n4915 : n4916;
  assign n4918 = pi19 ? n4914 : n4917;
  assign n4919 = pi18 ? n4911 : n4918;
  assign n4920 = pi22 ? n559 : n233;
  assign n4921 = pi21 ? n4920 : n233;
  assign n4922 = pi20 ? n4916 : n4921;
  assign n4923 = pi21 ? n4899 : n3411;
  assign n4924 = pi19 ? n4922 : n4923;
  assign n4925 = pi23 ? n233 : n4145;
  assign n4926 = pi22 ? n4925 : n706;
  assign n4927 = pi21 ? n4926 : n32;
  assign n4928 = pi20 ? n4927 : n32;
  assign n4929 = pi19 ? n4928 : n32;
  assign n4930 = pi18 ? n4924 : n4929;
  assign n4931 = pi17 ? n4919 : n4930;
  assign n4932 = pi16 ? n4898 : n4931;
  assign n4933 = pi15 ? n4890 : n4932;
  assign n4934 = pi20 ? n3299 : n2004;
  assign n4935 = pi19 ? n37 : n4934;
  assign n4936 = pi18 ? n374 : n4935;
  assign n4937 = pi17 ? n32 : n4936;
  assign n4938 = pi22 ? n583 : n335;
  assign n4939 = pi21 ? n4938 : n335;
  assign n4940 = pi20 ? n4939 : n335;
  assign n4941 = pi19 ? n4940 : n335;
  assign n4942 = pi18 ? n4941 : n335;
  assign n4943 = pi23 ? n335 : n4145;
  assign n4944 = pi22 ? n4943 : n32;
  assign n4945 = pi21 ? n4944 : n32;
  assign n4946 = pi20 ? n4945 : n32;
  assign n4947 = pi19 ? n4946 : n32;
  assign n4948 = pi18 ? n335 : n4947;
  assign n4949 = pi17 ? n4942 : n4948;
  assign n4950 = pi16 ? n4937 : n4949;
  assign n4951 = pi21 ? n2007 : n566;
  assign n4952 = pi21 ? n583 : n569;
  assign n4953 = pi20 ? n4951 : n4952;
  assign n4954 = pi21 ? n1943 : n569;
  assign n4955 = pi20 ? n4954 : n335;
  assign n4956 = pi19 ? n4953 : n4955;
  assign n4957 = pi18 ? n4956 : n335;
  assign n4958 = pi23 ? n335 : n2766;
  assign n4959 = pi22 ? n4958 : n32;
  assign n4960 = pi21 ? n4959 : n32;
  assign n4961 = pi20 ? n4960 : n32;
  assign n4962 = pi19 ? n4961 : n32;
  assign n4963 = pi18 ? n335 : n4962;
  assign n4964 = pi17 ? n4957 : n4963;
  assign n4965 = pi16 ? n439 : n4964;
  assign n4966 = pi15 ? n4950 : n4965;
  assign n4967 = pi14 ? n4933 : n4966;
  assign n4968 = pi13 ? n4859 : n4967;
  assign n4969 = pi12 ? n4797 : n4968;
  assign n4970 = pi11 ? n4612 : n4969;
  assign n4971 = pi21 ? n37 : n580;
  assign n4972 = pi20 ? n37 : n4971;
  assign n4973 = pi22 ? n566 : n583;
  assign n4974 = pi21 ? n4973 : n580;
  assign n4975 = pi22 ? n583 : n566;
  assign n4976 = pi21 ? n4973 : n4975;
  assign n4977 = pi20 ? n4974 : n4976;
  assign n4978 = pi19 ? n4972 : n4977;
  assign n4979 = pi20 ? n4976 : n2025;
  assign n4980 = pi21 ? n567 : n4938;
  assign n4981 = pi20 ? n4980 : n335;
  assign n4982 = pi19 ? n4979 : n4981;
  assign n4983 = pi18 ? n4978 : n4982;
  assign n4984 = pi20 ? n605 : n335;
  assign n4985 = pi19 ? n4984 : n335;
  assign n4986 = pi18 ? n4985 : n4962;
  assign n4987 = pi17 ? n4983 : n4986;
  assign n4988 = pi16 ? n439 : n4987;
  assign n4989 = pi21 ? n37 : n4975;
  assign n4990 = pi22 ? n335 : n566;
  assign n4991 = pi21 ? n335 : n4990;
  assign n4992 = pi20 ? n4989 : n4991;
  assign n4993 = pi19 ? n37 : n4992;
  assign n4994 = pi18 ? n37 : n4993;
  assign n4995 = pi21 ? n233 : n580;
  assign n4996 = pi21 ? n1943 : n567;
  assign n4997 = pi20 ? n4995 : n4996;
  assign n4998 = pi22 ? n566 : n233;
  assign n4999 = pi21 ? n570 : n4998;
  assign n5000 = pi21 ? n335 : n4998;
  assign n5001 = pi20 ? n4999 : n5000;
  assign n5002 = pi19 ? n4997 : n5001;
  assign n5003 = pi22 ? n1333 : n32;
  assign n5004 = pi21 ? n5003 : n32;
  assign n5005 = pi20 ? n5004 : n32;
  assign n5006 = pi19 ? n5005 : n32;
  assign n5007 = pi18 ? n5002 : n5006;
  assign n5008 = pi17 ? n4994 : n5007;
  assign n5009 = pi16 ? n439 : n5008;
  assign n5010 = pi15 ? n4988 : n5009;
  assign n5011 = pi23 ? n37 : n363;
  assign n5012 = pi22 ? n5011 : n37;
  assign n5013 = pi21 ? n37 : n5012;
  assign n5014 = pi22 ? n233 : n363;
  assign n5015 = pi22 ? n363 : n37;
  assign n5016 = pi21 ? n5014 : n5015;
  assign n5017 = pi20 ? n5013 : n5016;
  assign n5018 = pi19 ? n37 : n5017;
  assign n5019 = pi18 ? n37 : n5018;
  assign n5020 = pi21 ? n5014 : n233;
  assign n5021 = pi21 ? n2707 : n5014;
  assign n5022 = pi20 ? n5020 : n5021;
  assign n5023 = pi21 ? n2048 : n233;
  assign n5024 = pi20 ? n5023 : n233;
  assign n5025 = pi19 ? n5022 : n5024;
  assign n5026 = pi18 ? n5025 : n3342;
  assign n5027 = pi17 ? n5019 : n5026;
  assign n5028 = pi16 ? n439 : n5027;
  assign n5029 = pi20 ? n37 : n3393;
  assign n5030 = pi19 ? n37 : n5029;
  assign n5031 = pi18 ? n5030 : n2581;
  assign n5032 = pi17 ? n37 : n5031;
  assign n5033 = pi16 ? n439 : n5032;
  assign n5034 = pi15 ? n5028 : n5033;
  assign n5035 = pi14 ? n5010 : n5034;
  assign n5036 = pi20 ? n1921 : n2094;
  assign n5037 = pi19 ? n37 : n5036;
  assign n5038 = pi18 ? n5037 : n2581;
  assign n5039 = pi17 ? n37 : n5038;
  assign n5040 = pi16 ? n439 : n5039;
  assign n5041 = pi18 ? n2102 : n4112;
  assign n5042 = pi17 ? n37 : n5041;
  assign n5043 = pi16 ? n439 : n5042;
  assign n5044 = pi15 ? n5040 : n5043;
  assign n5045 = pi18 ? n2102 : n2640;
  assign n5046 = pi17 ? n37 : n5045;
  assign n5047 = pi16 ? n439 : n5046;
  assign n5048 = pi18 ? n2109 : n2640;
  assign n5049 = pi17 ? n37 : n5048;
  assign n5050 = pi16 ? n439 : n5049;
  assign n5051 = pi15 ? n5047 : n5050;
  assign n5052 = pi14 ? n5044 : n5051;
  assign n5053 = pi13 ? n5035 : n5052;
  assign n5054 = pi22 ? n363 : n157;
  assign n5055 = pi21 ? n37 : n5054;
  assign n5056 = pi20 ? n37 : n5055;
  assign n5057 = pi19 ? n37 : n5056;
  assign n5058 = pi18 ? n5057 : n2681;
  assign n5059 = pi17 ? n37 : n5058;
  assign n5060 = pi16 ? n439 : n5059;
  assign n5061 = pi23 ? n363 : n204;
  assign n5062 = pi22 ? n363 : n5061;
  assign n5063 = pi21 ? n37 : n5062;
  assign n5064 = pi20 ? n37 : n5063;
  assign n5065 = pi19 ? n37 : n5064;
  assign n5066 = pi18 ? n5065 : n2655;
  assign n5067 = pi17 ? n37 : n5066;
  assign n5068 = pi16 ? n439 : n5067;
  assign n5069 = pi15 ? n5060 : n5068;
  assign n5070 = pi22 ? n37 : n5061;
  assign n5071 = pi21 ? n37 : n5070;
  assign n5072 = pi20 ? n37 : n5071;
  assign n5073 = pi19 ? n37 : n5072;
  assign n5074 = pi18 ? n5073 : n2703;
  assign n5075 = pi17 ? n37 : n5074;
  assign n5076 = pi16 ? n439 : n5075;
  assign n5077 = pi21 ? n37 : n181;
  assign n5078 = pi20 ? n5077 : n2722;
  assign n5079 = pi19 ? n37 : n5078;
  assign n5080 = pi18 ? n5079 : n2703;
  assign n5081 = pi17 ? n37 : n5080;
  assign n5082 = pi16 ? n439 : n5081;
  assign n5083 = pi15 ? n5076 : n5082;
  assign n5084 = pi14 ? n5069 : n5083;
  assign n5085 = pi21 ? n99 : n685;
  assign n5086 = pi20 ? n99 : n5085;
  assign n5087 = pi19 ? n99 : n5086;
  assign n5088 = pi18 ? n5087 : n1824;
  assign n5089 = pi17 ? n99 : n5088;
  assign n5090 = pi16 ? n744 : n5089;
  assign n5091 = pi21 ? n767 : n685;
  assign n5092 = pi20 ? n99 : n5091;
  assign n5093 = pi19 ? n99 : n5092;
  assign n5094 = pi18 ? n5093 : n1824;
  assign n5095 = pi17 ? n99 : n5094;
  assign n5096 = pi16 ? n721 : n5095;
  assign n5097 = pi15 ? n5090 : n5096;
  assign n5098 = pi18 ? n5087 : n32;
  assign n5099 = pi17 ? n99 : n5098;
  assign n5100 = pi16 ? n721 : n5099;
  assign n5101 = pi22 ? n158 : n685;
  assign n5102 = pi21 ? n99 : n5101;
  assign n5103 = pi20 ? n99 : n5102;
  assign n5104 = pi19 ? n99 : n5103;
  assign n5105 = pi18 ? n5104 : n32;
  assign n5106 = pi17 ? n99 : n5105;
  assign n5107 = pi16 ? n721 : n5106;
  assign n5108 = pi15 ? n5100 : n5107;
  assign n5109 = pi14 ? n5097 : n5108;
  assign n5110 = pi13 ? n5084 : n5109;
  assign n5111 = pi12 ? n5053 : n5110;
  assign n5112 = pi16 ? n721 : n4187;
  assign n5113 = pi22 ? n685 : n1475;
  assign n5114 = pi21 ? n99 : n5113;
  assign n5115 = pi20 ? n99 : n5114;
  assign n5116 = pi19 ? n99 : n5115;
  assign n5117 = pi18 ? n5116 : n32;
  assign n5118 = pi17 ? n99 : n5117;
  assign n5119 = pi16 ? n721 : n5118;
  assign n5120 = pi15 ? n5112 : n5119;
  assign n5121 = pi20 ? n99 : n220;
  assign n5122 = pi19 ? n5121 : n99;
  assign n5123 = pi18 ? n719 : n5122;
  assign n5124 = pi17 ? n32 : n5123;
  assign n5125 = pi20 ? n2243 : n2208;
  assign n5126 = pi19 ? n99 : n5125;
  assign n5127 = pi18 ? n5126 : n32;
  assign n5128 = pi17 ? n99 : n5127;
  assign n5129 = pi16 ? n5124 : n5128;
  assign n5130 = pi21 ? n1505 : n1143;
  assign n5131 = pi20 ? n32 : n5130;
  assign n5132 = pi19 ? n32 : n5131;
  assign n5133 = pi20 ? n3888 : n220;
  assign n5134 = pi20 ? n2749 : n4202;
  assign n5135 = pi19 ? n5133 : n5134;
  assign n5136 = pi18 ? n5132 : n5135;
  assign n5137 = pi17 ? n32 : n5136;
  assign n5138 = pi20 ? n2174 : n3807;
  assign n5139 = pi19 ? n5138 : n99;
  assign n5140 = pi20 ? n99 : n2749;
  assign n5141 = pi20 ? n4202 : n2749;
  assign n5142 = pi19 ? n5140 : n5141;
  assign n5143 = pi18 ? n5139 : n5142;
  assign n5144 = pi20 ? n3506 : n2238;
  assign n5145 = pi22 ? n157 : n317;
  assign n5146 = pi21 ? n99 : n5145;
  assign n5147 = pi20 ? n157 : n5146;
  assign n5148 = pi19 ? n5144 : n5147;
  assign n5149 = pi18 ? n5148 : n32;
  assign n5150 = pi17 ? n5143 : n5149;
  assign n5151 = pi16 ? n5137 : n5150;
  assign n5152 = pi15 ? n5129 : n5151;
  assign n5153 = pi14 ? n5120 : n5152;
  assign n5154 = pi23 ? n961 : n157;
  assign n5155 = pi22 ? n5154 : n157;
  assign n5156 = pi21 ? n5155 : n157;
  assign n5157 = pi20 ? n32 : n5156;
  assign n5158 = pi19 ? n32 : n5157;
  assign n5159 = pi18 ? n5158 : n157;
  assign n5160 = pi17 ? n32 : n5159;
  assign n5161 = pi21 ? n157 : n5145;
  assign n5162 = pi20 ? n157 : n5161;
  assign n5163 = pi19 ? n157 : n5162;
  assign n5164 = pi18 ? n5163 : n32;
  assign n5165 = pi17 ? n157 : n5164;
  assign n5166 = pi16 ? n5160 : n5165;
  assign n5167 = pi23 ? n38 : n157;
  assign n5168 = pi22 ? n5167 : n157;
  assign n5169 = pi21 ? n5168 : n157;
  assign n5170 = pi20 ? n32 : n5169;
  assign n5171 = pi19 ? n32 : n5170;
  assign n5172 = pi20 ? n157 : n259;
  assign n5173 = pi19 ? n5172 : n157;
  assign n5174 = pi18 ? n5171 : n5173;
  assign n5175 = pi17 ? n32 : n5174;
  assign n5176 = pi22 ? n204 : n157;
  assign n5177 = pi21 ? n5176 : n204;
  assign n5178 = pi22 ? n316 : n317;
  assign n5179 = pi21 ? n157 : n5178;
  assign n5180 = pi20 ? n5177 : n5179;
  assign n5181 = pi19 ? n157 : n5180;
  assign n5182 = pi18 ? n5181 : n32;
  assign n5183 = pi17 ? n157 : n5182;
  assign n5184 = pi16 ? n5175 : n5183;
  assign n5185 = pi15 ? n5166 : n5184;
  assign n5186 = pi22 ? n909 : n204;
  assign n5187 = pi21 ? n5186 : n916;
  assign n5188 = pi20 ? n32 : n5187;
  assign n5189 = pi19 ? n32 : n5188;
  assign n5190 = pi20 ? n921 : n2318;
  assign n5191 = pi20 ? n2318 : n916;
  assign n5192 = pi19 ? n5190 : n5191;
  assign n5193 = pi18 ? n5189 : n5192;
  assign n5194 = pi17 ? n32 : n5193;
  assign n5195 = pi20 ? n1016 : n2316;
  assign n5196 = pi20 ? n204 : n921;
  assign n5197 = pi19 ? n5195 : n5196;
  assign n5198 = pi20 ? n204 : n916;
  assign n5199 = pi21 ? n921 : n204;
  assign n5200 = pi20 ? n5199 : n916;
  assign n5201 = pi19 ? n5198 : n5200;
  assign n5202 = pi18 ? n5197 : n5201;
  assign n5203 = pi20 ? n921 : n5199;
  assign n5204 = pi21 ? n204 : n921;
  assign n5205 = pi21 ? n316 : n5178;
  assign n5206 = pi20 ? n5204 : n5205;
  assign n5207 = pi19 ? n5203 : n5206;
  assign n5208 = pi18 ? n5207 : n32;
  assign n5209 = pi17 ? n5202 : n5208;
  assign n5210 = pi16 ? n5194 : n5209;
  assign n5211 = pi21 ? n2856 : n1793;
  assign n5212 = pi20 ? n32 : n5211;
  assign n5213 = pi19 ? n32 : n5212;
  assign n5214 = pi21 ? n2863 : n2869;
  assign n5215 = pi21 ? n2876 : n139;
  assign n5216 = pi20 ? n5214 : n5215;
  assign n5217 = pi21 ? n1793 : n919;
  assign n5218 = pi20 ? n5215 : n5217;
  assign n5219 = pi19 ? n5216 : n5218;
  assign n5220 = pi18 ? n5213 : n5219;
  assign n5221 = pi17 ? n32 : n5220;
  assign n5222 = pi21 ? n139 : n2876;
  assign n5223 = pi21 ? n919 : n4712;
  assign n5224 = pi20 ? n5222 : n5223;
  assign n5225 = pi20 ? n4712 : n921;
  assign n5226 = pi19 ? n5224 : n5225;
  assign n5227 = pi21 ? n916 : n919;
  assign n5228 = pi20 ? n2876 : n5227;
  assign n5229 = pi21 ? n921 : n2876;
  assign n5230 = pi20 ? n5229 : n5227;
  assign n5231 = pi19 ? n5228 : n5230;
  assign n5232 = pi18 ? n5226 : n5231;
  assign n5233 = pi21 ? n2863 : n204;
  assign n5234 = pi20 ? n921 : n5233;
  assign n5235 = pi22 ? n139 : n2299;
  assign n5236 = pi21 ? n5235 : n139;
  assign n5237 = pi20 ? n5236 : n5205;
  assign n5238 = pi19 ? n5234 : n5237;
  assign n5239 = pi18 ? n5238 : n32;
  assign n5240 = pi17 ? n5232 : n5239;
  assign n5241 = pi16 ? n5221 : n5240;
  assign n5242 = pi15 ? n5210 : n5241;
  assign n5243 = pi14 ? n5185 : n5242;
  assign n5244 = pi13 ? n5153 : n5243;
  assign n5245 = pi21 ? n316 : n3523;
  assign n5246 = pi20 ? n4437 : n5245;
  assign n5247 = pi19 ? n3578 : n5246;
  assign n5248 = pi18 ? n5247 : n32;
  assign n5249 = pi17 ? n139 : n5248;
  assign n5250 = pi16 ? n2810 : n5249;
  assign n5251 = pi22 ? n909 : n295;
  assign n5252 = pi21 ? n5251 : n297;
  assign n5253 = pi20 ? n32 : n5252;
  assign n5254 = pi19 ? n32 : n5253;
  assign n5255 = pi21 ? n1698 : n37;
  assign n5256 = pi20 ? n3932 : n5255;
  assign n5257 = pi21 ? n1531 : n37;
  assign n5258 = pi21 ? n297 : n1696;
  assign n5259 = pi20 ? n5257 : n5258;
  assign n5260 = pi19 ? n5256 : n5259;
  assign n5261 = pi18 ? n5254 : n5260;
  assign n5262 = pi17 ? n32 : n5261;
  assign n5263 = pi21 ? n3073 : n1529;
  assign n5264 = pi20 ? n5263 : n1719;
  assign n5265 = pi21 ? n1721 : n295;
  assign n5266 = pi20 ? n5265 : n2830;
  assign n5267 = pi19 ? n5264 : n5266;
  assign n5268 = pi20 ? n3913 : n2527;
  assign n5269 = pi21 ? n1696 : n1531;
  assign n5270 = pi20 ? n2513 : n5269;
  assign n5271 = pi19 ? n5268 : n5270;
  assign n5272 = pi18 ? n5267 : n5271;
  assign n5273 = pi21 ? n1211 : n139;
  assign n5274 = pi21 ? n1531 : n1785;
  assign n5275 = pi20 ? n5273 : n5274;
  assign n5276 = pi20 ? n316 : n5245;
  assign n5277 = pi19 ? n5275 : n5276;
  assign n5278 = pi18 ? n5277 : n32;
  assign n5279 = pi17 ? n5272 : n5278;
  assign n5280 = pi16 ? n5262 : n5279;
  assign n5281 = pi15 ? n5250 : n5280;
  assign n5282 = pi22 ? n909 : n316;
  assign n5283 = pi21 ? n5282 : n316;
  assign n5284 = pi20 ? n32 : n5283;
  assign n5285 = pi19 ? n32 : n5284;
  assign n5286 = pi21 ? n316 : n4020;
  assign n5287 = pi20 ? n316 : n5286;
  assign n5288 = pi20 ? n2353 : n316;
  assign n5289 = pi19 ? n5287 : n5288;
  assign n5290 = pi18 ? n5285 : n5289;
  assign n5291 = pi17 ? n32 : n5290;
  assign n5292 = pi19 ? n316 : n5276;
  assign n5293 = pi18 ? n5292 : n32;
  assign n5294 = pi17 ? n316 : n5293;
  assign n5295 = pi16 ? n5291 : n5294;
  assign n5296 = pi21 ? n4472 : n356;
  assign n5297 = pi20 ? n32 : n5296;
  assign n5298 = pi19 ? n32 : n5297;
  assign n5299 = pi21 ? n316 : n381;
  assign n5300 = pi20 ? n5299 : n1022;
  assign n5301 = pi20 ? n2353 : n975;
  assign n5302 = pi19 ? n5300 : n5301;
  assign n5303 = pi18 ? n5298 : n5302;
  assign n5304 = pi17 ? n32 : n5303;
  assign n5305 = pi20 ? n4437 : n316;
  assign n5306 = pi19 ? n5305 : n316;
  assign n5307 = pi18 ? n5306 : n316;
  assign n5308 = pi17 ? n5307 : n5293;
  assign n5309 = pi16 ? n5304 : n5308;
  assign n5310 = pi15 ? n5295 : n5309;
  assign n5311 = pi14 ? n5281 : n5310;
  assign n5312 = pi20 ? n1022 : n139;
  assign n5313 = pi19 ? n5312 : n139;
  assign n5314 = pi18 ? n1573 : n5313;
  assign n5315 = pi17 ? n32 : n5314;
  assign n5316 = pi19 ? n1820 : n316;
  assign n5317 = pi21 ? n316 : n356;
  assign n5318 = pi20 ? n4437 : n5317;
  assign n5319 = pi20 ? n975 : n1008;
  assign n5320 = pi19 ? n5318 : n5319;
  assign n5321 = pi18 ? n5316 : n5320;
  assign n5322 = pi19 ? n999 : n5276;
  assign n5323 = pi18 ? n5322 : n32;
  assign n5324 = pi17 ? n5321 : n5323;
  assign n5325 = pi16 ? n5315 : n5324;
  assign n5326 = pi21 ? n4472 : n3258;
  assign n5327 = pi20 ? n32 : n5326;
  assign n5328 = pi19 ? n32 : n5327;
  assign n5329 = pi21 ? n1027 : n37;
  assign n5330 = pi20 ? n5299 : n5329;
  assign n5331 = pi21 ? n3693 : n1018;
  assign n5332 = pi21 ? n335 : n1018;
  assign n5333 = pi20 ? n5331 : n5332;
  assign n5334 = pi19 ? n5330 : n5333;
  assign n5335 = pi18 ? n5328 : n5334;
  assign n5336 = pi17 ? n32 : n5335;
  assign n5337 = pi20 ? n3697 : n316;
  assign n5338 = pi20 ? n316 : n4002;
  assign n5339 = pi19 ? n5337 : n5338;
  assign n5340 = pi20 ? n2383 : n1019;
  assign n5341 = pi20 ? n316 : n1019;
  assign n5342 = pi19 ? n5340 : n5341;
  assign n5343 = pi18 ? n5339 : n5342;
  assign n5344 = pi20 ? n1018 : n2330;
  assign n5345 = pi19 ? n316 : n5344;
  assign n5346 = pi18 ? n5345 : n32;
  assign n5347 = pi17 ? n5343 : n5346;
  assign n5348 = pi16 ? n5336 : n5347;
  assign n5349 = pi15 ? n5325 : n5348;
  assign n5350 = pi22 ? n1591 : n204;
  assign n5351 = pi21 ? n5350 : n204;
  assign n5352 = pi20 ? n32 : n5351;
  assign n5353 = pi19 ? n32 : n5352;
  assign n5354 = pi18 ? n5353 : n204;
  assign n5355 = pi17 ? n32 : n5354;
  assign n5356 = pi21 ? n204 : n2637;
  assign n5357 = pi20 ? n204 : n5356;
  assign n5358 = pi19 ? n204 : n5357;
  assign n5359 = pi18 ? n5358 : n32;
  assign n5360 = pi17 ? n204 : n5359;
  assign n5361 = pi16 ? n5355 : n5360;
  assign n5362 = pi22 ? n2419 : n204;
  assign n5363 = pi21 ? n5362 : n204;
  assign n5364 = pi20 ? n32 : n5363;
  assign n5365 = pi19 ? n32 : n5364;
  assign n5366 = pi19 ? n204 : n1100;
  assign n5367 = pi18 ? n5365 : n5366;
  assign n5368 = pi17 ? n32 : n5367;
  assign n5369 = pi23 ? n2766 : n32;
  assign n5370 = pi22 ? n5369 : n32;
  assign n5371 = pi21 ? n204 : n5370;
  assign n5372 = pi20 ? n204 : n5371;
  assign n5373 = pi19 ? n204 : n5372;
  assign n5374 = pi18 ? n5373 : n32;
  assign n5375 = pi17 ? n204 : n5374;
  assign n5376 = pi16 ? n5368 : n5375;
  assign n5377 = pi15 ? n5361 : n5376;
  assign n5378 = pi14 ? n5349 : n5377;
  assign n5379 = pi13 ? n5311 : n5378;
  assign n5380 = pi12 ? n5244 : n5379;
  assign n5381 = pi11 ? n5111 : n5380;
  assign n5382 = pi10 ? n4970 : n5381;
  assign n5383 = pi09 ? n32 : n5382;
  assign n5384 = pi16 ? n3784 : n4524;
  assign n5385 = pi16 ? n70 : n4524;
  assign n5386 = pi15 ? n5384 : n5385;
  assign n5387 = pi20 ? n372 : n37;
  assign n5388 = pi19 ? n5387 : n37;
  assign n5389 = pi18 ? n32 : n5388;
  assign n5390 = pi17 ? n32 : n5389;
  assign n5391 = pi16 ? n5390 : n4524;
  assign n5392 = pi16 ? n73 : n4524;
  assign n5393 = pi15 ? n5391 : n5392;
  assign n5394 = pi14 ? n5386 : n5393;
  assign n5395 = pi15 ? n4525 : n4527;
  assign n5396 = pi21 ? n85 : n32;
  assign n5397 = pi20 ? n5396 : n32;
  assign n5398 = pi19 ? n5397 : n32;
  assign n5399 = pi18 ? n37 : n5398;
  assign n5400 = pi17 ? n37 : n5399;
  assign n5401 = pi16 ? n439 : n5400;
  assign n5402 = pi15 ? n4533 : n5401;
  assign n5403 = pi14 ? n5395 : n5402;
  assign n5404 = pi13 ? n5394 : n5403;
  assign n5405 = pi21 ? n2161 : n99;
  assign n5406 = pi19 ? n5405 : n99;
  assign n5407 = pi18 ? n184 : n5406;
  assign n5408 = pi17 ? n32 : n5407;
  assign n5409 = pi22 ? n4543 : n112;
  assign n5410 = pi21 ? n2161 : n5409;
  assign n5411 = pi20 ? n99 : n5410;
  assign n5412 = pi19 ? n99 : n5411;
  assign n5413 = pi21 ? n99 : n5409;
  assign n5414 = pi20 ? n5413 : n4549;
  assign n5415 = pi21 ? n4538 : n2164;
  assign n5416 = pi20 ? n5410 : n5415;
  assign n5417 = pi19 ? n5414 : n5416;
  assign n5418 = pi18 ? n5412 : n5417;
  assign n5419 = pi20 ? n5415 : n5405;
  assign n5420 = pi21 ? n99 : n2746;
  assign n5421 = pi20 ? n5420 : n99;
  assign n5422 = pi19 ? n5419 : n5421;
  assign n5423 = pi22 ? n99 : n47;
  assign n5424 = pi21 ? n5423 : n32;
  assign n5425 = pi20 ? n5424 : n32;
  assign n5426 = pi19 ? n5425 : n32;
  assign n5427 = pi18 ? n5422 : n5426;
  assign n5428 = pi17 ? n5418 : n5427;
  assign n5429 = pi16 ? n5408 : n5428;
  assign n5430 = pi21 ? n120 : n32;
  assign n5431 = pi20 ? n5430 : n32;
  assign n5432 = pi19 ? n5431 : n32;
  assign n5433 = pi18 ? n99 : n5432;
  assign n5434 = pi17 ? n99 : n5433;
  assign n5435 = pi16 ? n721 : n5434;
  assign n5436 = pi15 ? n5429 : n5435;
  assign n5437 = pi14 ? n5436 : n5435;
  assign n5438 = pi21 ? n141 : n32;
  assign n5439 = pi20 ? n5438 : n32;
  assign n5440 = pi19 ? n5439 : n32;
  assign n5441 = pi18 ? n99 : n5440;
  assign n5442 = pi17 ? n99 : n5441;
  assign n5443 = pi16 ? n801 : n5442;
  assign n5444 = pi22 ? n99 : n1344;
  assign n5445 = pi21 ? n5444 : n32;
  assign n5446 = pi20 ? n5445 : n32;
  assign n5447 = pi19 ? n5446 : n32;
  assign n5448 = pi18 ? n4586 : n5447;
  assign n5449 = pi17 ? n4585 : n5448;
  assign n5450 = pi16 ? n801 : n5449;
  assign n5451 = pi15 ? n5443 : n5450;
  assign n5452 = pi23 ? n685 : n99;
  assign n5453 = pi22 ? n99 : n5452;
  assign n5454 = pi21 ? n99 : n5453;
  assign n5455 = pi20 ? n99 : n5454;
  assign n5456 = pi19 ? n99 : n5455;
  assign n5457 = pi20 ? n5454 : n99;
  assign n5458 = pi22 ? n5452 : n99;
  assign n5459 = pi21 ? n5458 : n99;
  assign n5460 = pi20 ? n99 : n5459;
  assign n5461 = pi19 ? n5457 : n5460;
  assign n5462 = pi18 ? n5456 : n5461;
  assign n5463 = pi21 ? n5458 : n5453;
  assign n5464 = pi22 ? n3443 : n99;
  assign n5465 = pi21 ? n5464 : n99;
  assign n5466 = pi20 ? n5463 : n5465;
  assign n5467 = pi21 ? n99 : n3444;
  assign n5468 = pi20 ? n5467 : n99;
  assign n5469 = pi19 ? n5466 : n5468;
  assign n5470 = pi22 ? n99 : n759;
  assign n5471 = pi21 ? n5470 : n32;
  assign n5472 = pi20 ? n5471 : n32;
  assign n5473 = pi19 ? n5472 : n32;
  assign n5474 = pi18 ? n5469 : n5473;
  assign n5475 = pi17 ? n5462 : n5474;
  assign n5476 = pi16 ? n744 : n5475;
  assign n5477 = pi19 ? n4599 : n3481;
  assign n5478 = pi18 ? n4598 : n5477;
  assign n5479 = pi21 ? n2998 : n165;
  assign n5480 = pi20 ? n5479 : n169;
  assign n5481 = pi19 ? n5480 : n4604;
  assign n5482 = pi22 ? n99 : n1378;
  assign n5483 = pi21 ? n5482 : n32;
  assign n5484 = pi20 ? n5483 : n32;
  assign n5485 = pi19 ? n5484 : n32;
  assign n5486 = pi18 ? n5481 : n5485;
  assign n5487 = pi17 ? n5478 : n5486;
  assign n5488 = pi16 ? n1676 : n5487;
  assign n5489 = pi15 ? n5476 : n5488;
  assign n5490 = pi14 ? n5451 : n5489;
  assign n5491 = pi13 ? n5437 : n5490;
  assign n5492 = pi12 ? n5404 : n5491;
  assign n5493 = pi21 ? n1671 : n2164;
  assign n5494 = pi20 ? n32 : n5493;
  assign n5495 = pi19 ? n32 : n5494;
  assign n5496 = pi21 ? n2175 : n2168;
  assign n5497 = pi20 ? n2968 : n3814;
  assign n5498 = pi19 ? n5496 : n5497;
  assign n5499 = pi18 ? n5495 : n5498;
  assign n5500 = pi17 ? n32 : n5499;
  assign n5501 = pi21 ? n2160 : n112;
  assign n5502 = pi20 ? n3870 : n5501;
  assign n5503 = pi19 ? n5502 : n3824;
  assign n5504 = pi20 ? n3824 : n5501;
  assign n5505 = pi20 ? n5496 : n2169;
  assign n5506 = pi19 ? n5504 : n5505;
  assign n5507 = pi18 ? n5503 : n5506;
  assign n5508 = pi20 ? n2174 : n2163;
  assign n5509 = pi21 ? n2168 : n2162;
  assign n5510 = pi19 ? n5508 : n5509;
  assign n5511 = pi22 ? n2160 : n396;
  assign n5512 = pi21 ? n5511 : n32;
  assign n5513 = pi20 ? n5512 : n32;
  assign n5514 = pi19 ? n5513 : n32;
  assign n5515 = pi18 ? n5510 : n5514;
  assign n5516 = pi17 ? n5507 : n5515;
  assign n5517 = pi16 ? n5500 : n5516;
  assign n5518 = pi22 ? n157 : n295;
  assign n5519 = pi21 ? n180 : n5518;
  assign n5520 = pi20 ? n32 : n5519;
  assign n5521 = pi19 ? n32 : n5520;
  assign n5522 = pi22 ? n893 : n1043;
  assign n5523 = pi21 ? n5522 : n248;
  assign n5524 = pi22 ? n295 : n893;
  assign n5525 = pi21 ? n5524 : n1211;
  assign n5526 = pi21 ? n5518 : n5522;
  assign n5527 = pi20 ? n5525 : n5526;
  assign n5528 = pi19 ? n5523 : n5527;
  assign n5529 = pi18 ? n5521 : n5528;
  assign n5530 = pi17 ? n32 : n5529;
  assign n5531 = pi21 ? n248 : n5524;
  assign n5532 = pi21 ? n1211 : n5518;
  assign n5533 = pi20 ? n5531 : n5532;
  assign n5534 = pi21 ? n4652 : n5518;
  assign n5535 = pi21 ? n5522 : n157;
  assign n5536 = pi20 ? n5534 : n5535;
  assign n5537 = pi19 ? n5533 : n5536;
  assign n5538 = pi21 ? n139 : n5518;
  assign n5539 = pi20 ? n5535 : n5538;
  assign n5540 = pi22 ? n157 : n1043;
  assign n5541 = pi21 ? n5540 : n248;
  assign n5542 = pi20 ? n5523 : n5541;
  assign n5543 = pi19 ? n5539 : n5542;
  assign n5544 = pi18 ? n5537 : n5543;
  assign n5545 = pi21 ? n5540 : n157;
  assign n5546 = pi20 ? n5545 : n258;
  assign n5547 = pi21 ? n248 : n1526;
  assign n5548 = pi21 ? n248 : n1721;
  assign n5549 = pi20 ? n5547 : n5548;
  assign n5550 = pi19 ? n5546 : n5549;
  assign n5551 = pi22 ? n139 : n396;
  assign n5552 = pi21 ? n5551 : n32;
  assign n5553 = pi20 ? n5552 : n32;
  assign n5554 = pi19 ? n5553 : n32;
  assign n5555 = pi18 ? n5550 : n5554;
  assign n5556 = pi17 ? n5544 : n5555;
  assign n5557 = pi16 ? n5530 : n5556;
  assign n5558 = pi15 ? n5517 : n5557;
  assign n5559 = pi22 ? n204 : n295;
  assign n5560 = pi21 ? n180 : n5559;
  assign n5561 = pi20 ? n32 : n5560;
  assign n5562 = pi19 ? n32 : n5561;
  assign n5563 = pi21 ? n5522 : n916;
  assign n5564 = pi21 ? n5559 : n5522;
  assign n5565 = pi20 ? n5525 : n5564;
  assign n5566 = pi19 ? n5563 : n5565;
  assign n5567 = pi18 ? n5562 : n5566;
  assign n5568 = pi17 ? n32 : n5567;
  assign n5569 = pi21 ? n916 : n5524;
  assign n5570 = pi21 ? n1211 : n5559;
  assign n5571 = pi20 ? n5569 : n5570;
  assign n5572 = pi21 ? n4652 : n5559;
  assign n5573 = pi21 ? n5522 : n139;
  assign n5574 = pi20 ? n5572 : n5573;
  assign n5575 = pi19 ? n5571 : n5574;
  assign n5576 = pi21 ? n139 : n5559;
  assign n5577 = pi20 ? n5573 : n5576;
  assign n5578 = pi21 ? n1711 : n916;
  assign n5579 = pi20 ? n5563 : n5578;
  assign n5580 = pi19 ? n5577 : n5579;
  assign n5581 = pi18 ? n5575 : n5580;
  assign n5582 = pi20 ? n5578 : n139;
  assign n5583 = pi21 ? n916 : n1721;
  assign n5584 = pi19 ? n5582 : n5583;
  assign n5585 = pi21 ? n318 : n32;
  assign n5586 = pi20 ? n5585 : n32;
  assign n5587 = pi19 ? n5586 : n32;
  assign n5588 = pi18 ? n5584 : n5587;
  assign n5589 = pi17 ? n5581 : n5588;
  assign n5590 = pi16 ? n5568 : n5589;
  assign n5591 = pi21 ? n180 : n1531;
  assign n5592 = pi20 ? n32 : n5591;
  assign n5593 = pi19 ? n32 : n5592;
  assign n5594 = pi21 ? n1834 : n916;
  assign n5595 = pi21 ? n2585 : n1211;
  assign n5596 = pi21 ? n5559 : n1834;
  assign n5597 = pi20 ? n5595 : n5596;
  assign n5598 = pi19 ? n5594 : n5597;
  assign n5599 = pi18 ? n5593 : n5598;
  assign n5600 = pi17 ? n32 : n5599;
  assign n5601 = pi21 ? n916 : n2585;
  assign n5602 = pi20 ? n5601 : n5570;
  assign n5603 = pi21 ? n1834 : n1211;
  assign n5604 = pi19 ? n5602 : n5603;
  assign n5605 = pi20 ? n1707 : n2527;
  assign n5606 = pi21 ? n295 : n916;
  assign n5607 = pi20 ? n5594 : n5606;
  assign n5608 = pi19 ? n5605 : n5607;
  assign n5609 = pi18 ? n5604 : n5608;
  assign n5610 = pi20 ? n1714 : n3625;
  assign n5611 = pi19 ? n5610 : n1738;
  assign n5612 = pi24 ? n37 : n139;
  assign n5613 = pi23 ? n139 : n5612;
  assign n5614 = pi22 ? n5613 : n587;
  assign n5615 = pi21 ? n5614 : n32;
  assign n5616 = pi20 ? n5615 : n32;
  assign n5617 = pi19 ? n5616 : n32;
  assign n5618 = pi18 ? n5611 : n5617;
  assign n5619 = pi17 ? n5609 : n5618;
  assign n5620 = pi16 ? n5600 : n5619;
  assign n5621 = pi15 ? n5590 : n5620;
  assign n5622 = pi14 ? n5558 : n5621;
  assign n5623 = pi22 ? n139 : n587;
  assign n5624 = pi21 ? n5623 : n32;
  assign n5625 = pi20 ? n5624 : n32;
  assign n5626 = pi19 ? n5625 : n32;
  assign n5627 = pi18 ? n139 : n5626;
  assign n5628 = pi17 ? n139 : n5627;
  assign n5629 = pi16 ? n314 : n5628;
  assign n5630 = pi24 ? n363 : n32;
  assign n5631 = pi23 ? n5630 : n32;
  assign n5632 = pi22 ? n204 : n5631;
  assign n5633 = pi21 ? n5632 : n32;
  assign n5634 = pi20 ? n5633 : n32;
  assign n5635 = pi19 ? n5634 : n32;
  assign n5636 = pi18 ? n139 : n5635;
  assign n5637 = pi17 ? n139 : n5636;
  assign n5638 = pi16 ? n1773 : n5637;
  assign n5639 = pi15 ? n5629 : n5638;
  assign n5640 = pi22 ? n335 : n5631;
  assign n5641 = pi21 ? n5640 : n32;
  assign n5642 = pi20 ? n5641 : n32;
  assign n5643 = pi19 ? n5642 : n32;
  assign n5644 = pi18 ? n139 : n5643;
  assign n5645 = pi17 ? n139 : n5644;
  assign n5646 = pi16 ? n1773 : n5645;
  assign n5647 = pi21 ? n3986 : n346;
  assign n5648 = pi20 ? n32 : n5647;
  assign n5649 = pi19 ? n32 : n5648;
  assign n5650 = pi21 ? n4780 : n2319;
  assign n5651 = pi21 ? n354 : n1784;
  assign n5652 = pi21 ? n4020 : n4780;
  assign n5653 = pi20 ? n5651 : n5652;
  assign n5654 = pi19 ? n5650 : n5653;
  assign n5655 = pi18 ? n5649 : n5654;
  assign n5656 = pi17 ? n32 : n5655;
  assign n5657 = pi21 ? n2319 : n354;
  assign n5658 = pi21 ? n1784 : n4020;
  assign n5659 = pi20 ? n5657 : n5658;
  assign n5660 = pi21 ? n4780 : n346;
  assign n5661 = pi20 ? n5660 : n316;
  assign n5662 = pi19 ? n5659 : n5661;
  assign n5663 = pi18 ? n5662 : n4782;
  assign n5664 = pi21 ? n2319 : n4429;
  assign n5665 = pi20 ? n5657 : n5664;
  assign n5666 = pi19 ? n4785 : n5665;
  assign n5667 = pi21 ? n5178 : n32;
  assign n5668 = pi20 ? n5667 : n32;
  assign n5669 = pi19 ? n5668 : n32;
  assign n5670 = pi18 ? n5666 : n5669;
  assign n5671 = pi17 ? n5663 : n5670;
  assign n5672 = pi16 ? n5656 : n5671;
  assign n5673 = pi15 ? n5646 : n5672;
  assign n5674 = pi14 ? n5639 : n5673;
  assign n5675 = pi13 ? n5622 : n5674;
  assign n5676 = pi21 ? n4052 : n4015;
  assign n5677 = pi20 ? n5676 : n4054;
  assign n5678 = pi19 ? n5677 : n4059;
  assign n5679 = pi18 ? n3254 : n5678;
  assign n5680 = pi17 ? n32 : n5679;
  assign n5681 = pi21 ? n417 : n381;
  assign n5682 = pi20 ? n5681 : n4053;
  assign n5683 = pi19 ? n4065 : n5682;
  assign n5684 = pi20 ? n4053 : n3275;
  assign n5685 = pi21 ? n392 : n4015;
  assign n5686 = pi20 ? n5676 : n5685;
  assign n5687 = pi19 ? n5684 : n5686;
  assign n5688 = pi18 ? n5683 : n5687;
  assign n5689 = pi21 ? n384 : n316;
  assign n5690 = pi21 ? n384 : n3258;
  assign n5691 = pi20 ? n5689 : n5690;
  assign n5692 = pi19 ? n4810 : n5691;
  assign n5693 = pi18 ? n5692 : n5669;
  assign n5694 = pi17 ? n5688 : n5693;
  assign n5695 = pi16 ? n5680 : n5694;
  assign n5696 = pi21 ? n37 : n384;
  assign n5697 = pi20 ? n5696 : n37;
  assign n5698 = pi19 ? n5697 : n37;
  assign n5699 = pi18 ? n374 : n5698;
  assign n5700 = pi17 ? n32 : n5699;
  assign n5701 = pi18 ? n4820 : n5669;
  assign n5702 = pi17 ? n4818 : n5701;
  assign n5703 = pi16 ? n5700 : n5702;
  assign n5704 = pi15 ? n5695 : n5703;
  assign n5705 = pi22 ? n2401 : n383;
  assign n5706 = pi21 ? n37 : n5705;
  assign n5707 = pi21 ? n37 : n417;
  assign n5708 = pi20 ? n5706 : n5707;
  assign n5709 = pi21 ? n384 : n391;
  assign n5710 = pi20 ? n5709 : n3256;
  assign n5711 = pi19 ? n5708 : n5710;
  assign n5712 = pi18 ? n4827 : n5711;
  assign n5713 = pi17 ? n32 : n5712;
  assign n5714 = pi21 ? n417 : n384;
  assign n5715 = pi20 ? n5714 : n429;
  assign n5716 = pi21 ? n37 : n4052;
  assign n5717 = pi20 ? n3277 : n5716;
  assign n5718 = pi19 ? n5715 : n5717;
  assign n5719 = pi20 ? n5716 : n429;
  assign n5720 = pi20 ? n5707 : n418;
  assign n5721 = pi19 ? n5719 : n5720;
  assign n5722 = pi18 ? n5718 : n5721;
  assign n5723 = pi21 ? n391 : n384;
  assign n5724 = pi20 ? n426 : n5723;
  assign n5725 = pi19 ? n5724 : n5714;
  assign n5726 = pi22 ? n2401 : n532;
  assign n5727 = pi21 ? n5726 : n32;
  assign n5728 = pi20 ? n5727 : n32;
  assign n5729 = pi19 ? n5728 : n32;
  assign n5730 = pi18 ? n5725 : n5729;
  assign n5731 = pi17 ? n5722 : n5730;
  assign n5732 = pi16 ? n5713 : n5731;
  assign n5733 = pi21 ? n37 : n499;
  assign n5734 = pi20 ? n5733 : n37;
  assign n5735 = pi19 ? n5734 : n37;
  assign n5736 = pi18 ? n374 : n5735;
  assign n5737 = pi17 ? n32 : n5736;
  assign n5738 = pi16 ? n5737 : n4856;
  assign n5739 = pi15 ? n5732 : n5738;
  assign n5740 = pi14 ? n5704 : n5739;
  assign n5741 = pi21 ? n499 : n1309;
  assign n5742 = pi20 ? n5741 : n508;
  assign n5743 = pi19 ? n5742 : n4865;
  assign n5744 = pi18 ? n374 : n5743;
  assign n5745 = pi17 ? n32 : n5744;
  assign n5746 = pi22 ? n204 : n688;
  assign n5747 = pi21 ? n5746 : n32;
  assign n5748 = pi20 ? n5747 : n32;
  assign n5749 = pi19 ? n5748 : n32;
  assign n5750 = pi18 ? n4881 : n5749;
  assign n5751 = pi17 ? n4877 : n5750;
  assign n5752 = pi16 ? n5745 : n5751;
  assign n5753 = pi21 ? n3404 : n4893;
  assign n5754 = pi20 ? n37 : n5753;
  assign n5755 = pi19 ? n37 : n5754;
  assign n5756 = pi18 ? n374 : n5755;
  assign n5757 = pi17 ? n32 : n5756;
  assign n5758 = pi22 ? n233 : n706;
  assign n5759 = pi21 ? n5758 : n32;
  assign n5760 = pi20 ? n5759 : n32;
  assign n5761 = pi19 ? n5760 : n32;
  assign n5762 = pi18 ? n4924 : n5761;
  assign n5763 = pi17 ? n4919 : n5762;
  assign n5764 = pi16 ? n5757 : n5763;
  assign n5765 = pi15 ? n5752 : n5764;
  assign n5766 = pi21 ? n37 : n567;
  assign n5767 = pi20 ? n37 : n5766;
  assign n5768 = pi19 ? n37 : n5767;
  assign n5769 = pi18 ? n374 : n5768;
  assign n5770 = pi17 ? n32 : n5769;
  assign n5771 = pi22 ? n2060 : n32;
  assign n5772 = pi21 ? n5771 : n32;
  assign n5773 = pi20 ? n5772 : n32;
  assign n5774 = pi19 ? n5773 : n32;
  assign n5775 = pi18 ? n335 : n5774;
  assign n5776 = pi17 ? n4942 : n5775;
  assign n5777 = pi16 ? n5770 : n5776;
  assign n5778 = pi21 ? n584 : n569;
  assign n5779 = pi20 ? n4971 : n5778;
  assign n5780 = pi19 ? n5779 : n4955;
  assign n5781 = pi18 ? n5780 : n335;
  assign n5782 = pi23 ? n335 : n685;
  assign n5783 = pi22 ? n5782 : n32;
  assign n5784 = pi21 ? n5783 : n32;
  assign n5785 = pi20 ? n5784 : n32;
  assign n5786 = pi19 ? n5785 : n32;
  assign n5787 = pi18 ? n335 : n5786;
  assign n5788 = pi17 ? n5781 : n5787;
  assign n5789 = pi16 ? n439 : n5788;
  assign n5790 = pi15 ? n5777 : n5789;
  assign n5791 = pi14 ? n5765 : n5790;
  assign n5792 = pi13 ? n5740 : n5791;
  assign n5793 = pi12 ? n5675 : n5792;
  assign n5794 = pi11 ? n5492 : n5793;
  assign n5795 = pi19 ? n37 : n4981;
  assign n5796 = pi18 ? n37 : n5795;
  assign n5797 = pi18 ? n4985 : n4947;
  assign n5798 = pi17 ? n5796 : n5797;
  assign n5799 = pi16 ? n439 : n5798;
  assign n5800 = pi23 ? n335 : n2120;
  assign n5801 = pi22 ? n5800 : n32;
  assign n5802 = pi21 ? n5801 : n32;
  assign n5803 = pi20 ? n5802 : n32;
  assign n5804 = pi19 ? n5803 : n32;
  assign n5805 = pi18 ? n5002 : n5804;
  assign n5806 = pi17 ? n4994 : n5805;
  assign n5807 = pi16 ? n439 : n5806;
  assign n5808 = pi15 ? n5799 : n5807;
  assign n5809 = pi18 ? n5025 : n4104;
  assign n5810 = pi17 ? n5019 : n5809;
  assign n5811 = pi16 ? n439 : n5810;
  assign n5812 = pi23 ? n233 : n531;
  assign n5813 = pi22 ? n5812 : n32;
  assign n5814 = pi21 ? n5813 : n32;
  assign n5815 = pi20 ? n5814 : n32;
  assign n5816 = pi19 ? n5815 : n32;
  assign n5817 = pi18 ? n5030 : n5816;
  assign n5818 = pi17 ? n37 : n5817;
  assign n5819 = pi16 ? n439 : n5818;
  assign n5820 = pi15 ? n5811 : n5819;
  assign n5821 = pi14 ? n5808 : n5820;
  assign n5822 = pi18 ? n5037 : n4112;
  assign n5823 = pi17 ? n37 : n5822;
  assign n5824 = pi16 ? n439 : n5823;
  assign n5825 = pi15 ? n5824 : n5043;
  assign n5826 = pi18 ? n2102 : n4118;
  assign n5827 = pi17 ? n37 : n5826;
  assign n5828 = pi16 ? n439 : n5827;
  assign n5829 = pi22 ? n2192 : n32;
  assign n5830 = pi21 ? n5829 : n32;
  assign n5831 = pi20 ? n5830 : n32;
  assign n5832 = pi19 ? n5831 : n32;
  assign n5833 = pi18 ? n2109 : n5832;
  assign n5834 = pi17 ? n37 : n5833;
  assign n5835 = pi16 ? n439 : n5834;
  assign n5836 = pi15 ? n5828 : n5835;
  assign n5837 = pi14 ? n5825 : n5836;
  assign n5838 = pi13 ? n5821 : n5837;
  assign n5839 = pi18 ? n5057 : n2640;
  assign n5840 = pi17 ? n37 : n5839;
  assign n5841 = pi16 ? n439 : n5840;
  assign n5842 = pi15 ? n5841 : n5068;
  assign n5843 = pi18 ? n5073 : n2640;
  assign n5844 = pi17 ? n37 : n5843;
  assign n5845 = pi16 ? n439 : n5844;
  assign n5846 = pi18 ? n5079 : n2640;
  assign n5847 = pi17 ? n37 : n5846;
  assign n5848 = pi16 ? n439 : n5847;
  assign n5849 = pi15 ? n5845 : n5848;
  assign n5850 = pi14 ? n5842 : n5849;
  assign n5851 = pi18 ? n5087 : n2655;
  assign n5852 = pi17 ? n99 : n5851;
  assign n5853 = pi16 ? n721 : n5852;
  assign n5854 = pi18 ? n5093 : n2655;
  assign n5855 = pi17 ? n99 : n5854;
  assign n5856 = pi16 ? n744 : n5855;
  assign n5857 = pi15 ? n5853 : n5856;
  assign n5858 = pi18 ? n5104 : n1824;
  assign n5859 = pi17 ? n99 : n5858;
  assign n5860 = pi16 ? n744 : n5859;
  assign n5861 = pi15 ? n5090 : n5860;
  assign n5862 = pi14 ? n5857 : n5861;
  assign n5863 = pi13 ? n5850 : n5862;
  assign n5864 = pi12 ? n5838 : n5863;
  assign n5865 = pi16 ? n744 : n4187;
  assign n5866 = pi16 ? n744 : n5118;
  assign n5867 = pi15 ? n5865 : n5866;
  assign n5868 = pi18 ? n742 : n5122;
  assign n5869 = pi17 ? n32 : n5868;
  assign n5870 = pi16 ? n5869 : n5128;
  assign n5871 = pi22 ? n5167 : n158;
  assign n5872 = pi21 ? n5871 : n164;
  assign n5873 = pi20 ? n32 : n5872;
  assign n5874 = pi19 ? n32 : n5873;
  assign n5875 = pi22 ? n164 : n158;
  assign n5876 = pi21 ? n3010 : n5875;
  assign n5877 = pi22 ? n893 : n99;
  assign n5878 = pi21 ? n165 : n5877;
  assign n5879 = pi20 ? n5876 : n5878;
  assign n5880 = pi21 ? n165 : n168;
  assign n5881 = pi21 ? n164 : n168;
  assign n5882 = pi20 ? n5880 : n5881;
  assign n5883 = pi19 ? n5879 : n5882;
  assign n5884 = pi18 ? n5874 : n5883;
  assign n5885 = pi17 ? n32 : n5884;
  assign n5886 = pi21 ? n5875 : n3010;
  assign n5887 = pi21 ? n3013 : n3002;
  assign n5888 = pi20 ? n5886 : n5887;
  assign n5889 = pi21 ? n3002 : n777;
  assign n5890 = pi20 ? n5875 : n5889;
  assign n5891 = pi19 ? n5888 : n5890;
  assign n5892 = pi21 ? n165 : n3010;
  assign n5893 = pi21 ? n775 : n3013;
  assign n5894 = pi20 ? n5892 : n5893;
  assign n5895 = pi21 ? n168 : n3013;
  assign n5896 = pi20 ? n3011 : n5895;
  assign n5897 = pi19 ? n5894 : n5896;
  assign n5898 = pi18 ? n5891 : n5897;
  assign n5899 = pi22 ? n158 : n157;
  assign n5900 = pi21 ? n3002 : n5899;
  assign n5901 = pi21 ? n165 : n777;
  assign n5902 = pi20 ? n5900 : n5901;
  assign n5903 = pi19 ? n5902 : n5147;
  assign n5904 = pi18 ? n5903 : n32;
  assign n5905 = pi17 ? n5898 : n5904;
  assign n5906 = pi16 ? n5885 : n5905;
  assign n5907 = pi15 ? n5870 : n5906;
  assign n5908 = pi14 ? n5867 : n5907;
  assign n5909 = pi18 ? n5171 : n157;
  assign n5910 = pi17 ? n32 : n5909;
  assign n5911 = pi16 ? n5910 : n5165;
  assign n5912 = pi15 ? n5911 : n5184;
  assign n5913 = pi22 ? n962 : n918;
  assign n5914 = pi21 ? n5913 : n1793;
  assign n5915 = pi20 ? n32 : n5914;
  assign n5916 = pi19 ? n32 : n5915;
  assign n5917 = pi20 ? n2872 : n5215;
  assign n5918 = pi19 ? n5917 : n5218;
  assign n5919 = pi18 ? n5916 : n5918;
  assign n5920 = pi17 ? n32 : n5919;
  assign n5921 = pi21 ? n919 : n921;
  assign n5922 = pi20 ? n5222 : n5921;
  assign n5923 = pi21 ? n921 : n2863;
  assign n5924 = pi20 ? n921 : n5923;
  assign n5925 = pi19 ? n5922 : n5924;
  assign n5926 = pi21 ? n2876 : n916;
  assign n5927 = pi20 ? n5926 : n919;
  assign n5928 = pi20 ? n5229 : n919;
  assign n5929 = pi19 ? n5927 : n5928;
  assign n5930 = pi18 ? n5925 : n5929;
  assign n5931 = pi21 ? n2863 : n1039;
  assign n5932 = pi20 ? n5923 : n5931;
  assign n5933 = pi19 ? n5932 : n5237;
  assign n5934 = pi18 ? n5933 : n32;
  assign n5935 = pi17 ? n5930 : n5934;
  assign n5936 = pi16 ? n5920 : n5935;
  assign n5937 = pi15 ? n5210 : n5936;
  assign n5938 = pi14 ? n5912 : n5937;
  assign n5939 = pi13 ? n5908 : n5938;
  assign n5940 = pi22 ? n2401 : n706;
  assign n5941 = pi21 ? n316 : n5940;
  assign n5942 = pi20 ? n4437 : n5941;
  assign n5943 = pi19 ? n3578 : n5942;
  assign n5944 = pi18 ? n5943 : n32;
  assign n5945 = pi17 ? n139 : n5944;
  assign n5946 = pi16 ? n2810 : n5945;
  assign n5947 = pi22 ? n909 : n348;
  assign n5948 = pi21 ? n5947 : n4017;
  assign n5949 = pi20 ? n32 : n5948;
  assign n5950 = pi19 ? n32 : n5949;
  assign n5951 = pi21 ? n354 : n1774;
  assign n5952 = pi21 ? n392 : n390;
  assign n5953 = pi20 ? n5951 : n5952;
  assign n5954 = pi21 ? n1777 : n424;
  assign n5955 = pi21 ? n4017 : n424;
  assign n5956 = pi20 ? n5954 : n5955;
  assign n5957 = pi19 ? n5953 : n5956;
  assign n5958 = pi18 ? n5950 : n5957;
  assign n5959 = pi17 ? n32 : n5958;
  assign n5960 = pi21 ? n4424 : n4429;
  assign n5961 = pi21 ? n349 : n3617;
  assign n5962 = pi20 ? n5960 : n5961;
  assign n5963 = pi21 ? n356 : n4780;
  assign n5964 = pi20 ? n4020 : n5963;
  assign n5965 = pi19 ? n5962 : n5964;
  assign n5966 = pi21 ? n392 : n354;
  assign n5967 = pi21 ? n346 : n4421;
  assign n5968 = pi20 ? n5966 : n5967;
  assign n5969 = pi21 ? n3617 : n4014;
  assign n5970 = pi21 ? n424 : n4421;
  assign n5971 = pi20 ? n5969 : n5970;
  assign n5972 = pi19 ? n5968 : n5971;
  assign n5973 = pi18 ? n5965 : n5972;
  assign n5974 = pi20 ? n4433 : n4430;
  assign n5975 = pi19 ? n5974 : n5276;
  assign n5976 = pi18 ? n5975 : n32;
  assign n5977 = pi17 ? n5973 : n5976;
  assign n5978 = pi16 ? n5959 : n5977;
  assign n5979 = pi15 ? n5946 : n5978;
  assign n5980 = pi14 ? n5979 : n5310;
  assign n5981 = pi18 ? n329 : n5313;
  assign n5982 = pi17 ? n32 : n5981;
  assign n5983 = pi16 ? n5982 : n5324;
  assign n5984 = pi15 ? n5983 : n5348;
  assign n5985 = pi21 ? n4485 : n204;
  assign n5986 = pi20 ? n32 : n5985;
  assign n5987 = pi19 ? n32 : n5986;
  assign n5988 = pi18 ? n5987 : n204;
  assign n5989 = pi17 ? n32 : n5988;
  assign n5990 = pi21 ? n204 : n5829;
  assign n5991 = pi20 ? n204 : n5990;
  assign n5992 = pi19 ? n204 : n5991;
  assign n5993 = pi18 ? n5992 : n32;
  assign n5994 = pi17 ? n204 : n5993;
  assign n5995 = pi16 ? n5989 : n5994;
  assign n5996 = pi23 ? n714 : n335;
  assign n5997 = pi22 ? n5996 : n204;
  assign n5998 = pi21 ? n5997 : n204;
  assign n5999 = pi20 ? n32 : n5998;
  assign n6000 = pi19 ? n32 : n5999;
  assign n6001 = pi18 ? n6000 : n5366;
  assign n6002 = pi17 ? n32 : n6001;
  assign n6003 = pi21 ? n204 : n928;
  assign n6004 = pi20 ? n204 : n6003;
  assign n6005 = pi19 ? n204 : n6004;
  assign n6006 = pi18 ? n6005 : n32;
  assign n6007 = pi17 ? n204 : n6006;
  assign n6008 = pi16 ? n6002 : n6007;
  assign n6009 = pi15 ? n5995 : n6008;
  assign n6010 = pi14 ? n5984 : n6009;
  assign n6011 = pi13 ? n5980 : n6010;
  assign n6012 = pi12 ? n5939 : n6011;
  assign n6013 = pi11 ? n5864 : n6012;
  assign n6014 = pi10 ? n5794 : n6013;
  assign n6015 = pi09 ? n32 : n6014;
  assign n6016 = pi08 ? n5383 : n6015;
  assign n6017 = pi16 ? n3784 : n4532;
  assign n6018 = pi16 ? n70 : n4532;
  assign n6019 = pi15 ? n6017 : n6018;
  assign n6020 = pi16 ? n5390 : n4532;
  assign n6021 = pi16 ? n73 : n4532;
  assign n6022 = pi15 ? n6020 : n6021;
  assign n6023 = pi14 ? n6019 : n6022;
  assign n6024 = pi16 ? n83 : n5400;
  assign n6025 = pi16 ? n1130 : n5400;
  assign n6026 = pi15 ? n6024 : n6025;
  assign n6027 = pi23 ? n37 : n5630;
  assign n6028 = pi22 ? n37 : n6027;
  assign n6029 = pi21 ? n6028 : n32;
  assign n6030 = pi20 ? n6029 : n32;
  assign n6031 = pi19 ? n6030 : n32;
  assign n6032 = pi18 ? n37 : n6031;
  assign n6033 = pi17 ? n37 : n6032;
  assign n6034 = pi16 ? n2461 : n6033;
  assign n6035 = pi16 ? n439 : n6033;
  assign n6036 = pi15 ? n6034 : n6035;
  assign n6037 = pi14 ? n6026 : n6036;
  assign n6038 = pi13 ? n6023 : n6037;
  assign n6039 = pi20 ? n2167 : n3805;
  assign n6040 = pi19 ? n4616 : n6039;
  assign n6041 = pi18 ? n184 : n6040;
  assign n6042 = pi17 ? n32 : n6041;
  assign n6043 = pi21 ? n2164 : n2162;
  assign n6044 = pi21 ? n2161 : n112;
  assign n6045 = pi20 ? n6043 : n6044;
  assign n6046 = pi20 ? n5405 : n99;
  assign n6047 = pi19 ? n6045 : n6046;
  assign n6048 = pi18 ? n6047 : n99;
  assign n6049 = pi19 ? n99 : n2191;
  assign n6050 = pi21 ? n1168 : n32;
  assign n6051 = pi20 ? n6050 : n32;
  assign n6052 = pi19 ? n6051 : n32;
  assign n6053 = pi18 ? n6049 : n6052;
  assign n6054 = pi17 ? n6048 : n6053;
  assign n6055 = pi16 ? n6042 : n6054;
  assign n6056 = pi18 ? n99 : n6052;
  assign n6057 = pi17 ? n99 : n6056;
  assign n6058 = pi16 ? n201 : n6057;
  assign n6059 = pi15 ? n6055 : n6058;
  assign n6060 = pi21 ? n1186 : n32;
  assign n6061 = pi20 ? n6060 : n32;
  assign n6062 = pi19 ? n6061 : n32;
  assign n6063 = pi18 ? n99 : n6062;
  assign n6064 = pi17 ? n99 : n6063;
  assign n6065 = pi16 ? n801 : n6064;
  assign n6066 = pi16 ? n721 : n6064;
  assign n6067 = pi15 ? n6065 : n6066;
  assign n6068 = pi14 ? n6059 : n6067;
  assign n6069 = pi23 ? n139 : n624;
  assign n6070 = pi22 ? n99 : n6069;
  assign n6071 = pi21 ? n6070 : n32;
  assign n6072 = pi20 ? n6071 : n32;
  assign n6073 = pi19 ? n6072 : n32;
  assign n6074 = pi18 ? n99 : n6073;
  assign n6075 = pi17 ? n99 : n6074;
  assign n6076 = pi16 ? n721 : n6075;
  assign n6077 = pi23 ? n335 : n624;
  assign n6078 = pi22 ? n99 : n6077;
  assign n6079 = pi21 ? n6078 : n32;
  assign n6080 = pi20 ? n6079 : n32;
  assign n6081 = pi19 ? n6080 : n32;
  assign n6082 = pi18 ? n99 : n6081;
  assign n6083 = pi17 ? n99 : n6082;
  assign n6084 = pi16 ? n721 : n6083;
  assign n6085 = pi15 ? n6076 : n6084;
  assign n6086 = pi19 ? n99 : n5468;
  assign n6087 = pi21 ? n5464 : n5458;
  assign n6088 = pi20 ? n5465 : n6087;
  assign n6089 = pi22 ? n685 : n99;
  assign n6090 = pi21 ? n99 : n6089;
  assign n6091 = pi20 ? n99 : n6090;
  assign n6092 = pi19 ? n6088 : n6091;
  assign n6093 = pi18 ? n6086 : n6092;
  assign n6094 = pi22 ? n685 : n3443;
  assign n6095 = pi21 ? n99 : n6094;
  assign n6096 = pi22 ? n5452 : n3443;
  assign n6097 = pi21 ? n99 : n6096;
  assign n6098 = pi20 ? n6095 : n6097;
  assign n6099 = pi21 ? n5453 : n99;
  assign n6100 = pi19 ? n6098 : n6099;
  assign n6101 = pi21 ? n767 : n32;
  assign n6102 = pi20 ? n6101 : n32;
  assign n6103 = pi19 ? n6102 : n32;
  assign n6104 = pi18 ? n6100 : n6103;
  assign n6105 = pi17 ? n6093 : n6104;
  assign n6106 = pi16 ? n721 : n6105;
  assign n6107 = pi23 ? n714 : n157;
  assign n6108 = pi22 ? n6107 : n37;
  assign n6109 = pi21 ? n6108 : n157;
  assign n6110 = pi20 ? n32 : n6109;
  assign n6111 = pi19 ? n32 : n6110;
  assign n6112 = pi18 ? n6111 : n157;
  assign n6113 = pi17 ? n32 : n6112;
  assign n6114 = pi23 ? n157 : n1149;
  assign n6115 = pi22 ? n157 : n6114;
  assign n6116 = pi21 ? n6115 : n32;
  assign n6117 = pi20 ? n6116 : n32;
  assign n6118 = pi19 ? n6117 : n32;
  assign n6119 = pi18 ? n157 : n6118;
  assign n6120 = pi17 ? n157 : n6119;
  assign n6121 = pi16 ? n6113 : n6120;
  assign n6122 = pi15 ? n6106 : n6121;
  assign n6123 = pi14 ? n6085 : n6122;
  assign n6124 = pi13 ? n6068 : n6123;
  assign n6125 = pi12 ? n6038 : n6124;
  assign n6126 = pi22 ? n5167 : n37;
  assign n6127 = pi21 ? n6126 : n157;
  assign n6128 = pi20 ? n32 : n6127;
  assign n6129 = pi19 ? n32 : n6128;
  assign n6130 = pi18 ? n6129 : n157;
  assign n6131 = pi17 ? n32 : n6130;
  assign n6132 = pi22 ? n157 : n1484;
  assign n6133 = pi21 ? n6132 : n32;
  assign n6134 = pi20 ? n6133 : n32;
  assign n6135 = pi19 ? n6134 : n32;
  assign n6136 = pi18 ? n157 : n6135;
  assign n6137 = pi17 ? n157 : n6136;
  assign n6138 = pi16 ? n6131 : n6137;
  assign n6139 = pi21 ? n180 : n157;
  assign n6140 = pi20 ? n32 : n6139;
  assign n6141 = pi19 ? n32 : n6140;
  assign n6142 = pi18 ? n6141 : n157;
  assign n6143 = pi17 ? n32 : n6142;
  assign n6144 = pi19 ? n254 : n157;
  assign n6145 = pi18 ? n157 : n6144;
  assign n6146 = pi23 ? n157 : n395;
  assign n6147 = pi22 ? n157 : n6146;
  assign n6148 = pi21 ? n6147 : n32;
  assign n6149 = pi20 ? n6148 : n32;
  assign n6150 = pi19 ? n6149 : n32;
  assign n6151 = pi18 ? n5173 : n6150;
  assign n6152 = pi17 ? n6145 : n6151;
  assign n6153 = pi16 ? n6143 : n6152;
  assign n6154 = pi15 ? n6138 : n6153;
  assign n6155 = pi21 ? n180 : n204;
  assign n6156 = pi20 ? n32 : n6155;
  assign n6157 = pi19 ? n32 : n6156;
  assign n6158 = pi21 ? n204 : n916;
  assign n6159 = pi20 ? n5199 : n6158;
  assign n6160 = pi19 ? n204 : n6159;
  assign n6161 = pi18 ? n6157 : n6160;
  assign n6162 = pi17 ? n32 : n6161;
  assign n6163 = pi20 ? n5204 : n204;
  assign n6164 = pi20 ? n5921 : n1794;
  assign n6165 = pi19 ? n6163 : n6164;
  assign n6166 = pi20 ? n1794 : n5921;
  assign n6167 = pi21 ? n2869 : n916;
  assign n6168 = pi20 ? n1026 : n6167;
  assign n6169 = pi19 ? n6166 : n6168;
  assign n6170 = pi18 ? n6165 : n6169;
  assign n6171 = pi21 ? n2869 : n139;
  assign n6172 = pi21 ? n916 : n2869;
  assign n6173 = pi20 ? n6171 : n6172;
  assign n6174 = pi21 ? n2876 : n921;
  assign n6175 = pi20 ? n5215 : n6174;
  assign n6176 = pi19 ? n6173 : n6175;
  assign n6177 = pi22 ? n918 : n430;
  assign n6178 = pi21 ? n6177 : n32;
  assign n6179 = pi20 ? n6178 : n32;
  assign n6180 = pi19 ? n6179 : n32;
  assign n6181 = pi18 ? n6176 : n6180;
  assign n6182 = pi17 ? n6170 : n6181;
  assign n6183 = pi16 ? n6162 : n6182;
  assign n6184 = pi22 ? n139 : n2564;
  assign n6185 = pi21 ? n6184 : n32;
  assign n6186 = pi20 ? n6185 : n32;
  assign n6187 = pi19 ? n6186 : n32;
  assign n6188 = pi18 ? n139 : n6187;
  assign n6189 = pi17 ? n139 : n6188;
  assign n6190 = pi16 ? n314 : n6189;
  assign n6191 = pi15 ? n6183 : n6190;
  assign n6192 = pi14 ? n6154 : n6191;
  assign n6193 = pi16 ? n1773 : n6189;
  assign n6194 = pi22 ? n204 : n2564;
  assign n6195 = pi21 ? n6194 : n32;
  assign n6196 = pi20 ? n6195 : n32;
  assign n6197 = pi19 ? n6196 : n32;
  assign n6198 = pi18 ? n139 : n6197;
  assign n6199 = pi17 ? n139 : n6198;
  assign n6200 = pi16 ? n1773 : n6199;
  assign n6201 = pi15 ? n6193 : n6200;
  assign n6202 = pi20 ? n5273 : n2513;
  assign n6203 = pi19 ? n6202 : n2520;
  assign n6204 = pi18 ? n990 : n6203;
  assign n6205 = pi17 ? n32 : n6204;
  assign n6206 = pi20 ? n2510 : n2512;
  assign n6207 = pi19 ? n6206 : n5273;
  assign n6208 = pi21 ? n3617 : n139;
  assign n6209 = pi20 ? n6208 : n1008;
  assign n6210 = pi20 ? n2513 : n1531;
  assign n6211 = pi19 ? n6209 : n6210;
  assign n6212 = pi18 ? n6207 : n6211;
  assign n6213 = pi19 ? n1720 : n976;
  assign n6214 = pi21 ? n336 : n32;
  assign n6215 = pi20 ? n6214 : n32;
  assign n6216 = pi19 ? n6215 : n32;
  assign n6217 = pi18 ? n6213 : n6216;
  assign n6218 = pi17 ? n6212 : n6217;
  assign n6219 = pi16 ? n6205 : n6218;
  assign n6220 = pi21 ? n3986 : n316;
  assign n6221 = pi20 ? n32 : n6220;
  assign n6222 = pi19 ? n32 : n6221;
  assign n6223 = pi18 ? n6222 : n316;
  assign n6224 = pi17 ? n32 : n6223;
  assign n6225 = pi18 ? n316 : n5669;
  assign n6226 = pi17 ? n316 : n6225;
  assign n6227 = pi16 ? n6224 : n6226;
  assign n6228 = pi15 ? n6219 : n6227;
  assign n6229 = pi14 ? n6201 : n6228;
  assign n6230 = pi13 ? n6192 : n6229;
  assign n6231 = pi21 ? n180 : n316;
  assign n6232 = pi20 ? n32 : n6231;
  assign n6233 = pi19 ? n32 : n6232;
  assign n6234 = pi18 ? n6233 : n316;
  assign n6235 = pi17 ? n32 : n6234;
  assign n6236 = pi16 ? n6235 : n6226;
  assign n6237 = pi21 ? n180 : n424;
  assign n6238 = pi20 ? n32 : n6237;
  assign n6239 = pi19 ? n32 : n6238;
  assign n6240 = pi20 ? n5689 : n3697;
  assign n6241 = pi21 ? n316 : n3258;
  assign n6242 = pi20 ? n5299 : n6241;
  assign n6243 = pi19 ? n6240 : n6242;
  assign n6244 = pi18 ? n6239 : n6243;
  assign n6245 = pi17 ? n32 : n6244;
  assign n6246 = pi16 ? n6245 : n6226;
  assign n6247 = pi15 ? n6236 : n6246;
  assign n6248 = pi21 ? n180 : n1309;
  assign n6249 = pi20 ? n32 : n6248;
  assign n6250 = pi19 ? n32 : n6249;
  assign n6251 = pi20 ? n2634 : n508;
  assign n6252 = pi21 ? n516 : n1046;
  assign n6253 = pi20 ? n513 : n6252;
  assign n6254 = pi19 ? n6251 : n6253;
  assign n6255 = pi18 ? n6250 : n6254;
  assign n6256 = pi17 ? n32 : n6255;
  assign n6257 = pi18 ? n204 : n6197;
  assign n6258 = pi17 ? n204 : n6257;
  assign n6259 = pi16 ? n6256 : n6258;
  assign n6260 = pi21 ? n1313 : n499;
  assign n6261 = pi20 ? n37 : n6260;
  assign n6262 = pi19 ? n37 : n6261;
  assign n6263 = pi18 ? n374 : n6262;
  assign n6264 = pi17 ? n32 : n6263;
  assign n6265 = pi21 ? n455 : n204;
  assign n6266 = pi20 ? n6265 : n1057;
  assign n6267 = pi19 ? n6266 : n1919;
  assign n6268 = pi20 ? n1582 : n204;
  assign n6269 = pi18 ? n6267 : n6268;
  assign n6270 = pi22 ? n204 : n664;
  assign n6271 = pi21 ? n6270 : n32;
  assign n6272 = pi20 ? n6271 : n32;
  assign n6273 = pi19 ? n6272 : n32;
  assign n6274 = pi18 ? n204 : n6273;
  assign n6275 = pi17 ? n6269 : n6274;
  assign n6276 = pi16 ? n6264 : n6275;
  assign n6277 = pi15 ? n6259 : n6276;
  assign n6278 = pi14 ? n6247 : n6277;
  assign n6279 = pi21 ? n37 : n559;
  assign n6280 = pi21 ? n4891 : n3409;
  assign n6281 = pi20 ? n6279 : n6280;
  assign n6282 = pi21 ? n4893 : n3409;
  assign n6283 = pi20 ? n6282 : n4916;
  assign n6284 = pi19 ? n6281 : n6283;
  assign n6285 = pi21 ? n4908 : n4899;
  assign n6286 = pi21 ? n4893 : n4899;
  assign n6287 = pi20 ? n6285 : n6286;
  assign n6288 = pi19 ? n4915 : n6287;
  assign n6289 = pi18 ? n6284 : n6288;
  assign n6290 = pi21 ? n4908 : n4900;
  assign n6291 = pi20 ? n4916 : n6290;
  assign n6292 = pi21 ? n4902 : n4900;
  assign n6293 = pi19 ? n6291 : n6292;
  assign n6294 = pi22 ? n2060 : n1407;
  assign n6295 = pi21 ? n6294 : n32;
  assign n6296 = pi20 ? n6295 : n32;
  assign n6297 = pi19 ? n6296 : n32;
  assign n6298 = pi18 ? n6293 : n6297;
  assign n6299 = pi17 ? n6289 : n6298;
  assign n6300 = pi16 ? n439 : n6299;
  assign n6301 = pi21 ? n2007 : n580;
  assign n6302 = pi20 ? n37 : n6301;
  assign n6303 = pi21 ? n583 : n566;
  assign n6304 = pi21 ? n4938 : n580;
  assign n6305 = pi20 ? n6303 : n6304;
  assign n6306 = pi19 ? n6302 : n6305;
  assign n6307 = pi20 ? n581 : n604;
  assign n6308 = pi19 ? n6307 : n581;
  assign n6309 = pi18 ? n6306 : n6308;
  assign n6310 = pi20 ? n4991 : n1893;
  assign n6311 = pi21 ? n569 : n567;
  assign n6312 = pi21 ? n580 : n567;
  assign n6313 = pi20 ? n6311 : n6312;
  assign n6314 = pi19 ? n6310 : n6313;
  assign n6315 = pi22 ? n2060 : n317;
  assign n6316 = pi21 ? n6315 : n32;
  assign n6317 = pi20 ? n6316 : n32;
  assign n6318 = pi19 ? n6317 : n32;
  assign n6319 = pi18 ? n6314 : n6318;
  assign n6320 = pi17 ? n6309 : n6319;
  assign n6321 = pi16 ? n439 : n6320;
  assign n6322 = pi15 ? n6300 : n6321;
  assign n6323 = pi20 ? n4971 : n3292;
  assign n6324 = pi21 ? n567 : n570;
  assign n6325 = pi20 ? n37 : n6324;
  assign n6326 = pi19 ? n6323 : n6325;
  assign n6327 = pi18 ? n37 : n6326;
  assign n6328 = pi20 ? n647 : n1893;
  assign n6329 = pi20 ? n569 : n605;
  assign n6330 = pi19 ? n6328 : n6329;
  assign n6331 = pi22 ? n2060 : n688;
  assign n6332 = pi21 ? n6331 : n32;
  assign n6333 = pi20 ? n6332 : n32;
  assign n6334 = pi19 ? n6333 : n32;
  assign n6335 = pi18 ? n6330 : n6334;
  assign n6336 = pi17 ? n6327 : n6335;
  assign n6337 = pi16 ? n439 : n6336;
  assign n6338 = pi19 ? n37 : n3332;
  assign n6339 = pi18 ? n37 : n6338;
  assign n6340 = pi20 ? n647 : n37;
  assign n6341 = pi20 ? n649 : n605;
  assign n6342 = pi19 ? n6340 : n6341;
  assign n6343 = pi22 ? n5782 : n706;
  assign n6344 = pi21 ? n6343 : n32;
  assign n6345 = pi20 ? n6344 : n32;
  assign n6346 = pi19 ? n6345 : n32;
  assign n6347 = pi18 ? n6342 : n6346;
  assign n6348 = pi17 ? n6339 : n6347;
  assign n6349 = pi16 ? n439 : n6348;
  assign n6350 = pi15 ? n6337 : n6349;
  assign n6351 = pi14 ? n6322 : n6350;
  assign n6352 = pi13 ? n6278 : n6351;
  assign n6353 = pi12 ? n6230 : n6352;
  assign n6354 = pi11 ? n6125 : n6353;
  assign n6355 = pi20 ? n37 : n2049;
  assign n6356 = pi19 ? n37 : n6355;
  assign n6357 = pi18 ? n37 : n6356;
  assign n6358 = pi21 ? n233 : n37;
  assign n6359 = pi20 ? n6358 : n37;
  assign n6360 = pi21 ? n37 : n3409;
  assign n6361 = pi22 ? n233 : n335;
  assign n6362 = pi21 ? n6361 : n233;
  assign n6363 = pi20 ? n6360 : n6362;
  assign n6364 = pi19 ? n6359 : n6363;
  assign n6365 = pi23 ? n233 : n685;
  assign n6366 = pi22 ? n6365 : n706;
  assign n6367 = pi21 ? n6366 : n32;
  assign n6368 = pi20 ? n6367 : n32;
  assign n6369 = pi19 ? n6368 : n32;
  assign n6370 = pi18 ? n6364 : n6369;
  assign n6371 = pi17 ? n6357 : n6370;
  assign n6372 = pi16 ? n439 : n6371;
  assign n6373 = pi20 ? n37 : n639;
  assign n6374 = pi19 ? n37 : n6373;
  assign n6375 = pi18 ? n37 : n6374;
  assign n6376 = pi22 ? n335 : n233;
  assign n6377 = pi21 ? n335 : n6376;
  assign n6378 = pi20 ? n2094 : n6377;
  assign n6379 = pi19 ? n6359 : n6378;
  assign n6380 = pi23 ? n335 : n316;
  assign n6381 = pi22 ? n6380 : n32;
  assign n6382 = pi21 ? n6381 : n32;
  assign n6383 = pi20 ? n6382 : n32;
  assign n6384 = pi19 ? n6383 : n32;
  assign n6385 = pi18 ? n6379 : n6384;
  assign n6386 = pi17 ? n6375 : n6385;
  assign n6387 = pi16 ? n439 : n6386;
  assign n6388 = pi15 ? n6372 : n6387;
  assign n6389 = pi21 ? n4891 : n37;
  assign n6390 = pi20 ? n6389 : n37;
  assign n6391 = pi20 ? n2094 : n233;
  assign n6392 = pi19 ? n6390 : n6391;
  assign n6393 = pi23 ? n363 : n2120;
  assign n6394 = pi22 ? n6393 : n32;
  assign n6395 = pi21 ? n6394 : n32;
  assign n6396 = pi20 ? n6395 : n32;
  assign n6397 = pi19 ? n6396 : n32;
  assign n6398 = pi18 ? n6392 : n6397;
  assign n6399 = pi17 ? n2115 : n6398;
  assign n6400 = pi16 ? n439 : n6399;
  assign n6401 = pi22 ? n37 : n5011;
  assign n6402 = pi21 ? n37 : n6401;
  assign n6403 = pi20 ? n37 : n6402;
  assign n6404 = pi19 ? n37 : n6403;
  assign n6405 = pi23 ? n363 : n624;
  assign n6406 = pi22 ? n6405 : n32;
  assign n6407 = pi21 ? n6406 : n32;
  assign n6408 = pi20 ? n6407 : n32;
  assign n6409 = pi19 ? n6408 : n32;
  assign n6410 = pi18 ? n6404 : n6409;
  assign n6411 = pi17 ? n37 : n6410;
  assign n6412 = pi16 ? n439 : n6411;
  assign n6413 = pi15 ? n6400 : n6412;
  assign n6414 = pi14 ? n6388 : n6413;
  assign n6415 = pi23 ? n233 : n687;
  assign n6416 = pi22 ? n6415 : n32;
  assign n6417 = pi21 ? n6416 : n32;
  assign n6418 = pi20 ? n6417 : n32;
  assign n6419 = pi19 ? n6418 : n32;
  assign n6420 = pi18 ? n2102 : n6419;
  assign n6421 = pi17 ? n37 : n6420;
  assign n6422 = pi16 ? n439 : n6421;
  assign n6423 = pi15 ? n6422 : n5835;
  assign n6424 = pi14 ? n5043 : n6423;
  assign n6425 = pi13 ? n6414 : n6424;
  assign n6426 = pi22 ? n363 : n893;
  assign n6427 = pi21 ? n37 : n6426;
  assign n6428 = pi20 ? n37 : n6427;
  assign n6429 = pi19 ? n37 : n6428;
  assign n6430 = pi18 ? n6429 : n2640;
  assign n6431 = pi17 ? n37 : n6430;
  assign n6432 = pi16 ? n439 : n6431;
  assign n6433 = pi22 ? n37 : n893;
  assign n6434 = pi21 ? n37 : n6433;
  assign n6435 = pi20 ? n37 : n6434;
  assign n6436 = pi19 ? n37 : n6435;
  assign n6437 = pi18 ? n6436 : n2640;
  assign n6438 = pi17 ? n37 : n6437;
  assign n6439 = pi16 ? n439 : n6438;
  assign n6440 = pi15 ? n6432 : n6439;
  assign n6441 = pi22 ? n37 : n3961;
  assign n6442 = pi21 ? n37 : n6441;
  assign n6443 = pi20 ? n37 : n6442;
  assign n6444 = pi19 ? n37 : n6443;
  assign n6445 = pi18 ? n6444 : n2640;
  assign n6446 = pi17 ? n37 : n6445;
  assign n6447 = pi16 ? n439 : n6446;
  assign n6448 = pi21 ? n722 : n2721;
  assign n6449 = pi20 ? n99 : n6448;
  assign n6450 = pi19 ? n99 : n6449;
  assign n6451 = pi18 ? n6450 : n2640;
  assign n6452 = pi17 ? n99 : n6451;
  assign n6453 = pi16 ? n744 : n6452;
  assign n6454 = pi15 ? n6447 : n6453;
  assign n6455 = pi14 ? n6440 : n6454;
  assign n6456 = pi16 ? n744 : n5852;
  assign n6457 = pi15 ? n6456 : n5856;
  assign n6458 = pi18 ? n5087 : n2703;
  assign n6459 = pi17 ? n99 : n6458;
  assign n6460 = pi16 ? n744 : n6459;
  assign n6461 = pi22 ? n157 : n685;
  assign n6462 = pi21 ? n99 : n6461;
  assign n6463 = pi20 ? n99 : n6462;
  assign n6464 = pi19 ? n99 : n6463;
  assign n6465 = pi18 ? n6464 : n2703;
  assign n6466 = pi17 ? n99 : n6465;
  assign n6467 = pi16 ? n744 : n6466;
  assign n6468 = pi15 ? n6460 : n6467;
  assign n6469 = pi14 ? n6457 : n6468;
  assign n6470 = pi13 ? n6455 : n6469;
  assign n6471 = pi12 ? n6425 : n6470;
  assign n6472 = pi22 ? n738 : n112;
  assign n6473 = pi21 ? n6472 : n2746;
  assign n6474 = pi20 ? n32 : n6473;
  assign n6475 = pi19 ? n32 : n6474;
  assign n6476 = pi20 ? n2749 : n2174;
  assign n6477 = pi21 ? n181 : n2164;
  assign n6478 = pi20 ? n6477 : n2962;
  assign n6479 = pi19 ? n6476 : n6478;
  assign n6480 = pi18 ? n6475 : n6479;
  assign n6481 = pi17 ? n32 : n6480;
  assign n6482 = pi20 ? n2752 : n99;
  assign n6483 = pi20 ? n2164 : n99;
  assign n6484 = pi19 ? n6482 : n6483;
  assign n6485 = pi20 ? n3812 : n99;
  assign n6486 = pi20 ? n99 : n3888;
  assign n6487 = pi19 ? n6485 : n6486;
  assign n6488 = pi18 ? n6484 : n6487;
  assign n6489 = pi20 ? n99 : n2191;
  assign n6490 = pi21 ? n168 : n777;
  assign n6491 = pi21 ? n775 : n685;
  assign n6492 = pi20 ? n6490 : n6491;
  assign n6493 = pi19 ? n6489 : n6492;
  assign n6494 = pi18 ? n6493 : n1824;
  assign n6495 = pi17 ? n6488 : n6494;
  assign n6496 = pi16 ? n6481 : n6495;
  assign n6497 = pi21 ? n716 : n157;
  assign n6498 = pi20 ? n32 : n6497;
  assign n6499 = pi19 ? n32 : n6498;
  assign n6500 = pi21 ? n777 : n775;
  assign n6501 = pi20 ? n6500 : n157;
  assign n6502 = pi21 ? n2998 : n157;
  assign n6503 = pi21 ? n775 : n777;
  assign n6504 = pi20 ? n6502 : n6503;
  assign n6505 = pi19 ? n6501 : n6504;
  assign n6506 = pi18 ? n6499 : n6505;
  assign n6507 = pi17 ? n32 : n6506;
  assign n6508 = pi21 ? n157 : n777;
  assign n6509 = pi20 ? n6508 : n157;
  assign n6510 = pi19 ? n6509 : n157;
  assign n6511 = pi18 ? n6510 : n157;
  assign n6512 = pi20 ? n157 : n775;
  assign n6513 = pi20 ? n6508 : n5114;
  assign n6514 = pi19 ? n6512 : n6513;
  assign n6515 = pi18 ? n6514 : n1824;
  assign n6516 = pi17 ? n6511 : n6515;
  assign n6517 = pi16 ? n6507 : n6516;
  assign n6518 = pi15 ? n6496 : n6517;
  assign n6519 = pi22 ? n715 : n157;
  assign n6520 = pi21 ? n6519 : n775;
  assign n6521 = pi20 ? n32 : n6520;
  assign n6522 = pi19 ? n32 : n6521;
  assign n6523 = pi21 ? n775 : n157;
  assign n6524 = pi20 ? n787 : n6523;
  assign n6525 = pi19 ? n6509 : n6524;
  assign n6526 = pi18 ? n6522 : n6525;
  assign n6527 = pi17 ? n32 : n6526;
  assign n6528 = pi20 ? n157 : n6500;
  assign n6529 = pi20 ? n157 : n6523;
  assign n6530 = pi19 ? n6528 : n6529;
  assign n6531 = pi20 ? n157 : n787;
  assign n6532 = pi20 ? n6523 : n157;
  assign n6533 = pi19 ? n6531 : n6532;
  assign n6534 = pi18 ? n6530 : n6533;
  assign n6535 = pi22 ? n157 : n396;
  assign n6536 = pi21 ? n777 : n6535;
  assign n6537 = pi20 ? n6523 : n6536;
  assign n6538 = pi19 ? n6532 : n6537;
  assign n6539 = pi18 ? n6538 : n32;
  assign n6540 = pi17 ? n6534 : n6539;
  assign n6541 = pi16 ? n6527 : n6540;
  assign n6542 = pi20 ? n99 : n787;
  assign n6543 = pi21 ? n157 : n6535;
  assign n6544 = pi20 ? n157 : n6543;
  assign n6545 = pi19 ? n6542 : n6544;
  assign n6546 = pi18 ? n6545 : n32;
  assign n6547 = pi17 ? n99 : n6546;
  assign n6548 = pi16 ? n744 : n6547;
  assign n6549 = pi15 ? n6541 : n6548;
  assign n6550 = pi14 ? n6518 : n6549;
  assign n6551 = pi22 ? n909 : n157;
  assign n6552 = pi21 ? n6551 : n157;
  assign n6553 = pi20 ? n32 : n6552;
  assign n6554 = pi19 ? n32 : n6553;
  assign n6555 = pi18 ? n6554 : n157;
  assign n6556 = pi17 ? n32 : n6555;
  assign n6557 = pi19 ? n157 : n6544;
  assign n6558 = pi18 ? n6557 : n32;
  assign n6559 = pi17 ? n157 : n6558;
  assign n6560 = pi16 ? n6556 : n6559;
  assign n6561 = pi21 ? n204 : n397;
  assign n6562 = pi20 ? n5199 : n6561;
  assign n6563 = pi19 ? n2317 : n6562;
  assign n6564 = pi18 ? n6563 : n32;
  assign n6565 = pi17 ? n139 : n6564;
  assign n6566 = pi16 ? n915 : n6565;
  assign n6567 = pi15 ? n6560 : n6566;
  assign n6568 = pi21 ? n139 : n921;
  assign n6569 = pi20 ? n6568 : n927;
  assign n6570 = pi19 ? n6569 : n139;
  assign n6571 = pi18 ? n913 : n6570;
  assign n6572 = pi17 ? n32 : n6571;
  assign n6573 = pi20 ? n1026 : n6568;
  assign n6574 = pi20 ? n916 : n139;
  assign n6575 = pi19 ? n6573 : n6574;
  assign n6576 = pi20 ? n927 : n139;
  assign n6577 = pi21 ? n921 : n916;
  assign n6578 = pi20 ? n6577 : n139;
  assign n6579 = pi19 ? n6576 : n6578;
  assign n6580 = pi18 ? n6575 : n6579;
  assign n6581 = pi20 ? n922 : n1016;
  assign n6582 = pi21 ? n316 : n397;
  assign n6583 = pi20 ? n5204 : n6582;
  assign n6584 = pi19 ? n6581 : n6583;
  assign n6585 = pi18 ? n6584 : n32;
  assign n6586 = pi17 ? n6580 : n6585;
  assign n6587 = pi16 ? n6572 : n6586;
  assign n6588 = pi22 ? n909 : n1043;
  assign n6589 = pi21 ? n6588 : n139;
  assign n6590 = pi20 ? n32 : n6589;
  assign n6591 = pi19 ? n32 : n6590;
  assign n6592 = pi20 ? n139 : n2830;
  assign n6593 = pi19 ? n6592 : n1719;
  assign n6594 = pi18 ? n6591 : n6593;
  assign n6595 = pi17 ? n32 : n6594;
  assign n6596 = pi20 ? n2521 : n139;
  assign n6597 = pi19 ? n6596 : n3582;
  assign n6598 = pi19 ? n1720 : n139;
  assign n6599 = pi18 ? n6597 : n6598;
  assign n6600 = pi20 ? n350 : n6582;
  assign n6601 = pi19 ? n139 : n6600;
  assign n6602 = pi18 ? n6601 : n32;
  assign n6603 = pi17 ? n6599 : n6602;
  assign n6604 = pi16 ? n6595 : n6603;
  assign n6605 = pi15 ? n6587 : n6604;
  assign n6606 = pi14 ? n6567 : n6605;
  assign n6607 = pi13 ? n6550 : n6606;
  assign n6608 = pi23 ? n38 : n316;
  assign n6609 = pi22 ? n6608 : n37;
  assign n6610 = pi21 ? n6609 : n316;
  assign n6611 = pi20 ? n32 : n6610;
  assign n6612 = pi19 ? n32 : n6611;
  assign n6613 = pi21 ? n316 : n4015;
  assign n6614 = pi20 ? n6613 : n316;
  assign n6615 = pi19 ? n316 : n6614;
  assign n6616 = pi18 ? n6612 : n6615;
  assign n6617 = pi17 ? n32 : n6616;
  assign n6618 = pi20 ? n316 : n5205;
  assign n6619 = pi19 ? n316 : n6618;
  assign n6620 = pi18 ? n6619 : n32;
  assign n6621 = pi17 ? n316 : n6620;
  assign n6622 = pi16 ? n6617 : n6621;
  assign n6623 = pi20 ? n3697 : n3702;
  assign n6624 = pi21 ? n3258 : n4015;
  assign n6625 = pi21 ? n3258 : n37;
  assign n6626 = pi20 ? n6624 : n6625;
  assign n6627 = pi19 ? n6623 : n6626;
  assign n6628 = pi18 ? n3254 : n6627;
  assign n6629 = pi17 ? n32 : n6628;
  assign n6630 = pi20 ? n6241 : n316;
  assign n6631 = pi19 ? n6630 : n316;
  assign n6632 = pi18 ? n6631 : n316;
  assign n6633 = pi17 ? n6632 : n6620;
  assign n6634 = pi16 ? n6629 : n6633;
  assign n6635 = pi15 ? n6622 : n6634;
  assign n6636 = pi21 ? n326 : n346;
  assign n6637 = pi20 ? n32 : n6636;
  assign n6638 = pi19 ? n32 : n6637;
  assign n6639 = pi20 ? n4437 : n1001;
  assign n6640 = pi21 ? n297 : n4015;
  assign n6641 = pi20 ? n6640 : n1022;
  assign n6642 = pi19 ? n6639 : n6641;
  assign n6643 = pi18 ? n6638 : n6642;
  assign n6644 = pi17 ? n32 : n6643;
  assign n6645 = pi20 ? n5317 : n316;
  assign n6646 = pi19 ? n6645 : n316;
  assign n6647 = pi18 ? n6646 : n316;
  assign n6648 = pi17 ? n6647 : n6620;
  assign n6649 = pi16 ? n6644 : n6648;
  assign n6650 = pi21 ? n139 : n2863;
  assign n6651 = pi20 ? n6650 : n139;
  assign n6652 = pi19 ? n6651 : n139;
  assign n6653 = pi18 ? n913 : n6652;
  assign n6654 = pi17 ? n32 : n6653;
  assign n6655 = pi20 ? n139 : n976;
  assign n6656 = pi21 ? n3188 : n356;
  assign n6657 = pi20 ? n3188 : n6656;
  assign n6658 = pi19 ? n6655 : n6657;
  assign n6659 = pi21 ? n4383 : n139;
  assign n6660 = pi21 ? n3189 : n1810;
  assign n6661 = pi20 ? n6659 : n6660;
  assign n6662 = pi20 ? n1008 : n6660;
  assign n6663 = pi19 ? n6661 : n6662;
  assign n6664 = pi18 ? n6658 : n6663;
  assign n6665 = pi20 ? n1008 : n2383;
  assign n6666 = pi19 ? n6665 : n6618;
  assign n6667 = pi18 ? n6666 : n32;
  assign n6668 = pi17 ? n6664 : n6667;
  assign n6669 = pi16 ? n6654 : n6668;
  assign n6670 = pi15 ? n6649 : n6669;
  assign n6671 = pi14 ? n6635 : n6670;
  assign n6672 = pi21 ? n2497 : n4725;
  assign n6673 = pi20 ? n32 : n6672;
  assign n6674 = pi19 ? n32 : n6673;
  assign n6675 = pi21 ? n1531 : n921;
  assign n6676 = pi22 ? n295 : n204;
  assign n6677 = pi21 ? n6676 : n919;
  assign n6678 = pi20 ? n6675 : n6677;
  assign n6679 = pi21 ? n1696 : n919;
  assign n6680 = pi21 ? n921 : n1531;
  assign n6681 = pi20 ? n6679 : n6680;
  assign n6682 = pi19 ? n6678 : n6681;
  assign n6683 = pi18 ? n6674 : n6682;
  assign n6684 = pi17 ? n32 : n6683;
  assign n6685 = pi21 ? n921 : n1847;
  assign n6686 = pi20 ? n6685 : n4360;
  assign n6687 = pi21 ? n916 : n2876;
  assign n6688 = pi20 ? n6687 : n5926;
  assign n6689 = pi19 ? n6686 : n6688;
  assign n6690 = pi20 ? n5227 : n921;
  assign n6691 = pi21 ? n2864 : n919;
  assign n6692 = pi22 ? n1038 : n918;
  assign n6693 = pi21 ? n6692 : n921;
  assign n6694 = pi20 ? n6691 : n6693;
  assign n6695 = pi19 ? n6690 : n6694;
  assign n6696 = pi18 ? n6689 : n6695;
  assign n6697 = pi21 ? n3207 : n316;
  assign n6698 = pi20 ? n6691 : n6697;
  assign n6699 = pi19 ? n6698 : n6618;
  assign n6700 = pi18 ? n6699 : n32;
  assign n6701 = pi17 ? n6696 : n6700;
  assign n6702 = pi16 ? n6684 : n6701;
  assign n6703 = pi21 ? n555 : n476;
  assign n6704 = pi20 ? n32 : n6703;
  assign n6705 = pi19 ? n32 : n6704;
  assign n6706 = pi22 ? n37 : n448;
  assign n6707 = pi22 ? n450 : n37;
  assign n6708 = pi21 ? n6706 : n6707;
  assign n6709 = pi21 ? n1940 : n1949;
  assign n6710 = pi20 ? n6708 : n6709;
  assign n6711 = pi21 ? n570 : n1949;
  assign n6712 = pi21 ? n335 : n6706;
  assign n6713 = pi20 ? n6711 : n6712;
  assign n6714 = pi19 ? n6710 : n6713;
  assign n6715 = pi18 ? n6705 : n6714;
  assign n6716 = pi17 ? n32 : n6715;
  assign n6717 = pi21 ? n476 : n335;
  assign n6718 = pi21 ? n1949 : n476;
  assign n6719 = pi20 ? n6717 : n6718;
  assign n6720 = pi22 ? n204 : n450;
  assign n6721 = pi21 ? n6720 : n1083;
  assign n6722 = pi20 ? n6720 : n6721;
  assign n6723 = pi19 ? n6719 : n6722;
  assign n6724 = pi21 ? n1083 : n1949;
  assign n6725 = pi21 ? n1949 : n1079;
  assign n6726 = pi20 ? n6724 : n6725;
  assign n6727 = pi21 ? n476 : n1083;
  assign n6728 = pi20 ? n6727 : n6725;
  assign n6729 = pi19 ? n6726 : n6728;
  assign n6730 = pi18 ? n6723 : n6729;
  assign n6731 = pi23 ? n316 : n335;
  assign n6732 = pi22 ? n6731 : n6380;
  assign n6733 = pi21 ? n1083 : n6732;
  assign n6734 = pi20 ? n6727 : n6733;
  assign n6735 = pi22 ? n335 : n2401;
  assign n6736 = pi21 ? n6735 : n4101;
  assign n6737 = pi20 ? n204 : n6736;
  assign n6738 = pi19 ? n6734 : n6737;
  assign n6739 = pi18 ? n6738 : n32;
  assign n6740 = pi17 ? n6730 : n6739;
  assign n6741 = pi16 ? n6716 : n6740;
  assign n6742 = pi15 ? n6702 : n6741;
  assign n6743 = pi21 ? n204 : n760;
  assign n6744 = pi20 ? n204 : n6743;
  assign n6745 = pi19 ? n204 : n6744;
  assign n6746 = pi18 ? n6745 : n32;
  assign n6747 = pi17 ? n204 : n6746;
  assign n6748 = pi16 ? n5355 : n6747;
  assign n6749 = pi20 ? n1089 : n204;
  assign n6750 = pi19 ? n204 : n6749;
  assign n6751 = pi18 ? n5353 : n6750;
  assign n6752 = pi17 ? n32 : n6751;
  assign n6753 = pi16 ? n6752 : n5994;
  assign n6754 = pi15 ? n6748 : n6753;
  assign n6755 = pi14 ? n6742 : n6754;
  assign n6756 = pi13 ? n6671 : n6755;
  assign n6757 = pi12 ? n6607 : n6756;
  assign n6758 = pi11 ? n6471 : n6757;
  assign n6759 = pi10 ? n6354 : n6758;
  assign n6760 = pi09 ? n32 : n6759;
  assign n6761 = pi21 ? n37 : n32;
  assign n6762 = pi20 ? n6761 : n32;
  assign n6763 = pi19 ? n6762 : n32;
  assign n6764 = pi18 ? n37 : n6763;
  assign n6765 = pi17 ? n37 : n6764;
  assign n6766 = pi16 ? n70 : n6765;
  assign n6767 = pi15 ? n32 : n6766;
  assign n6768 = pi14 ? n32 : n6767;
  assign n6769 = pi13 ? n32 : n6768;
  assign n6770 = pi12 ? n32 : n6769;
  assign n6771 = pi11 ? n32 : n6770;
  assign n6772 = pi10 ? n32 : n6771;
  assign n6773 = pi16 ? n5390 : n5400;
  assign n6774 = pi23 ? n37 : n102;
  assign n6775 = pi22 ? n37 : n6774;
  assign n6776 = pi21 ? n6775 : n32;
  assign n6777 = pi20 ? n6776 : n32;
  assign n6778 = pi19 ? n6777 : n32;
  assign n6779 = pi18 ? n37 : n6778;
  assign n6780 = pi17 ? n37 : n6779;
  assign n6781 = pi16 ? n73 : n6780;
  assign n6782 = pi15 ? n6773 : n6781;
  assign n6783 = pi21 ? n32 : n40;
  assign n6784 = pi20 ? n32 : n6783;
  assign n6785 = pi19 ? n32 : n6784;
  assign n6786 = pi18 ? n6785 : n37;
  assign n6787 = pi17 ? n32 : n6786;
  assign n6788 = pi16 ? n6787 : n5400;
  assign n6789 = pi22 ? n37 : n1762;
  assign n6790 = pi21 ? n6789 : n32;
  assign n6791 = pi20 ? n6790 : n32;
  assign n6792 = pi19 ? n6791 : n32;
  assign n6793 = pi18 ? n37 : n6792;
  assign n6794 = pi17 ? n37 : n6793;
  assign n6795 = pi16 ? n83 : n6794;
  assign n6796 = pi15 ? n6788 : n6795;
  assign n6797 = pi14 ? n6782 : n6796;
  assign n6798 = pi23 ? n37 : n586;
  assign n6799 = pi22 ? n37 : n6798;
  assign n6800 = pi21 ? n6799 : n32;
  assign n6801 = pi20 ? n6800 : n32;
  assign n6802 = pi19 ? n6801 : n32;
  assign n6803 = pi18 ? n37 : n6802;
  assign n6804 = pi17 ? n37 : n6803;
  assign n6805 = pi16 ? n2461 : n6804;
  assign n6806 = pi15 ? n6025 : n6805;
  assign n6807 = pi21 ? n6401 : n32;
  assign n6808 = pi20 ? n6807 : n32;
  assign n6809 = pi19 ? n6808 : n32;
  assign n6810 = pi18 ? n37 : n6809;
  assign n6811 = pi17 ? n37 : n6810;
  assign n6812 = pi16 ? n439 : n6811;
  assign n6813 = pi14 ? n6806 : n6812;
  assign n6814 = pi13 ? n6797 : n6813;
  assign n6815 = pi21 ? n159 : n32;
  assign n6816 = pi20 ? n6815 : n32;
  assign n6817 = pi19 ? n6816 : n32;
  assign n6818 = pi18 ? n99 : n6817;
  assign n6819 = pi17 ? n99 : n6818;
  assign n6820 = pi16 ? n721 : n6819;
  assign n6821 = pi16 ? n201 : n6819;
  assign n6822 = pi15 ? n6820 : n6821;
  assign n6823 = pi22 ? n99 : n3961;
  assign n6824 = pi21 ? n6823 : n32;
  assign n6825 = pi20 ? n6824 : n32;
  assign n6826 = pi19 ? n6825 : n32;
  assign n6827 = pi18 ? n99 : n6826;
  assign n6828 = pi17 ? n99 : n6827;
  assign n6829 = pi16 ? n801 : n6828;
  assign n6830 = pi16 ? n744 : n6828;
  assign n6831 = pi15 ? n6829 : n6830;
  assign n6832 = pi14 ? n6822 : n6831;
  assign n6833 = pi23 ? n139 : n233;
  assign n6834 = pi22 ? n99 : n6833;
  assign n6835 = pi21 ? n6834 : n32;
  assign n6836 = pi20 ? n6835 : n32;
  assign n6837 = pi19 ? n6836 : n32;
  assign n6838 = pi18 ? n99 : n6837;
  assign n6839 = pi17 ? n99 : n6838;
  assign n6840 = pi16 ? n744 : n6839;
  assign n6841 = pi19 ? n5459 : n99;
  assign n6842 = pi18 ? n742 : n6841;
  assign n6843 = pi17 ? n32 : n6842;
  assign n6844 = pi21 ? n3444 : n5453;
  assign n6845 = pi22 ? n3443 : n5452;
  assign n6846 = pi21 ? n6096 : n6845;
  assign n6847 = pi20 ? n6844 : n6846;
  assign n6848 = pi19 ? n99 : n6847;
  assign n6849 = pi21 ? n6096 : n5453;
  assign n6850 = pi20 ? n6846 : n6849;
  assign n6851 = pi21 ? n6096 : n5464;
  assign n6852 = pi19 ? n6850 : n6851;
  assign n6853 = pi18 ? n6848 : n6852;
  assign n6854 = pi21 ? n6094 : n5453;
  assign n6855 = pi20 ? n6846 : n6854;
  assign n6856 = pi21 ? n5464 : n767;
  assign n6857 = pi21 ? n5464 : n3444;
  assign n6858 = pi20 ? n6856 : n6857;
  assign n6859 = pi19 ? n6855 : n6858;
  assign n6860 = pi22 ? n3443 : n2060;
  assign n6861 = pi21 ? n6860 : n32;
  assign n6862 = pi20 ? n6861 : n32;
  assign n6863 = pi19 ? n6862 : n32;
  assign n6864 = pi18 ? n6859 : n6863;
  assign n6865 = pi17 ? n6853 : n6864;
  assign n6866 = pi16 ? n6843 : n6865;
  assign n6867 = pi15 ? n6840 : n6866;
  assign n6868 = pi20 ? n5405 : n2191;
  assign n6869 = pi19 ? n6868 : n6091;
  assign n6870 = pi18 ? n6086 : n6869;
  assign n6871 = pi20 ? n6095 : n99;
  assign n6872 = pi19 ? n6871 : n3888;
  assign n6873 = pi21 ? n3444 : n32;
  assign n6874 = pi20 ? n6873 : n32;
  assign n6875 = pi19 ? n6874 : n32;
  assign n6876 = pi18 ? n6872 : n6875;
  assign n6877 = pi17 ? n6870 : n6876;
  assign n6878 = pi16 ? n744 : n6877;
  assign n6879 = pi22 ? n4263 : n37;
  assign n6880 = pi21 ? n6879 : n157;
  assign n6881 = pi20 ? n32 : n6880;
  assign n6882 = pi19 ? n32 : n6881;
  assign n6883 = pi18 ? n6882 : n157;
  assign n6884 = pi17 ? n32 : n6883;
  assign n6885 = pi16 ? n6884 : n6137;
  assign n6886 = pi15 ? n6878 : n6885;
  assign n6887 = pi14 ? n6867 : n6886;
  assign n6888 = pi13 ? n6832 : n6887;
  assign n6889 = pi12 ? n6814 : n6888;
  assign n6890 = pi23 ? n4262 : n37;
  assign n6891 = pi22 ? n6890 : n37;
  assign n6892 = pi21 ? n6891 : n157;
  assign n6893 = pi20 ? n32 : n6892;
  assign n6894 = pi19 ? n32 : n6893;
  assign n6895 = pi18 ? n6894 : n157;
  assign n6896 = pi17 ? n32 : n6895;
  assign n6897 = pi22 ? n157 : n1511;
  assign n6898 = pi21 ? n6897 : n32;
  assign n6899 = pi20 ? n6898 : n32;
  assign n6900 = pi19 ? n6899 : n32;
  assign n6901 = pi18 ? n5173 : n6900;
  assign n6902 = pi17 ? n6145 : n6901;
  assign n6903 = pi16 ? n6896 : n6902;
  assign n6904 = pi15 ? n6885 : n6903;
  assign n6905 = pi14 ? n6904 : n6191;
  assign n6906 = pi21 ? n180 : n349;
  assign n6907 = pi20 ? n32 : n6906;
  assign n6908 = pi19 ? n32 : n6907;
  assign n6909 = pi21 ? n1784 : n349;
  assign n6910 = pi21 ? n4429 : n3617;
  assign n6911 = pi21 ? n348 : n1784;
  assign n6912 = pi20 ? n6910 : n6911;
  assign n6913 = pi19 ? n6909 : n6912;
  assign n6914 = pi18 ? n6908 : n6913;
  assign n6915 = pi17 ? n32 : n6914;
  assign n6916 = pi21 ? n349 : n4429;
  assign n6917 = pi21 ? n3617 : n348;
  assign n6918 = pi20 ? n6916 : n6917;
  assign n6919 = pi21 ? n3617 : n349;
  assign n6920 = pi21 ? n1784 : n139;
  assign n6921 = pi20 ? n6919 : n6920;
  assign n6922 = pi19 ? n6918 : n6921;
  assign n6923 = pi21 ? n139 : n4020;
  assign n6924 = pi20 ? n6920 : n6923;
  assign n6925 = pi21 ? n1777 : n349;
  assign n6926 = pi20 ? n6909 : n6925;
  assign n6927 = pi19 ? n6924 : n6926;
  assign n6928 = pi18 ? n6922 : n6927;
  assign n6929 = pi20 ? n6925 : n139;
  assign n6930 = pi21 ? n346 : n359;
  assign n6931 = pi19 ? n6929 : n6930;
  assign n6932 = pi18 ? n6931 : n6216;
  assign n6933 = pi17 ? n6928 : n6932;
  assign n6934 = pi16 ? n6915 : n6933;
  assign n6935 = pi21 ? n397 : n32;
  assign n6936 = pi20 ? n6935 : n32;
  assign n6937 = pi19 ? n6936 : n32;
  assign n6938 = pi18 ? n316 : n6937;
  assign n6939 = pi17 ? n316 : n6938;
  assign n6940 = pi16 ? n6224 : n6939;
  assign n6941 = pi15 ? n6934 : n6940;
  assign n6942 = pi14 ? n6201 : n6941;
  assign n6943 = pi13 ? n6905 : n6942;
  assign n6944 = pi16 ? n6235 : n6939;
  assign n6945 = pi16 ? n6245 : n6939;
  assign n6946 = pi15 ? n6944 : n6945;
  assign n6947 = pi21 ? n37 : n506;
  assign n6948 = pi20 ? n37 : n6947;
  assign n6949 = pi20 ? n2616 : n6252;
  assign n6950 = pi19 ? n6948 : n6949;
  assign n6951 = pi18 ? n374 : n6950;
  assign n6952 = pi17 ? n32 : n6951;
  assign n6953 = pi16 ? n6952 : n6258;
  assign n6954 = pi16 ? n439 : n6275;
  assign n6955 = pi15 ? n6953 : n6954;
  assign n6956 = pi14 ? n6946 : n6955;
  assign n6957 = pi20 ? n1921 : n6280;
  assign n6958 = pi19 ? n6957 : n6283;
  assign n6959 = pi18 ? n6958 : n6288;
  assign n6960 = pi24 ? n335 : n233;
  assign n6961 = pi23 ? n335 : n6960;
  assign n6962 = pi22 ? n6961 : n4146;
  assign n6963 = pi21 ? n6962 : n32;
  assign n6964 = pi20 ? n6963 : n32;
  assign n6965 = pi19 ? n6964 : n32;
  assign n6966 = pi18 ? n6293 : n6965;
  assign n6967 = pi17 ? n6959 : n6966;
  assign n6968 = pi16 ? n439 : n6967;
  assign n6969 = pi21 ? n569 : n580;
  assign n6970 = pi20 ? n3289 : n6969;
  assign n6971 = pi19 ? n37 : n6970;
  assign n6972 = pi18 ? n6971 : n6308;
  assign n6973 = pi22 ? n2060 : n3396;
  assign n6974 = pi21 ? n6973 : n32;
  assign n6975 = pi20 ? n6974 : n32;
  assign n6976 = pi19 ? n6975 : n32;
  assign n6977 = pi18 ? n6314 : n6976;
  assign n6978 = pi17 ? n6972 : n6977;
  assign n6979 = pi16 ? n439 : n6978;
  assign n6980 = pi15 ? n6968 : n6979;
  assign n6981 = pi19 ? n37 : n6325;
  assign n6982 = pi18 ? n37 : n6981;
  assign n6983 = pi22 ? n2060 : n625;
  assign n6984 = pi21 ? n6983 : n32;
  assign n6985 = pi20 ? n6984 : n32;
  assign n6986 = pi19 ? n6985 : n32;
  assign n6987 = pi18 ? n6330 : n6986;
  assign n6988 = pi17 ? n6982 : n6987;
  assign n6989 = pi16 ? n439 : n6988;
  assign n6990 = pi22 ? n5782 : n688;
  assign n6991 = pi21 ? n6990 : n32;
  assign n6992 = pi20 ? n6991 : n32;
  assign n6993 = pi19 ? n6992 : n32;
  assign n6994 = pi18 ? n6342 : n6993;
  assign n6995 = pi17 ? n6339 : n6994;
  assign n6996 = pi16 ? n439 : n6995;
  assign n6997 = pi15 ? n6989 : n6996;
  assign n6998 = pi14 ? n6980 : n6997;
  assign n6999 = pi13 ? n6956 : n6998;
  assign n7000 = pi12 ? n6943 : n6999;
  assign n7001 = pi11 ? n6889 : n7000;
  assign n7002 = pi22 ? n6365 : n688;
  assign n7003 = pi21 ? n7002 : n32;
  assign n7004 = pi20 ? n7003 : n32;
  assign n7005 = pi19 ? n7004 : n32;
  assign n7006 = pi18 ? n6364 : n7005;
  assign n7007 = pi17 ? n6357 : n7006;
  assign n7008 = pi16 ? n439 : n7007;
  assign n7009 = pi22 ? n6380 : n706;
  assign n7010 = pi21 ? n7009 : n32;
  assign n7011 = pi20 ? n7010 : n32;
  assign n7012 = pi19 ? n7011 : n32;
  assign n7013 = pi18 ? n6379 : n7012;
  assign n7014 = pi17 ? n6375 : n7013;
  assign n7015 = pi16 ? n439 : n7014;
  assign n7016 = pi15 ? n7008 : n7015;
  assign n7017 = pi22 ? n673 : n32;
  assign n7018 = pi21 ? n7017 : n32;
  assign n7019 = pi20 ? n7018 : n32;
  assign n7020 = pi19 ? n7019 : n32;
  assign n7021 = pi18 ? n6392 : n7020;
  assign n7022 = pi17 ? n2115 : n7021;
  assign n7023 = pi16 ? n439 : n7022;
  assign n7024 = pi23 ? n37 : n1432;
  assign n7025 = pi22 ? n37 : n7024;
  assign n7026 = pi21 ? n37 : n7025;
  assign n7027 = pi20 ? n37 : n7026;
  assign n7028 = pi19 ? n37 : n7027;
  assign n7029 = pi18 ? n7028 : n7020;
  assign n7030 = pi17 ? n37 : n7029;
  assign n7031 = pi16 ? n439 : n7030;
  assign n7032 = pi15 ? n7023 : n7031;
  assign n7033 = pi14 ? n7016 : n7032;
  assign n7034 = pi22 ? n233 : n32;
  assign n7035 = pi21 ? n7034 : n32;
  assign n7036 = pi20 ? n7035 : n32;
  assign n7037 = pi19 ? n7036 : n32;
  assign n7038 = pi18 ? n2102 : n7037;
  assign n7039 = pi17 ? n37 : n7038;
  assign n7040 = pi16 ? n439 : n7039;
  assign n7041 = pi22 ? n6365 : n32;
  assign n7042 = pi21 ? n7041 : n32;
  assign n7043 = pi20 ? n7042 : n32;
  assign n7044 = pi19 ? n7043 : n32;
  assign n7045 = pi18 ? n2102 : n7044;
  assign n7046 = pi17 ? n37 : n7045;
  assign n7047 = pi16 ? n439 : n7046;
  assign n7048 = pi22 ? n1475 : n32;
  assign n7049 = pi21 ? n7048 : n32;
  assign n7050 = pi20 ? n7049 : n32;
  assign n7051 = pi19 ? n7050 : n32;
  assign n7052 = pi18 ? n2109 : n7051;
  assign n7053 = pi17 ? n37 : n7052;
  assign n7054 = pi16 ? n439 : n7053;
  assign n7055 = pi15 ? n7047 : n7054;
  assign n7056 = pi14 ? n7040 : n7055;
  assign n7057 = pi13 ? n7033 : n7056;
  assign n7058 = pi18 ? n6429 : n4118;
  assign n7059 = pi17 ? n37 : n7058;
  assign n7060 = pi16 ? n439 : n7059;
  assign n7061 = pi18 ? n6436 : n4118;
  assign n7062 = pi17 ? n37 : n7061;
  assign n7063 = pi16 ? n439 : n7062;
  assign n7064 = pi15 ? n7060 : n7063;
  assign n7065 = pi18 ? n6444 : n4118;
  assign n7066 = pi17 ? n37 : n7065;
  assign n7067 = pi16 ? n439 : n7066;
  assign n7068 = pi18 ? n6450 : n4118;
  assign n7069 = pi17 ? n99 : n7068;
  assign n7070 = pi16 ? n721 : n7069;
  assign n7071 = pi15 ? n7067 : n7070;
  assign n7072 = pi14 ? n7064 : n7071;
  assign n7073 = pi18 ? n5087 : n5832;
  assign n7074 = pi17 ? n99 : n7073;
  assign n7075 = pi16 ? n721 : n7074;
  assign n7076 = pi18 ? n5093 : n2640;
  assign n7077 = pi17 ? n99 : n7076;
  assign n7078 = pi16 ? n721 : n7077;
  assign n7079 = pi15 ? n7075 : n7078;
  assign n7080 = pi15 ? n5853 : n6467;
  assign n7081 = pi14 ? n7079 : n7080;
  assign n7082 = pi13 ? n7072 : n7081;
  assign n7083 = pi12 ? n7057 : n7082;
  assign n7084 = pi22 ? n738 : n164;
  assign n7085 = pi21 ? n7084 : n5875;
  assign n7086 = pi20 ? n32 : n7085;
  assign n7087 = pi19 ? n32 : n7086;
  assign n7088 = pi21 ? n165 : n775;
  assign n7089 = pi20 ? n7088 : n3011;
  assign n7090 = pi21 ? n775 : n3010;
  assign n7091 = pi21 ? n3013 : n165;
  assign n7092 = pi20 ? n7090 : n7091;
  assign n7093 = pi19 ? n7089 : n7092;
  assign n7094 = pi18 ? n7087 : n7093;
  assign n7095 = pi17 ? n32 : n7094;
  assign n7096 = pi21 ? n3013 : n164;
  assign n7097 = pi21 ? n168 : n5875;
  assign n7098 = pi20 ? n7096 : n7097;
  assign n7099 = pi21 ? n777 : n3002;
  assign n7100 = pi20 ? n7099 : n5889;
  assign n7101 = pi19 ? n7098 : n7100;
  assign n7102 = pi21 ? n5899 : n3010;
  assign n7103 = pi20 ? n7102 : n5893;
  assign n7104 = pi21 ? n5875 : n165;
  assign n7105 = pi21 ? n3010 : n3013;
  assign n7106 = pi20 ? n7104 : n7105;
  assign n7107 = pi19 ? n7103 : n7106;
  assign n7108 = pi18 ? n7101 : n7107;
  assign n7109 = pi21 ? n3010 : n5877;
  assign n7110 = pi20 ? n7104 : n7109;
  assign n7111 = pi21 ? n5899 : n777;
  assign n7112 = pi20 ? n7111 : n6491;
  assign n7113 = pi19 ? n7110 : n7112;
  assign n7114 = pi18 ? n7113 : n1824;
  assign n7115 = pi17 ? n7108 : n7114;
  assign n7116 = pi16 ? n7095 : n7115;
  assign n7117 = pi21 ? n739 : n157;
  assign n7118 = pi20 ? n32 : n7117;
  assign n7119 = pi19 ? n32 : n7118;
  assign n7120 = pi18 ? n7119 : n6505;
  assign n7121 = pi17 ? n32 : n7120;
  assign n7122 = pi20 ? n6508 : n2769;
  assign n7123 = pi19 ? n6512 : n7122;
  assign n7124 = pi18 ? n7123 : n32;
  assign n7125 = pi17 ? n6511 : n7124;
  assign n7126 = pi16 ? n7121 : n7125;
  assign n7127 = pi15 ? n7116 : n7126;
  assign n7128 = pi22 ? n738 : n157;
  assign n7129 = pi21 ? n7128 : n775;
  assign n7130 = pi20 ? n32 : n7129;
  assign n7131 = pi19 ? n32 : n7130;
  assign n7132 = pi18 ? n7131 : n6525;
  assign n7133 = pi17 ? n32 : n7132;
  assign n7134 = pi16 ? n7133 : n6540;
  assign n7135 = pi15 ? n7134 : n6548;
  assign n7136 = pi14 ? n7127 : n7135;
  assign n7137 = pi22 ? n316 : n2834;
  assign n7138 = pi21 ? n204 : n7137;
  assign n7139 = pi20 ? n5199 : n7138;
  assign n7140 = pi19 ? n2317 : n7139;
  assign n7141 = pi18 ? n7140 : n32;
  assign n7142 = pi17 ? n139 : n7141;
  assign n7143 = pi16 ? n915 : n7142;
  assign n7144 = pi15 ? n6560 : n7143;
  assign n7145 = pi23 ? n3690 : n139;
  assign n7146 = pi22 ? n7145 : n1784;
  assign n7147 = pi21 ? n7146 : n3617;
  assign n7148 = pi20 ? n32 : n7147;
  assign n7149 = pi19 ? n32 : n7148;
  assign n7150 = pi21 ? n4429 : n4421;
  assign n7151 = pi21 ? n1784 : n354;
  assign n7152 = pi20 ? n7150 : n7151;
  assign n7153 = pi21 ? n4421 : n346;
  assign n7154 = pi21 ? n4421 : n4429;
  assign n7155 = pi20 ? n7153 : n7154;
  assign n7156 = pi19 ? n7152 : n7155;
  assign n7157 = pi18 ? n7149 : n7156;
  assign n7158 = pi17 ? n32 : n7157;
  assign n7159 = pi21 ? n4421 : n4780;
  assign n7160 = pi20 ? n7159 : n5961;
  assign n7161 = pi21 ? n4429 : n4780;
  assign n7162 = pi21 ? n4780 : n4429;
  assign n7163 = pi20 ? n7161 : n7162;
  assign n7164 = pi19 ? n7160 : n7163;
  assign n7165 = pi20 ? n354 : n4421;
  assign n7166 = pi21 ? n356 : n4429;
  assign n7167 = pi20 ? n7166 : n5967;
  assign n7168 = pi19 ? n7165 : n7167;
  assign n7169 = pi18 ? n7164 : n7168;
  assign n7170 = pi21 ? n346 : n349;
  assign n7171 = pi20 ? n7166 : n7170;
  assign n7172 = pi20 ? n6930 : n5205;
  assign n7173 = pi19 ? n7171 : n7172;
  assign n7174 = pi18 ? n7173 : n32;
  assign n7175 = pi17 ? n7169 : n7174;
  assign n7176 = pi16 ? n7158 : n7175;
  assign n7177 = pi15 ? n6587 : n7176;
  assign n7178 = pi14 ? n7144 : n7177;
  assign n7179 = pi13 ? n7136 : n7178;
  assign n7180 = pi19 ? n6655 : n356;
  assign n7181 = pi21 ? n346 : n1531;
  assign n7182 = pi20 ? n3625 : n7181;
  assign n7183 = pi21 ? n3189 : n1531;
  assign n7184 = pi20 ? n1008 : n7183;
  assign n7185 = pi19 ? n7182 : n7184;
  assign n7186 = pi18 ? n7180 : n7185;
  assign n7187 = pi21 ? n3189 : n316;
  assign n7188 = pi20 ? n1008 : n7187;
  assign n7189 = pi19 ? n7188 : n6618;
  assign n7190 = pi18 ? n7189 : n32;
  assign n7191 = pi17 ? n7186 : n7190;
  assign n7192 = pi16 ? n915 : n7191;
  assign n7193 = pi15 ? n6649 : n7192;
  assign n7194 = pi14 ? n6635 : n7193;
  assign n7195 = pi22 ? n37 : n1038;
  assign n7196 = pi21 ? n296 : n7195;
  assign n7197 = pi20 ? n32 : n7196;
  assign n7198 = pi19 ? n32 : n7197;
  assign n7199 = pi21 ? n295 : n5559;
  assign n7200 = pi20 ? n7199 : n6677;
  assign n7201 = pi21 ? n921 : n295;
  assign n7202 = pi20 ? n6679 : n7201;
  assign n7203 = pi19 ? n7200 : n7202;
  assign n7204 = pi18 ? n7198 : n7203;
  assign n7205 = pi17 ? n32 : n7204;
  assign n7206 = pi22 ? n918 : n37;
  assign n7207 = pi21 ? n921 : n7206;
  assign n7208 = pi22 ? n1038 : n295;
  assign n7209 = pi21 ? n7208 : n4343;
  assign n7210 = pi20 ? n7207 : n7209;
  assign n7211 = pi21 ? n6676 : n2876;
  assign n7212 = pi21 ? n2876 : n6676;
  assign n7213 = pi20 ? n7211 : n7212;
  assign n7214 = pi19 ? n7210 : n7213;
  assign n7215 = pi21 ? n5559 : n921;
  assign n7216 = pi20 ? n5227 : n7215;
  assign n7217 = pi22 ? n295 : n455;
  assign n7218 = pi21 ? n4343 : n7217;
  assign n7219 = pi20 ? n7218 : n6693;
  assign n7220 = pi19 ? n7216 : n7219;
  assign n7221 = pi18 ? n7214 : n7220;
  assign n7222 = pi20 ? n7218 : n6697;
  assign n7223 = pi19 ? n7222 : n5276;
  assign n7224 = pi18 ? n7223 : n32;
  assign n7225 = pi17 ? n7221 : n7224;
  assign n7226 = pi16 ? n7205 : n7225;
  assign n7227 = pi21 ? n6706 : n570;
  assign n7228 = pi20 ? n7227 : n6709;
  assign n7229 = pi19 ? n7228 : n6713;
  assign n7230 = pi18 ? n6705 : n7229;
  assign n7231 = pi17 ? n32 : n7230;
  assign n7232 = pi19 ? n6719 : n1083;
  assign n7233 = pi21 ? n1929 : n1949;
  assign n7234 = pi21 ? n1079 : n476;
  assign n7235 = pi20 ? n7233 : n7234;
  assign n7236 = pi20 ? n6727 : n6718;
  assign n7237 = pi19 ? n7235 : n7236;
  assign n7238 = pi18 ? n7232 : n7237;
  assign n7239 = pi22 ? n6731 : n566;
  assign n7240 = pi21 ? n1929 : n7239;
  assign n7241 = pi20 ? n6727 : n7240;
  assign n7242 = pi22 ? n335 : n448;
  assign n7243 = pi23 ? n4882 : n316;
  assign n7244 = pi22 ? n7243 : n32;
  assign n7245 = pi21 ? n7242 : n7244;
  assign n7246 = pi20 ? n204 : n7245;
  assign n7247 = pi19 ? n7241 : n7246;
  assign n7248 = pi18 ? n7247 : n32;
  assign n7249 = pi17 ? n7238 : n7248;
  assign n7250 = pi16 ? n7231 : n7249;
  assign n7251 = pi15 ? n7226 : n7250;
  assign n7252 = pi23 ? n1598 : n2766;
  assign n7253 = pi22 ? n7252 : n32;
  assign n7254 = pi21 ? n204 : n7253;
  assign n7255 = pi20 ? n204 : n7254;
  assign n7256 = pi19 ? n204 : n7255;
  assign n7257 = pi18 ? n7256 : n32;
  assign n7258 = pi17 ? n204 : n7257;
  assign n7259 = pi16 ? n5989 : n7258;
  assign n7260 = pi18 ? n5987 : n6750;
  assign n7261 = pi17 ? n32 : n7260;
  assign n7262 = pi23 ? n1598 : n395;
  assign n7263 = pi22 ? n7262 : n32;
  assign n7264 = pi21 ? n204 : n7263;
  assign n7265 = pi20 ? n204 : n7264;
  assign n7266 = pi19 ? n204 : n7265;
  assign n7267 = pi18 ? n7266 : n32;
  assign n7268 = pi17 ? n204 : n7267;
  assign n7269 = pi16 ? n7261 : n7268;
  assign n7270 = pi15 ? n7259 : n7269;
  assign n7271 = pi14 ? n7251 : n7270;
  assign n7272 = pi13 ? n7194 : n7271;
  assign n7273 = pi12 ? n7179 : n7272;
  assign n7274 = pi11 ? n7083 : n7273;
  assign n7275 = pi10 ? n7001 : n7274;
  assign n7276 = pi09 ? n6772 : n7275;
  assign n7277 = pi08 ? n6760 : n7276;
  assign n7278 = pi07 ? n6016 : n7277;
  assign n7279 = pi06 ? n4511 : n7278;
  assign n7280 = pi05 ? n1616 : n7279;
  assign n7281 = pi04 ? n32 : n7280;
  assign n7282 = pi21 ? n37 : n2933;
  assign n7283 = pi20 ? n7282 : n32;
  assign n7284 = pi19 ? n7283 : n32;
  assign n7285 = pi18 ? n37 : n7284;
  assign n7286 = pi17 ? n37 : n7285;
  assign n7287 = pi16 ? n70 : n7286;
  assign n7288 = pi15 ? n32 : n7287;
  assign n7289 = pi14 ? n32 : n7288;
  assign n7290 = pi13 ? n32 : n7289;
  assign n7291 = pi12 ? n32 : n7290;
  assign n7292 = pi11 ? n32 : n7291;
  assign n7293 = pi10 ? n32 : n7292;
  assign n7294 = pi21 ? n1618 : n32;
  assign n7295 = pi20 ? n7294 : n32;
  assign n7296 = pi19 ? n7295 : n32;
  assign n7297 = pi18 ? n37 : n7296;
  assign n7298 = pi17 ? n37 : n7297;
  assign n7299 = pi16 ? n5390 : n7298;
  assign n7300 = pi21 ? n99 : n32;
  assign n7301 = pi20 ? n7300 : n32;
  assign n7302 = pi19 ? n7301 : n32;
  assign n7303 = pi18 ? n37 : n7302;
  assign n7304 = pi17 ? n37 : n7303;
  assign n7305 = pi16 ? n73 : n7304;
  assign n7306 = pi15 ? n7299 : n7305;
  assign n7307 = pi16 ? n6787 : n7298;
  assign n7308 = pi21 ? n139 : n32;
  assign n7309 = pi20 ? n7308 : n32;
  assign n7310 = pi19 ? n7309 : n32;
  assign n7311 = pi18 ? n37 : n7310;
  assign n7312 = pi17 ? n37 : n7311;
  assign n7313 = pi16 ? n83 : n7312;
  assign n7314 = pi15 ? n7307 : n7313;
  assign n7315 = pi14 ? n7306 : n7314;
  assign n7316 = pi21 ? n584 : n32;
  assign n7317 = pi20 ? n7316 : n32;
  assign n7318 = pi19 ? n7317 : n32;
  assign n7319 = pi18 ? n37 : n7318;
  assign n7320 = pi17 ? n37 : n7319;
  assign n7321 = pi16 ? n1130 : n7320;
  assign n7322 = pi21 ? n5012 : n37;
  assign n7323 = pi19 ? n7322 : n37;
  assign n7324 = pi18 ? n2459 : n7323;
  assign n7325 = pi17 ? n32 : n7324;
  assign n7326 = pi23 ? n363 : n37;
  assign n7327 = pi22 ? n37 : n7326;
  assign n7328 = pi21 ? n5011 : n7327;
  assign n7329 = pi20 ? n37 : n7328;
  assign n7330 = pi19 ? n37 : n7329;
  assign n7331 = pi21 ? n6401 : n7327;
  assign n7332 = pi21 ? n37 : n7327;
  assign n7333 = pi20 ? n7331 : n7332;
  assign n7334 = pi22 ? n7326 : n37;
  assign n7335 = pi21 ? n7334 : n7327;
  assign n7336 = pi20 ? n7328 : n7335;
  assign n7337 = pi19 ? n7333 : n7336;
  assign n7338 = pi18 ? n7330 : n7337;
  assign n7339 = pi20 ? n7335 : n7322;
  assign n7340 = pi20 ? n6402 : n37;
  assign n7341 = pi19 ? n7339 : n7340;
  assign n7342 = pi18 ? n7341 : n6809;
  assign n7343 = pi17 ? n7338 : n7342;
  assign n7344 = pi16 ? n7325 : n7343;
  assign n7345 = pi15 ? n7321 : n7344;
  assign n7346 = pi21 ? n37 : n2164;
  assign n7347 = pi20 ? n7346 : n3039;
  assign n7348 = pi20 ? n3032 : n2970;
  assign n7349 = pi19 ? n7347 : n7348;
  assign n7350 = pi18 ? n184 : n7349;
  assign n7351 = pi17 ? n32 : n7350;
  assign n7352 = pi20 ? n3033 : n3038;
  assign n7353 = pi22 ? n99 : n7326;
  assign n7354 = pi21 ? n37 : n7353;
  assign n7355 = pi20 ? n226 : n7354;
  assign n7356 = pi19 ? n7352 : n7355;
  assign n7357 = pi21 ? n218 : n7353;
  assign n7358 = pi20 ? n7357 : n4625;
  assign n7359 = pi21 ? n2998 : n218;
  assign n7360 = pi20 ? n3039 : n7359;
  assign n7361 = pi19 ? n7358 : n7360;
  assign n7362 = pi18 ? n7356 : n7361;
  assign n7363 = pi21 ? n2998 : n4551;
  assign n7364 = pi22 ? n5011 : n99;
  assign n7365 = pi21 ? n7364 : n99;
  assign n7366 = pi20 ? n7363 : n7365;
  assign n7367 = pi22 ? n112 : n5011;
  assign n7368 = pi21 ? n99 : n7367;
  assign n7369 = pi20 ? n7368 : n2191;
  assign n7370 = pi19 ? n7366 : n7369;
  assign n7371 = pi18 ? n7370 : n6817;
  assign n7372 = pi17 ? n7362 : n7371;
  assign n7373 = pi16 ? n7351 : n7372;
  assign n7374 = pi15 ? n6812 : n7373;
  assign n7375 = pi14 ? n7345 : n7374;
  assign n7376 = pi13 ? n7315 : n7375;
  assign n7377 = pi23 ? n99 : n170;
  assign n7378 = pi22 ? n99 : n7377;
  assign n7379 = pi21 ? n7378 : n32;
  assign n7380 = pi20 ? n7379 : n32;
  assign n7381 = pi19 ? n7380 : n32;
  assign n7382 = pi18 ? n99 : n7381;
  assign n7383 = pi17 ? n99 : n7382;
  assign n7384 = pi16 ? n721 : n7383;
  assign n7385 = pi15 ? n6820 : n7384;
  assign n7386 = pi21 ? n1683 : n32;
  assign n7387 = pi20 ? n7386 : n32;
  assign n7388 = pi19 ? n7387 : n32;
  assign n7389 = pi18 ? n99 : n7388;
  assign n7390 = pi17 ? n99 : n7389;
  assign n7391 = pi16 ? n721 : n7390;
  assign n7392 = pi14 ? n7385 : n7391;
  assign n7393 = pi24 ? n139 : n233;
  assign n7394 = pi23 ? n99 : n7393;
  assign n7395 = pi22 ? n99 : n7394;
  assign n7396 = pi21 ? n7395 : n32;
  assign n7397 = pi20 ? n7396 : n32;
  assign n7398 = pi19 ? n7397 : n32;
  assign n7399 = pi18 ? n99 : n7398;
  assign n7400 = pi17 ? n99 : n7399;
  assign n7401 = pi16 ? n721 : n7400;
  assign n7402 = pi21 ? n685 : n5464;
  assign n7403 = pi20 ? n7402 : n685;
  assign n7404 = pi19 ? n7403 : n685;
  assign n7405 = pi18 ? n719 : n7404;
  assign n7406 = pi17 ? n32 : n7405;
  assign n7407 = pi21 ? n685 : n2700;
  assign n7408 = pi20 ? n7407 : n32;
  assign n7409 = pi19 ? n7408 : n32;
  assign n7410 = pi18 ? n685 : n7409;
  assign n7411 = pi17 ? n685 : n7410;
  assign n7412 = pi16 ? n7406 : n7411;
  assign n7413 = pi15 ? n7401 : n7412;
  assign n7414 = pi22 ? n6107 : n157;
  assign n7415 = pi21 ? n7414 : n157;
  assign n7416 = pi20 ? n32 : n7415;
  assign n7417 = pi19 ? n32 : n7416;
  assign n7418 = pi18 ? n7417 : n157;
  assign n7419 = pi17 ? n32 : n7418;
  assign n7420 = pi24 ? n363 : n685;
  assign n7421 = pi23 ? n157 : n7420;
  assign n7422 = pi22 ? n157 : n7421;
  assign n7423 = pi21 ? n7422 : n32;
  assign n7424 = pi20 ? n7423 : n32;
  assign n7425 = pi19 ? n7424 : n32;
  assign n7426 = pi18 ? n157 : n7425;
  assign n7427 = pi17 ? n157 : n7426;
  assign n7428 = pi16 ? n7419 : n7427;
  assign n7429 = pi22 ? n316 : n157;
  assign n7430 = pi21 ? n7429 : n157;
  assign n7431 = pi19 ? n7430 : n157;
  assign n7432 = pi18 ? n157 : n7431;
  assign n7433 = pi21 ? n7429 : n3562;
  assign n7434 = pi20 ? n157 : n7433;
  assign n7435 = pi21 ? n157 : n3562;
  assign n7436 = pi20 ? n7435 : n157;
  assign n7437 = pi19 ? n7434 : n7436;
  assign n7438 = pi21 ? n6132 : n1009;
  assign n7439 = pi20 ? n7438 : n32;
  assign n7440 = pi19 ? n7439 : n32;
  assign n7441 = pi18 ? n7437 : n7440;
  assign n7442 = pi17 ? n7432 : n7441;
  assign n7443 = pi16 ? n6143 : n7442;
  assign n7444 = pi15 ? n7428 : n7443;
  assign n7445 = pi14 ? n7413 : n7444;
  assign n7446 = pi13 ? n7392 : n7445;
  assign n7447 = pi12 ? n7376 : n7446;
  assign n7448 = pi18 ? n157 : n7440;
  assign n7449 = pi17 ? n157 : n7448;
  assign n7450 = pi16 ? n6143 : n7449;
  assign n7451 = pi21 ? n296 : n204;
  assign n7452 = pi20 ? n32 : n7451;
  assign n7453 = pi19 ? n32 : n7452;
  assign n7454 = pi20 ? n204 : n6158;
  assign n7455 = pi19 ? n7454 : n6163;
  assign n7456 = pi18 ? n7453 : n7455;
  assign n7457 = pi17 ? n32 : n7456;
  assign n7458 = pi20 ? n2316 : n5199;
  assign n7459 = pi20 ? n6577 : n2318;
  assign n7460 = pi19 ? n7458 : n7459;
  assign n7461 = pi20 ? n2318 : n5199;
  assign n7462 = pi20 ? n6158 : n916;
  assign n7463 = pi19 ? n7461 : n7462;
  assign n7464 = pi18 ? n7460 : n7463;
  assign n7465 = pi20 ? n916 : n1016;
  assign n7466 = pi21 ? n916 : n921;
  assign n7467 = pi19 ? n7465 : n7466;
  assign n7468 = pi22 ? n139 : n1484;
  assign n7469 = pi21 ? n7468 : n32;
  assign n7470 = pi20 ? n7469 : n32;
  assign n7471 = pi19 ? n7470 : n32;
  assign n7472 = pi18 ? n7467 : n7471;
  assign n7473 = pi17 ? n7464 : n7472;
  assign n7474 = pi16 ? n7457 : n7473;
  assign n7475 = pi15 ? n7450 : n7474;
  assign n7476 = pi21 ? n1039 : n919;
  assign n7477 = pi21 ? n2864 : n921;
  assign n7478 = pi21 ? n918 : n1039;
  assign n7479 = pi20 ? n7477 : n7478;
  assign n7480 = pi19 ? n7476 : n7479;
  assign n7481 = pi18 ? n990 : n7480;
  assign n7482 = pi17 ? n32 : n7481;
  assign n7483 = pi21 ? n919 : n2864;
  assign n7484 = pi21 ? n921 : n918;
  assign n7485 = pi20 ? n7483 : n7484;
  assign n7486 = pi20 ? n6171 : n139;
  assign n7487 = pi19 ? n7485 : n7486;
  assign n7488 = pi20 ? n139 : n6659;
  assign n7489 = pi19 ? n7488 : n139;
  assign n7490 = pi18 ? n7487 : n7489;
  assign n7491 = pi21 ? n139 : n1832;
  assign n7492 = pi20 ? n139 : n7491;
  assign n7493 = pi21 ? n919 : n2863;
  assign n7494 = pi20 ? n920 : n7493;
  assign n7495 = pi19 ? n7492 : n7494;
  assign n7496 = pi21 ? n1785 : n32;
  assign n7497 = pi20 ? n7496 : n32;
  assign n7498 = pi19 ? n7497 : n32;
  assign n7499 = pi18 ? n7495 : n7498;
  assign n7500 = pi17 ? n7490 : n7499;
  assign n7501 = pi16 ? n7482 : n7500;
  assign n7502 = pi21 ? n1218 : n32;
  assign n7503 = pi20 ? n7502 : n32;
  assign n7504 = pi19 ? n7503 : n32;
  assign n7505 = pi18 ? n139 : n7504;
  assign n7506 = pi17 ? n139 : n7505;
  assign n7507 = pi16 ? n1773 : n7506;
  assign n7508 = pi15 ? n7501 : n7507;
  assign n7509 = pi14 ? n7475 : n7508;
  assign n7510 = pi16 ? n331 : n7506;
  assign n7511 = pi18 ? n990 : n967;
  assign n7512 = pi17 ? n32 : n7511;
  assign n7513 = pi23 ? n335 : n531;
  assign n7514 = pi22 ? n139 : n7513;
  assign n7515 = pi21 ? n7514 : n32;
  assign n7516 = pi20 ? n7515 : n32;
  assign n7517 = pi19 ? n7516 : n32;
  assign n7518 = pi18 ? n139 : n7517;
  assign n7519 = pi17 ? n139 : n7518;
  assign n7520 = pi16 ? n7512 : n7519;
  assign n7521 = pi15 ? n7510 : n7520;
  assign n7522 = pi21 ? n180 : n4052;
  assign n7523 = pi20 ? n32 : n7522;
  assign n7524 = pi19 ? n32 : n7523;
  assign n7525 = pi20 ? n4837 : n393;
  assign n7526 = pi21 ? n3118 : n424;
  assign n7527 = pi20 ? n7526 : n425;
  assign n7528 = pi19 ? n7525 : n7527;
  assign n7529 = pi18 ? n7524 : n7528;
  assign n7530 = pi17 ? n32 : n7529;
  assign n7531 = pi21 ? n349 : n4780;
  assign n7532 = pi20 ? n5652 : n7531;
  assign n7533 = pi19 ? n316 : n7532;
  assign n7534 = pi21 ? n349 : n354;
  assign n7535 = pi21 ? n4421 : n354;
  assign n7536 = pi20 ? n7534 : n7535;
  assign n7537 = pi19 ? n7531 : n7536;
  assign n7538 = pi18 ? n7533 : n7537;
  assign n7539 = pi21 ? n354 : n3617;
  assign n7540 = pi20 ? n7159 : n7539;
  assign n7541 = pi21 ? n316 : n4421;
  assign n7542 = pi20 ? n7541 : n5286;
  assign n7543 = pi19 ? n7540 : n7542;
  assign n7544 = pi22 ? n348 : n7513;
  assign n7545 = pi21 ? n7544 : n32;
  assign n7546 = pi20 ? n7545 : n32;
  assign n7547 = pi19 ? n7546 : n32;
  assign n7548 = pi18 ? n7543 : n7547;
  assign n7549 = pi17 ? n7538 : n7548;
  assign n7550 = pi16 ? n7530 : n7549;
  assign n7551 = pi20 ? n37 : n408;
  assign n7552 = pi21 ? n392 : n952;
  assign n7553 = pi20 ? n7552 : n316;
  assign n7554 = pi19 ? n7551 : n7553;
  assign n7555 = pi18 ? n374 : n7554;
  assign n7556 = pi17 ? n32 : n7555;
  assign n7557 = pi20 ? n316 : n4437;
  assign n7558 = pi19 ? n316 : n7557;
  assign n7559 = pi19 ? n5305 : n4437;
  assign n7560 = pi18 ? n7558 : n7559;
  assign n7561 = pi18 ? n5306 : n6937;
  assign n7562 = pi17 ? n7560 : n7561;
  assign n7563 = pi16 ? n7556 : n7562;
  assign n7564 = pi15 ? n7550 : n7563;
  assign n7565 = pi14 ? n7521 : n7564;
  assign n7566 = pi13 ? n7509 : n7565;
  assign n7567 = pi20 ? n4831 : n4038;
  assign n7568 = pi19 ? n37 : n7567;
  assign n7569 = pi18 ? n374 : n7568;
  assign n7570 = pi17 ? n32 : n7569;
  assign n7571 = pi21 ? n424 : n316;
  assign n7572 = pi20 ? n7571 : n316;
  assign n7573 = pi21 ? n1091 : n316;
  assign n7574 = pi20 ? n316 : n7573;
  assign n7575 = pi19 ? n7572 : n7574;
  assign n7576 = pi20 ? n7573 : n316;
  assign n7577 = pi19 ? n7576 : n7573;
  assign n7578 = pi18 ? n7575 : n7577;
  assign n7579 = pi20 ? n7573 : n4437;
  assign n7580 = pi19 ? n7579 : n316;
  assign n7581 = pi18 ? n7580 : n6937;
  assign n7582 = pi17 ? n7578 : n7581;
  assign n7583 = pi16 ? n7570 : n7582;
  assign n7584 = pi20 ? n2019 : n5766;
  assign n7585 = pi19 ? n37 : n7584;
  assign n7586 = pi20 ? n5766 : n638;
  assign n7587 = pi21 ? n2007 : n569;
  assign n7588 = pi20 ? n649 : n7587;
  assign n7589 = pi19 ? n7586 : n7588;
  assign n7590 = pi18 ? n7585 : n7589;
  assign n7591 = pi21 ? n2007 : n335;
  assign n7592 = pi20 ? n7591 : n2019;
  assign n7593 = pi21 ? n574 : n570;
  assign n7594 = pi21 ? n574 : n2007;
  assign n7595 = pi20 ? n7593 : n7594;
  assign n7596 = pi19 ? n7592 : n7595;
  assign n7597 = pi22 ? n335 : n3174;
  assign n7598 = pi21 ? n7597 : n32;
  assign n7599 = pi20 ? n7598 : n32;
  assign n7600 = pi19 ? n7599 : n32;
  assign n7601 = pi18 ? n7596 : n7600;
  assign n7602 = pi17 ? n7590 : n7601;
  assign n7603 = pi16 ? n439 : n7602;
  assign n7604 = pi15 ? n7583 : n7603;
  assign n7605 = pi20 ? n37 : n507;
  assign n7606 = pi22 ? n455 : n583;
  assign n7607 = pi21 ? n499 : n7606;
  assign n7608 = pi21 ? n570 : n516;
  assign n7609 = pi20 ? n7607 : n7608;
  assign n7610 = pi19 ? n7605 : n7609;
  assign n7611 = pi20 ? n6711 : n1941;
  assign n7612 = pi21 ? n335 : n476;
  assign n7613 = pi21 ? n1083 : n476;
  assign n7614 = pi20 ? n7612 : n7613;
  assign n7615 = pi19 ? n7611 : n7614;
  assign n7616 = pi18 ? n7610 : n7615;
  assign n7617 = pi20 ? n1099 : n1988;
  assign n7618 = pi21 ? n476 : n474;
  assign n7619 = pi20 ? n1954 : n7618;
  assign n7620 = pi19 ? n7617 : n7619;
  assign n7621 = pi22 ? n204 : n3174;
  assign n7622 = pi21 ? n7621 : n32;
  assign n7623 = pi20 ? n7622 : n32;
  assign n7624 = pi19 ? n7623 : n32;
  assign n7625 = pi18 ? n7620 : n7624;
  assign n7626 = pi17 ? n7616 : n7625;
  assign n7627 = pi16 ? n439 : n7626;
  assign n7628 = pi19 ? n37 : n6948;
  assign n7629 = pi20 ? n6947 : n1583;
  assign n7630 = pi20 ? n1912 : n4864;
  assign n7631 = pi19 ? n7629 : n7630;
  assign n7632 = pi18 ? n7628 : n7631;
  assign n7633 = pi20 ? n1063 : n204;
  assign n7634 = pi21 ? n1046 : n1056;
  assign n7635 = pi20 ? n7634 : n4864;
  assign n7636 = pi19 ? n7633 : n7635;
  assign n7637 = pi22 ? n204 : n1388;
  assign n7638 = pi21 ? n7637 : n32;
  assign n7639 = pi20 ? n7638 : n32;
  assign n7640 = pi19 ? n7639 : n32;
  assign n7641 = pi18 ? n7636 : n7640;
  assign n7642 = pi17 ? n7632 : n7641;
  assign n7643 = pi16 ? n439 : n7642;
  assign n7644 = pi15 ? n7627 : n7643;
  assign n7645 = pi14 ? n7604 : n7644;
  assign n7646 = pi21 ? n37 : n2007;
  assign n7647 = pi21 ? n4973 : n566;
  assign n7648 = pi20 ? n7646 : n7647;
  assign n7649 = pi21 ? n1943 : n4975;
  assign n7650 = pi21 ? n4973 : n4990;
  assign n7651 = pi20 ? n7649 : n7650;
  assign n7652 = pi19 ? n7648 : n7651;
  assign n7653 = pi18 ? n37 : n7652;
  assign n7654 = pi20 ? n581 : n4996;
  assign n7655 = pi21 ? n4975 : n567;
  assign n7656 = pi20 ? n7655 : n335;
  assign n7657 = pi19 ? n7654 : n7656;
  assign n7658 = pi22 ? n335 : n6415;
  assign n7659 = pi21 ? n7658 : n32;
  assign n7660 = pi20 ? n7659 : n32;
  assign n7661 = pi19 ? n7660 : n32;
  assign n7662 = pi18 ? n7657 : n7661;
  assign n7663 = pi17 ? n7653 : n7662;
  assign n7664 = pi16 ? n439 : n7663;
  assign n7665 = pi20 ? n575 : n37;
  assign n7666 = pi20 ? n649 : n2008;
  assign n7667 = pi19 ? n7665 : n7666;
  assign n7668 = pi22 ? n335 : n2192;
  assign n7669 = pi21 ? n7668 : n32;
  assign n7670 = pi20 ? n7669 : n32;
  assign n7671 = pi19 ? n7670 : n32;
  assign n7672 = pi18 ? n7667 : n7671;
  assign n7673 = pi17 ? n37 : n7672;
  assign n7674 = pi16 ? n439 : n7673;
  assign n7675 = pi15 ? n7664 : n7674;
  assign n7676 = pi20 ? n37 : n649;
  assign n7677 = pi19 ? n37 : n7676;
  assign n7678 = pi22 ? n335 : n3396;
  assign n7679 = pi21 ? n7678 : n32;
  assign n7680 = pi20 ? n7679 : n32;
  assign n7681 = pi19 ? n7680 : n32;
  assign n7682 = pi18 ? n7677 : n7681;
  assign n7683 = pi17 ? n37 : n7682;
  assign n7684 = pi16 ? n439 : n7683;
  assign n7685 = pi20 ? n37 : n577;
  assign n7686 = pi19 ? n37 : n7685;
  assign n7687 = pi18 ? n7686 : n6216;
  assign n7688 = pi17 ? n37 : n7687;
  assign n7689 = pi16 ? n439 : n7688;
  assign n7690 = pi15 ? n7684 : n7689;
  assign n7691 = pi14 ? n7675 : n7690;
  assign n7692 = pi13 ? n7645 : n7691;
  assign n7693 = pi12 ? n7566 : n7692;
  assign n7694 = pi11 ? n7447 : n7693;
  assign n7695 = pi20 ? n642 : n37;
  assign n7696 = pi20 ? n37 : n6377;
  assign n7697 = pi19 ? n7695 : n7696;
  assign n7698 = pi18 ? n7697 : n5761;
  assign n7699 = pi17 ? n37 : n7698;
  assign n7700 = pi16 ? n439 : n7699;
  assign n7701 = pi18 ? n2114 : n5761;
  assign n7702 = pi17 ? n37 : n7701;
  assign n7703 = pi16 ? n439 : n7702;
  assign n7704 = pi15 ? n7700 : n7703;
  assign n7705 = pi21 ? n2091 : n233;
  assign n7706 = pi20 ? n37 : n7705;
  assign n7707 = pi19 ? n37 : n7706;
  assign n7708 = pi18 ? n7707 : n7037;
  assign n7709 = pi17 ? n37 : n7708;
  assign n7710 = pi16 ? n439 : n7709;
  assign n7711 = pi18 ? n37 : n7037;
  assign n7712 = pi17 ? n37 : n7711;
  assign n7713 = pi16 ? n439 : n7712;
  assign n7714 = pi15 ? n7710 : n7713;
  assign n7715 = pi14 ? n7704 : n7714;
  assign n7716 = pi21 ? n37 : n4891;
  assign n7717 = pi20 ? n37 : n7716;
  assign n7718 = pi19 ? n37 : n7717;
  assign n7719 = pi18 ? n7718 : n7037;
  assign n7720 = pi17 ? n37 : n7719;
  assign n7721 = pi16 ? n439 : n7720;
  assign n7722 = pi15 ? n7040 : n7721;
  assign n7723 = pi22 ? n685 : n32;
  assign n7724 = pi21 ? n7723 : n32;
  assign n7725 = pi20 ? n7724 : n32;
  assign n7726 = pi19 ? n7725 : n32;
  assign n7727 = pi18 ? n2109 : n7726;
  assign n7728 = pi17 ? n37 : n7727;
  assign n7729 = pi16 ? n439 : n7728;
  assign n7730 = pi21 ? n37 : n363;
  assign n7731 = pi20 ? n37 : n7730;
  assign n7732 = pi19 ? n37 : n7731;
  assign n7733 = pi21 ? n1485 : n32;
  assign n7734 = pi20 ? n7733 : n32;
  assign n7735 = pi19 ? n7734 : n32;
  assign n7736 = pi18 ? n7732 : n7735;
  assign n7737 = pi17 ? n37 : n7736;
  assign n7738 = pi16 ? n439 : n7737;
  assign n7739 = pi15 ? n7729 : n7738;
  assign n7740 = pi14 ? n7722 : n7739;
  assign n7741 = pi13 ? n7715 : n7740;
  assign n7742 = pi18 ? n5030 : n3322;
  assign n7743 = pi17 ? n37 : n7742;
  assign n7744 = pi16 ? n439 : n7743;
  assign n7745 = pi21 ? n99 : n37;
  assign n7746 = pi20 ? n99 : n7745;
  assign n7747 = pi21 ? n181 : n218;
  assign n7748 = pi21 ? n218 : n3392;
  assign n7749 = pi20 ? n7747 : n7748;
  assign n7750 = pi19 ? n7746 : n7749;
  assign n7751 = pi18 ? n7750 : n6419;
  assign n7752 = pi17 ? n99 : n7751;
  assign n7753 = pi16 ? n801 : n7752;
  assign n7754 = pi21 ? n99 : n767;
  assign n7755 = pi20 ? n99 : n7754;
  assign n7756 = pi19 ? n99 : n7755;
  assign n7757 = pi18 ? n7756 : n3342;
  assign n7758 = pi17 ? n99 : n7757;
  assign n7759 = pi16 ? n744 : n7758;
  assign n7760 = pi15 ? n7753 : n7759;
  assign n7761 = pi14 ? n7744 : n7760;
  assign n7762 = pi16 ? n744 : n7074;
  assign n7763 = pi20 ? n99 : n6491;
  assign n7764 = pi19 ? n99 : n7763;
  assign n7765 = pi18 ? n7764 : n2640;
  assign n7766 = pi17 ? n99 : n7765;
  assign n7767 = pi16 ? n744 : n7766;
  assign n7768 = pi15 ? n7762 : n7767;
  assign n7769 = pi21 ? n739 : n2161;
  assign n7770 = pi20 ? n32 : n7769;
  assign n7771 = pi19 ? n32 : n7770;
  assign n7772 = pi18 ? n7771 : n6049;
  assign n7773 = pi17 ? n32 : n7772;
  assign n7774 = pi20 ? n2749 : n5405;
  assign n7775 = pi19 ? n5421 : n7774;
  assign n7776 = pi20 ? n2191 : n99;
  assign n7777 = pi19 ? n7776 : n99;
  assign n7778 = pi18 ? n7775 : n7777;
  assign n7779 = pi21 ? n99 : n2998;
  assign n7780 = pi23 ? n685 : n157;
  assign n7781 = pi22 ? n157 : n7780;
  assign n7782 = pi21 ? n7781 : n685;
  assign n7783 = pi20 ? n7779 : n7782;
  assign n7784 = pi19 ? n99 : n7783;
  assign n7785 = pi18 ? n7784 : n2640;
  assign n7786 = pi17 ? n7778 : n7785;
  assign n7787 = pi16 ? n7773 : n7786;
  assign n7788 = pi22 ? n4263 : n157;
  assign n7789 = pi21 ? n7788 : n157;
  assign n7790 = pi20 ? n32 : n7789;
  assign n7791 = pi19 ? n32 : n7790;
  assign n7792 = pi18 ? n7791 : n157;
  assign n7793 = pi17 ? n32 : n7792;
  assign n7794 = pi21 ? n157 : n767;
  assign n7795 = pi20 ? n157 : n7794;
  assign n7796 = pi19 ? n157 : n7795;
  assign n7797 = pi18 ? n7796 : n2655;
  assign n7798 = pi17 ? n157 : n7797;
  assign n7799 = pi16 ? n7793 : n7798;
  assign n7800 = pi15 ? n7787 : n7799;
  assign n7801 = pi14 ? n7768 : n7800;
  assign n7802 = pi13 ? n7761 : n7801;
  assign n7803 = pi12 ? n7741 : n7802;
  assign n7804 = pi21 ? n7788 : n165;
  assign n7805 = pi20 ? n32 : n7804;
  assign n7806 = pi19 ? n32 : n7805;
  assign n7807 = pi21 ? n775 : n3002;
  assign n7808 = pi20 ? n6508 : n7807;
  assign n7809 = pi21 ? n165 : n159;
  assign n7810 = pi21 ? n165 : n3013;
  assign n7811 = pi20 ? n7809 : n7810;
  assign n7812 = pi19 ? n7808 : n7811;
  assign n7813 = pi18 ? n7806 : n7812;
  assign n7814 = pi17 ? n32 : n7813;
  assign n7815 = pi22 ? n157 : n164;
  assign n7816 = pi21 ? n3002 : n7815;
  assign n7817 = pi20 ? n7088 : n7816;
  assign n7818 = pi21 ? n157 : n775;
  assign n7819 = pi20 ? n7818 : n6523;
  assign n7820 = pi19 ? n7817 : n7819;
  assign n7821 = pi21 ? n777 : n7815;
  assign n7822 = pi20 ? n3002 : n7821;
  assign n7823 = pi21 ? n7815 : n157;
  assign n7824 = pi21 ? n3002 : n165;
  assign n7825 = pi20 ? n7823 : n7824;
  assign n7826 = pi19 ? n7822 : n7825;
  assign n7827 = pi18 ? n7820 : n7826;
  assign n7828 = pi20 ? n7823 : n5889;
  assign n7829 = pi21 ? n157 : n685;
  assign n7830 = pi20 ? n157 : n7829;
  assign n7831 = pi19 ? n7828 : n7830;
  assign n7832 = pi21 ? n5370 : n32;
  assign n7833 = pi20 ? n7832 : n32;
  assign n7834 = pi19 ? n7833 : n32;
  assign n7835 = pi18 ? n7831 : n7834;
  assign n7836 = pi17 ? n7827 : n7835;
  assign n7837 = pi16 ? n7814 : n7836;
  assign n7838 = pi21 ? n157 : n6132;
  assign n7839 = pi20 ? n157 : n7838;
  assign n7840 = pi19 ? n99 : n7839;
  assign n7841 = pi18 ? n7840 : n1824;
  assign n7842 = pi17 ? n99 : n7841;
  assign n7843 = pi16 ? n721 : n7842;
  assign n7844 = pi15 ? n7837 : n7843;
  assign n7845 = pi20 ? n99 : n2243;
  assign n7846 = pi19 ? n7845 : n7839;
  assign n7847 = pi18 ? n7846 : n32;
  assign n7848 = pi17 ? n99 : n7847;
  assign n7849 = pi16 ? n721 : n7848;
  assign n7850 = pi21 ? n139 : n157;
  assign n7851 = pi20 ? n139 : n7850;
  assign n7852 = pi19 ? n7851 : n7839;
  assign n7853 = pi18 ? n7852 : n32;
  assign n7854 = pi17 ? n139 : n7853;
  assign n7855 = pi16 ? n2291 : n7854;
  assign n7856 = pi15 ? n7849 : n7855;
  assign n7857 = pi14 ? n7844 : n7856;
  assign n7858 = pi21 ? n204 : n1027;
  assign n7859 = pi20 ? n204 : n7858;
  assign n7860 = pi19 ? n7851 : n7859;
  assign n7861 = pi18 ? n7860 : n32;
  assign n7862 = pi17 ? n139 : n7861;
  assign n7863 = pi16 ? n2291 : n7862;
  assign n7864 = pi19 ? n139 : n2521;
  assign n7865 = pi18 ? n966 : n7864;
  assign n7866 = pi17 ? n32 : n7865;
  assign n7867 = pi20 ? n2365 : n139;
  assign n7868 = pi19 ? n3626 : n7867;
  assign n7869 = pi18 ? n7868 : n139;
  assign n7870 = pi20 ? n139 : n2872;
  assign n7871 = pi21 ? n921 : n349;
  assign n7872 = pi20 ? n7871 : n316;
  assign n7873 = pi19 ? n7870 : n7872;
  assign n7874 = pi18 ? n7873 : n32;
  assign n7875 = pi17 ? n7869 : n7874;
  assign n7876 = pi16 ? n7866 : n7875;
  assign n7877 = pi15 ? n7863 : n7876;
  assign n7878 = pi22 ? n6608 : n316;
  assign n7879 = pi21 ? n7878 : n316;
  assign n7880 = pi20 ? n32 : n7879;
  assign n7881 = pi19 ? n32 : n7880;
  assign n7882 = pi18 ? n7881 : n316;
  assign n7883 = pi17 ? n32 : n7882;
  assign n7884 = pi18 ? n316 : n32;
  assign n7885 = pi17 ? n316 : n7884;
  assign n7886 = pi16 ? n7883 : n7885;
  assign n7887 = pi19 ? n316 : n6645;
  assign n7888 = pi18 ? n7881 : n7887;
  assign n7889 = pi17 ? n32 : n7888;
  assign n7890 = pi22 ? n316 : n3338;
  assign n7891 = pi21 ? n316 : n7890;
  assign n7892 = pi20 ? n316 : n7891;
  assign n7893 = pi19 ? n316 : n7892;
  assign n7894 = pi18 ? n7893 : n32;
  assign n7895 = pi17 ? n316 : n7894;
  assign n7896 = pi16 ? n7889 : n7895;
  assign n7897 = pi15 ? n7886 : n7896;
  assign n7898 = pi14 ? n7877 : n7897;
  assign n7899 = pi13 ? n7857 : n7898;
  assign n7900 = pi21 ? n316 : n37;
  assign n7901 = pi20 ? n7900 : n316;
  assign n7902 = pi19 ? n316 : n7901;
  assign n7903 = pi18 ? n7881 : n7902;
  assign n7904 = pi17 ? n32 : n7903;
  assign n7905 = pi16 ? n7904 : n7895;
  assign n7906 = pi21 ? n2391 : n316;
  assign n7907 = pi20 ? n32 : n7906;
  assign n7908 = pi19 ? n32 : n7907;
  assign n7909 = pi21 ? n204 : n316;
  assign n7910 = pi20 ? n7900 : n7909;
  assign n7911 = pi19 ? n316 : n7910;
  assign n7912 = pi18 ? n7908 : n7911;
  assign n7913 = pi17 ? n32 : n7912;
  assign n7914 = pi20 ? n316 : n6582;
  assign n7915 = pi19 ? n316 : n7914;
  assign n7916 = pi18 ? n7915 : n32;
  assign n7917 = pi17 ? n316 : n7916;
  assign n7918 = pi16 ? n7913 : n7917;
  assign n7919 = pi15 ? n7905 : n7918;
  assign n7920 = pi19 ? n1820 : n7914;
  assign n7921 = pi18 ? n7920 : n32;
  assign n7922 = pi17 ? n139 : n7921;
  assign n7923 = pi16 ? n915 : n7922;
  assign n7924 = pi21 ? n963 : n297;
  assign n7925 = pi20 ? n32 : n7924;
  assign n7926 = pi19 ? n32 : n7925;
  assign n7927 = pi19 ? n139 : n1806;
  assign n7928 = pi18 ? n7926 : n7927;
  assign n7929 = pi17 ? n32 : n7928;
  assign n7930 = pi20 ? n347 : n5205;
  assign n7931 = pi19 ? n139 : n7930;
  assign n7932 = pi18 ? n7931 : n32;
  assign n7933 = pi17 ? n139 : n7932;
  assign n7934 = pi16 ? n7929 : n7933;
  assign n7935 = pi15 ? n7923 : n7934;
  assign n7936 = pi14 ? n7919 : n7935;
  assign n7937 = pi23 ? n38 : n335;
  assign n7938 = pi22 ? n7937 : n335;
  assign n7939 = pi21 ? n7938 : n335;
  assign n7940 = pi20 ? n32 : n7939;
  assign n7941 = pi19 ? n32 : n7940;
  assign n7942 = pi18 ? n7941 : n335;
  assign n7943 = pi17 ? n32 : n7942;
  assign n7944 = pi20 ? n335 : n3311;
  assign n7945 = pi21 ? n1079 : n3693;
  assign n7946 = pi21 ? n1018 : n5178;
  assign n7947 = pi20 ? n7945 : n7946;
  assign n7948 = pi19 ? n7944 : n7947;
  assign n7949 = pi18 ? n7948 : n32;
  assign n7950 = pi17 ? n335 : n7949;
  assign n7951 = pi16 ? n7943 : n7950;
  assign n7952 = pi21 ? n204 : n7723;
  assign n7953 = pi20 ? n3311 : n7952;
  assign n7954 = pi19 ? n335 : n7953;
  assign n7955 = pi18 ? n7954 : n32;
  assign n7956 = pi17 ? n335 : n7955;
  assign n7957 = pi16 ? n2425 : n7956;
  assign n7958 = pi15 ? n7951 : n7957;
  assign n7959 = pi23 ? n1590 : n204;
  assign n7960 = pi22 ? n7959 : n204;
  assign n7961 = pi21 ? n7960 : n204;
  assign n7962 = pi20 ? n32 : n7961;
  assign n7963 = pi19 ? n32 : n7962;
  assign n7964 = pi21 ? n204 : n1079;
  assign n7965 = pi20 ? n7964 : n204;
  assign n7966 = pi19 ? n204 : n7965;
  assign n7967 = pi18 ? n7963 : n7966;
  assign n7968 = pi17 ? n32 : n7967;
  assign n7969 = pi21 ? n204 : n2300;
  assign n7970 = pi20 ? n204 : n7969;
  assign n7971 = pi19 ? n204 : n7970;
  assign n7972 = pi18 ? n7971 : n32;
  assign n7973 = pi17 ? n204 : n7972;
  assign n7974 = pi16 ? n7968 : n7973;
  assign n7975 = pi23 ? n1590 : n233;
  assign n7976 = pi22 ? n7975 : n335;
  assign n7977 = pi21 ? n7976 : n233;
  assign n7978 = pi20 ? n32 : n7977;
  assign n7979 = pi19 ? n32 : n7978;
  assign n7980 = pi21 ? n233 : n335;
  assign n7981 = pi20 ? n7980 : n233;
  assign n7982 = pi19 ? n233 : n7981;
  assign n7983 = pi18 ? n7979 : n7982;
  assign n7984 = pi17 ? n32 : n7983;
  assign n7985 = pi20 ? n233 : n7980;
  assign n7986 = pi22 ? n335 : n363;
  assign n7987 = pi21 ? n7986 : n2320;
  assign n7988 = pi20 ? n6377 : n7987;
  assign n7989 = pi19 ? n7985 : n7988;
  assign n7990 = pi18 ? n7989 : n32;
  assign n7991 = pi17 ? n233 : n7990;
  assign n7992 = pi16 ? n7984 : n7991;
  assign n7993 = pi15 ? n7974 : n7992;
  assign n7994 = pi14 ? n7958 : n7993;
  assign n7995 = pi13 ? n7936 : n7994;
  assign n7996 = pi12 ? n7899 : n7995;
  assign n7997 = pi11 ? n7803 : n7996;
  assign n7998 = pi10 ? n7694 : n7997;
  assign n7999 = pi09 ? n7293 : n7998;
  assign n8000 = pi16 ? n5390 : n7286;
  assign n8001 = pi16 ? n73 : n7286;
  assign n8002 = pi15 ? n8000 : n8001;
  assign n8003 = pi14 ? n32 : n8002;
  assign n8004 = pi13 ? n32 : n8003;
  assign n8005 = pi12 ? n32 : n8004;
  assign n8006 = pi11 ? n32 : n8005;
  assign n8007 = pi10 ? n32 : n8006;
  assign n8008 = pi22 ? n103 : n32;
  assign n8009 = pi21 ? n2957 : n8008;
  assign n8010 = pi20 ? n8009 : n32;
  assign n8011 = pi19 ? n8010 : n32;
  assign n8012 = pi18 ? n37 : n8011;
  assign n8013 = pi17 ? n37 : n8012;
  assign n8014 = pi16 ? n6787 : n8013;
  assign n8015 = pi22 ? n261 : n32;
  assign n8016 = pi21 ? n99 : n8015;
  assign n8017 = pi20 ? n8016 : n32;
  assign n8018 = pi19 ? n8017 : n32;
  assign n8019 = pi18 ? n37 : n8018;
  assign n8020 = pi17 ? n37 : n8019;
  assign n8021 = pi16 ? n83 : n8020;
  assign n8022 = pi15 ? n8014 : n8021;
  assign n8023 = pi21 ? n32 : n56;
  assign n8024 = pi20 ? n32 : n8023;
  assign n8025 = pi19 ? n32 : n8024;
  assign n8026 = pi18 ? n8025 : n37;
  assign n8027 = pi17 ? n32 : n8026;
  assign n8028 = pi21 ? n3073 : n32;
  assign n8029 = pi20 ? n8028 : n32;
  assign n8030 = pi19 ? n8029 : n32;
  assign n8031 = pi18 ? n37 : n8030;
  assign n8032 = pi17 ? n37 : n8031;
  assign n8033 = pi16 ? n8027 : n8032;
  assign n8034 = pi16 ? n1130 : n7312;
  assign n8035 = pi15 ? n8033 : n8034;
  assign n8036 = pi14 ? n8022 : n8035;
  assign n8037 = pi16 ? n2461 : n7320;
  assign n8038 = pi21 ? n7334 : n37;
  assign n8039 = pi20 ? n37 : n8038;
  assign n8040 = pi19 ? n37 : n8039;
  assign n8041 = pi18 ? n37 : n8040;
  assign n8042 = pi20 ? n8038 : n37;
  assign n8043 = pi19 ? n8042 : n37;
  assign n8044 = pi22 ? n5631 : n32;
  assign n8045 = pi21 ? n6401 : n8044;
  assign n8046 = pi20 ? n8045 : n32;
  assign n8047 = pi19 ? n8046 : n32;
  assign n8048 = pi18 ? n8043 : n8047;
  assign n8049 = pi17 ? n8041 : n8048;
  assign n8050 = pi16 ? n439 : n8049;
  assign n8051 = pi15 ? n8037 : n8050;
  assign n8052 = pi18 ? n37 : n8047;
  assign n8053 = pi17 ? n37 : n8052;
  assign n8054 = pi16 ? n439 : n8053;
  assign n8055 = pi21 ? n180 : n2161;
  assign n8056 = pi20 ? n32 : n8055;
  assign n8057 = pi19 ? n32 : n8056;
  assign n8058 = pi21 ? n112 : n2746;
  assign n8059 = pi20 ? n3879 : n8058;
  assign n8060 = pi21 ? n2164 : n1143;
  assign n8061 = pi20 ? n8060 : n6044;
  assign n8062 = pi19 ? n8059 : n8061;
  assign n8063 = pi18 ? n8057 : n8062;
  assign n8064 = pi17 ? n32 : n8063;
  assign n8065 = pi20 ? n4616 : n3506;
  assign n8066 = pi20 ? n4202 : n8058;
  assign n8067 = pi19 ? n8065 : n8066;
  assign n8068 = pi20 ? n4619 : n99;
  assign n8069 = pi21 ? n2998 : n2746;
  assign n8070 = pi20 ? n8058 : n8069;
  assign n8071 = pi19 ? n8068 : n8070;
  assign n8072 = pi18 ? n8067 : n8071;
  assign n8073 = pi20 ? n2999 : n4202;
  assign n8074 = pi20 ? n4625 : n99;
  assign n8075 = pi19 ? n8073 : n8074;
  assign n8076 = pi21 ? n159 : n2469;
  assign n8077 = pi20 ? n8076 : n32;
  assign n8078 = pi19 ? n8077 : n32;
  assign n8079 = pi18 ? n8075 : n8078;
  assign n8080 = pi17 ? n8072 : n8079;
  assign n8081 = pi16 ? n8064 : n8080;
  assign n8082 = pi15 ? n8054 : n8081;
  assign n8083 = pi14 ? n8051 : n8082;
  assign n8084 = pi13 ? n8036 : n8083;
  assign n8085 = pi18 ? n99 : n8078;
  assign n8086 = pi17 ? n99 : n8085;
  assign n8087 = pi16 ? n744 : n8086;
  assign n8088 = pi21 ? n99 : n2469;
  assign n8089 = pi20 ? n8088 : n32;
  assign n8090 = pi19 ? n8089 : n32;
  assign n8091 = pi18 ? n99 : n8090;
  assign n8092 = pi17 ? n99 : n8091;
  assign n8093 = pi16 ? n744 : n8092;
  assign n8094 = pi15 ? n8087 : n8093;
  assign n8095 = pi21 ? n99 : n2553;
  assign n8096 = pi20 ? n8095 : n32;
  assign n8097 = pi19 ? n8096 : n32;
  assign n8098 = pi18 ? n99 : n8097;
  assign n8099 = pi17 ? n99 : n8098;
  assign n8100 = pi16 ? n744 : n8099;
  assign n8101 = pi14 ? n8094 : n8100;
  assign n8102 = pi21 ? n746 : n2678;
  assign n8103 = pi20 ? n8102 : n32;
  assign n8104 = pi19 ? n8103 : n32;
  assign n8105 = pi18 ? n99 : n8104;
  assign n8106 = pi17 ? n99 : n8105;
  assign n8107 = pi16 ? n744 : n8106;
  assign n8108 = pi18 ? n742 : n7404;
  assign n8109 = pi17 ? n32 : n8108;
  assign n8110 = pi16 ? n8109 : n7411;
  assign n8111 = pi15 ? n8107 : n8110;
  assign n8112 = pi21 ? n157 : n2700;
  assign n8113 = pi20 ? n8112 : n32;
  assign n8114 = pi19 ? n8113 : n32;
  assign n8115 = pi18 ? n157 : n8114;
  assign n8116 = pi17 ? n157 : n8115;
  assign n8117 = pi16 ? n7793 : n8116;
  assign n8118 = pi23 ? n157 : n842;
  assign n8119 = pi22 ? n157 : n8118;
  assign n8120 = pi21 ? n8119 : n1009;
  assign n8121 = pi20 ? n8120 : n32;
  assign n8122 = pi19 ? n8121 : n32;
  assign n8123 = pi18 ? n7437 : n8122;
  assign n8124 = pi17 ? n7432 : n8123;
  assign n8125 = pi16 ? n6143 : n8124;
  assign n8126 = pi15 ? n8117 : n8125;
  assign n8127 = pi14 ? n8111 : n8126;
  assign n8128 = pi13 ? n8101 : n8127;
  assign n8129 = pi12 ? n8084 : n8128;
  assign n8130 = pi18 ? n157 : n8122;
  assign n8131 = pi17 ? n157 : n8130;
  assign n8132 = pi16 ? n6143 : n8131;
  assign n8133 = pi24 ? n204 : n316;
  assign n8134 = pi23 ? n157 : n8133;
  assign n8135 = pi22 ? n139 : n8134;
  assign n8136 = pi21 ? n8135 : n32;
  assign n8137 = pi20 ? n8136 : n32;
  assign n8138 = pi19 ? n8137 : n32;
  assign n8139 = pi18 ? n7467 : n8138;
  assign n8140 = pi17 ? n7464 : n8139;
  assign n8141 = pi16 ? n7457 : n8140;
  assign n8142 = pi15 ? n8132 : n8141;
  assign n8143 = pi22 ? n55 : n1043;
  assign n8144 = pi21 ? n8143 : n139;
  assign n8145 = pi20 ? n32 : n8144;
  assign n8146 = pi19 ? n32 : n8145;
  assign n8147 = pi20 ? n5227 : n927;
  assign n8148 = pi21 ? n2863 : n921;
  assign n8149 = pi21 ? n919 : n916;
  assign n8150 = pi20 ? n8148 : n8149;
  assign n8151 = pi19 ? n8147 : n8150;
  assign n8152 = pi18 ? n8146 : n8151;
  assign n8153 = pi17 ? n32 : n8152;
  assign n8154 = pi21 ? n921 : n919;
  assign n8155 = pi20 ? n6650 : n8154;
  assign n8156 = pi19 ? n8155 : n139;
  assign n8157 = pi18 ? n8156 : n3627;
  assign n8158 = pi20 ? n139 : n6650;
  assign n8159 = pi19 ? n2551 : n8158;
  assign n8160 = pi24 ? n139 : n316;
  assign n8161 = pi23 ? n139 : n8160;
  assign n8162 = pi22 ? n139 : n8161;
  assign n8163 = pi21 ? n8162 : n32;
  assign n8164 = pi20 ? n8163 : n32;
  assign n8165 = pi19 ? n8164 : n32;
  assign n8166 = pi18 ? n8159 : n8165;
  assign n8167 = pi17 ? n8157 : n8166;
  assign n8168 = pi16 ? n8153 : n8167;
  assign n8169 = pi18 ? n8146 : n139;
  assign n8170 = pi17 ? n32 : n8169;
  assign n8171 = pi16 ? n8170 : n7506;
  assign n8172 = pi15 ? n8168 : n8171;
  assign n8173 = pi14 ? n8142 : n8172;
  assign n8174 = pi23 ? n139 : n586;
  assign n8175 = pi22 ? n139 : n8174;
  assign n8176 = pi21 ? n8175 : n32;
  assign n8177 = pi20 ? n8176 : n32;
  assign n8178 = pi19 ? n8177 : n32;
  assign n8179 = pi18 ? n139 : n8178;
  assign n8180 = pi17 ? n139 : n8179;
  assign n8181 = pi16 ? n915 : n8180;
  assign n8182 = pi18 ? n2500 : n967;
  assign n8183 = pi17 ? n32 : n8182;
  assign n8184 = pi24 ? n139 : n335;
  assign n8185 = pi23 ? n8184 : n531;
  assign n8186 = pi22 ? n139 : n8185;
  assign n8187 = pi21 ? n8186 : n32;
  assign n8188 = pi20 ? n8187 : n32;
  assign n8189 = pi19 ? n8188 : n32;
  assign n8190 = pi18 ? n139 : n8189;
  assign n8191 = pi17 ? n139 : n8190;
  assign n8192 = pi16 ? n8183 : n8191;
  assign n8193 = pi15 ? n8181 : n8192;
  assign n8194 = pi20 ? n5709 : n3275;
  assign n8195 = pi19 ? n37 : n8194;
  assign n8196 = pi18 ? n374 : n8195;
  assign n8197 = pi17 ? n32 : n8196;
  assign n8198 = pi23 ? n335 : n5630;
  assign n8199 = pi22 ? n348 : n8198;
  assign n8200 = pi21 ? n8199 : n32;
  assign n8201 = pi20 ? n8200 : n32;
  assign n8202 = pi19 ? n8201 : n32;
  assign n8203 = pi18 ? n7543 : n8202;
  assign n8204 = pi17 ? n7538 : n8203;
  assign n8205 = pi16 ? n8197 : n8204;
  assign n8206 = pi21 ? n180 : n3668;
  assign n8207 = pi20 ? n32 : n8206;
  assign n8208 = pi19 ? n32 : n8207;
  assign n8209 = pi21 ? n37 : n1698;
  assign n8210 = pi21 ? n37 : n952;
  assign n8211 = pi20 ? n8209 : n8210;
  assign n8212 = pi19 ? n8211 : n7553;
  assign n8213 = pi18 ? n8208 : n8212;
  assign n8214 = pi17 ? n32 : n8213;
  assign n8215 = pi21 ? n1246 : n32;
  assign n8216 = pi20 ? n8215 : n32;
  assign n8217 = pi19 ? n8216 : n32;
  assign n8218 = pi18 ? n5306 : n8217;
  assign n8219 = pi17 ? n7560 : n8218;
  assign n8220 = pi16 ? n8214 : n8219;
  assign n8221 = pi15 ? n8205 : n8220;
  assign n8222 = pi14 ? n8193 : n8221;
  assign n8223 = pi13 ? n8173 : n8222;
  assign n8224 = pi20 ? n37 : n5714;
  assign n8225 = pi19 ? n37 : n8224;
  assign n8226 = pi18 ? n374 : n8225;
  assign n8227 = pi17 ? n32 : n8226;
  assign n8228 = pi23 ? n316 : n1149;
  assign n8229 = pi22 ? n316 : n8228;
  assign n8230 = pi21 ? n8229 : n32;
  assign n8231 = pi20 ? n8230 : n32;
  assign n8232 = pi19 ? n8231 : n32;
  assign n8233 = pi18 ? n7580 : n8232;
  assign n8234 = pi17 ? n7578 : n8233;
  assign n8235 = pi16 ? n8227 : n8234;
  assign n8236 = pi15 ? n8235 : n7603;
  assign n8237 = pi20 ? n37 : n1315;
  assign n8238 = pi20 ? n5741 : n7608;
  assign n8239 = pi19 ? n8237 : n8238;
  assign n8240 = pi18 ? n8239 : n7615;
  assign n8241 = pi17 ? n8240 : n7625;
  assign n8242 = pi16 ? n439 : n8241;
  assign n8243 = pi18 ? n37 : n7631;
  assign n8244 = pi17 ? n8243 : n7641;
  assign n8245 = pi16 ? n439 : n8244;
  assign n8246 = pi15 ? n8242 : n8245;
  assign n8247 = pi14 ? n8236 : n8246;
  assign n8248 = pi20 ? n647 : n4974;
  assign n8249 = pi20 ? n2008 : n335;
  assign n8250 = pi19 ? n8248 : n8249;
  assign n8251 = pi18 ? n8250 : n7661;
  assign n8252 = pi17 ? n6375 : n8251;
  assign n8253 = pi16 ? n439 : n8252;
  assign n8254 = pi20 ? n4971 : n2008;
  assign n8255 = pi19 ? n7665 : n8254;
  assign n8256 = pi18 ? n8255 : n7671;
  assign n8257 = pi17 ? n37 : n8256;
  assign n8258 = pi16 ? n439 : n8257;
  assign n8259 = pi15 ? n8253 : n8258;
  assign n8260 = pi22 ? n335 : n1407;
  assign n8261 = pi21 ? n8260 : n32;
  assign n8262 = pi20 ? n8261 : n32;
  assign n8263 = pi19 ? n8262 : n32;
  assign n8264 = pi18 ? n7677 : n8263;
  assign n8265 = pi17 ? n37 : n8264;
  assign n8266 = pi16 ? n439 : n8265;
  assign n8267 = pi15 ? n8266 : n7689;
  assign n8268 = pi14 ? n8259 : n8267;
  assign n8269 = pi13 ? n8247 : n8268;
  assign n8270 = pi12 ? n8223 : n8269;
  assign n8271 = pi11 ? n8129 : n8270;
  assign n8272 = pi22 ? n233 : n3396;
  assign n8273 = pi21 ? n8272 : n32;
  assign n8274 = pi20 ? n8273 : n32;
  assign n8275 = pi19 ? n8274 : n32;
  assign n8276 = pi18 ? n7697 : n8275;
  assign n8277 = pi17 ? n37 : n8276;
  assign n8278 = pi16 ? n439 : n8277;
  assign n8279 = pi18 ? n2114 : n8275;
  assign n8280 = pi17 ? n37 : n8279;
  assign n8281 = pi16 ? n439 : n8280;
  assign n8282 = pi15 ? n8278 : n8281;
  assign n8283 = pi18 ? n7707 : n4854;
  assign n8284 = pi17 ? n37 : n8283;
  assign n8285 = pi16 ? n439 : n8284;
  assign n8286 = pi15 ? n8285 : n4857;
  assign n8287 = pi14 ? n8282 : n8286;
  assign n8288 = pi18 ? n2102 : n4854;
  assign n8289 = pi17 ? n37 : n8288;
  assign n8290 = pi16 ? n439 : n8289;
  assign n8291 = pi18 ? n7718 : n4854;
  assign n8292 = pi17 ? n37 : n8291;
  assign n8293 = pi16 ? n439 : n8292;
  assign n8294 = pi15 ? n8290 : n8293;
  assign n8295 = pi21 ? n696 : n32;
  assign n8296 = pi20 ? n8295 : n32;
  assign n8297 = pi19 ? n8296 : n32;
  assign n8298 = pi18 ? n2109 : n8297;
  assign n8299 = pi17 ? n37 : n8298;
  assign n8300 = pi16 ? n439 : n8299;
  assign n8301 = pi21 ? n2245 : n32;
  assign n8302 = pi20 ? n8301 : n32;
  assign n8303 = pi19 ? n8302 : n32;
  assign n8304 = pi18 ? n7732 : n8303;
  assign n8305 = pi17 ? n37 : n8304;
  assign n8306 = pi16 ? n439 : n8305;
  assign n8307 = pi15 ? n8300 : n8306;
  assign n8308 = pi14 ? n8294 : n8307;
  assign n8309 = pi13 ? n8287 : n8308;
  assign n8310 = pi24 ? n363 : n157;
  assign n8311 = pi23 ? n8310 : n685;
  assign n8312 = pi22 ? n8311 : n32;
  assign n8313 = pi21 ? n8312 : n32;
  assign n8314 = pi20 ? n8313 : n32;
  assign n8315 = pi19 ? n8314 : n32;
  assign n8316 = pi18 ? n5030 : n8315;
  assign n8317 = pi17 ? n37 : n8316;
  assign n8318 = pi16 ? n439 : n8317;
  assign n8319 = pi24 ? n363 : n204;
  assign n8320 = pi23 ? n8319 : n685;
  assign n8321 = pi22 ? n8320 : n32;
  assign n8322 = pi21 ? n8321 : n32;
  assign n8323 = pi20 ? n8322 : n32;
  assign n8324 = pi19 ? n8323 : n32;
  assign n8325 = pi18 ? n7750 : n8324;
  assign n8326 = pi17 ? n99 : n8325;
  assign n8327 = pi16 ? n801 : n8326;
  assign n8328 = pi23 ? n778 : n316;
  assign n8329 = pi22 ? n8328 : n32;
  assign n8330 = pi21 ? n8329 : n32;
  assign n8331 = pi20 ? n8330 : n32;
  assign n8332 = pi19 ? n8331 : n32;
  assign n8333 = pi18 ? n7756 : n8332;
  assign n8334 = pi17 ? n99 : n8333;
  assign n8335 = pi16 ? n721 : n8334;
  assign n8336 = pi15 ? n8327 : n8335;
  assign n8337 = pi14 ? n8318 : n8336;
  assign n8338 = pi18 ? n5087 : n7051;
  assign n8339 = pi17 ? n99 : n8338;
  assign n8340 = pi16 ? n721 : n8339;
  assign n8341 = pi22 ? n157 : n3443;
  assign n8342 = pi21 ? n8341 : n685;
  assign n8343 = pi20 ? n99 : n8342;
  assign n8344 = pi19 ? n99 : n8343;
  assign n8345 = pi18 ? n8344 : n5832;
  assign n8346 = pi17 ? n99 : n8345;
  assign n8347 = pi16 ? n721 : n8346;
  assign n8348 = pi15 ? n8340 : n8347;
  assign n8349 = pi22 ? n715 : n164;
  assign n8350 = pi21 ? n8349 : n158;
  assign n8351 = pi20 ? n32 : n8350;
  assign n8352 = pi19 ? n32 : n8351;
  assign n8353 = pi21 ? n165 : n158;
  assign n8354 = pi20 ? n8353 : n5886;
  assign n8355 = pi21 ? n3013 : n2998;
  assign n8356 = pi20 ? n8355 : n7096;
  assign n8357 = pi19 ? n8354 : n8356;
  assign n8358 = pi18 ? n8352 : n8357;
  assign n8359 = pi17 ? n32 : n8358;
  assign n8360 = pi21 ? n158 : n3002;
  assign n8361 = pi20 ? n8360 : n7097;
  assign n8362 = pi21 ? n165 : n5899;
  assign n8363 = pi20 ? n8362 : n7102;
  assign n8364 = pi19 ? n8361 : n8363;
  assign n8365 = pi21 ? n3010 : n7815;
  assign n8366 = pi21 ? n3013 : n5875;
  assign n8367 = pi20 ? n8365 : n8366;
  assign n8368 = pi20 ? n7824 : n5895;
  assign n8369 = pi19 ? n8367 : n8368;
  assign n8370 = pi18 ? n8364 : n8369;
  assign n8371 = pi21 ? n168 : n775;
  assign n8372 = pi20 ? n7824 : n8371;
  assign n8373 = pi21 ? n2998 : n775;
  assign n8374 = pi20 ? n8373 : n7829;
  assign n8375 = pi19 ? n8372 : n8374;
  assign n8376 = pi18 ? n8375 : n5832;
  assign n8377 = pi17 ? n8370 : n8376;
  assign n8378 = pi16 ? n8359 : n8377;
  assign n8379 = pi16 ? n5910 : n7798;
  assign n8380 = pi15 ? n8378 : n8379;
  assign n8381 = pi14 ? n8348 : n8380;
  assign n8382 = pi13 ? n8337 : n8381;
  assign n8383 = pi12 ? n8309 : n8382;
  assign n8384 = pi21 ? n7128 : n165;
  assign n8385 = pi20 ? n32 : n8384;
  assign n8386 = pi19 ? n32 : n8385;
  assign n8387 = pi20 ? n7824 : n7807;
  assign n8388 = pi19 ? n8387 : n7811;
  assign n8389 = pi18 ? n8386 : n8388;
  assign n8390 = pi17 ? n32 : n8389;
  assign n8391 = pi21 ? n164 : n775;
  assign n8392 = pi20 ? n7088 : n8391;
  assign n8393 = pi21 ? n2998 : n3002;
  assign n8394 = pi20 ? n3004 : n8393;
  assign n8395 = pi19 ? n8392 : n8394;
  assign n8396 = pi20 ? n777 : n7088;
  assign n8397 = pi20 ? n7807 : n165;
  assign n8398 = pi19 ? n8396 : n8397;
  assign n8399 = pi18 ? n8395 : n8398;
  assign n8400 = pi20 ? n7807 : n5901;
  assign n8401 = pi19 ? n8400 : n7830;
  assign n8402 = pi18 ? n8401 : n2655;
  assign n8403 = pi17 ? n8399 : n8402;
  assign n8404 = pi16 ? n8390 : n8403;
  assign n8405 = pi16 ? n744 : n7842;
  assign n8406 = pi15 ? n8404 : n8405;
  assign n8407 = pi16 ? n744 : n7848;
  assign n8408 = pi16 ? n915 : n7854;
  assign n8409 = pi15 ? n8407 : n8408;
  assign n8410 = pi14 ? n8406 : n8409;
  assign n8411 = pi16 ? n915 : n7862;
  assign n8412 = pi22 ? n909 : n1784;
  assign n8413 = pi21 ? n8412 : n139;
  assign n8414 = pi20 ? n32 : n8413;
  assign n8415 = pi19 ? n32 : n8414;
  assign n8416 = pi21 ? n3617 : n1785;
  assign n8417 = pi20 ? n4767 : n8416;
  assign n8418 = pi19 ? n8417 : n5961;
  assign n8419 = pi18 ? n8415 : n8418;
  assign n8420 = pi17 ? n32 : n8419;
  assign n8421 = pi21 ? n139 : n3617;
  assign n8422 = pi20 ? n8421 : n4411;
  assign n8423 = pi21 ? n4429 : n346;
  assign n8424 = pi20 ? n8423 : n4429;
  assign n8425 = pi19 ? n8422 : n8424;
  assign n8426 = pi20 ? n346 : n5961;
  assign n8427 = pi20 ? n7166 : n4422;
  assign n8428 = pi19 ? n8426 : n8427;
  assign n8429 = pi18 ? n8425 : n8428;
  assign n8430 = pi20 ? n4433 : n4422;
  assign n8431 = pi22 ? n204 : n348;
  assign n8432 = pi21 ? n8431 : n346;
  assign n8433 = pi20 ? n8432 : n316;
  assign n8434 = pi19 ? n8430 : n8433;
  assign n8435 = pi18 ? n8434 : n32;
  assign n8436 = pi17 ? n8429 : n8435;
  assign n8437 = pi16 ? n8420 : n8436;
  assign n8438 = pi15 ? n8411 : n8437;
  assign n8439 = pi23 ? n3690 : n316;
  assign n8440 = pi22 ? n8439 : n316;
  assign n8441 = pi21 ? n8440 : n316;
  assign n8442 = pi20 ? n32 : n8441;
  assign n8443 = pi19 ? n32 : n8442;
  assign n8444 = pi18 ? n8443 : n316;
  assign n8445 = pi17 ? n32 : n8444;
  assign n8446 = pi16 ? n8445 : n7885;
  assign n8447 = pi23 ? n961 : n316;
  assign n8448 = pi22 ? n8447 : n316;
  assign n8449 = pi21 ? n8448 : n316;
  assign n8450 = pi20 ? n32 : n8449;
  assign n8451 = pi19 ? n32 : n8450;
  assign n8452 = pi18 ? n8451 : n7887;
  assign n8453 = pi17 ? n32 : n8452;
  assign n8454 = pi22 ? n316 : n1388;
  assign n8455 = pi21 ? n316 : n8454;
  assign n8456 = pi20 ? n316 : n8455;
  assign n8457 = pi19 ? n316 : n8456;
  assign n8458 = pi18 ? n8457 : n32;
  assign n8459 = pi17 ? n316 : n8458;
  assign n8460 = pi16 ? n8453 : n8459;
  assign n8461 = pi15 ? n8446 : n8460;
  assign n8462 = pi14 ? n8438 : n8461;
  assign n8463 = pi13 ? n8410 : n8462;
  assign n8464 = pi22 ? n316 : n6415;
  assign n8465 = pi21 ? n316 : n8464;
  assign n8466 = pi20 ? n316 : n8465;
  assign n8467 = pi19 ? n316 : n8466;
  assign n8468 = pi18 ? n8467 : n32;
  assign n8469 = pi17 ? n316 : n8468;
  assign n8470 = pi16 ? n7904 : n8469;
  assign n8471 = pi15 ? n8470 : n7918;
  assign n8472 = pi21 ? n910 : n297;
  assign n8473 = pi20 ? n32 : n8472;
  assign n8474 = pi19 ? n32 : n8473;
  assign n8475 = pi18 ? n8474 : n7927;
  assign n8476 = pi17 ? n32 : n8475;
  assign n8477 = pi16 ? n8476 : n7933;
  assign n8478 = pi15 ? n7923 : n8477;
  assign n8479 = pi14 ? n8471 : n8478;
  assign n8480 = pi21 ? n476 : n3693;
  assign n8481 = pi20 ? n8480 : n7946;
  assign n8482 = pi19 ? n7944 : n8481;
  assign n8483 = pi18 ? n8482 : n32;
  assign n8484 = pi17 ? n335 : n8483;
  assign n8485 = pi16 ? n7943 : n8484;
  assign n8486 = pi22 ? n685 : n706;
  assign n8487 = pi21 ? n204 : n8486;
  assign n8488 = pi20 ? n3311 : n8487;
  assign n8489 = pi19 ? n335 : n8488;
  assign n8490 = pi18 ? n8489 : n32;
  assign n8491 = pi17 ? n335 : n8490;
  assign n8492 = pi16 ? n7943 : n8491;
  assign n8493 = pi15 ? n8485 : n8492;
  assign n8494 = pi22 ? n2895 : n204;
  assign n8495 = pi21 ? n8494 : n204;
  assign n8496 = pi20 ? n32 : n8495;
  assign n8497 = pi19 ? n32 : n8496;
  assign n8498 = pi18 ? n8497 : n7966;
  assign n8499 = pi17 ? n32 : n8498;
  assign n8500 = pi16 ? n8499 : n7973;
  assign n8501 = pi23 ? n714 : n233;
  assign n8502 = pi22 ? n8501 : n335;
  assign n8503 = pi21 ? n8502 : n233;
  assign n8504 = pi20 ? n32 : n8503;
  assign n8505 = pi19 ? n32 : n8504;
  assign n8506 = pi18 ? n8505 : n7982;
  assign n8507 = pi17 ? n32 : n8506;
  assign n8508 = pi16 ? n8507 : n7991;
  assign n8509 = pi15 ? n8500 : n8508;
  assign n8510 = pi14 ? n8493 : n8509;
  assign n8511 = pi13 ? n8479 : n8510;
  assign n8512 = pi12 ? n8463 : n8511;
  assign n8513 = pi11 ? n8383 : n8512;
  assign n8514 = pi10 ? n8271 : n8513;
  assign n8515 = pi09 ? n8007 : n8514;
  assign n8516 = pi08 ? n7999 : n8515;
  assign n8517 = pi21 ? n37 : n2946;
  assign n8518 = pi20 ? n8517 : n32;
  assign n8519 = pi19 ? n8518 : n32;
  assign n8520 = pi18 ? n37 : n8519;
  assign n8521 = pi17 ? n37 : n8520;
  assign n8522 = pi16 ? n5390 : n8521;
  assign n8523 = pi16 ? n73 : n8521;
  assign n8524 = pi15 ? n8522 : n8523;
  assign n8525 = pi14 ? n32 : n8524;
  assign n8526 = pi13 ? n32 : n8525;
  assign n8527 = pi12 ? n32 : n8526;
  assign n8528 = pi11 ? n32 : n8527;
  assign n8529 = pi10 ? n32 : n8528;
  assign n8530 = pi21 ? n37 : n2989;
  assign n8531 = pi20 ? n8530 : n32;
  assign n8532 = pi19 ? n8531 : n32;
  assign n8533 = pi18 ? n37 : n8532;
  assign n8534 = pi17 ? n37 : n8533;
  assign n8535 = pi16 ? n6787 : n8534;
  assign n8536 = pi21 ? n99 : n3022;
  assign n8537 = pi20 ? n8536 : n32;
  assign n8538 = pi19 ? n8537 : n32;
  assign n8539 = pi18 ? n37 : n8538;
  assign n8540 = pi17 ? n37 : n8539;
  assign n8541 = pi16 ? n83 : n8540;
  assign n8542 = pi15 ? n8535 : n8541;
  assign n8543 = pi21 ? n37 : n8015;
  assign n8544 = pi20 ? n8543 : n32;
  assign n8545 = pi19 ? n8544 : n32;
  assign n8546 = pi18 ? n37 : n8545;
  assign n8547 = pi17 ? n37 : n8546;
  assign n8548 = pi16 ? n8027 : n8547;
  assign n8549 = pi21 ? n139 : n8015;
  assign n8550 = pi20 ? n8549 : n32;
  assign n8551 = pi19 ? n8550 : n32;
  assign n8552 = pi18 ? n37 : n8551;
  assign n8553 = pi17 ? n37 : n8552;
  assign n8554 = pi16 ? n1130 : n8553;
  assign n8555 = pi15 ? n8548 : n8554;
  assign n8556 = pi14 ? n8542 : n8555;
  assign n8557 = pi22 ? n587 : n32;
  assign n8558 = pi21 ? n37 : n8557;
  assign n8559 = pi20 ? n8558 : n32;
  assign n8560 = pi19 ? n8559 : n32;
  assign n8561 = pi18 ? n37 : n8560;
  assign n8562 = pi17 ? n37 : n8561;
  assign n8563 = pi16 ? n2461 : n8562;
  assign n8564 = pi20 ? n37 : n7322;
  assign n8565 = pi19 ? n8564 : n37;
  assign n8566 = pi18 ? n37 : n8565;
  assign n8567 = pi22 ? n7326 : n5011;
  assign n8568 = pi21 ? n37 : n8567;
  assign n8569 = pi20 ? n37 : n8568;
  assign n8570 = pi19 ? n8569 : n37;
  assign n8571 = pi21 ? n37 : n8044;
  assign n8572 = pi20 ? n8571 : n32;
  assign n8573 = pi19 ? n8572 : n32;
  assign n8574 = pi18 ? n8570 : n8573;
  assign n8575 = pi17 ? n8566 : n8574;
  assign n8576 = pi16 ? n439 : n8575;
  assign n8577 = pi15 ? n8563 : n8576;
  assign n8578 = pi20 ? n99 : n169;
  assign n8579 = pi19 ? n8578 : n99;
  assign n8580 = pi18 ? n99 : n8579;
  assign n8581 = pi21 ? n99 : n5875;
  assign n8582 = pi20 ? n99 : n8581;
  assign n8583 = pi19 ? n8582 : n99;
  assign n8584 = pi18 ? n8583 : n8090;
  assign n8585 = pi17 ? n8580 : n8584;
  assign n8586 = pi16 ? n721 : n8585;
  assign n8587 = pi15 ? n8576 : n8586;
  assign n8588 = pi14 ? n8577 : n8587;
  assign n8589 = pi13 ? n8556 : n8588;
  assign n8590 = pi16 ? n721 : n8092;
  assign n8591 = pi15 ? n8586 : n8590;
  assign n8592 = pi16 ? n721 : n8099;
  assign n8593 = pi21 ? n716 : n165;
  assign n8594 = pi20 ? n32 : n8593;
  assign n8595 = pi19 ? n32 : n8594;
  assign n8596 = pi18 ? n8595 : n99;
  assign n8597 = pi17 ? n32 : n8596;
  assign n8598 = pi21 ? n99 : n2678;
  assign n8599 = pi20 ? n8598 : n32;
  assign n8600 = pi19 ? n8599 : n32;
  assign n8601 = pi18 ? n99 : n8600;
  assign n8602 = pi17 ? n99 : n8601;
  assign n8603 = pi16 ? n8597 : n8602;
  assign n8604 = pi15 ? n8592 : n8603;
  assign n8605 = pi14 ? n8591 : n8604;
  assign n8606 = pi21 ? n4237 : n2678;
  assign n8607 = pi20 ? n8606 : n32;
  assign n8608 = pi19 ? n8607 : n32;
  assign n8609 = pi18 ? n99 : n8608;
  assign n8610 = pi17 ? n99 : n8609;
  assign n8611 = pi16 ? n721 : n8610;
  assign n8612 = pi21 ? n1657 : n2700;
  assign n8613 = pi20 ? n8612 : n32;
  assign n8614 = pi19 ? n8613 : n32;
  assign n8615 = pi18 ? n99 : n8614;
  assign n8616 = pi17 ? n99 : n8615;
  assign n8617 = pi16 ? n801 : n8616;
  assign n8618 = pi15 ? n8611 : n8617;
  assign n8619 = pi18 ? n6499 : n157;
  assign n8620 = pi17 ? n32 : n8619;
  assign n8621 = pi16 ? n8620 : n8116;
  assign n8622 = pi21 ? n6132 : n3562;
  assign n8623 = pi23 ? n316 : n157;
  assign n8624 = pi22 ? n157 : n8623;
  assign n8625 = pi21 ? n157 : n8624;
  assign n8626 = pi20 ? n8622 : n8625;
  assign n8627 = pi19 ? n157 : n8626;
  assign n8628 = pi21 ? n7429 : n8624;
  assign n8629 = pi22 ? n316 : n1484;
  assign n8630 = pi21 ? n8629 : n157;
  assign n8631 = pi20 ? n8628 : n8630;
  assign n8632 = pi22 ? n8623 : n316;
  assign n8633 = pi21 ? n8632 : n157;
  assign n8634 = pi20 ? n157 : n8633;
  assign n8635 = pi19 ? n8631 : n8634;
  assign n8636 = pi18 ? n8627 : n8635;
  assign n8637 = pi21 ? n8632 : n3562;
  assign n8638 = pi21 ? n8629 : n8632;
  assign n8639 = pi20 ? n8637 : n8638;
  assign n8640 = pi22 ? n1484 : n157;
  assign n8641 = pi21 ? n8640 : n3562;
  assign n8642 = pi19 ? n8639 : n8641;
  assign n8643 = pi22 ? n1484 : n316;
  assign n8644 = pi21 ? n8643 : n928;
  assign n8645 = pi20 ? n8644 : n32;
  assign n8646 = pi19 ? n8645 : n32;
  assign n8647 = pi18 ? n8642 : n8646;
  assign n8648 = pi17 ? n8636 : n8647;
  assign n8649 = pi16 ? n6143 : n8648;
  assign n8650 = pi15 ? n8621 : n8649;
  assign n8651 = pi14 ? n8618 : n8650;
  assign n8652 = pi13 ? n8605 : n8651;
  assign n8653 = pi12 ? n8589 : n8652;
  assign n8654 = pi22 ? n37 : n889;
  assign n8655 = pi21 ? n180 : n8654;
  assign n8656 = pi20 ? n32 : n8655;
  assign n8657 = pi19 ? n32 : n8656;
  assign n8658 = pi22 ? n893 : n157;
  assign n8659 = pi21 ? n8658 : n8654;
  assign n8660 = pi21 ? n8658 : n890;
  assign n8661 = pi20 ? n8659 : n8660;
  assign n8662 = pi21 ? n4320 : n258;
  assign n8663 = pi21 ? n852 : n8658;
  assign n8664 = pi20 ? n8662 : n8663;
  assign n8665 = pi19 ? n8661 : n8664;
  assign n8666 = pi18 ? n8657 : n8665;
  assign n8667 = pi17 ? n32 : n8666;
  assign n8668 = pi21 ? n858 : n4320;
  assign n8669 = pi21 ? n258 : n852;
  assign n8670 = pi20 ? n8668 : n8669;
  assign n8671 = pi22 ? n893 : n1784;
  assign n8672 = pi21 ? n8671 : n349;
  assign n8673 = pi21 ? n8658 : n349;
  assign n8674 = pi20 ? n8672 : n8673;
  assign n8675 = pi19 ? n8670 : n8674;
  assign n8676 = pi22 ? n8623 : n157;
  assign n8677 = pi21 ? n8676 : n349;
  assign n8678 = pi22 ? n889 : n852;
  assign n8679 = pi21 ? n4780 : n8678;
  assign n8680 = pi20 ? n8677 : n8679;
  assign n8681 = pi21 ? n8658 : n858;
  assign n8682 = pi21 ? n354 : n858;
  assign n8683 = pi20 ? n8681 : n8682;
  assign n8684 = pi19 ? n8680 : n8683;
  assign n8685 = pi18 ? n8675 : n8684;
  assign n8686 = pi21 ? n354 : n349;
  assign n8687 = pi22 ? n383 : n1784;
  assign n8688 = pi21 ? n8687 : n354;
  assign n8689 = pi20 ? n8686 : n8688;
  assign n8690 = pi22 ? n1784 : n889;
  assign n8691 = pi22 ? n852 : n383;
  assign n8692 = pi21 ? n8690 : n8691;
  assign n8693 = pi22 ? n1784 : n852;
  assign n8694 = pi21 ? n8693 : n8691;
  assign n8695 = pi20 ? n8692 : n8694;
  assign n8696 = pi19 ? n8689 : n8695;
  assign n8697 = pi22 ? n1784 : n1484;
  assign n8698 = pi21 ? n8697 : n928;
  assign n8699 = pi20 ? n8698 : n32;
  assign n8700 = pi19 ? n8699 : n32;
  assign n8701 = pi18 ? n8696 : n8700;
  assign n8702 = pi17 ? n8685 : n8701;
  assign n8703 = pi16 ? n8667 : n8702;
  assign n8704 = pi21 ? n180 : n1696;
  assign n8705 = pi20 ? n32 : n8704;
  assign n8706 = pi19 ? n32 : n8705;
  assign n8707 = pi21 ? n37 : n1696;
  assign n8708 = pi21 ? n1056 : n820;
  assign n8709 = pi20 ? n8707 : n8708;
  assign n8710 = pi21 ? n297 : n921;
  assign n8711 = pi20 ? n8710 : n1026;
  assign n8712 = pi19 ? n8709 : n8711;
  assign n8713 = pi18 ? n8706 : n8712;
  assign n8714 = pi17 ? n32 : n8713;
  assign n8715 = pi19 ? n926 : n139;
  assign n8716 = pi20 ? n139 : n360;
  assign n8717 = pi19 ? n8716 : n139;
  assign n8718 = pi18 ? n8715 : n8717;
  assign n8719 = pi21 ? n1785 : n349;
  assign n8720 = pi20 ? n139 : n8719;
  assign n8721 = pi19 ? n8720 : n6208;
  assign n8722 = pi21 ? n1785 : n1009;
  assign n8723 = pi20 ? n8722 : n32;
  assign n8724 = pi19 ? n8723 : n32;
  assign n8725 = pi18 ? n8721 : n8724;
  assign n8726 = pi17 ? n8718 : n8725;
  assign n8727 = pi16 ? n8714 : n8726;
  assign n8728 = pi15 ? n8703 : n8727;
  assign n8729 = pi21 ? n3073 : n375;
  assign n8730 = pi20 ? n37 : n8729;
  assign n8731 = pi21 ? n1711 : n1721;
  assign n8732 = pi20 ? n8731 : n942;
  assign n8733 = pi19 ? n8730 : n8732;
  assign n8734 = pi18 ? n374 : n8733;
  assign n8735 = pi17 ? n32 : n8734;
  assign n8736 = pi19 ? n1804 : n139;
  assign n8737 = pi18 ? n8736 : n139;
  assign n8738 = pi19 ? n940 : n3578;
  assign n8739 = pi18 ? n8738 : n8724;
  assign n8740 = pi17 ? n8737 : n8739;
  assign n8741 = pi16 ? n8735 : n8740;
  assign n8742 = pi21 ? n37 : n3073;
  assign n8743 = pi20 ? n37 : n8742;
  assign n8744 = pi20 ? n1705 : n1707;
  assign n8745 = pi19 ? n8743 : n8744;
  assign n8746 = pi18 ? n374 : n8745;
  assign n8747 = pi17 ? n32 : n8746;
  assign n8748 = pi21 ? n1793 : n32;
  assign n8749 = pi20 ? n8748 : n32;
  assign n8750 = pi19 ? n8749 : n32;
  assign n8751 = pi18 ? n139 : n8750;
  assign n8752 = pi17 ? n139 : n8751;
  assign n8753 = pi16 ? n8747 : n8752;
  assign n8754 = pi15 ? n8741 : n8753;
  assign n8755 = pi14 ? n8728 : n8754;
  assign n8756 = pi20 ? n37 : n1694;
  assign n8757 = pi19 ? n37 : n8756;
  assign n8758 = pi18 ? n374 : n8757;
  assign n8759 = pi17 ? n32 : n8758;
  assign n8760 = pi20 ? n1708 : n139;
  assign n8761 = pi19 ? n8760 : n139;
  assign n8762 = pi18 ? n8761 : n139;
  assign n8763 = pi17 ? n8762 : n8751;
  assign n8764 = pi16 ? n8759 : n8763;
  assign n8765 = pi20 ? n3096 : n139;
  assign n8766 = pi19 ? n8765 : n139;
  assign n8767 = pi18 ? n8766 : n139;
  assign n8768 = pi21 ? n916 : n32;
  assign n8769 = pi20 ? n8768 : n32;
  assign n8770 = pi19 ? n8769 : n32;
  assign n8771 = pi18 ? n139 : n8770;
  assign n8772 = pi17 ? n8767 : n8771;
  assign n8773 = pi16 ? n439 : n8772;
  assign n8774 = pi15 ? n8764 : n8773;
  assign n8775 = pi21 ? n37 : n295;
  assign n8776 = pi20 ? n8775 : n1747;
  assign n8777 = pi19 ? n8776 : n139;
  assign n8778 = pi18 ? n8777 : n139;
  assign n8779 = pi18 ? n139 : n7498;
  assign n8780 = pi17 ? n8778 : n8779;
  assign n8781 = pi16 ? n439 : n8780;
  assign n8782 = pi21 ? n1696 : n346;
  assign n8783 = pi20 ? n37 : n8782;
  assign n8784 = pi22 ? n1043 : n316;
  assign n8785 = pi21 ? n1529 : n8784;
  assign n8786 = pi21 ? n139 : n8784;
  assign n8787 = pi20 ? n8785 : n8786;
  assign n8788 = pi19 ? n8783 : n8787;
  assign n8789 = pi18 ? n8788 : n347;
  assign n8790 = pi20 ? n347 : n1008;
  assign n8791 = pi20 ? n356 : n5317;
  assign n8792 = pi19 ? n8790 : n8791;
  assign n8793 = pi21 ? n346 : n32;
  assign n8794 = pi20 ? n8793 : n32;
  assign n8795 = pi19 ? n8794 : n32;
  assign n8796 = pi18 ? n8792 : n8795;
  assign n8797 = pi17 ? n8789 : n8796;
  assign n8798 = pi16 ? n439 : n8797;
  assign n8799 = pi15 ? n8781 : n8798;
  assign n8800 = pi14 ? n8774 : n8799;
  assign n8801 = pi13 ? n8755 : n8800;
  assign n8802 = pi20 ? n37 : n3299;
  assign n8803 = pi21 ? n37 : n4973;
  assign n8804 = pi20 ? n8803 : n2008;
  assign n8805 = pi19 ? n8802 : n8804;
  assign n8806 = pi21 ? n4975 : n335;
  assign n8807 = pi20 ? n1893 : n8806;
  assign n8808 = pi19 ? n8807 : n335;
  assign n8809 = pi18 ? n8805 : n8808;
  assign n8810 = pi21 ? n1079 : n32;
  assign n8811 = pi20 ? n8810 : n32;
  assign n8812 = pi19 ? n8811 : n32;
  assign n8813 = pi18 ? n335 : n8812;
  assign n8814 = pi17 ? n8809 : n8813;
  assign n8815 = pi16 ? n439 : n8814;
  assign n8816 = pi21 ? n570 : n580;
  assign n8817 = pi20 ? n4971 : n8816;
  assign n8818 = pi19 ? n37 : n8817;
  assign n8819 = pi18 ? n37 : n8818;
  assign n8820 = pi21 ? n4975 : n1943;
  assign n8821 = pi20 ? n604 : n8820;
  assign n8822 = pi21 ? n574 : n1943;
  assign n8823 = pi21 ? n566 : n1943;
  assign n8824 = pi20 ? n8822 : n8823;
  assign n8825 = pi19 ? n8821 : n8824;
  assign n8826 = pi18 ? n8825 : n8812;
  assign n8827 = pi17 ? n8819 : n8826;
  assign n8828 = pi16 ? n439 : n8827;
  assign n8829 = pi15 ? n8815 : n8828;
  assign n8830 = pi21 ? n583 : n506;
  assign n8831 = pi19 ? n4972 : n8830;
  assign n8832 = pi18 ? n37 : n8831;
  assign n8833 = pi22 ? n583 : n456;
  assign n8834 = pi22 ? n566 : n455;
  assign n8835 = pi21 ? n8833 : n8834;
  assign n8836 = pi21 ? n2007 : n4973;
  assign n8837 = pi20 ? n8835 : n8836;
  assign n8838 = pi21 ? n580 : n7606;
  assign n8839 = pi21 ? n37 : n1083;
  assign n8840 = pi20 ? n8838 : n8839;
  assign n8841 = pi19 ? n8837 : n8840;
  assign n8842 = pi22 ? n204 : n4079;
  assign n8843 = pi21 ? n8842 : n32;
  assign n8844 = pi20 ? n8843 : n32;
  assign n8845 = pi19 ? n8844 : n32;
  assign n8846 = pi18 ? n8841 : n8845;
  assign n8847 = pi17 ? n8832 : n8846;
  assign n8848 = pi16 ? n439 : n8847;
  assign n8849 = pi21 ? n6376 : n32;
  assign n8850 = pi20 ? n8849 : n32;
  assign n8851 = pi19 ? n8850 : n32;
  assign n8852 = pi18 ? n37 : n8851;
  assign n8853 = pi17 ? n37 : n8852;
  assign n8854 = pi16 ? n439 : n8853;
  assign n8855 = pi15 ? n8848 : n8854;
  assign n8856 = pi14 ? n8829 : n8855;
  assign n8857 = pi21 ? n584 : n335;
  assign n8858 = pi20 ? n37 : n8857;
  assign n8859 = pi19 ? n37 : n8858;
  assign n8860 = pi22 ? n335 : n6365;
  assign n8861 = pi21 ? n8860 : n32;
  assign n8862 = pi20 ? n8861 : n32;
  assign n8863 = pi19 ? n8862 : n32;
  assign n8864 = pi18 ? n8859 : n8863;
  assign n8865 = pi17 ? n37 : n8864;
  assign n8866 = pi16 ? n439 : n8865;
  assign n8867 = pi20 ? n37 : n5778;
  assign n8868 = pi19 ? n37 : n8867;
  assign n8869 = pi22 ? n335 : n1070;
  assign n8870 = pi21 ? n8869 : n32;
  assign n8871 = pi20 ? n8870 : n32;
  assign n8872 = pi19 ? n8871 : n32;
  assign n8873 = pi18 ? n8868 : n8872;
  assign n8874 = pi17 ? n37 : n8873;
  assign n8875 = pi16 ? n439 : n8874;
  assign n8876 = pi15 ? n8866 : n8875;
  assign n8877 = pi18 ? n8868 : n7671;
  assign n8878 = pi17 ? n37 : n8877;
  assign n8879 = pi16 ? n439 : n8878;
  assign n8880 = pi23 ? n1590 : n37;
  assign n8881 = pi22 ? n8880 : n37;
  assign n8882 = pi21 ? n8881 : n37;
  assign n8883 = pi20 ? n32 : n8882;
  assign n8884 = pi19 ? n32 : n8883;
  assign n8885 = pi20 ? n3335 : n577;
  assign n8886 = pi19 ? n642 : n8885;
  assign n8887 = pi18 ? n8884 : n8886;
  assign n8888 = pi17 ? n32 : n8887;
  assign n8889 = pi20 ? n569 : n638;
  assign n8890 = pi19 ? n8889 : n571;
  assign n8891 = pi20 ? n610 : n604;
  assign n8892 = pi19 ? n8891 : n612;
  assign n8893 = pi18 ? n8890 : n8892;
  assign n8894 = pi20 ? n649 : n610;
  assign n8895 = pi19 ? n8894 : n7685;
  assign n8896 = pi18 ? n8895 : n7671;
  assign n8897 = pi17 ? n8893 : n8896;
  assign n8898 = pi16 ? n8888 : n8897;
  assign n8899 = pi15 ? n8879 : n8898;
  assign n8900 = pi14 ? n8876 : n8899;
  assign n8901 = pi13 ? n8856 : n8900;
  assign n8902 = pi12 ? n8801 : n8901;
  assign n8903 = pi11 ? n8653 : n8902;
  assign n8904 = pi20 ? n604 : n569;
  assign n8905 = pi19 ? n642 : n8904;
  assign n8906 = pi18 ? n374 : n8905;
  assign n8907 = pi17 ? n32 : n8906;
  assign n8908 = pi20 ? n3335 : n642;
  assign n8909 = pi20 ? n570 : n571;
  assign n8910 = pi19 ? n8908 : n8909;
  assign n8911 = pi19 ? n335 : n4984;
  assign n8912 = pi18 ? n8910 : n8911;
  assign n8913 = pi20 ? n647 : n639;
  assign n8914 = pi20 ? n335 : n6377;
  assign n8915 = pi19 ? n8913 : n8914;
  assign n8916 = pi22 ? n233 : n317;
  assign n8917 = pi21 ? n8916 : n32;
  assign n8918 = pi20 ? n8917 : n32;
  assign n8919 = pi19 ? n8918 : n32;
  assign n8920 = pi18 ? n8915 : n8919;
  assign n8921 = pi17 ? n8912 : n8920;
  assign n8922 = pi16 ? n8907 : n8921;
  assign n8923 = pi18 ? n2102 : n8919;
  assign n8924 = pi17 ? n37 : n8923;
  assign n8925 = pi16 ? n439 : n8924;
  assign n8926 = pi15 ? n8922 : n8925;
  assign n8927 = pi21 ? n37 : n233;
  assign n8928 = pi20 ? n37 : n8927;
  assign n8929 = pi19 ? n37 : n8928;
  assign n8930 = pi22 ? n233 : n5631;
  assign n8931 = pi21 ? n8930 : n32;
  assign n8932 = pi20 ? n8931 : n32;
  assign n8933 = pi19 ? n8932 : n32;
  assign n8934 = pi18 ? n8929 : n8933;
  assign n8935 = pi17 ? n37 : n8934;
  assign n8936 = pi16 ? n439 : n8935;
  assign n8937 = pi22 ? n233 : n2468;
  assign n8938 = pi21 ? n8937 : n32;
  assign n8939 = pi20 ? n8938 : n32;
  assign n8940 = pi19 ? n8939 : n32;
  assign n8941 = pi18 ? n37 : n8940;
  assign n8942 = pi17 ? n37 : n8941;
  assign n8943 = pi16 ? n439 : n8942;
  assign n8944 = pi15 ? n8936 : n8943;
  assign n8945 = pi14 ? n8926 : n8944;
  assign n8946 = pi22 ? n233 : n532;
  assign n8947 = pi21 ? n8946 : n32;
  assign n8948 = pi20 ? n8947 : n32;
  assign n8949 = pi19 ? n8948 : n32;
  assign n8950 = pi18 ? n2102 : n8949;
  assign n8951 = pi17 ? n37 : n8950;
  assign n8952 = pi16 ? n439 : n8951;
  assign n8953 = pi15 ? n8952 : n4857;
  assign n8954 = pi18 ? n37 : n8297;
  assign n8955 = pi17 ? n37 : n8954;
  assign n8956 = pi16 ? n439 : n8955;
  assign n8957 = pi22 ? n686 : n706;
  assign n8958 = pi21 ? n8957 : n32;
  assign n8959 = pi20 ? n8958 : n32;
  assign n8960 = pi19 ? n8959 : n32;
  assign n8961 = pi18 ? n7732 : n8960;
  assign n8962 = pi17 ? n37 : n8961;
  assign n8963 = pi16 ? n439 : n8962;
  assign n8964 = pi15 ? n8956 : n8963;
  assign n8965 = pi14 ? n8953 : n8964;
  assign n8966 = pi13 ? n8945 : n8965;
  assign n8967 = pi21 ? n2256 : n32;
  assign n8968 = pi20 ? n8967 : n32;
  assign n8969 = pi19 ? n8968 : n32;
  assign n8970 = pi18 ? n6404 : n8969;
  assign n8971 = pi17 ? n37 : n8970;
  assign n8972 = pi16 ? n439 : n8971;
  assign n8973 = pi18 ? n6404 : n7726;
  assign n8974 = pi17 ? n37 : n8973;
  assign n8975 = pi16 ? n439 : n8974;
  assign n8976 = pi15 ? n8972 : n8975;
  assign n8977 = pi22 ? n4537 : n158;
  assign n8978 = pi21 ? n99 : n8977;
  assign n8979 = pi20 ? n99 : n8978;
  assign n8980 = pi19 ? n99 : n8979;
  assign n8981 = pi18 ? n8980 : n7726;
  assign n8982 = pi17 ? n99 : n8981;
  assign n8983 = pi16 ? n744 : n8982;
  assign n8984 = pi18 ? n7756 : n3212;
  assign n8985 = pi17 ? n99 : n8984;
  assign n8986 = pi16 ? n744 : n8985;
  assign n8987 = pi15 ? n8983 : n8986;
  assign n8988 = pi14 ? n8976 : n8987;
  assign n8989 = pi22 ? n2767 : n32;
  assign n8990 = pi21 ? n8989 : n32;
  assign n8991 = pi20 ? n8990 : n32;
  assign n8992 = pi19 ? n8991 : n32;
  assign n8993 = pi18 ? n5087 : n8992;
  assign n8994 = pi17 ? n99 : n8993;
  assign n8995 = pi16 ? n744 : n8994;
  assign n8996 = pi20 ? n157 : n6491;
  assign n8997 = pi19 ? n157 : n8996;
  assign n8998 = pi18 ? n8997 : n4118;
  assign n8999 = pi17 ? n157 : n8998;
  assign n9000 = pi16 ? n5910 : n8999;
  assign n9001 = pi15 ? n8995 : n9000;
  assign n9002 = pi20 ? n157 : n278;
  assign n9003 = pi19 ? n157 : n9002;
  assign n9004 = pi18 ? n5171 : n9003;
  assign n9005 = pi17 ? n32 : n9004;
  assign n9006 = pi16 ? n9005 : n8999;
  assign n9007 = pi21 ? n7815 : n3002;
  assign n9008 = pi20 ? n7096 : n9007;
  assign n9009 = pi19 ? n9008 : n7088;
  assign n9010 = pi18 ? n5874 : n9009;
  assign n9011 = pi17 ? n32 : n9010;
  assign n9012 = pi20 ? n8391 : n3011;
  assign n9013 = pi21 ? n157 : n3002;
  assign n9014 = pi19 ? n9012 : n9013;
  assign n9015 = pi21 ? n3002 : n157;
  assign n9016 = pi20 ? n9015 : n7815;
  assign n9017 = pi20 ? n157 : n7816;
  assign n9018 = pi19 ? n9016 : n9017;
  assign n9019 = pi18 ? n9014 : n9018;
  assign n9020 = pi20 ? n6523 : n7816;
  assign n9021 = pi21 ? n157 : n6461;
  assign n9022 = pi20 ? n157 : n9021;
  assign n9023 = pi19 ? n9020 : n9022;
  assign n9024 = pi18 ? n9023 : n5832;
  assign n9025 = pi17 ? n9019 : n9024;
  assign n9026 = pi16 ? n9011 : n9025;
  assign n9027 = pi15 ? n9006 : n9026;
  assign n9028 = pi14 ? n9001 : n9027;
  assign n9029 = pi13 ? n8988 : n9028;
  assign n9030 = pi12 ? n8966 : n9029;
  assign n9031 = pi19 ? n99 : n7795;
  assign n9032 = pi18 ? n9031 : n5832;
  assign n9033 = pi17 ? n99 : n9032;
  assign n9034 = pi16 ? n721 : n9033;
  assign n9035 = pi20 ? n157 : n7435;
  assign n9036 = pi19 ? n99 : n9035;
  assign n9037 = pi18 ? n9036 : n2655;
  assign n9038 = pi17 ? n99 : n9037;
  assign n9039 = pi16 ? n721 : n9038;
  assign n9040 = pi15 ? n9034 : n9039;
  assign n9041 = pi18 ? n9036 : n1824;
  assign n9042 = pi17 ? n99 : n9041;
  assign n9043 = pi16 ? n721 : n9042;
  assign n9044 = pi21 ? n157 : n8119;
  assign n9045 = pi20 ? n157 : n9044;
  assign n9046 = pi19 ? n139 : n9045;
  assign n9047 = pi18 ? n9046 : n1824;
  assign n9048 = pi17 ? n139 : n9047;
  assign n9049 = pi16 ? n915 : n9048;
  assign n9050 = pi15 ? n9043 : n9049;
  assign n9051 = pi14 ? n9040 : n9050;
  assign n9052 = pi19 ? n139 : n7859;
  assign n9053 = pi18 ? n9052 : n1824;
  assign n9054 = pi17 ? n139 : n9053;
  assign n9055 = pi16 ? n915 : n9054;
  assign n9056 = pi21 ? n910 : n349;
  assign n9057 = pi20 ? n32 : n9056;
  assign n9058 = pi19 ? n32 : n9057;
  assign n9059 = pi20 ? n3172 : n6930;
  assign n9060 = pi20 ? n1001 : n1008;
  assign n9061 = pi19 ? n9059 : n9060;
  assign n9062 = pi18 ? n9058 : n9061;
  assign n9063 = pi17 ? n32 : n9062;
  assign n9064 = pi20 ? n360 : n1022;
  assign n9065 = pi21 ? n316 : n346;
  assign n9066 = pi20 ? n9065 : n316;
  assign n9067 = pi19 ? n9064 : n9066;
  assign n9068 = pi20 ? n316 : n2353;
  assign n9069 = pi19 ? n316 : n9068;
  assign n9070 = pi18 ? n9067 : n9069;
  assign n9071 = pi20 ? n4437 : n2353;
  assign n9072 = pi19 ? n9071 : n316;
  assign n9073 = pi18 ? n9072 : n1824;
  assign n9074 = pi17 ? n9070 : n9073;
  assign n9075 = pi16 ? n9063 : n9074;
  assign n9076 = pi15 ? n9055 : n9075;
  assign n9077 = pi18 ? n7881 : n9069;
  assign n9078 = pi17 ? n32 : n9077;
  assign n9079 = pi18 ? n316 : n1824;
  assign n9080 = pi17 ? n316 : n9079;
  assign n9081 = pi16 ? n9078 : n9080;
  assign n9082 = pi21 ? n1785 : n316;
  assign n9083 = pi20 ? n316 : n9082;
  assign n9084 = pi19 ? n316 : n9083;
  assign n9085 = pi18 ? n5285 : n9084;
  assign n9086 = pi17 ? n32 : n9085;
  assign n9087 = pi16 ? n9086 : n7885;
  assign n9088 = pi15 ? n9081 : n9087;
  assign n9089 = pi14 ? n9076 : n9088;
  assign n9090 = pi13 ? n9051 : n9089;
  assign n9091 = pi21 ? n4472 : n316;
  assign n9092 = pi20 ? n32 : n9091;
  assign n9093 = pi19 ? n32 : n9092;
  assign n9094 = pi20 ? n6241 : n3255;
  assign n9095 = pi19 ? n316 : n9094;
  assign n9096 = pi18 ? n9093 : n9095;
  assign n9097 = pi17 ? n32 : n9096;
  assign n9098 = pi16 ? n9097 : n7885;
  assign n9099 = pi21 ? n1037 : n316;
  assign n9100 = pi20 ? n32 : n9099;
  assign n9101 = pi19 ? n32 : n9100;
  assign n9102 = pi21 ? n316 : n820;
  assign n9103 = pi21 ? n297 : n316;
  assign n9104 = pi20 ? n9102 : n9103;
  assign n9105 = pi19 ? n316 : n9104;
  assign n9106 = pi18 ? n9101 : n9105;
  assign n9107 = pi17 ? n32 : n9106;
  assign n9108 = pi16 ? n9107 : n7885;
  assign n9109 = pi15 ? n9098 : n9108;
  assign n9110 = pi20 ? n139 : n316;
  assign n9111 = pi19 ? n139 : n9110;
  assign n9112 = pi18 ? n9111 : n32;
  assign n9113 = pi17 ? n139 : n9112;
  assign n9114 = pi16 ? n915 : n9113;
  assign n9115 = pi21 ? n296 : n570;
  assign n9116 = pi20 ? n32 : n9115;
  assign n9117 = pi19 ? n32 : n9116;
  assign n9118 = pi21 ? n3073 : n570;
  assign n9119 = pi22 ? n295 : n335;
  assign n9120 = pi21 ? n9119 : n3073;
  assign n9121 = pi20 ? n9118 : n9120;
  assign n9122 = pi22 ? n335 : n139;
  assign n9123 = pi23 ? n335 : n139;
  assign n9124 = pi22 ? n9123 : n37;
  assign n9125 = pi21 ? n9122 : n9124;
  assign n9126 = pi22 ? n9123 : n335;
  assign n9127 = pi21 ? n297 : n9126;
  assign n9128 = pi20 ? n9125 : n9127;
  assign n9129 = pi19 ? n9121 : n9128;
  assign n9130 = pi18 ? n9117 : n9129;
  assign n9131 = pi17 ? n32 : n9130;
  assign n9132 = pi21 ? n820 : n9119;
  assign n9133 = pi22 ? n139 : n566;
  assign n9134 = pi21 ? n9133 : n9119;
  assign n9135 = pi20 ? n9132 : n9134;
  assign n9136 = pi22 ? n1043 : n9123;
  assign n9137 = pi21 ? n9136 : n9122;
  assign n9138 = pi22 ? n335 : n9123;
  assign n9139 = pi20 ? n9137 : n9138;
  assign n9140 = pi19 ? n9135 : n9139;
  assign n9141 = pi21 ? n9122 : n9126;
  assign n9142 = pi20 ? n9122 : n9141;
  assign n9143 = pi22 ? n139 : n335;
  assign n9144 = pi22 ? n139 : n9123;
  assign n9145 = pi21 ? n9143 : n9144;
  assign n9146 = pi22 ? n335 : n1043;
  assign n9147 = pi21 ? n9146 : n9126;
  assign n9148 = pi20 ? n9145 : n9147;
  assign n9149 = pi19 ? n9142 : n9148;
  assign n9150 = pi18 ? n9140 : n9149;
  assign n9151 = pi21 ? n9126 : n9144;
  assign n9152 = pi20 ? n9151 : n9147;
  assign n9153 = pi22 ? n9123 : n316;
  assign n9154 = pi20 ? n9153 : n6582;
  assign n9155 = pi19 ? n9152 : n9154;
  assign n9156 = pi18 ? n9155 : n32;
  assign n9157 = pi17 ? n9150 : n9156;
  assign n9158 = pi16 ? n9131 : n9157;
  assign n9159 = pi15 ? n9114 : n9158;
  assign n9160 = pi14 ? n9109 : n9159;
  assign n9161 = pi20 ? n4991 : n335;
  assign n9162 = pi19 ? n335 : n9161;
  assign n9163 = pi18 ? n602 : n9162;
  assign n9164 = pi17 ? n32 : n9163;
  assign n9165 = pi22 ? n4079 : n5369;
  assign n9166 = pi21 ? n1079 : n9165;
  assign n9167 = pi20 ? n335 : n9166;
  assign n9168 = pi19 ? n335 : n9167;
  assign n9169 = pi18 ? n9168 : n32;
  assign n9170 = pi17 ? n335 : n9169;
  assign n9171 = pi16 ? n9164 : n9170;
  assign n9172 = pi22 ? n3762 : n688;
  assign n9173 = pi21 ? n204 : n9172;
  assign n9174 = pi20 ? n335 : n9173;
  assign n9175 = pi19 ? n335 : n9174;
  assign n9176 = pi18 ? n9175 : n32;
  assign n9177 = pi17 ? n335 : n9176;
  assign n9178 = pi16 ? n2035 : n9177;
  assign n9179 = pi15 ? n9171 : n9178;
  assign n9180 = pi21 ? n204 : n335;
  assign n9181 = pi21 ? n3759 : n204;
  assign n9182 = pi20 ? n9180 : n9181;
  assign n9183 = pi19 ? n204 : n9182;
  assign n9184 = pi18 ? n5987 : n9183;
  assign n9185 = pi17 ? n32 : n9184;
  assign n9186 = pi22 ? n3762 : n706;
  assign n9187 = pi21 ? n204 : n9186;
  assign n9188 = pi20 ? n204 : n9187;
  assign n9189 = pi19 ? n204 : n9188;
  assign n9190 = pi18 ? n9189 : n32;
  assign n9191 = pi17 ? n204 : n9190;
  assign n9192 = pi16 ? n9185 : n9191;
  assign n9193 = pi21 ? n1078 : n233;
  assign n9194 = pi20 ? n32 : n9193;
  assign n9195 = pi19 ? n32 : n9194;
  assign n9196 = pi22 ? n99 : n233;
  assign n9197 = pi21 ? n9196 : n233;
  assign n9198 = pi20 ? n7980 : n9197;
  assign n9199 = pi19 ? n233 : n9198;
  assign n9200 = pi18 ? n9195 : n9199;
  assign n9201 = pi17 ? n32 : n9200;
  assign n9202 = pi22 ? n1070 : n706;
  assign n9203 = pi21 ? n335 : n9202;
  assign n9204 = pi20 ? n335 : n9203;
  assign n9205 = pi19 ? n7985 : n9204;
  assign n9206 = pi18 ? n9205 : n32;
  assign n9207 = pi17 ? n233 : n9206;
  assign n9208 = pi16 ? n9201 : n9207;
  assign n9209 = pi15 ? n9192 : n9208;
  assign n9210 = pi14 ? n9179 : n9209;
  assign n9211 = pi13 ? n9160 : n9210;
  assign n9212 = pi12 ? n9090 : n9211;
  assign n9213 = pi11 ? n9030 : n9212;
  assign n9214 = pi10 ? n8903 : n9213;
  assign n9215 = pi09 ? n8529 : n9214;
  assign n9216 = pi15 ? n32 : n8523;
  assign n9217 = pi16 ? n6787 : n8521;
  assign n9218 = pi16 ? n83 : n8521;
  assign n9219 = pi15 ? n9217 : n9218;
  assign n9220 = pi14 ? n9216 : n9219;
  assign n9221 = pi13 ? n32 : n9220;
  assign n9222 = pi12 ? n32 : n9221;
  assign n9223 = pi11 ? n32 : n9222;
  assign n9224 = pi10 ? n32 : n9223;
  assign n9225 = pi16 ? n8027 : n8534;
  assign n9226 = pi16 ? n1130 : n8540;
  assign n9227 = pi15 ? n9225 : n9226;
  assign n9228 = pi21 ? n32 : n3779;
  assign n9229 = pi20 ? n32 : n9228;
  assign n9230 = pi19 ? n32 : n9229;
  assign n9231 = pi18 ? n9230 : n37;
  assign n9232 = pi17 ? n32 : n9231;
  assign n9233 = pi16 ? n9232 : n8547;
  assign n9234 = pi16 ? n2461 : n8553;
  assign n9235 = pi15 ? n9233 : n9234;
  assign n9236 = pi14 ? n9227 : n9235;
  assign n9237 = pi16 ? n439 : n8562;
  assign n9238 = pi22 ? n1370 : n32;
  assign n9239 = pi21 ? n37 : n9238;
  assign n9240 = pi20 ? n9239 : n32;
  assign n9241 = pi19 ? n9240 : n32;
  assign n9242 = pi18 ? n8570 : n9241;
  assign n9243 = pi17 ? n8566 : n9242;
  assign n9244 = pi16 ? n439 : n9243;
  assign n9245 = pi15 ? n9237 : n9244;
  assign n9246 = pi22 ? n1378 : n32;
  assign n9247 = pi21 ? n99 : n9246;
  assign n9248 = pi20 ? n9247 : n32;
  assign n9249 = pi19 ? n9248 : n32;
  assign n9250 = pi18 ? n8583 : n9249;
  assign n9251 = pi17 ? n8580 : n9250;
  assign n9252 = pi16 ? n744 : n9251;
  assign n9253 = pi15 ? n9244 : n9252;
  assign n9254 = pi14 ? n9245 : n9253;
  assign n9255 = pi13 ? n9236 : n9254;
  assign n9256 = pi21 ? n99 : n2565;
  assign n9257 = pi20 ? n9256 : n32;
  assign n9258 = pi19 ? n9257 : n32;
  assign n9259 = pi18 ? n99 : n9258;
  assign n9260 = pi17 ? n99 : n9259;
  assign n9261 = pi16 ? n744 : n9260;
  assign n9262 = pi15 ? n9252 : n9261;
  assign n9263 = pi21 ? n739 : n165;
  assign n9264 = pi20 ? n32 : n9263;
  assign n9265 = pi19 ? n32 : n9264;
  assign n9266 = pi18 ? n9265 : n99;
  assign n9267 = pi17 ? n32 : n9266;
  assign n9268 = pi22 ? n235 : n32;
  assign n9269 = pi21 ? n99 : n9268;
  assign n9270 = pi20 ? n9269 : n32;
  assign n9271 = pi19 ? n9270 : n32;
  assign n9272 = pi18 ? n99 : n9271;
  assign n9273 = pi17 ? n99 : n9272;
  assign n9274 = pi16 ? n9267 : n9273;
  assign n9275 = pi15 ? n9261 : n9274;
  assign n9276 = pi14 ? n9262 : n9275;
  assign n9277 = pi21 ? n4237 : n2578;
  assign n9278 = pi20 ? n9277 : n32;
  assign n9279 = pi19 ? n9278 : n32;
  assign n9280 = pi18 ? n99 : n9279;
  assign n9281 = pi17 ? n99 : n9280;
  assign n9282 = pi16 ? n744 : n9281;
  assign n9283 = pi21 ? n99 : n2637;
  assign n9284 = pi20 ? n9283 : n32;
  assign n9285 = pi19 ? n9284 : n32;
  assign n9286 = pi18 ? n99 : n9285;
  assign n9287 = pi17 ? n99 : n9286;
  assign n9288 = pi16 ? n801 : n9287;
  assign n9289 = pi15 ? n9282 : n9288;
  assign n9290 = pi18 ? n7119 : n157;
  assign n9291 = pi17 ? n32 : n9290;
  assign n9292 = pi23 ? n778 : n32;
  assign n9293 = pi22 ? n9292 : n32;
  assign n9294 = pi21 ? n157 : n9293;
  assign n9295 = pi20 ? n9294 : n32;
  assign n9296 = pi19 ? n9295 : n32;
  assign n9297 = pi18 ? n157 : n9296;
  assign n9298 = pi17 ? n157 : n9297;
  assign n9299 = pi16 ? n9291 : n9298;
  assign n9300 = pi15 ? n9299 : n8649;
  assign n9301 = pi14 ? n9289 : n9300;
  assign n9302 = pi13 ? n9276 : n9301;
  assign n9303 = pi12 ? n9255 : n9302;
  assign n9304 = pi21 ? n244 : n8654;
  assign n9305 = pi21 ? n1526 : n1711;
  assign n9306 = pi20 ? n9304 : n9305;
  assign n9307 = pi22 ? n852 : n295;
  assign n9308 = pi21 ? n9307 : n258;
  assign n9309 = pi21 ? n858 : n1526;
  assign n9310 = pi20 ? n9308 : n9309;
  assign n9311 = pi19 ? n9306 : n9310;
  assign n9312 = pi18 ? n8657 : n9311;
  assign n9313 = pi17 ? n32 : n9312;
  assign n9314 = pi21 ? n139 : n9307;
  assign n9315 = pi20 ? n9314 : n869;
  assign n9316 = pi22 ? n295 : n1784;
  assign n9317 = pi21 ? n9316 : n349;
  assign n9318 = pi21 ? n1526 : n139;
  assign n9319 = pi20 ? n9317 : n9318;
  assign n9320 = pi19 ? n9315 : n9319;
  assign n9321 = pi22 ? n348 : n157;
  assign n9322 = pi21 ? n9321 : n139;
  assign n9323 = pi22 ? n1043 : n852;
  assign n9324 = pi21 ? n4429 : n9323;
  assign n9325 = pi20 ? n9322 : n9324;
  assign n9326 = pi21 ? n354 : n139;
  assign n9327 = pi20 ? n9318 : n9326;
  assign n9328 = pi19 ? n9325 : n9327;
  assign n9329 = pi18 ? n9320 : n9328;
  assign n9330 = pi20 ? n8686 : n9317;
  assign n9331 = pi22 ? n1784 : n1043;
  assign n9332 = pi21 ? n9331 : n9307;
  assign n9333 = pi21 ? n3617 : n9307;
  assign n9334 = pi20 ? n9332 : n9333;
  assign n9335 = pi19 ? n9330 : n9334;
  assign n9336 = pi21 ? n1784 : n928;
  assign n9337 = pi20 ? n9336 : n32;
  assign n9338 = pi19 ? n9337 : n32;
  assign n9339 = pi18 ? n9335 : n9338;
  assign n9340 = pi17 ? n9329 : n9339;
  assign n9341 = pi16 ? n9313 : n9340;
  assign n9342 = pi20 ? n37 : n8708;
  assign n9343 = pi19 ? n9342 : n8711;
  assign n9344 = pi18 ? n374 : n9343;
  assign n9345 = pi17 ? n32 : n9344;
  assign n9346 = pi16 ? n9345 : n8726;
  assign n9347 = pi15 ? n9341 : n9346;
  assign n9348 = pi21 ? n1711 : n297;
  assign n9349 = pi20 ? n9348 : n942;
  assign n9350 = pi19 ? n37 : n9349;
  assign n9351 = pi18 ? n374 : n9350;
  assign n9352 = pi17 ? n32 : n9351;
  assign n9353 = pi16 ? n9352 : n8740;
  assign n9354 = pi21 ? n37 : n3668;
  assign n9355 = pi20 ? n9354 : n1694;
  assign n9356 = pi19 ? n37 : n9355;
  assign n9357 = pi18 ? n374 : n9356;
  assign n9358 = pi17 ? n32 : n9357;
  assign n9359 = pi16 ? n9358 : n8752;
  assign n9360 = pi15 ? n9353 : n9359;
  assign n9361 = pi14 ? n9347 : n9360;
  assign n9362 = pi17 ? n8767 : n8751;
  assign n9363 = pi16 ? n439 : n9362;
  assign n9364 = pi15 ? n9363 : n8773;
  assign n9365 = pi20 ? n8742 : n1761;
  assign n9366 = pi19 ? n9365 : n139;
  assign n9367 = pi18 ? n9366 : n139;
  assign n9368 = pi17 ? n9367 : n8779;
  assign n9369 = pi16 ? n439 : n9368;
  assign n9370 = pi21 ? n37 : n8784;
  assign n9371 = pi20 ? n37 : n9370;
  assign n9372 = pi21 ? n375 : n8784;
  assign n9373 = pi20 ? n9372 : n8786;
  assign n9374 = pi19 ? n9371 : n9373;
  assign n9375 = pi18 ? n9374 : n347;
  assign n9376 = pi17 ? n9375 : n8796;
  assign n9377 = pi16 ? n439 : n9376;
  assign n9378 = pi15 ? n9369 : n9377;
  assign n9379 = pi14 ? n9364 : n9378;
  assign n9380 = pi13 ? n9361 : n9379;
  assign n9381 = pi19 ? n37 : n4972;
  assign n9382 = pi20 ? n8816 : n7591;
  assign n9383 = pi19 ? n9382 : n335;
  assign n9384 = pi18 ? n9381 : n9383;
  assign n9385 = pi17 ? n9384 : n8813;
  assign n9386 = pi16 ? n439 : n9385;
  assign n9387 = pi15 ? n9386 : n8828;
  assign n9388 = pi20 ? n37 : n8839;
  assign n9389 = pi19 ? n37 : n9388;
  assign n9390 = pi21 ? n204 : n32;
  assign n9391 = pi20 ? n9390 : n32;
  assign n9392 = pi19 ? n9391 : n32;
  assign n9393 = pi18 ? n9389 : n9392;
  assign n9394 = pi17 ? n37 : n9393;
  assign n9395 = pi16 ? n439 : n9394;
  assign n9396 = pi15 ? n9395 : n8854;
  assign n9397 = pi14 ? n9387 : n9396;
  assign n9398 = pi22 ? n335 : n4925;
  assign n9399 = pi21 ? n9398 : n32;
  assign n9400 = pi20 ? n9399 : n32;
  assign n9401 = pi19 ? n9400 : n32;
  assign n9402 = pi18 ? n8859 : n9401;
  assign n9403 = pi17 ? n37 : n9402;
  assign n9404 = pi16 ? n439 : n9403;
  assign n9405 = pi22 ? n335 : n2121;
  assign n9406 = pi21 ? n9405 : n32;
  assign n9407 = pi20 ? n9406 : n32;
  assign n9408 = pi19 ? n9407 : n32;
  assign n9409 = pi18 ? n8868 : n9408;
  assign n9410 = pi17 ? n37 : n9409;
  assign n9411 = pi16 ? n439 : n9410;
  assign n9412 = pi15 ? n9404 : n9411;
  assign n9413 = pi22 ? n335 : n759;
  assign n9414 = pi21 ? n9413 : n32;
  assign n9415 = pi20 ? n9414 : n32;
  assign n9416 = pi19 ? n9415 : n32;
  assign n9417 = pi18 ? n7677 : n9416;
  assign n9418 = pi17 ? n37 : n9417;
  assign n9419 = pi16 ? n439 : n9418;
  assign n9420 = pi18 ? n374 : n8886;
  assign n9421 = pi17 ? n32 : n9420;
  assign n9422 = pi18 ? n8895 : n9416;
  assign n9423 = pi17 ? n8893 : n9422;
  assign n9424 = pi16 ? n9421 : n9423;
  assign n9425 = pi15 ? n9419 : n9424;
  assign n9426 = pi14 ? n9412 : n9425;
  assign n9427 = pi13 ? n9397 : n9426;
  assign n9428 = pi12 ? n9380 : n9427;
  assign n9429 = pi11 ? n9303 : n9428;
  assign n9430 = pi22 ? n233 : n3338;
  assign n9431 = pi21 ? n9430 : n32;
  assign n9432 = pi20 ? n9431 : n32;
  assign n9433 = pi19 ? n9432 : n32;
  assign n9434 = pi18 ? n8915 : n9433;
  assign n9435 = pi17 ? n8912 : n9434;
  assign n9436 = pi16 ? n8907 : n9435;
  assign n9437 = pi18 ? n2102 : n9433;
  assign n9438 = pi17 ? n37 : n9437;
  assign n9439 = pi16 ? n439 : n9438;
  assign n9440 = pi15 ? n9436 : n9439;
  assign n9441 = pi21 ? n665 : n32;
  assign n9442 = pi20 ? n9441 : n32;
  assign n9443 = pi19 ? n9442 : n32;
  assign n9444 = pi18 ? n8929 : n9443;
  assign n9445 = pi17 ? n37 : n9444;
  assign n9446 = pi16 ? n439 : n9445;
  assign n9447 = pi18 ? n37 : n9443;
  assign n9448 = pi17 ? n37 : n9447;
  assign n9449 = pi16 ? n439 : n9448;
  assign n9450 = pi15 ? n9446 : n9449;
  assign n9451 = pi14 ? n9440 : n9450;
  assign n9452 = pi18 ? n2102 : n9443;
  assign n9453 = pi17 ? n37 : n9452;
  assign n9454 = pi16 ? n439 : n9453;
  assign n9455 = pi15 ? n9454 : n9449;
  assign n9456 = pi21 ? n1423 : n32;
  assign n9457 = pi20 ? n9456 : n32;
  assign n9458 = pi19 ? n9457 : n32;
  assign n9459 = pi18 ? n37 : n9458;
  assign n9460 = pi17 ? n37 : n9459;
  assign n9461 = pi16 ? n439 : n9460;
  assign n9462 = pi22 ? n686 : n317;
  assign n9463 = pi21 ? n9462 : n32;
  assign n9464 = pi20 ? n9463 : n32;
  assign n9465 = pi19 ? n9464 : n32;
  assign n9466 = pi18 ? n7732 : n9465;
  assign n9467 = pi17 ? n37 : n9466;
  assign n9468 = pi16 ? n439 : n9467;
  assign n9469 = pi15 ? n9461 : n9468;
  assign n9470 = pi14 ? n9455 : n9469;
  assign n9471 = pi13 ? n9451 : n9470;
  assign n9472 = pi21 ? n689 : n32;
  assign n9473 = pi20 ? n9472 : n32;
  assign n9474 = pi19 ? n9473 : n32;
  assign n9475 = pi18 ? n6404 : n9474;
  assign n9476 = pi17 ? n37 : n9475;
  assign n9477 = pi16 ? n439 : n9476;
  assign n9478 = pi18 ? n6404 : n8297;
  assign n9479 = pi17 ? n37 : n9478;
  assign n9480 = pi16 ? n439 : n9479;
  assign n9481 = pi15 ? n9477 : n9480;
  assign n9482 = pi21 ? n8486 : n32;
  assign n9483 = pi20 ? n9482 : n32;
  assign n9484 = pi19 ? n9483 : n32;
  assign n9485 = pi18 ? n1667 : n9484;
  assign n9486 = pi17 ? n99 : n9485;
  assign n9487 = pi16 ? n744 : n9486;
  assign n9488 = pi18 ? n7756 : n4010;
  assign n9489 = pi17 ? n99 : n9488;
  assign n9490 = pi16 ? n744 : n9489;
  assign n9491 = pi15 ? n9487 : n9490;
  assign n9492 = pi14 ? n9481 : n9491;
  assign n9493 = pi18 ? n5087 : n7726;
  assign n9494 = pi17 ? n99 : n9493;
  assign n9495 = pi16 ? n744 : n9494;
  assign n9496 = pi18 ? n8997 : n7051;
  assign n9497 = pi17 ? n157 : n9496;
  assign n9498 = pi16 ? n7793 : n9497;
  assign n9499 = pi15 ? n9495 : n9498;
  assign n9500 = pi16 ? n9005 : n9497;
  assign n9501 = pi21 ? n5871 : n165;
  assign n9502 = pi20 ? n32 : n9501;
  assign n9503 = pi19 ? n32 : n9502;
  assign n9504 = pi20 ? n7091 : n7807;
  assign n9505 = pi19 ? n9504 : n7088;
  assign n9506 = pi18 ? n9503 : n9505;
  assign n9507 = pi17 ? n32 : n9506;
  assign n9508 = pi20 ? n8391 : n3004;
  assign n9509 = pi20 ? n7824 : n6508;
  assign n9510 = pi19 ? n9508 : n9509;
  assign n9511 = pi21 ? n165 : n7815;
  assign n9512 = pi21 ? n7815 : n775;
  assign n9513 = pi20 ? n9511 : n9512;
  assign n9514 = pi20 ? n3002 : n7088;
  assign n9515 = pi19 ? n9513 : n9514;
  assign n9516 = pi18 ? n9510 : n9515;
  assign n9517 = pi20 ? n7807 : n7088;
  assign n9518 = pi19 ? n9517 : n9022;
  assign n9519 = pi18 ? n9518 : n5832;
  assign n9520 = pi17 ? n9516 : n9519;
  assign n9521 = pi16 ? n9507 : n9520;
  assign n9522 = pi15 ? n9500 : n9521;
  assign n9523 = pi14 ? n9499 : n9522;
  assign n9524 = pi13 ? n9492 : n9523;
  assign n9525 = pi12 ? n9471 : n9524;
  assign n9526 = pi16 ? n744 : n9033;
  assign n9527 = pi16 ? n744 : n9038;
  assign n9528 = pi15 ? n9526 : n9527;
  assign n9529 = pi18 ? n9036 : n2681;
  assign n9530 = pi17 ? n99 : n9529;
  assign n9531 = pi16 ? n744 : n9530;
  assign n9532 = pi18 ? n2277 : n2703;
  assign n9533 = pi17 ? n139 : n9532;
  assign n9534 = pi16 ? n915 : n9533;
  assign n9535 = pi15 ? n9531 : n9534;
  assign n9536 = pi14 ? n9528 : n9535;
  assign n9537 = pi21 ? n359 : n356;
  assign n9538 = pi20 ? n1001 : n9537;
  assign n9539 = pi19 ? n9059 : n9538;
  assign n9540 = pi18 ? n9058 : n9539;
  assign n9541 = pi17 ? n32 : n9540;
  assign n9542 = pi16 ? n9541 : n9074;
  assign n9543 = pi15 ? n9055 : n9542;
  assign n9544 = pi21 ? n354 : n316;
  assign n9545 = pi20 ? n316 : n9544;
  assign n9546 = pi19 ? n316 : n9545;
  assign n9547 = pi18 ? n7881 : n9546;
  assign n9548 = pi17 ? n32 : n9547;
  assign n9549 = pi16 ? n9548 : n9080;
  assign n9550 = pi15 ? n9549 : n9087;
  assign n9551 = pi14 ? n9543 : n9550;
  assign n9552 = pi13 ? n9536 : n9551;
  assign n9553 = pi16 ? n2291 : n9113;
  assign n9554 = pi21 ? n180 : n570;
  assign n9555 = pi20 ? n32 : n9554;
  assign n9556 = pi19 ? n32 : n9555;
  assign n9557 = pi20 ? n639 : n9120;
  assign n9558 = pi19 ? n9557 : n9128;
  assign n9559 = pi18 ? n9556 : n9558;
  assign n9560 = pi17 ? n32 : n9559;
  assign n9561 = pi21 ? n9133 : n569;
  assign n9562 = pi20 ? n9132 : n9561;
  assign n9563 = pi22 ? n335 : n295;
  assign n9564 = pi21 ? n580 : n9563;
  assign n9565 = pi20 ? n9564 : n9138;
  assign n9566 = pi19 ? n9562 : n9565;
  assign n9567 = pi21 ? n9563 : n9122;
  assign n9568 = pi20 ? n9567 : n9141;
  assign n9569 = pi21 ? n9119 : n9133;
  assign n9570 = pi20 ? n9569 : n1893;
  assign n9571 = pi19 ? n9568 : n9570;
  assign n9572 = pi18 ? n9566 : n9571;
  assign n9573 = pi21 ? n9126 : n9133;
  assign n9574 = pi20 ? n9573 : n1893;
  assign n9575 = pi22 ? n566 : n316;
  assign n9576 = pi21 ? n9575 : n9153;
  assign n9577 = pi20 ? n9576 : n316;
  assign n9578 = pi19 ? n9574 : n9577;
  assign n9579 = pi18 ? n9578 : n32;
  assign n9580 = pi17 ? n9572 : n9579;
  assign n9581 = pi16 ? n9560 : n9580;
  assign n9582 = pi15 ? n9553 : n9581;
  assign n9583 = pi14 ? n9109 : n9582;
  assign n9584 = pi22 ? n4079 : n396;
  assign n9585 = pi21 ? n1079 : n9584;
  assign n9586 = pi20 ? n335 : n9585;
  assign n9587 = pi19 ? n335 : n9586;
  assign n9588 = pi18 ? n9587 : n32;
  assign n9589 = pi17 ? n335 : n9588;
  assign n9590 = pi16 ? n9164 : n9589;
  assign n9591 = pi22 ? n3762 : n5369;
  assign n9592 = pi21 ? n204 : n9591;
  assign n9593 = pi20 ? n335 : n9592;
  assign n9594 = pi19 ? n335 : n9593;
  assign n9595 = pi18 ? n9594 : n32;
  assign n9596 = pi17 ? n335 : n9595;
  assign n9597 = pi16 ? n2035 : n9596;
  assign n9598 = pi15 ? n9590 : n9597;
  assign n9599 = pi14 ? n9598 : n9209;
  assign n9600 = pi13 ? n9583 : n9599;
  assign n9601 = pi12 ? n9552 : n9600;
  assign n9602 = pi11 ? n9525 : n9601;
  assign n9603 = pi10 ? n9429 : n9602;
  assign n9604 = pi09 ? n9224 : n9603;
  assign n9605 = pi08 ? n9215 : n9604;
  assign n9606 = pi07 ? n8516 : n9605;
  assign n9607 = pi21 ? n37 : n3791;
  assign n9608 = pi20 ? n9607 : n32;
  assign n9609 = pi19 ? n9608 : n32;
  assign n9610 = pi18 ? n37 : n9609;
  assign n9611 = pi17 ? n37 : n9610;
  assign n9612 = pi16 ? n73 : n9611;
  assign n9613 = pi15 ? n32 : n9612;
  assign n9614 = pi16 ? n6787 : n9611;
  assign n9615 = pi16 ? n83 : n9611;
  assign n9616 = pi15 ? n9614 : n9615;
  assign n9617 = pi14 ? n9613 : n9616;
  assign n9618 = pi13 ? n32 : n9617;
  assign n9619 = pi12 ? n32 : n9618;
  assign n9620 = pi11 ? n32 : n9619;
  assign n9621 = pi10 ? n32 : n9620;
  assign n9622 = pi21 ? n37 : n3832;
  assign n9623 = pi20 ? n9622 : n32;
  assign n9624 = pi19 ? n9623 : n32;
  assign n9625 = pi18 ? n37 : n9624;
  assign n9626 = pi17 ? n37 : n9625;
  assign n9627 = pi16 ? n8027 : n9626;
  assign n9628 = pi23 ? n99 : n260;
  assign n9629 = pi22 ? n9628 : n32;
  assign n9630 = pi21 ? n37 : n9629;
  assign n9631 = pi20 ? n9630 : n32;
  assign n9632 = pi19 ? n9631 : n32;
  assign n9633 = pi18 ? n37 : n9632;
  assign n9634 = pi17 ? n37 : n9633;
  assign n9635 = pi16 ? n1130 : n9634;
  assign n9636 = pi15 ? n9627 : n9635;
  assign n9637 = pi21 ? n37 : n3022;
  assign n9638 = pi20 ? n9637 : n32;
  assign n9639 = pi19 ? n9638 : n32;
  assign n9640 = pi18 ? n37 : n9639;
  assign n9641 = pi17 ? n37 : n9640;
  assign n9642 = pi16 ? n9232 : n9641;
  assign n9643 = pi16 ? n2461 : n9641;
  assign n9644 = pi15 ? n9642 : n9643;
  assign n9645 = pi14 ? n9636 : n9644;
  assign n9646 = pi23 ? n1342 : n32;
  assign n9647 = pi22 ? n9646 : n32;
  assign n9648 = pi21 ? n37 : n9647;
  assign n9649 = pi20 ? n9648 : n32;
  assign n9650 = pi19 ? n9649 : n32;
  assign n9651 = pi18 ? n37 : n9650;
  assign n9652 = pi17 ? n37 : n9651;
  assign n9653 = pi16 ? n439 : n9652;
  assign n9654 = pi21 ? n5015 : n7327;
  assign n9655 = pi20 ? n7331 : n9654;
  assign n9656 = pi19 ? n37 : n9655;
  assign n9657 = pi22 ? n363 : n5011;
  assign n9658 = pi21 ? n9657 : n37;
  assign n9659 = pi20 ? n9654 : n9658;
  assign n9660 = pi21 ? n5015 : n37;
  assign n9661 = pi21 ? n8567 : n37;
  assign n9662 = pi20 ? n9660 : n9661;
  assign n9663 = pi19 ? n9659 : n9662;
  assign n9664 = pi18 ? n9656 : n9663;
  assign n9665 = pi21 ? n8567 : n7327;
  assign n9666 = pi22 ? n7326 : n363;
  assign n9667 = pi21 ? n9657 : n9666;
  assign n9668 = pi20 ? n9665 : n9667;
  assign n9669 = pi21 ? n5012 : n3392;
  assign n9670 = pi21 ? n5012 : n6401;
  assign n9671 = pi20 ? n9669 : n9670;
  assign n9672 = pi19 ? n9668 : n9671;
  assign n9673 = pi21 ? n5012 : n9238;
  assign n9674 = pi20 ? n9673 : n32;
  assign n9675 = pi19 ? n9674 : n32;
  assign n9676 = pi18 ? n9672 : n9675;
  assign n9677 = pi17 ? n9664 : n9676;
  assign n9678 = pi16 ? n439 : n9677;
  assign n9679 = pi15 ? n9653 : n9678;
  assign n9680 = pi21 ? n99 : n9238;
  assign n9681 = pi20 ? n9680 : n32;
  assign n9682 = pi19 ? n9681 : n32;
  assign n9683 = pi18 ? n99 : n9682;
  assign n9684 = pi17 ? n99 : n9683;
  assign n9685 = pi16 ? n721 : n9684;
  assign n9686 = pi21 ? n159 : n165;
  assign n9687 = pi21 ? n775 : n165;
  assign n9688 = pi20 ? n9686 : n9687;
  assign n9689 = pi19 ? n99 : n9688;
  assign n9690 = pi20 ? n9687 : n3014;
  assign n9691 = pi21 ? n5875 : n99;
  assign n9692 = pi20 ? n802 : n9691;
  assign n9693 = pi19 ? n9690 : n9692;
  assign n9694 = pi18 ? n9689 : n9693;
  assign n9695 = pi20 ? n7104 : n5887;
  assign n9696 = pi21 ? n168 : n159;
  assign n9697 = pi20 ? n6490 : n9696;
  assign n9698 = pi19 ? n9695 : n9697;
  assign n9699 = pi21 ? n168 : n9246;
  assign n9700 = pi20 ? n9699 : n32;
  assign n9701 = pi19 ? n9700 : n32;
  assign n9702 = pi18 ? n9698 : n9701;
  assign n9703 = pi17 ? n9694 : n9702;
  assign n9704 = pi16 ? n721 : n9703;
  assign n9705 = pi15 ? n9685 : n9704;
  assign n9706 = pi14 ? n9679 : n9705;
  assign n9707 = pi13 ? n9645 : n9706;
  assign n9708 = pi20 ? n9686 : n166;
  assign n9709 = pi19 ? n99 : n9708;
  assign n9710 = pi20 ? n99 : n9691;
  assign n9711 = pi19 ? n9690 : n9710;
  assign n9712 = pi18 ? n9709 : n9711;
  assign n9713 = pi17 ? n9712 : n9702;
  assign n9714 = pi16 ? n721 : n9713;
  assign n9715 = pi20 ? n99 : n802;
  assign n9716 = pi19 ? n9715 : n99;
  assign n9717 = pi18 ? n719 : n9716;
  assign n9718 = pi17 ? n32 : n9717;
  assign n9719 = pi16 ? n9718 : n9260;
  assign n9720 = pi15 ? n9714 : n9719;
  assign n9721 = pi16 ? n801 : n9260;
  assign n9722 = pi21 ? n796 : n168;
  assign n9723 = pi20 ? n32 : n9722;
  assign n9724 = pi19 ? n32 : n9723;
  assign n9725 = pi18 ? n9724 : n99;
  assign n9726 = pi17 ? n32 : n9725;
  assign n9727 = pi21 ? n99 : n2578;
  assign n9728 = pi20 ? n9727 : n32;
  assign n9729 = pi19 ? n9728 : n32;
  assign n9730 = pi18 ? n99 : n9729;
  assign n9731 = pi17 ? n99 : n9730;
  assign n9732 = pi16 ? n9726 : n9731;
  assign n9733 = pi15 ? n9721 : n9732;
  assign n9734 = pi14 ? n9720 : n9733;
  assign n9735 = pi16 ? n744 : n9731;
  assign n9736 = pi15 ? n9735 : n9288;
  assign n9737 = pi21 ? n180 : n775;
  assign n9738 = pi20 ? n32 : n9737;
  assign n9739 = pi19 ? n32 : n9738;
  assign n9740 = pi20 ? n6500 : n99;
  assign n9741 = pi19 ? n9740 : n99;
  assign n9742 = pi18 ? n9739 : n9741;
  assign n9743 = pi17 ? n32 : n9742;
  assign n9744 = pi16 ? n9743 : n9287;
  assign n9745 = pi21 ? n381 : n384;
  assign n9746 = pi20 ? n37 : n9745;
  assign n9747 = pi21 ? n3562 : n316;
  assign n9748 = pi20 ? n7571 : n9747;
  assign n9749 = pi19 ? n9746 : n9748;
  assign n9750 = pi18 ? n374 : n9749;
  assign n9751 = pi17 ? n32 : n9750;
  assign n9752 = pi21 ? n7429 : n316;
  assign n9753 = pi20 ? n9752 : n316;
  assign n9754 = pi19 ? n9753 : n316;
  assign n9755 = pi18 ? n9754 : n316;
  assign n9756 = pi20 ? n2330 : n32;
  assign n9757 = pi19 ? n9756 : n32;
  assign n9758 = pi18 ? n316 : n9757;
  assign n9759 = pi17 ? n9755 : n9758;
  assign n9760 = pi16 ? n9751 : n9759;
  assign n9761 = pi15 ? n9744 : n9760;
  assign n9762 = pi14 ? n9736 : n9761;
  assign n9763 = pi13 ? n9734 : n9762;
  assign n9764 = pi12 ? n9707 : n9763;
  assign n9765 = pi20 ? n37 : n942;
  assign n9766 = pi19 ? n37 : n9765;
  assign n9767 = pi18 ? n374 : n9766;
  assign n9768 = pi17 ? n32 : n9767;
  assign n9769 = pi20 ? n942 : n139;
  assign n9770 = pi19 ? n9769 : n139;
  assign n9771 = pi18 ? n9770 : n8717;
  assign n9772 = pi20 ? n139 : n7170;
  assign n9773 = pi21 ? n356 : n139;
  assign n9774 = pi19 ? n9772 : n9773;
  assign n9775 = pi21 ? n139 : n882;
  assign n9776 = pi20 ? n9775 : n32;
  assign n9777 = pi19 ? n9776 : n32;
  assign n9778 = pi18 ? n9774 : n9777;
  assign n9779 = pi17 ? n9771 : n9778;
  assign n9780 = pi16 ? n9768 : n9779;
  assign n9781 = pi18 ? n8766 : n8717;
  assign n9782 = pi21 ? n139 : n928;
  assign n9783 = pi20 ? n9782 : n32;
  assign n9784 = pi19 ? n9783 : n32;
  assign n9785 = pi18 ? n9774 : n9784;
  assign n9786 = pi17 ? n9781 : n9785;
  assign n9787 = pi16 ? n439 : n9786;
  assign n9788 = pi15 ? n9780 : n9787;
  assign n9789 = pi20 ? n3656 : n139;
  assign n9790 = pi19 ? n9789 : n139;
  assign n9791 = pi18 ? n9790 : n139;
  assign n9792 = pi18 ? n139 : n9784;
  assign n9793 = pi17 ? n9791 : n9792;
  assign n9794 = pi16 ? n439 : n9793;
  assign n9795 = pi20 ? n37 : n139;
  assign n9796 = pi19 ? n9795 : n139;
  assign n9797 = pi18 ? n9796 : n139;
  assign n9798 = pi21 ? n139 : n2553;
  assign n9799 = pi20 ? n9798 : n32;
  assign n9800 = pi19 ? n9799 : n32;
  assign n9801 = pi18 ? n139 : n9800;
  assign n9802 = pi17 ? n9797 : n9801;
  assign n9803 = pi16 ? n439 : n9802;
  assign n9804 = pi15 ? n9794 : n9803;
  assign n9805 = pi14 ? n9788 : n9804;
  assign n9806 = pi19 ? n37 : n2374;
  assign n9807 = pi18 ? n9806 : n139;
  assign n9808 = pi21 ? n139 : n8557;
  assign n9809 = pi20 ? n9808 : n32;
  assign n9810 = pi19 ? n9809 : n32;
  assign n9811 = pi18 ? n139 : n9810;
  assign n9812 = pi17 ? n9807 : n9811;
  assign n9813 = pi16 ? n439 : n9812;
  assign n9814 = pi20 ? n37 : n3096;
  assign n9815 = pi19 ? n9814 : n139;
  assign n9816 = pi18 ? n37 : n9815;
  assign n9817 = pi21 ? n9143 : n2553;
  assign n9818 = pi20 ? n9817 : n32;
  assign n9819 = pi19 ? n9818 : n32;
  assign n9820 = pi18 ? n139 : n9819;
  assign n9821 = pi17 ? n9816 : n9820;
  assign n9822 = pi16 ? n439 : n9821;
  assign n9823 = pi15 ? n9813 : n9822;
  assign n9824 = pi20 ? n37 : n3086;
  assign n9825 = pi19 ? n9824 : n139;
  assign n9826 = pi18 ? n37 : n9825;
  assign n9827 = pi23 ? n139 : n335;
  assign n9828 = pi22 ? n139 : n9827;
  assign n9829 = pi21 ? n9828 : n2553;
  assign n9830 = pi20 ? n9829 : n32;
  assign n9831 = pi19 ? n9830 : n32;
  assign n9832 = pi18 ? n139 : n9831;
  assign n9833 = pi17 ? n9826 : n9832;
  assign n9834 = pi16 ? n439 : n9833;
  assign n9835 = pi22 ? n295 : n9123;
  assign n9836 = pi22 ? n335 : n9827;
  assign n9837 = pi21 ? n9835 : n9836;
  assign n9838 = pi21 ? n9144 : n9836;
  assign n9839 = pi20 ? n9837 : n9838;
  assign n9840 = pi19 ? n37 : n9839;
  assign n9841 = pi18 ? n37 : n9840;
  assign n9842 = pi21 ? n9144 : n921;
  assign n9843 = pi20 ? n9842 : n9151;
  assign n9844 = pi21 ? n9836 : n9144;
  assign n9845 = pi19 ? n9843 : n9844;
  assign n9846 = pi22 ? n335 : n364;
  assign n9847 = pi21 ? n9846 : n2553;
  assign n9848 = pi20 ? n9847 : n32;
  assign n9849 = pi19 ? n9848 : n32;
  assign n9850 = pi18 ? n9845 : n9849;
  assign n9851 = pi17 ? n9841 : n9850;
  assign n9852 = pi16 ? n439 : n9851;
  assign n9853 = pi15 ? n9834 : n9852;
  assign n9854 = pi14 ? n9823 : n9853;
  assign n9855 = pi13 ? n9805 : n9854;
  assign n9856 = pi19 ? n37 : n335;
  assign n9857 = pi18 ? n37 : n9856;
  assign n9858 = pi21 ? n1079 : n2553;
  assign n9859 = pi20 ? n9858 : n32;
  assign n9860 = pi19 ? n9859 : n32;
  assign n9861 = pi18 ? n335 : n9860;
  assign n9862 = pi17 ? n9857 : n9861;
  assign n9863 = pi16 ? n439 : n9862;
  assign n9864 = pi21 ? n1056 : n2553;
  assign n9865 = pi20 ? n9864 : n32;
  assign n9866 = pi19 ? n9865 : n32;
  assign n9867 = pi18 ? n37 : n9866;
  assign n9868 = pi17 ? n37 : n9867;
  assign n9869 = pi16 ? n439 : n9868;
  assign n9870 = pi15 ? n9863 : n9869;
  assign n9871 = pi22 ? n456 : n233;
  assign n9872 = pi21 ? n9871 : n2678;
  assign n9873 = pi20 ? n9872 : n32;
  assign n9874 = pi19 ? n9873 : n32;
  assign n9875 = pi18 ? n37 : n9874;
  assign n9876 = pi17 ? n37 : n9875;
  assign n9877 = pi16 ? n439 : n9876;
  assign n9878 = pi21 ? n2091 : n2678;
  assign n9879 = pi20 ? n9878 : n32;
  assign n9880 = pi19 ? n9879 : n32;
  assign n9881 = pi18 ? n37 : n9880;
  assign n9882 = pi17 ? n37 : n9881;
  assign n9883 = pi16 ? n439 : n9882;
  assign n9884 = pi15 ? n9877 : n9883;
  assign n9885 = pi14 ? n9870 : n9884;
  assign n9886 = pi22 ? n335 : n5782;
  assign n9887 = pi21 ? n9886 : n2700;
  assign n9888 = pi20 ? n9887 : n32;
  assign n9889 = pi19 ? n9888 : n32;
  assign n9890 = pi18 ? n37 : n9889;
  assign n9891 = pi17 ? n37 : n9890;
  assign n9892 = pi16 ? n439 : n9891;
  assign n9893 = pi21 ? n9886 : n1009;
  assign n9894 = pi20 ? n9893 : n32;
  assign n9895 = pi19 ? n9894 : n32;
  assign n9896 = pi18 ? n37 : n9895;
  assign n9897 = pi17 ? n37 : n9896;
  assign n9898 = pi16 ? n439 : n9897;
  assign n9899 = pi15 ? n9892 : n9898;
  assign n9900 = pi22 ? n335 : n6380;
  assign n9901 = pi21 ? n9900 : n32;
  assign n9902 = pi20 ? n9901 : n32;
  assign n9903 = pi19 ? n9902 : n32;
  assign n9904 = pi18 ? n37 : n9903;
  assign n9905 = pi17 ? n37 : n9904;
  assign n9906 = pi16 ? n439 : n9905;
  assign n9907 = pi14 ? n9899 : n9906;
  assign n9908 = pi13 ? n9885 : n9907;
  assign n9909 = pi12 ? n9855 : n9908;
  assign n9910 = pi11 ? n9764 : n9909;
  assign n9911 = pi20 ? n7646 : n3292;
  assign n9912 = pi21 ? n37 : n574;
  assign n9913 = pi20 ? n9912 : n37;
  assign n9914 = pi19 ? n9911 : n9913;
  assign n9915 = pi18 ? n37 : n9914;
  assign n9916 = pi20 ? n37 : n584;
  assign n9917 = pi19 ? n37 : n9916;
  assign n9918 = pi22 ? n233 : n3124;
  assign n9919 = pi21 ? n9918 : n32;
  assign n9920 = pi20 ? n9919 : n32;
  assign n9921 = pi19 ? n9920 : n32;
  assign n9922 = pi18 ? n9917 : n9921;
  assign n9923 = pi17 ? n9915 : n9922;
  assign n9924 = pi16 ? n439 : n9923;
  assign n9925 = pi22 ? n363 : n3124;
  assign n9926 = pi21 ? n9925 : n32;
  assign n9927 = pi20 ? n9926 : n32;
  assign n9928 = pi19 ? n9927 : n32;
  assign n9929 = pi18 ? n37 : n9928;
  assign n9930 = pi17 ? n37 : n9929;
  assign n9931 = pi16 ? n439 : n9930;
  assign n9932 = pi15 ? n9924 : n9931;
  assign n9933 = pi22 ? n5011 : n664;
  assign n9934 = pi21 ? n9933 : n32;
  assign n9935 = pi20 ? n9934 : n32;
  assign n9936 = pi19 ? n9935 : n32;
  assign n9937 = pi18 ? n37 : n9936;
  assign n9938 = pi17 ? n37 : n9937;
  assign n9939 = pi16 ? n439 : n9938;
  assign n9940 = pi15 ? n9939 : n9449;
  assign n9941 = pi14 ? n9932 : n9940;
  assign n9942 = pi22 ? n363 : n664;
  assign n9943 = pi21 ? n9942 : n32;
  assign n9944 = pi20 ? n9943 : n32;
  assign n9945 = pi19 ? n9944 : n32;
  assign n9946 = pi18 ? n37 : n9945;
  assign n9947 = pi17 ? n37 : n9946;
  assign n9948 = pi16 ? n439 : n9947;
  assign n9949 = pi21 ? n1408 : n32;
  assign n9950 = pi20 ? n9949 : n32;
  assign n9951 = pi19 ? n9950 : n32;
  assign n9952 = pi18 ? n37 : n9951;
  assign n9953 = pi17 ? n37 : n9952;
  assign n9954 = pi16 ? n439 : n9953;
  assign n9955 = pi15 ? n9948 : n9954;
  assign n9956 = pi22 ? n157 : n1407;
  assign n9957 = pi21 ? n9956 : n32;
  assign n9958 = pi20 ? n9957 : n32;
  assign n9959 = pi19 ? n9958 : n32;
  assign n9960 = pi18 ? n37 : n9959;
  assign n9961 = pi17 ? n37 : n9960;
  assign n9962 = pi16 ? n439 : n9961;
  assign n9963 = pi21 ? n2230 : n32;
  assign n9964 = pi20 ? n9963 : n32;
  assign n9965 = pi19 ? n9964 : n32;
  assign n9966 = pi18 ? n37 : n9965;
  assign n9967 = pi17 ? n37 : n9966;
  assign n9968 = pi16 ? n439 : n9967;
  assign n9969 = pi15 ? n9962 : n9968;
  assign n9970 = pi14 ? n9955 : n9969;
  assign n9971 = pi13 ? n9941 : n9970;
  assign n9972 = pi20 ? n99 : n37;
  assign n9973 = pi19 ? n99 : n9972;
  assign n9974 = pi18 ? n9973 : n5749;
  assign n9975 = pi17 ? n99 : n9974;
  assign n9976 = pi16 ? n201 : n9975;
  assign n9977 = pi19 ? n99 : n5121;
  assign n9978 = pi18 ? n9977 : n9474;
  assign n9979 = pi17 ? n99 : n9978;
  assign n9980 = pi16 ? n801 : n9979;
  assign n9981 = pi15 ? n9976 : n9980;
  assign n9982 = pi18 ? n99 : n9484;
  assign n9983 = pi17 ? n99 : n9982;
  assign n9984 = pi16 ? n721 : n9983;
  assign n9985 = pi19 ? n99 : n7845;
  assign n9986 = pi18 ? n9985 : n9484;
  assign n9987 = pi17 ? n99 : n9986;
  assign n9988 = pi16 ? n721 : n9987;
  assign n9989 = pi15 ? n9984 : n9988;
  assign n9990 = pi14 ? n9981 : n9989;
  assign n9991 = pi16 ? n721 : n9494;
  assign n9992 = pi19 ? n157 : n9022;
  assign n9993 = pi18 ? n9992 : n7726;
  assign n9994 = pi17 ? n157 : n9993;
  assign n9995 = pi16 ? n5910 : n9994;
  assign n9996 = pi15 ? n9991 : n9995;
  assign n9997 = pi21 ? n157 : n159;
  assign n9998 = pi20 ? n99 : n9997;
  assign n9999 = pi19 ? n99 : n9998;
  assign n10000 = pi18 ? n9999 : n3212;
  assign n10001 = pi17 ? n99 : n10000;
  assign n10002 = pi16 ? n744 : n10001;
  assign n10003 = pi15 ? n9995 : n10002;
  assign n10004 = pi14 ? n9996 : n10003;
  assign n10005 = pi13 ? n9990 : n10004;
  assign n10006 = pi12 ? n9971 : n10005;
  assign n10007 = pi18 ? n1667 : n3212;
  assign n10008 = pi17 ? n99 : n10007;
  assign n10009 = pi16 ? n744 : n10008;
  assign n10010 = pi19 ? n99 : n2242;
  assign n10011 = pi21 ? n882 : n32;
  assign n10012 = pi20 ? n10011 : n32;
  assign n10013 = pi19 ? n10012 : n32;
  assign n10014 = pi18 ? n10010 : n10013;
  assign n10015 = pi17 ? n99 : n10014;
  assign n10016 = pi16 ? n721 : n10015;
  assign n10017 = pi15 ? n10009 : n10016;
  assign n10018 = pi18 ? n2277 : n2655;
  assign n10019 = pi17 ? n139 : n10018;
  assign n10020 = pi16 ? n915 : n10019;
  assign n10021 = pi22 ? n157 : n204;
  assign n10022 = pi21 ? n248 : n10021;
  assign n10023 = pi20 ? n10022 : n7858;
  assign n10024 = pi19 ? n139 : n10023;
  assign n10025 = pi18 ? n10024 : n2655;
  assign n10026 = pi17 ? n139 : n10025;
  assign n10027 = pi16 ? n1575 : n10026;
  assign n10028 = pi15 ? n10020 : n10027;
  assign n10029 = pi14 ? n10017 : n10028;
  assign n10030 = pi19 ? n139 : n3578;
  assign n10031 = pi18 ? n1573 : n10030;
  assign n10032 = pi17 ? n32 : n10031;
  assign n10033 = pi21 ? n139 : n1027;
  assign n10034 = pi20 ? n139 : n10033;
  assign n10035 = pi19 ? n139 : n10034;
  assign n10036 = pi18 ? n10035 : n2655;
  assign n10037 = pi17 ? n139 : n10036;
  assign n10038 = pi16 ? n10032 : n10037;
  assign n10039 = pi20 ? n316 : n9065;
  assign n10040 = pi19 ? n316 : n10039;
  assign n10041 = pi18 ? n8451 : n10040;
  assign n10042 = pi17 ? n32 : n10041;
  assign n10043 = pi18 ? n316 : n2655;
  assign n10044 = pi17 ? n316 : n10043;
  assign n10045 = pi16 ? n10042 : n10044;
  assign n10046 = pi15 ? n10038 : n10045;
  assign n10047 = pi16 ? n7883 : n10044;
  assign n10048 = pi21 ? n4020 : n346;
  assign n10049 = pi20 ? n316 : n10048;
  assign n10050 = pi19 ? n316 : n10049;
  assign n10051 = pi18 ? n7881 : n10050;
  assign n10052 = pi17 ? n32 : n10051;
  assign n10053 = pi16 ? n10052 : n9080;
  assign n10054 = pi15 ? n10047 : n10053;
  assign n10055 = pi14 ? n10046 : n10054;
  assign n10056 = pi13 ? n10029 : n10055;
  assign n10057 = pi22 ? n6608 : n139;
  assign n10058 = pi21 ? n10057 : n316;
  assign n10059 = pi20 ? n32 : n10058;
  assign n10060 = pi19 ? n32 : n10059;
  assign n10061 = pi20 ? n316 : n4804;
  assign n10062 = pi19 ? n316 : n10061;
  assign n10063 = pi18 ? n10060 : n10062;
  assign n10064 = pi17 ? n32 : n10063;
  assign n10065 = pi16 ? n10064 : n9080;
  assign n10066 = pi21 ? n910 : n316;
  assign n10067 = pi20 ? n32 : n10066;
  assign n10068 = pi19 ? n32 : n10067;
  assign n10069 = pi20 ? n316 : n139;
  assign n10070 = pi19 ? n316 : n10069;
  assign n10071 = pi18 ? n10068 : n10070;
  assign n10072 = pi17 ? n32 : n10071;
  assign n10073 = pi19 ? n999 : n316;
  assign n10074 = pi18 ? n10073 : n316;
  assign n10075 = pi17 ? n10074 : n9079;
  assign n10076 = pi16 ? n10072 : n10075;
  assign n10077 = pi15 ? n10065 : n10076;
  assign n10078 = pi19 ? n139 : n2352;
  assign n10079 = pi18 ? n10078 : n1824;
  assign n10080 = pi17 ? n139 : n10079;
  assign n10081 = pi16 ? n915 : n10080;
  assign n10082 = pi22 ? n6380 : n335;
  assign n10083 = pi21 ? n335 : n10082;
  assign n10084 = pi22 ? n6380 : n316;
  assign n10085 = pi21 ? n2427 : n10084;
  assign n10086 = pi20 ? n10083 : n10085;
  assign n10087 = pi19 ? n335 : n10086;
  assign n10088 = pi18 ? n10087 : n32;
  assign n10089 = pi17 ? n335 : n10088;
  assign n10090 = pi16 ? n2035 : n10089;
  assign n10091 = pi15 ? n10081 : n10090;
  assign n10092 = pi14 ? n10077 : n10091;
  assign n10093 = pi21 ? n335 : n4938;
  assign n10094 = pi20 ? n335 : n10093;
  assign n10095 = pi19 ? n335 : n10094;
  assign n10096 = pi18 ? n7941 : n10095;
  assign n10097 = pi17 ? n32 : n10096;
  assign n10098 = pi23 ? n4145 : n395;
  assign n10099 = pi22 ? n204 : n10098;
  assign n10100 = pi21 ? n335 : n10099;
  assign n10101 = pi20 ? n335 : n10100;
  assign n10102 = pi19 ? n335 : n10101;
  assign n10103 = pi18 ? n10102 : n32;
  assign n10104 = pi17 ? n335 : n10103;
  assign n10105 = pi16 ? n10097 : n10104;
  assign n10106 = pi22 ? n204 : n1407;
  assign n10107 = pi21 ? n335 : n10106;
  assign n10108 = pi20 ? n335 : n10107;
  assign n10109 = pi19 ? n335 : n10108;
  assign n10110 = pi18 ? n10109 : n32;
  assign n10111 = pi17 ? n335 : n10110;
  assign n10112 = pi16 ? n2035 : n10111;
  assign n10113 = pi15 ? n10105 : n10112;
  assign n10114 = pi21 ? n1078 : n335;
  assign n10115 = pi20 ? n32 : n10114;
  assign n10116 = pi19 ? n32 : n10115;
  assign n10117 = pi18 ? n10116 : n335;
  assign n10118 = pi17 ? n32 : n10117;
  assign n10119 = pi22 ? n233 : n5369;
  assign n10120 = pi21 ? n335 : n10119;
  assign n10121 = pi20 ? n335 : n10120;
  assign n10122 = pi19 ? n335 : n10121;
  assign n10123 = pi18 ? n10122 : n32;
  assign n10124 = pi17 ? n335 : n10123;
  assign n10125 = pi16 ? n10118 : n10124;
  assign n10126 = pi21 ? n335 : n8916;
  assign n10127 = pi20 ? n335 : n10126;
  assign n10128 = pi19 ? n335 : n10127;
  assign n10129 = pi18 ? n10128 : n32;
  assign n10130 = pi17 ? n335 : n10129;
  assign n10131 = pi16 ? n10118 : n10130;
  assign n10132 = pi15 ? n10125 : n10131;
  assign n10133 = pi14 ? n10113 : n10132;
  assign n10134 = pi13 ? n10092 : n10133;
  assign n10135 = pi12 ? n10056 : n10134;
  assign n10136 = pi11 ? n10006 : n10135;
  assign n10137 = pi10 ? n9910 : n10136;
  assign n10138 = pi09 ? n9621 : n10137;
  assign n10139 = pi15 ? n32 : n9614;
  assign n10140 = pi16 ? n8027 : n9611;
  assign n10141 = pi15 ? n9615 : n10140;
  assign n10142 = pi14 ? n10139 : n10141;
  assign n10143 = pi13 ? n32 : n10142;
  assign n10144 = pi12 ? n32 : n10143;
  assign n10145 = pi11 ? n32 : n10144;
  assign n10146 = pi10 ? n32 : n10145;
  assign n10147 = pi16 ? n1130 : n9626;
  assign n10148 = pi16 ? n9232 : n9634;
  assign n10149 = pi15 ? n10147 : n10148;
  assign n10150 = pi21 ? n32 : n180;
  assign n10151 = pi20 ? n32 : n10150;
  assign n10152 = pi19 ? n32 : n10151;
  assign n10153 = pi18 ? n10152 : n37;
  assign n10154 = pi17 ? n32 : n10153;
  assign n10155 = pi16 ? n10154 : n9641;
  assign n10156 = pi15 ? n9643 : n10155;
  assign n10157 = pi14 ? n10149 : n10156;
  assign n10158 = pi21 ? n37 : n3066;
  assign n10159 = pi20 ? n10158 : n32;
  assign n10160 = pi19 ? n10159 : n32;
  assign n10161 = pi18 ? n37 : n10160;
  assign n10162 = pi17 ? n37 : n10161;
  assign n10163 = pi16 ? n439 : n10162;
  assign n10164 = pi23 ? n363 : n5630;
  assign n10165 = pi22 ? n10164 : n32;
  assign n10166 = pi21 ? n5012 : n10165;
  assign n10167 = pi20 ? n10166 : n32;
  assign n10168 = pi19 ? n10167 : n32;
  assign n10169 = pi18 ? n9672 : n10168;
  assign n10170 = pi17 ? n9664 : n10169;
  assign n10171 = pi16 ? n439 : n10170;
  assign n10172 = pi15 ? n10163 : n10171;
  assign n10173 = pi16 ? n744 : n9684;
  assign n10174 = pi22 ? n6114 : n32;
  assign n10175 = pi21 ? n168 : n10174;
  assign n10176 = pi20 ? n10175 : n32;
  assign n10177 = pi19 ? n10176 : n32;
  assign n10178 = pi18 ? n9698 : n10177;
  assign n10179 = pi17 ? n9694 : n10178;
  assign n10180 = pi16 ? n744 : n10179;
  assign n10181 = pi15 ? n10173 : n10180;
  assign n10182 = pi14 ? n10172 : n10181;
  assign n10183 = pi13 ? n10157 : n10182;
  assign n10184 = pi17 ? n9712 : n10178;
  assign n10185 = pi16 ? n744 : n10184;
  assign n10186 = pi18 ? n742 : n9716;
  assign n10187 = pi17 ? n32 : n10186;
  assign n10188 = pi22 ? n1185 : n32;
  assign n10189 = pi21 ? n99 : n10188;
  assign n10190 = pi20 ? n10189 : n32;
  assign n10191 = pi19 ? n10190 : n32;
  assign n10192 = pi18 ? n99 : n10191;
  assign n10193 = pi17 ? n99 : n10192;
  assign n10194 = pi16 ? n10187 : n10193;
  assign n10195 = pi15 ? n10185 : n10194;
  assign n10196 = pi21 ? n99 : n3175;
  assign n10197 = pi20 ? n10196 : n32;
  assign n10198 = pi19 ? n10197 : n32;
  assign n10199 = pi18 ? n99 : n10198;
  assign n10200 = pi17 ? n99 : n10199;
  assign n10201 = pi16 ? n801 : n10200;
  assign n10202 = pi21 ? n99 : n4109;
  assign n10203 = pi20 ? n10202 : n32;
  assign n10204 = pi19 ? n10203 : n32;
  assign n10205 = pi18 ? n99 : n10204;
  assign n10206 = pi17 ? n99 : n10205;
  assign n10207 = pi16 ? n9726 : n10206;
  assign n10208 = pi15 ? n10201 : n10207;
  assign n10209 = pi14 ? n10195 : n10208;
  assign n10210 = pi16 ? n721 : n10206;
  assign n10211 = pi21 ? n99 : n760;
  assign n10212 = pi20 ? n10211 : n32;
  assign n10213 = pi19 ? n10212 : n32;
  assign n10214 = pi18 ? n99 : n10213;
  assign n10215 = pi17 ? n99 : n10214;
  assign n10216 = pi16 ? n801 : n10215;
  assign n10217 = pi15 ? n10210 : n10216;
  assign n10218 = pi16 ? n9743 : n10215;
  assign n10219 = pi15 ? n10218 : n9760;
  assign n10220 = pi14 ? n10217 : n10219;
  assign n10221 = pi13 ? n10209 : n10220;
  assign n10222 = pi12 ? n10183 : n10221;
  assign n10223 = pi17 ? n9797 : n9811;
  assign n10224 = pi16 ? n439 : n10223;
  assign n10225 = pi15 ? n9794 : n10224;
  assign n10226 = pi14 ? n9788 : n10225;
  assign n10227 = pi21 ? n9143 : n8044;
  assign n10228 = pi20 ? n10227 : n32;
  assign n10229 = pi19 ? n10228 : n32;
  assign n10230 = pi18 ? n139 : n10229;
  assign n10231 = pi17 ? n9816 : n10230;
  assign n10232 = pi16 ? n439 : n10231;
  assign n10233 = pi15 ? n9813 : n10232;
  assign n10234 = pi22 ? n295 : n566;
  assign n10235 = pi21 ? n10234 : n9836;
  assign n10236 = pi19 ? n37 : n10235;
  assign n10237 = pi18 ? n37 : n10236;
  assign n10238 = pi21 ? n10234 : n5559;
  assign n10239 = pi20 ? n10238 : n9151;
  assign n10240 = pi21 ? n9836 : n9835;
  assign n10241 = pi19 ? n10239 : n10240;
  assign n10242 = pi18 ? n10241 : n9849;
  assign n10243 = pi17 ? n10237 : n10242;
  assign n10244 = pi16 ? n439 : n10243;
  assign n10245 = pi15 ? n9834 : n10244;
  assign n10246 = pi14 ? n10233 : n10245;
  assign n10247 = pi13 ? n10226 : n10246;
  assign n10248 = pi14 ? n9870 : n9883;
  assign n10249 = pi21 ? n2061 : n2700;
  assign n10250 = pi20 ? n10249 : n32;
  assign n10251 = pi19 ? n10250 : n32;
  assign n10252 = pi18 ? n37 : n10251;
  assign n10253 = pi17 ? n37 : n10252;
  assign n10254 = pi16 ? n439 : n10253;
  assign n10255 = pi21 ? n2061 : n1009;
  assign n10256 = pi20 ? n10255 : n32;
  assign n10257 = pi19 ? n10256 : n32;
  assign n10258 = pi18 ? n37 : n10257;
  assign n10259 = pi17 ? n37 : n10258;
  assign n10260 = pi16 ? n439 : n10259;
  assign n10261 = pi15 ? n10254 : n10260;
  assign n10262 = pi21 ? n9886 : n32;
  assign n10263 = pi20 ? n10262 : n32;
  assign n10264 = pi19 ? n10263 : n32;
  assign n10265 = pi18 ? n37 : n10264;
  assign n10266 = pi17 ? n37 : n10265;
  assign n10267 = pi16 ? n439 : n10266;
  assign n10268 = pi14 ? n10261 : n10267;
  assign n10269 = pi13 ? n10248 : n10268;
  assign n10270 = pi12 ? n10247 : n10269;
  assign n10271 = pi11 ? n10222 : n10270;
  assign n10272 = pi20 ? n7646 : n37;
  assign n10273 = pi19 ? n10272 : n37;
  assign n10274 = pi18 ? n37 : n10273;
  assign n10275 = pi22 ? n233 : n705;
  assign n10276 = pi21 ? n10275 : n32;
  assign n10277 = pi20 ? n10276 : n32;
  assign n10278 = pi19 ? n10277 : n32;
  assign n10279 = pi18 ? n37 : n10278;
  assign n10280 = pi17 ? n10274 : n10279;
  assign n10281 = pi16 ? n439 : n10280;
  assign n10282 = pi22 ? n363 : n705;
  assign n10283 = pi21 ? n10282 : n32;
  assign n10284 = pi20 ? n10283 : n32;
  assign n10285 = pi19 ? n10284 : n32;
  assign n10286 = pi18 ? n37 : n10285;
  assign n10287 = pi17 ? n37 : n10286;
  assign n10288 = pi16 ? n439 : n10287;
  assign n10289 = pi15 ? n10281 : n10288;
  assign n10290 = pi22 ? n5011 : n1388;
  assign n10291 = pi21 ? n10290 : n32;
  assign n10292 = pi20 ? n10291 : n32;
  assign n10293 = pi19 ? n10292 : n32;
  assign n10294 = pi18 ? n37 : n10293;
  assign n10295 = pi17 ? n37 : n10294;
  assign n10296 = pi16 ? n439 : n10295;
  assign n10297 = pi21 ? n1389 : n32;
  assign n10298 = pi20 ? n10297 : n32;
  assign n10299 = pi19 ? n10298 : n32;
  assign n10300 = pi18 ? n37 : n10299;
  assign n10301 = pi17 ? n37 : n10300;
  assign n10302 = pi16 ? n439 : n10301;
  assign n10303 = pi15 ? n10296 : n10302;
  assign n10304 = pi14 ? n10289 : n10303;
  assign n10305 = pi21 ? n2132 : n32;
  assign n10306 = pi20 ? n10305 : n32;
  assign n10307 = pi19 ? n10306 : n32;
  assign n10308 = pi18 ? n37 : n10307;
  assign n10309 = pi17 ? n37 : n10308;
  assign n10310 = pi16 ? n439 : n10309;
  assign n10311 = pi21 ? n2139 : n32;
  assign n10312 = pi20 ? n10311 : n32;
  assign n10313 = pi19 ? n10312 : n32;
  assign n10314 = pi18 ? n37 : n10313;
  assign n10315 = pi17 ? n37 : n10314;
  assign n10316 = pi16 ? n439 : n10315;
  assign n10317 = pi15 ? n10310 : n10316;
  assign n10318 = pi22 ? n157 : n759;
  assign n10319 = pi21 ? n10318 : n32;
  assign n10320 = pi20 ? n10319 : n32;
  assign n10321 = pi19 ? n10320 : n32;
  assign n10322 = pi18 ? n37 : n10321;
  assign n10323 = pi17 ? n37 : n10322;
  assign n10324 = pi16 ? n439 : n10323;
  assign n10325 = pi22 ? n685 : n396;
  assign n10326 = pi21 ? n10325 : n32;
  assign n10327 = pi20 ? n10326 : n32;
  assign n10328 = pi19 ? n10327 : n32;
  assign n10329 = pi18 ? n37 : n10328;
  assign n10330 = pi17 ? n37 : n10329;
  assign n10331 = pi16 ? n439 : n10330;
  assign n10332 = pi15 ? n10324 : n10331;
  assign n10333 = pi14 ? n10317 : n10332;
  assign n10334 = pi13 ? n10304 : n10333;
  assign n10335 = pi21 ? n10106 : n32;
  assign n10336 = pi20 ? n10335 : n32;
  assign n10337 = pi19 ? n10336 : n32;
  assign n10338 = pi18 ? n9973 : n10337;
  assign n10339 = pi17 ? n99 : n10338;
  assign n10340 = pi16 ? n201 : n10339;
  assign n10341 = pi23 ? n363 : n8319;
  assign n10342 = pi22 ? n10341 : n1407;
  assign n10343 = pi21 ? n10342 : n32;
  assign n10344 = pi20 ? n10343 : n32;
  assign n10345 = pi19 ? n10344 : n32;
  assign n10346 = pi18 ? n9977 : n10345;
  assign n10347 = pi17 ? n99 : n10346;
  assign n10348 = pi16 ? n801 : n10347;
  assign n10349 = pi15 ? n10340 : n10348;
  assign n10350 = pi22 ? n685 : n5369;
  assign n10351 = pi21 ? n10350 : n32;
  assign n10352 = pi20 ? n10351 : n32;
  assign n10353 = pi19 ? n10352 : n32;
  assign n10354 = pi18 ? n99 : n10353;
  assign n10355 = pi17 ? n99 : n10354;
  assign n10356 = pi16 ? n744 : n10355;
  assign n10357 = pi18 ? n9985 : n9965;
  assign n10358 = pi17 ? n99 : n10357;
  assign n10359 = pi16 ? n744 : n10358;
  assign n10360 = pi15 ? n10356 : n10359;
  assign n10361 = pi14 ? n10349 : n10360;
  assign n10362 = pi18 ? n5087 : n8297;
  assign n10363 = pi17 ? n99 : n10362;
  assign n10364 = pi16 ? n744 : n10363;
  assign n10365 = pi18 ? n9992 : n9484;
  assign n10366 = pi17 ? n157 : n10365;
  assign n10367 = pi16 ? n7793 : n10366;
  assign n10368 = pi15 ? n10364 : n10367;
  assign n10369 = pi15 ? n10367 : n10002;
  assign n10370 = pi14 ? n10368 : n10369;
  assign n10371 = pi13 ? n10361 : n10370;
  assign n10372 = pi12 ? n10334 : n10371;
  assign n10373 = pi16 ? n744 : n10015;
  assign n10374 = pi15 ? n10009 : n10373;
  assign n10375 = pi16 ? n331 : n10026;
  assign n10376 = pi15 ? n10020 : n10375;
  assign n10377 = pi14 ? n10374 : n10376;
  assign n10378 = pi18 ? n329 : n10030;
  assign n10379 = pi17 ? n32 : n10378;
  assign n10380 = pi16 ? n10379 : n10037;
  assign n10381 = pi18 ? n7881 : n10040;
  assign n10382 = pi17 ? n32 : n10381;
  assign n10383 = pi16 ? n10382 : n10044;
  assign n10384 = pi15 ? n10380 : n10383;
  assign n10385 = pi18 ? n316 : n2703;
  assign n10386 = pi17 ? n316 : n10385;
  assign n10387 = pi16 ? n10052 : n10386;
  assign n10388 = pi15 ? n10047 : n10387;
  assign n10389 = pi14 ? n10384 : n10388;
  assign n10390 = pi13 ? n10377 : n10389;
  assign n10391 = pi16 ? n10064 : n10386;
  assign n10392 = pi15 ? n10391 : n10076;
  assign n10393 = pi16 ? n2291 : n10080;
  assign n10394 = pi22 ? n8880 : n335;
  assign n10395 = pi21 ? n10394 : n335;
  assign n10396 = pi20 ? n32 : n10395;
  assign n10397 = pi19 ? n32 : n10396;
  assign n10398 = pi18 ? n10397 : n335;
  assign n10399 = pi17 ? n32 : n10398;
  assign n10400 = pi23 ? n335 : n363;
  assign n10401 = pi22 ? n10400 : n316;
  assign n10402 = pi21 ? n1578 : n10401;
  assign n10403 = pi20 ? n10083 : n10402;
  assign n10404 = pi19 ? n335 : n10403;
  assign n10405 = pi18 ? n10404 : n32;
  assign n10406 = pi17 ? n335 : n10405;
  assign n10407 = pi16 ? n10399 : n10406;
  assign n10408 = pi15 ? n10393 : n10407;
  assign n10409 = pi14 ? n10392 : n10408;
  assign n10410 = pi22 ? n204 : n1475;
  assign n10411 = pi21 ? n335 : n10410;
  assign n10412 = pi20 ? n335 : n10411;
  assign n10413 = pi19 ? n335 : n10412;
  assign n10414 = pi18 ? n10413 : n32;
  assign n10415 = pi17 ? n335 : n10414;
  assign n10416 = pi16 ? n10097 : n10415;
  assign n10417 = pi22 ? n204 : n2192;
  assign n10418 = pi21 ? n335 : n10417;
  assign n10419 = pi20 ? n335 : n10418;
  assign n10420 = pi19 ? n335 : n10419;
  assign n10421 = pi18 ? n10420 : n32;
  assign n10422 = pi17 ? n335 : n10421;
  assign n10423 = pi16 ? n2035 : n10422;
  assign n10424 = pi15 ? n10416 : n10423;
  assign n10425 = pi14 ? n10424 : n10131;
  assign n10426 = pi13 ? n10409 : n10425;
  assign n10427 = pi12 ? n10390 : n10426;
  assign n10428 = pi11 ? n10372 : n10427;
  assign n10429 = pi10 ? n10271 : n10428;
  assign n10430 = pi09 ? n10146 : n10429;
  assign n10431 = pi08 ? n10138 : n10430;
  assign n10432 = pi21 ? n37 : n4519;
  assign n10433 = pi20 ? n10432 : n32;
  assign n10434 = pi19 ? n10433 : n32;
  assign n10435 = pi18 ? n37 : n10434;
  assign n10436 = pi17 ? n37 : n10435;
  assign n10437 = pi16 ? n6787 : n10436;
  assign n10438 = pi15 ? n32 : n10437;
  assign n10439 = pi16 ? n83 : n10436;
  assign n10440 = pi16 ? n8027 : n10436;
  assign n10441 = pi15 ? n10439 : n10440;
  assign n10442 = pi14 ? n10438 : n10441;
  assign n10443 = pi13 ? n32 : n10442;
  assign n10444 = pi12 ? n32 : n10443;
  assign n10445 = pi11 ? n32 : n10444;
  assign n10446 = pi10 ? n32 : n10445;
  assign n10447 = pi21 ? n37 : n4559;
  assign n10448 = pi20 ? n10447 : n32;
  assign n10449 = pi19 ? n10448 : n32;
  assign n10450 = pi18 ? n37 : n10449;
  assign n10451 = pi17 ? n37 : n10450;
  assign n10452 = pi16 ? n1130 : n10451;
  assign n10453 = pi22 ? n139 : n32;
  assign n10454 = pi21 ? n37 : n10453;
  assign n10455 = pi20 ? n10454 : n32;
  assign n10456 = pi19 ? n10455 : n32;
  assign n10457 = pi18 ? n37 : n10456;
  assign n10458 = pi17 ? n37 : n10457;
  assign n10459 = pi16 ? n9232 : n10458;
  assign n10460 = pi15 ? n10452 : n10459;
  assign n10461 = pi22 ? n1762 : n32;
  assign n10462 = pi21 ? n37 : n10461;
  assign n10463 = pi20 ? n10462 : n32;
  assign n10464 = pi19 ? n10463 : n32;
  assign n10465 = pi18 ? n37 : n10464;
  assign n10466 = pi17 ? n37 : n10465;
  assign n10467 = pi16 ? n2461 : n10466;
  assign n10468 = pi16 ? n10154 : n10466;
  assign n10469 = pi15 ? n10467 : n10468;
  assign n10470 = pi14 ? n10460 : n10469;
  assign n10471 = pi22 ? n6798 : n32;
  assign n10472 = pi21 ? n37 : n10471;
  assign n10473 = pi20 ? n10472 : n32;
  assign n10474 = pi19 ? n10473 : n32;
  assign n10475 = pi18 ? n37 : n10474;
  assign n10476 = pi17 ? n37 : n10475;
  assign n10477 = pi16 ? n439 : n10476;
  assign n10478 = pi21 ? n6401 : n5012;
  assign n10479 = pi20 ? n37 : n10478;
  assign n10480 = pi21 ? n9666 : n5011;
  assign n10481 = pi21 ? n7327 : n9657;
  assign n10482 = pi20 ? n10480 : n10481;
  assign n10483 = pi19 ? n10479 : n10482;
  assign n10484 = pi18 ? n374 : n10483;
  assign n10485 = pi17 ? n32 : n10484;
  assign n10486 = pi21 ? n5012 : n9666;
  assign n10487 = pi20 ? n10486 : n7328;
  assign n10488 = pi22 ? n5011 : n363;
  assign n10489 = pi21 ? n9657 : n10488;
  assign n10490 = pi22 ? n363 : n7326;
  assign n10491 = pi21 ? n363 : n10490;
  assign n10492 = pi20 ? n10489 : n10491;
  assign n10493 = pi19 ? n10487 : n10492;
  assign n10494 = pi21 ? n9657 : n3392;
  assign n10495 = pi20 ? n10491 : n10494;
  assign n10496 = pi21 ? n363 : n5015;
  assign n10497 = pi21 ? n9666 : n5015;
  assign n10498 = pi20 ? n10496 : n10497;
  assign n10499 = pi19 ? n10495 : n10498;
  assign n10500 = pi18 ? n10493 : n10499;
  assign n10501 = pi21 ? n9666 : n363;
  assign n10502 = pi20 ? n10501 : n9667;
  assign n10503 = pi21 ? n5012 : n363;
  assign n10504 = pi20 ? n10503 : n10486;
  assign n10505 = pi19 ? n10502 : n10504;
  assign n10506 = pi18 ? n10505 : n10168;
  assign n10507 = pi17 ? n10500 : n10506;
  assign n10508 = pi16 ? n10485 : n10507;
  assign n10509 = pi15 ? n10477 : n10508;
  assign n10510 = pi23 ? n99 : n5630;
  assign n10511 = pi22 ? n10510 : n32;
  assign n10512 = pi21 ? n99 : n10511;
  assign n10513 = pi20 ? n10512 : n32;
  assign n10514 = pi19 ? n10513 : n32;
  assign n10515 = pi18 ? n99 : n10514;
  assign n10516 = pi17 ? n99 : n10515;
  assign n10517 = pi16 ? n721 : n10516;
  assign n10518 = pi21 ? n159 : n168;
  assign n10519 = pi20 ? n99 : n10518;
  assign n10520 = pi21 ? n3002 : n158;
  assign n10521 = pi20 ? n10520 : n7810;
  assign n10522 = pi19 ? n10519 : n10521;
  assign n10523 = pi18 ? n719 : n10522;
  assign n10524 = pi17 ? n32 : n10523;
  assign n10525 = pi21 ? n168 : n3002;
  assign n10526 = pi21 ? n158 : n165;
  assign n10527 = pi20 ? n10525 : n10526;
  assign n10528 = pi21 ? n3013 : n5899;
  assign n10529 = pi21 ? n157 : n7815;
  assign n10530 = pi20 ? n10528 : n10529;
  assign n10531 = pi19 ? n10527 : n10530;
  assign n10532 = pi21 ? n3013 : n777;
  assign n10533 = pi20 ? n10529 : n10532;
  assign n10534 = pi21 ? n3002 : n775;
  assign n10535 = pi20 ? n7818 : n10534;
  assign n10536 = pi19 ? n10533 : n10535;
  assign n10537 = pi18 ? n10531 : n10536;
  assign n10538 = pi20 ? n9015 : n5887;
  assign n10539 = pi21 ? n168 : n157;
  assign n10540 = pi20 ? n10539 : n10525;
  assign n10541 = pi19 ? n10538 : n10540;
  assign n10542 = pi18 ? n10541 : n10177;
  assign n10543 = pi17 ? n10537 : n10542;
  assign n10544 = pi16 ? n10524 : n10543;
  assign n10545 = pi15 ? n10517 : n10544;
  assign n10546 = pi14 ? n10509 : n10545;
  assign n10547 = pi13 ? n10470 : n10546;
  assign n10548 = pi20 ? n10518 : n776;
  assign n10549 = pi19 ? n99 : n10548;
  assign n10550 = pi20 ? n775 : n3014;
  assign n10551 = pi20 ? n99 : n3003;
  assign n10552 = pi19 ? n10550 : n10551;
  assign n10553 = pi18 ? n10549 : n10552;
  assign n10554 = pi20 ? n10534 : n10532;
  assign n10555 = pi19 ? n10554 : n6490;
  assign n10556 = pi18 ? n10555 : n10177;
  assign n10557 = pi17 ? n10553 : n10556;
  assign n10558 = pi16 ? n801 : n10557;
  assign n10559 = pi18 ? n799 : n9716;
  assign n10560 = pi17 ? n32 : n10559;
  assign n10561 = pi16 ? n10560 : n10193;
  assign n10562 = pi15 ? n10558 : n10561;
  assign n10563 = pi16 ? n744 : n10193;
  assign n10564 = pi23 ? n99 : n624;
  assign n10565 = pi22 ? n10564 : n32;
  assign n10566 = pi21 ? n99 : n10565;
  assign n10567 = pi20 ? n10566 : n32;
  assign n10568 = pi19 ? n10567 : n32;
  assign n10569 = pi18 ? n99 : n10568;
  assign n10570 = pi17 ? n99 : n10569;
  assign n10571 = pi16 ? n9726 : n10570;
  assign n10572 = pi15 ? n10563 : n10571;
  assign n10573 = pi14 ? n10562 : n10572;
  assign n10574 = pi21 ? n99 : n748;
  assign n10575 = pi20 ? n10574 : n32;
  assign n10576 = pi19 ? n10575 : n32;
  assign n10577 = pi18 ? n99 : n10576;
  assign n10578 = pi17 ? n99 : n10577;
  assign n10579 = pi16 ? n9726 : n10578;
  assign n10580 = pi21 ? n99 : n1512;
  assign n10581 = pi20 ? n10580 : n32;
  assign n10582 = pi19 ? n10581 : n32;
  assign n10583 = pi18 ? n99 : n10582;
  assign n10584 = pi17 ? n99 : n10583;
  assign n10585 = pi16 ? n801 : n10584;
  assign n10586 = pi15 ? n10579 : n10585;
  assign n10587 = pi21 ? n37 : n383;
  assign n10588 = pi20 ? n37 : n10587;
  assign n10589 = pi21 ? n391 : n316;
  assign n10590 = pi21 ? n3118 : n316;
  assign n10591 = pi20 ? n10589 : n10590;
  assign n10592 = pi19 ? n10588 : n10591;
  assign n10593 = pi18 ? n374 : n10592;
  assign n10594 = pi17 ? n32 : n10593;
  assign n10595 = pi20 ? n3619 : n32;
  assign n10596 = pi19 ? n10595 : n32;
  assign n10597 = pi18 ? n316 : n10596;
  assign n10598 = pi17 ? n316 : n10597;
  assign n10599 = pi16 ? n10594 : n10598;
  assign n10600 = pi20 ? n37 : n413;
  assign n10601 = pi19 ? n37 : n10600;
  assign n10602 = pi18 ? n374 : n10601;
  assign n10603 = pi17 ? n32 : n10602;
  assign n10604 = pi19 ? n4810 : n316;
  assign n10605 = pi18 ? n10604 : n316;
  assign n10606 = pi17 ? n10605 : n10597;
  assign n10607 = pi16 ? n10603 : n10606;
  assign n10608 = pi15 ? n10599 : n10607;
  assign n10609 = pi14 ? n10586 : n10608;
  assign n10610 = pi13 ? n10573 : n10609;
  assign n10611 = pi12 ? n10547 : n10610;
  assign n10612 = pi18 ? n9770 : n3163;
  assign n10613 = pi20 ? n139 : n5961;
  assign n10614 = pi19 ? n10613 : n360;
  assign n10615 = pi21 ? n139 : n2320;
  assign n10616 = pi20 ? n10615 : n32;
  assign n10617 = pi19 ? n10616 : n32;
  assign n10618 = pi18 ? n10614 : n10617;
  assign n10619 = pi17 ? n10612 : n10618;
  assign n10620 = pi16 ? n439 : n10619;
  assign n10621 = pi20 ? n3086 : n942;
  assign n10622 = pi19 ? n10621 : n139;
  assign n10623 = pi20 ? n1778 : n942;
  assign n10624 = pi19 ? n10623 : n139;
  assign n10625 = pi18 ? n10622 : n10624;
  assign n10626 = pi18 ? n10614 : n9777;
  assign n10627 = pi17 ? n10625 : n10626;
  assign n10628 = pi16 ? n439 : n10627;
  assign n10629 = pi15 ? n10620 : n10628;
  assign n10630 = pi20 ? n3086 : n1761;
  assign n10631 = pi19 ? n10630 : n139;
  assign n10632 = pi18 ? n10631 : n139;
  assign n10633 = pi23 ? n139 : n395;
  assign n10634 = pi22 ? n10633 : n32;
  assign n10635 = pi21 ? n139 : n10634;
  assign n10636 = pi20 ? n10635 : n32;
  assign n10637 = pi19 ? n10636 : n32;
  assign n10638 = pi18 ? n139 : n10637;
  assign n10639 = pi17 ? n10632 : n10638;
  assign n10640 = pi16 ? n439 : n10639;
  assign n10641 = pi20 ? n37 : n3090;
  assign n10642 = pi19 ? n10641 : n139;
  assign n10643 = pi18 ? n10642 : n139;
  assign n10644 = pi21 ? n139 : n2565;
  assign n10645 = pi20 ? n10644 : n32;
  assign n10646 = pi19 ? n10645 : n32;
  assign n10647 = pi18 ? n139 : n10646;
  assign n10648 = pi17 ? n10643 : n10647;
  assign n10649 = pi16 ? n439 : n10648;
  assign n10650 = pi15 ? n10640 : n10649;
  assign n10651 = pi14 ? n10629 : n10650;
  assign n10652 = pi19 ? n9765 : n139;
  assign n10653 = pi18 ? n37 : n10652;
  assign n10654 = pi17 ? n10653 : n10647;
  assign n10655 = pi16 ? n439 : n10654;
  assign n10656 = pi17 ? n9816 : n10647;
  assign n10657 = pi16 ? n439 : n10656;
  assign n10658 = pi15 ? n10655 : n10657;
  assign n10659 = pi19 ? n9824 : n9769;
  assign n10660 = pi18 ? n37 : n10659;
  assign n10661 = pi17 ? n10660 : n10647;
  assign n10662 = pi16 ? n439 : n10661;
  assign n10663 = pi22 ? n335 : n455;
  assign n10664 = pi21 ? n37 : n10663;
  assign n10665 = pi20 ? n639 : n10664;
  assign n10666 = pi19 ? n37 : n10665;
  assign n10667 = pi18 ? n37 : n10666;
  assign n10668 = pi20 ? n204 : n4870;
  assign n10669 = pi21 ? n570 : n204;
  assign n10670 = pi20 ? n642 : n10669;
  assign n10671 = pi19 ? n10668 : n10670;
  assign n10672 = pi21 ? n1079 : n2565;
  assign n10673 = pi20 ? n10672 : n32;
  assign n10674 = pi19 ? n10673 : n32;
  assign n10675 = pi18 ? n10671 : n10674;
  assign n10676 = pi17 ? n10667 : n10675;
  assign n10677 = pi16 ? n439 : n10676;
  assign n10678 = pi15 ? n10662 : n10677;
  assign n10679 = pi14 ? n10658 : n10678;
  assign n10680 = pi13 ? n10651 : n10679;
  assign n10681 = pi20 ? n577 : n335;
  assign n10682 = pi19 ? n37 : n10681;
  assign n10683 = pi18 ? n37 : n10682;
  assign n10684 = pi22 ? n335 : n10400;
  assign n10685 = pi21 ? n10684 : n2565;
  assign n10686 = pi20 ? n10685 : n32;
  assign n10687 = pi19 ? n10686 : n32;
  assign n10688 = pi18 ? n335 : n10687;
  assign n10689 = pi17 ? n10683 : n10688;
  assign n10690 = pi16 ? n439 : n10689;
  assign n10691 = pi21 ? n6433 : n2565;
  assign n10692 = pi20 ? n10691 : n32;
  assign n10693 = pi19 ? n10692 : n32;
  assign n10694 = pi18 ? n37 : n10693;
  assign n10695 = pi17 ? n37 : n10694;
  assign n10696 = pi16 ? n439 : n10695;
  assign n10697 = pi15 ? n10690 : n10696;
  assign n10698 = pi21 ? n1313 : n2578;
  assign n10699 = pi20 ? n10698 : n32;
  assign n10700 = pi19 ? n10699 : n32;
  assign n10701 = pi18 ? n37 : n10700;
  assign n10702 = pi17 ? n37 : n10701;
  assign n10703 = pi16 ? n439 : n10702;
  assign n10704 = pi21 ? n6441 : n2578;
  assign n10705 = pi20 ? n10704 : n32;
  assign n10706 = pi19 ? n10705 : n32;
  assign n10707 = pi18 ? n37 : n10706;
  assign n10708 = pi17 ? n37 : n10707;
  assign n10709 = pi16 ? n439 : n10708;
  assign n10710 = pi15 ? n10703 : n10709;
  assign n10711 = pi14 ? n10697 : n10710;
  assign n10712 = pi23 ? n99 : n6960;
  assign n10713 = pi22 ? n37 : n10712;
  assign n10714 = pi21 ? n10713 : n2637;
  assign n10715 = pi20 ? n10714 : n32;
  assign n10716 = pi19 ? n10715 : n32;
  assign n10717 = pi18 ? n37 : n10716;
  assign n10718 = pi17 ? n37 : n10717;
  assign n10719 = pi16 ? n439 : n10718;
  assign n10720 = pi23 ? n139 : n6960;
  assign n10721 = pi22 ? n37 : n10720;
  assign n10722 = pi21 ? n10721 : n5370;
  assign n10723 = pi20 ? n10722 : n32;
  assign n10724 = pi19 ? n10723 : n32;
  assign n10725 = pi18 ? n37 : n10724;
  assign n10726 = pi17 ? n37 : n10725;
  assign n10727 = pi16 ? n439 : n10726;
  assign n10728 = pi15 ? n10719 : n10727;
  assign n10729 = pi24 ? n335 : n685;
  assign n10730 = pi23 ? n335 : n10729;
  assign n10731 = pi22 ? n37 : n10730;
  assign n10732 = pi21 ? n10731 : n1009;
  assign n10733 = pi20 ? n10732 : n32;
  assign n10734 = pi19 ? n10733 : n32;
  assign n10735 = pi18 ? n37 : n10734;
  assign n10736 = pi17 ? n37 : n10735;
  assign n10737 = pi16 ? n439 : n10736;
  assign n10738 = pi22 ? n335 : n10730;
  assign n10739 = pi21 ? n10738 : n1009;
  assign n10740 = pi20 ? n10739 : n32;
  assign n10741 = pi19 ? n10740 : n32;
  assign n10742 = pi18 ? n37 : n10741;
  assign n10743 = pi17 ? n37 : n10742;
  assign n10744 = pi16 ? n439 : n10743;
  assign n10745 = pi15 ? n10737 : n10744;
  assign n10746 = pi14 ? n10728 : n10745;
  assign n10747 = pi13 ? n10711 : n10746;
  assign n10748 = pi12 ? n10680 : n10747;
  assign n10749 = pi11 ? n10611 : n10748;
  assign n10750 = pi24 ? n363 : n316;
  assign n10751 = pi23 ? n363 : n10750;
  assign n10752 = pi22 ? n99 : n10751;
  assign n10753 = pi21 ? n10752 : n32;
  assign n10754 = pi20 ? n10753 : n32;
  assign n10755 = pi19 ? n10754 : n32;
  assign n10756 = pi18 ? n37 : n10755;
  assign n10757 = pi17 ? n37 : n10756;
  assign n10758 = pi16 ? n439 : n10757;
  assign n10759 = pi23 ? n233 : n10750;
  assign n10760 = pi22 ? n363 : n10759;
  assign n10761 = pi21 ? n10760 : n32;
  assign n10762 = pi20 ? n10761 : n32;
  assign n10763 = pi19 ? n10762 : n32;
  assign n10764 = pi18 ? n37 : n10763;
  assign n10765 = pi17 ? n37 : n10764;
  assign n10766 = pi16 ? n439 : n10765;
  assign n10767 = pi15 ? n10758 : n10766;
  assign n10768 = pi23 ? n233 : n1149;
  assign n10769 = pi22 ? n7024 : n10768;
  assign n10770 = pi21 ? n10769 : n32;
  assign n10771 = pi20 ? n10770 : n32;
  assign n10772 = pi19 ? n10771 : n32;
  assign n10773 = pi18 ? n37 : n10772;
  assign n10774 = pi17 ? n37 : n10773;
  assign n10775 = pi16 ? n439 : n10774;
  assign n10776 = pi14 ? n10767 : n10775;
  assign n10777 = pi22 ? n5011 : n730;
  assign n10778 = pi21 ? n10777 : n32;
  assign n10779 = pi20 ? n10778 : n32;
  assign n10780 = pi19 ? n10779 : n32;
  assign n10781 = pi18 ? n37 : n10780;
  assign n10782 = pi17 ? n37 : n10781;
  assign n10783 = pi16 ? n439 : n10782;
  assign n10784 = pi23 ? n685 : n624;
  assign n10785 = pi22 ? n363 : n10784;
  assign n10786 = pi21 ? n10785 : n32;
  assign n10787 = pi20 ? n10786 : n32;
  assign n10788 = pi19 ? n10787 : n32;
  assign n10789 = pi18 ? n37 : n10788;
  assign n10790 = pi17 ? n37 : n10789;
  assign n10791 = pi16 ? n439 : n10790;
  assign n10792 = pi15 ? n10783 : n10791;
  assign n10793 = pi22 ? n3944 : n2192;
  assign n10794 = pi21 ? n10793 : n32;
  assign n10795 = pi20 ? n10794 : n32;
  assign n10796 = pi19 ? n10795 : n32;
  assign n10797 = pi18 ? n37 : n10796;
  assign n10798 = pi17 ? n37 : n10797;
  assign n10799 = pi16 ? n439 : n10798;
  assign n10800 = pi15 ? n10316 : n10799;
  assign n10801 = pi14 ? n10792 : n10800;
  assign n10802 = pi13 ? n10776 : n10801;
  assign n10803 = pi18 ? n9973 : n9959;
  assign n10804 = pi17 ? n99 : n10803;
  assign n10805 = pi16 ? n201 : n10804;
  assign n10806 = pi21 ? n99 : n4538;
  assign n10807 = pi20 ? n99 : n10806;
  assign n10808 = pi19 ? n99 : n10807;
  assign n10809 = pi18 ? n10808 : n10337;
  assign n10810 = pi17 ? n99 : n10809;
  assign n10811 = pi16 ? n744 : n10810;
  assign n10812 = pi15 ? n10805 : n10811;
  assign n10813 = pi18 ? n99 : n9458;
  assign n10814 = pi17 ? n99 : n10813;
  assign n10815 = pi16 ? n721 : n10814;
  assign n10816 = pi16 ? n721 : n10358;
  assign n10817 = pi15 ? n10815 : n10816;
  assign n10818 = pi14 ? n10812 : n10817;
  assign n10819 = pi18 ? n5087 : n10353;
  assign n10820 = pi17 ? n99 : n10819;
  assign n10821 = pi16 ? n721 : n10820;
  assign n10822 = pi18 ? n9992 : n8297;
  assign n10823 = pi17 ? n157 : n10822;
  assign n10824 = pi16 ? n5910 : n10823;
  assign n10825 = pi15 ? n10821 : n10824;
  assign n10826 = pi21 ? n157 : n4237;
  assign n10827 = pi20 ? n99 : n10826;
  assign n10828 = pi19 ? n99 : n10827;
  assign n10829 = pi18 ? n10828 : n4010;
  assign n10830 = pi17 ? n99 : n10829;
  assign n10831 = pi16 ? n744 : n10830;
  assign n10832 = pi15 ? n10824 : n10831;
  assign n10833 = pi14 ? n10825 : n10832;
  assign n10834 = pi13 ? n10818 : n10833;
  assign n10835 = pi12 ? n10802 : n10834;
  assign n10836 = pi21 ? n99 : n4237;
  assign n10837 = pi20 ? n99 : n10836;
  assign n10838 = pi19 ? n99 : n10837;
  assign n10839 = pi18 ? n10838 : n4010;
  assign n10840 = pi17 ? n99 : n10839;
  assign n10841 = pi16 ? n744 : n10840;
  assign n10842 = pi18 ? n10010 : n3212;
  assign n10843 = pi17 ? n99 : n10842;
  assign n10844 = pi16 ? n721 : n10843;
  assign n10845 = pi15 ? n10841 : n10844;
  assign n10846 = pi18 ? n9046 : n10013;
  assign n10847 = pi17 ? n139 : n10846;
  assign n10848 = pi16 ? n915 : n10847;
  assign n10849 = pi20 ? n1026 : n7858;
  assign n10850 = pi19 ? n139 : n10849;
  assign n10851 = pi18 ? n10850 : n10013;
  assign n10852 = pi17 ? n139 : n10851;
  assign n10853 = pi16 ? n2291 : n10852;
  assign n10854 = pi15 ? n10848 : n10853;
  assign n10855 = pi14 ? n10845 : n10854;
  assign n10856 = pi21 ? n963 : n1721;
  assign n10857 = pi20 ? n32 : n10856;
  assign n10858 = pi19 ? n32 : n10857;
  assign n10859 = pi20 ? n1719 : n5269;
  assign n10860 = pi19 ? n2512 : n10859;
  assign n10861 = pi18 ? n10858 : n10860;
  assign n10862 = pi17 ? n32 : n10861;
  assign n10863 = pi20 ? n2527 : n992;
  assign n10864 = pi20 ? n5273 : n992;
  assign n10865 = pi19 ? n10863 : n10864;
  assign n10866 = pi21 ? n1531 : n1698;
  assign n10867 = pi20 ? n139 : n10866;
  assign n10868 = pi20 ? n942 : n2543;
  assign n10869 = pi19 ? n10867 : n10868;
  assign n10870 = pi18 ? n10865 : n10869;
  assign n10871 = pi20 ? n2830 : n2518;
  assign n10872 = pi19 ? n10871 : n10034;
  assign n10873 = pi18 ? n10872 : n10013;
  assign n10874 = pi17 ? n10870 : n10873;
  assign n10875 = pi16 ? n10862 : n10874;
  assign n10876 = pi22 ? n1519 : n316;
  assign n10877 = pi21 ? n10876 : n316;
  assign n10878 = pi20 ? n32 : n10877;
  assign n10879 = pi19 ? n32 : n10878;
  assign n10880 = pi19 ? n316 : n5287;
  assign n10881 = pi18 ? n10879 : n10880;
  assign n10882 = pi17 ? n32 : n10881;
  assign n10883 = pi20 ? n4778 : n316;
  assign n10884 = pi19 ? n10883 : n316;
  assign n10885 = pi18 ? n10884 : n316;
  assign n10886 = pi18 ? n316 : n10013;
  assign n10887 = pi17 ? n10885 : n10886;
  assign n10888 = pi16 ? n10882 : n10887;
  assign n10889 = pi15 ? n10875 : n10888;
  assign n10890 = pi17 ? n316 : n10886;
  assign n10891 = pi16 ? n7883 : n10890;
  assign n10892 = pi20 ? n316 : n5317;
  assign n10893 = pi19 ? n316 : n10892;
  assign n10894 = pi18 ? n5285 : n10893;
  assign n10895 = pi17 ? n32 : n10894;
  assign n10896 = pi17 ? n10885 : n10043;
  assign n10897 = pi16 ? n10895 : n10896;
  assign n10898 = pi15 ? n10891 : n10897;
  assign n10899 = pi14 ? n10889 : n10898;
  assign n10900 = pi13 ? n10855 : n10899;
  assign n10901 = pi21 ? n326 : n316;
  assign n10902 = pi20 ? n32 : n10901;
  assign n10903 = pi19 ? n32 : n10902;
  assign n10904 = pi21 ? n356 : n37;
  assign n10905 = pi20 ? n316 : n10904;
  assign n10906 = pi19 ? n316 : n10905;
  assign n10907 = pi18 ? n10903 : n10906;
  assign n10908 = pi17 ? n32 : n10907;
  assign n10909 = pi19 ? n5288 : n316;
  assign n10910 = pi18 ? n10909 : n316;
  assign n10911 = pi17 ? n10910 : n10043;
  assign n10912 = pi16 ? n10908 : n10911;
  assign n10913 = pi18 ? n10903 : n10070;
  assign n10914 = pi17 ? n32 : n10913;
  assign n10915 = pi17 ? n10074 : n10043;
  assign n10916 = pi16 ? n10914 : n10915;
  assign n10917 = pi15 ? n10912 : n10916;
  assign n10918 = pi21 ? n910 : n1211;
  assign n10919 = pi20 ? n32 : n10918;
  assign n10920 = pi19 ? n32 : n10919;
  assign n10921 = pi21 ? n9146 : n9143;
  assign n10922 = pi21 ? n9144 : n297;
  assign n10923 = pi20 ? n10921 : n10922;
  assign n10924 = pi19 ? n2521 : n10923;
  assign n10925 = pi18 ? n10920 : n10924;
  assign n10926 = pi17 ? n32 : n10925;
  assign n10927 = pi21 ? n9144 : n9122;
  assign n10928 = pi21 ? n139 : n9122;
  assign n10929 = pi20 ? n10927 : n10928;
  assign n10930 = pi22 ? n9123 : n139;
  assign n10931 = pi21 ? n10930 : n139;
  assign n10932 = pi21 ? n1721 : n9143;
  assign n10933 = pi20 ? n10931 : n10932;
  assign n10934 = pi19 ? n10929 : n10933;
  assign n10935 = pi20 ? n9126 : n9143;
  assign n10936 = pi21 ? n9122 : n10930;
  assign n10937 = pi20 ? n10927 : n10936;
  assign n10938 = pi19 ? n10935 : n10937;
  assign n10939 = pi18 ? n10934 : n10938;
  assign n10940 = pi21 ? n1531 : n9144;
  assign n10941 = pi20 ? n10940 : n10936;
  assign n10942 = pi21 ? n3188 : n316;
  assign n10943 = pi20 ? n10940 : n10942;
  assign n10944 = pi19 ? n10941 : n10943;
  assign n10945 = pi18 ? n10944 : n2655;
  assign n10946 = pi17 ? n10939 : n10945;
  assign n10947 = pi16 ? n10926 : n10946;
  assign n10948 = pi22 ? n448 : n685;
  assign n10949 = pi21 ? n1079 : n10948;
  assign n10950 = pi20 ? n335 : n10949;
  assign n10951 = pi19 ? n335 : n10950;
  assign n10952 = pi18 ? n10951 : n1824;
  assign n10953 = pi17 ? n335 : n10952;
  assign n10954 = pi16 ? n2035 : n10953;
  assign n10955 = pi15 ? n10947 : n10954;
  assign n10956 = pi14 ? n10917 : n10955;
  assign n10957 = pi20 ? n335 : n647;
  assign n10958 = pi19 ? n335 : n10957;
  assign n10959 = pi18 ? n7941 : n10958;
  assign n10960 = pi17 ? n32 : n10959;
  assign n10961 = pi21 ? n335 : n1071;
  assign n10962 = pi20 ? n335 : n10961;
  assign n10963 = pi19 ? n335 : n10962;
  assign n10964 = pi18 ? n10963 : n32;
  assign n10965 = pi17 ? n335 : n10964;
  assign n10966 = pi16 ? n10960 : n10965;
  assign n10967 = pi22 ? n3935 : n2192;
  assign n10968 = pi21 ? n335 : n10967;
  assign n10969 = pi20 ? n335 : n10968;
  assign n10970 = pi19 ? n335 : n10969;
  assign n10971 = pi18 ? n10970 : n32;
  assign n10972 = pi17 ? n335 : n10971;
  assign n10973 = pi16 ? n7943 : n10972;
  assign n10974 = pi15 ? n10966 : n10973;
  assign n10975 = pi22 ? n5996 : n335;
  assign n10976 = pi21 ? n10975 : n335;
  assign n10977 = pi20 ? n32 : n10976;
  assign n10978 = pi19 ? n32 : n10977;
  assign n10979 = pi18 ? n10978 : n335;
  assign n10980 = pi17 ? n32 : n10979;
  assign n10981 = pi22 ? n233 : n2192;
  assign n10982 = pi21 ? n335 : n10981;
  assign n10983 = pi20 ? n335 : n10982;
  assign n10984 = pi19 ? n335 : n10983;
  assign n10985 = pi18 ? n10984 : n32;
  assign n10986 = pi17 ? n335 : n10985;
  assign n10987 = pi16 ? n10980 : n10986;
  assign n10988 = pi16 ? n10980 : n10130;
  assign n10989 = pi15 ? n10987 : n10988;
  assign n10990 = pi14 ? n10974 : n10989;
  assign n10991 = pi13 ? n10956 : n10990;
  assign n10992 = pi12 ? n10900 : n10991;
  assign n10993 = pi11 ? n10835 : n10992;
  assign n10994 = pi10 ? n10749 : n10993;
  assign n10995 = pi09 ? n10446 : n10994;
  assign n10996 = pi15 ? n32 : n10439;
  assign n10997 = pi16 ? n1130 : n10436;
  assign n10998 = pi15 ? n10440 : n10997;
  assign n10999 = pi14 ? n10996 : n10998;
  assign n11000 = pi13 ? n32 : n10999;
  assign n11001 = pi12 ? n32 : n11000;
  assign n11002 = pi11 ? n32 : n11001;
  assign n11003 = pi10 ? n32 : n11002;
  assign n11004 = pi16 ? n9232 : n10451;
  assign n11005 = pi16 ? n2461 : n10458;
  assign n11006 = pi15 ? n11004 : n11005;
  assign n11007 = pi21 ? n32 : n37;
  assign n11008 = pi20 ? n32 : n11007;
  assign n11009 = pi19 ? n32 : n11008;
  assign n11010 = pi18 ? n11009 : n37;
  assign n11011 = pi17 ? n32 : n11010;
  assign n11012 = pi16 ? n11011 : n10476;
  assign n11013 = pi15 ? n10468 : n11012;
  assign n11014 = pi14 ? n11006 : n11013;
  assign n11015 = pi22 ? n363 : n32;
  assign n11016 = pi21 ? n5012 : n11015;
  assign n11017 = pi20 ? n11016 : n32;
  assign n11018 = pi19 ? n11017 : n32;
  assign n11019 = pi18 ? n10505 : n11018;
  assign n11020 = pi17 ? n10500 : n11019;
  assign n11021 = pi16 ? n10485 : n11020;
  assign n11022 = pi15 ? n10477 : n11021;
  assign n11023 = pi16 ? n744 : n10516;
  assign n11024 = pi18 ? n742 : n10522;
  assign n11025 = pi17 ? n32 : n11024;
  assign n11026 = pi22 ? n157 : n32;
  assign n11027 = pi21 ? n168 : n11026;
  assign n11028 = pi20 ? n11027 : n32;
  assign n11029 = pi19 ? n11028 : n32;
  assign n11030 = pi18 ? n10541 : n11029;
  assign n11031 = pi17 ? n10537 : n11030;
  assign n11032 = pi16 ? n11025 : n11031;
  assign n11033 = pi15 ? n11023 : n11032;
  assign n11034 = pi14 ? n11022 : n11033;
  assign n11035 = pi13 ? n11014 : n11034;
  assign n11036 = pi18 ? n10555 : n11029;
  assign n11037 = pi17 ? n10553 : n11036;
  assign n11038 = pi16 ? n801 : n11037;
  assign n11039 = pi21 ? n99 : n3962;
  assign n11040 = pi20 ? n11039 : n32;
  assign n11041 = pi19 ? n11040 : n32;
  assign n11042 = pi18 ? n99 : n11041;
  assign n11043 = pi17 ? n99 : n11042;
  assign n11044 = pi16 ? n10560 : n11043;
  assign n11045 = pi15 ? n11038 : n11044;
  assign n11046 = pi16 ? n721 : n11043;
  assign n11047 = pi23 ? n99 : n233;
  assign n11048 = pi22 ? n11047 : n32;
  assign n11049 = pi21 ? n99 : n11048;
  assign n11050 = pi20 ? n11049 : n32;
  assign n11051 = pi19 ? n11050 : n32;
  assign n11052 = pi18 ? n99 : n11051;
  assign n11053 = pi17 ? n99 : n11052;
  assign n11054 = pi16 ? n9726 : n11053;
  assign n11055 = pi15 ? n11046 : n11054;
  assign n11056 = pi14 ? n11045 : n11055;
  assign n11057 = pi22 ? n1457 : n32;
  assign n11058 = pi21 ? n99 : n11057;
  assign n11059 = pi20 ? n11058 : n32;
  assign n11060 = pi19 ? n11059 : n32;
  assign n11061 = pi18 ? n99 : n11060;
  assign n11062 = pi17 ? n99 : n11061;
  assign n11063 = pi16 ? n9726 : n11062;
  assign n11064 = pi21 ? n99 : n2256;
  assign n11065 = pi20 ? n11064 : n32;
  assign n11066 = pi19 ? n11065 : n32;
  assign n11067 = pi18 ? n99 : n11066;
  assign n11068 = pi17 ? n99 : n11067;
  assign n11069 = pi16 ? n801 : n11068;
  assign n11070 = pi15 ? n11063 : n11069;
  assign n11071 = pi21 ? n37 : n428;
  assign n11072 = pi20 ? n37 : n11071;
  assign n11073 = pi21 ? n37 : n424;
  assign n11074 = pi20 ? n11073 : n5689;
  assign n11075 = pi19 ? n11072 : n11074;
  assign n11076 = pi18 ? n374 : n11075;
  assign n11077 = pi17 ? n32 : n11076;
  assign n11078 = pi16 ? n11077 : n10598;
  assign n11079 = pi15 ? n11078 : n10607;
  assign n11080 = pi14 ? n11070 : n11079;
  assign n11081 = pi13 ? n11056 : n11080;
  assign n11082 = pi12 ? n11035 : n11081;
  assign n11083 = pi22 ? n1784 : n32;
  assign n11084 = pi21 ? n139 : n11083;
  assign n11085 = pi20 ? n11084 : n32;
  assign n11086 = pi19 ? n11085 : n32;
  assign n11087 = pi18 ? n10614 : n11086;
  assign n11088 = pi17 ? n10612 : n11087;
  assign n11089 = pi16 ? n439 : n11088;
  assign n11090 = pi18 ? n10614 : n10637;
  assign n11091 = pi17 ? n10625 : n11090;
  assign n11092 = pi16 ? n439 : n11091;
  assign n11093 = pi15 ? n11089 : n11092;
  assign n11094 = pi21 ? n139 : n5003;
  assign n11095 = pi20 ? n11094 : n32;
  assign n11096 = pi19 ? n11095 : n32;
  assign n11097 = pi18 ? n139 : n11096;
  assign n11098 = pi17 ? n10632 : n11097;
  assign n11099 = pi16 ? n439 : n11098;
  assign n11100 = pi21 ? n139 : n3066;
  assign n11101 = pi20 ? n11100 : n32;
  assign n11102 = pi19 ? n11101 : n32;
  assign n11103 = pi18 ? n139 : n11102;
  assign n11104 = pi17 ? n10643 : n11103;
  assign n11105 = pi16 ? n439 : n11104;
  assign n11106 = pi15 ? n11099 : n11105;
  assign n11107 = pi14 ? n11093 : n11106;
  assign n11108 = pi13 ? n11107 : n10679;
  assign n11109 = pi23 ? n335 : n1432;
  assign n11110 = pi22 ? n335 : n11109;
  assign n11111 = pi21 ? n11110 : n2565;
  assign n11112 = pi20 ? n11111 : n32;
  assign n11113 = pi19 ? n11112 : n32;
  assign n11114 = pi18 ? n335 : n11113;
  assign n11115 = pi17 ? n10683 : n11114;
  assign n11116 = pi16 ? n439 : n11115;
  assign n11117 = pi24 ? n37 : n204;
  assign n11118 = pi23 ? n37 : n11117;
  assign n11119 = pi22 ? n37 : n11118;
  assign n11120 = pi21 ? n11119 : n2565;
  assign n11121 = pi20 ? n11120 : n32;
  assign n11122 = pi19 ? n11121 : n32;
  assign n11123 = pi18 ? n37 : n11122;
  assign n11124 = pi17 ? n37 : n11123;
  assign n11125 = pi16 ? n439 : n11124;
  assign n11126 = pi15 ? n11116 : n11125;
  assign n11127 = pi24 ? n37 : n233;
  assign n11128 = pi23 ? n37 : n11127;
  assign n11129 = pi22 ? n37 : n11128;
  assign n11130 = pi21 ? n11129 : n2578;
  assign n11131 = pi20 ? n11130 : n32;
  assign n11132 = pi19 ? n11131 : n32;
  assign n11133 = pi18 ? n37 : n11132;
  assign n11134 = pi17 ? n37 : n11133;
  assign n11135 = pi16 ? n439 : n11134;
  assign n11136 = pi23 ? n99 : n234;
  assign n11137 = pi22 ? n37 : n11136;
  assign n11138 = pi21 ? n11137 : n2578;
  assign n11139 = pi20 ? n11138 : n32;
  assign n11140 = pi19 ? n11139 : n32;
  assign n11141 = pi18 ? n37 : n11140;
  assign n11142 = pi17 ? n37 : n11141;
  assign n11143 = pi16 ? n439 : n11142;
  assign n11144 = pi15 ? n11135 : n11143;
  assign n11145 = pi14 ? n11126 : n11144;
  assign n11146 = pi22 ? n37 : n11047;
  assign n11147 = pi21 ? n11146 : n2637;
  assign n11148 = pi20 ? n11147 : n32;
  assign n11149 = pi19 ? n11148 : n32;
  assign n11150 = pi18 ? n37 : n11149;
  assign n11151 = pi17 ? n37 : n11150;
  assign n11152 = pi16 ? n439 : n11151;
  assign n11153 = pi22 ? n37 : n6833;
  assign n11154 = pi21 ? n11153 : n2678;
  assign n11155 = pi20 ? n11154 : n32;
  assign n11156 = pi19 ? n11155 : n32;
  assign n11157 = pi18 ? n37 : n11156;
  assign n11158 = pi17 ? n37 : n11157;
  assign n11159 = pi16 ? n439 : n11158;
  assign n11160 = pi15 ? n11152 : n11159;
  assign n11161 = pi21 ? n2074 : n2700;
  assign n11162 = pi20 ? n11161 : n32;
  assign n11163 = pi19 ? n11162 : n32;
  assign n11164 = pi18 ? n37 : n11163;
  assign n11165 = pi17 ? n37 : n11164;
  assign n11166 = pi16 ? n439 : n11165;
  assign n11167 = pi21 ? n2061 : n928;
  assign n11168 = pi20 ? n11167 : n32;
  assign n11169 = pi19 ? n11168 : n32;
  assign n11170 = pi18 ? n37 : n11169;
  assign n11171 = pi17 ? n37 : n11170;
  assign n11172 = pi16 ? n439 : n11171;
  assign n11173 = pi15 ? n11166 : n11172;
  assign n11174 = pi14 ? n11160 : n11173;
  assign n11175 = pi13 ? n11145 : n11174;
  assign n11176 = pi12 ? n11108 : n11175;
  assign n11177 = pi11 ? n11082 : n11176;
  assign n11178 = pi22 ? n99 : n673;
  assign n11179 = pi21 ? n11178 : n1009;
  assign n11180 = pi20 ? n11179 : n32;
  assign n11181 = pi19 ? n11180 : n32;
  assign n11182 = pi18 ? n37 : n11181;
  assign n11183 = pi17 ? n37 : n11182;
  assign n11184 = pi16 ? n439 : n11183;
  assign n11185 = pi21 ? n2707 : n1009;
  assign n11186 = pi20 ? n11185 : n32;
  assign n11187 = pi19 ? n11186 : n32;
  assign n11188 = pi18 ? n37 : n11187;
  assign n11189 = pi17 ? n37 : n11188;
  assign n11190 = pi16 ? n439 : n11189;
  assign n11191 = pi15 ? n11184 : n11190;
  assign n11192 = pi22 ? n295 : n233;
  assign n11193 = pi21 ? n11192 : n32;
  assign n11194 = pi20 ? n11193 : n32;
  assign n11195 = pi19 ? n11194 : n32;
  assign n11196 = pi18 ? n37 : n11195;
  assign n11197 = pi17 ? n37 : n11196;
  assign n11198 = pi16 ? n439 : n11197;
  assign n11199 = pi22 ? n583 : n233;
  assign n11200 = pi21 ? n11199 : n32;
  assign n11201 = pi20 ? n11200 : n32;
  assign n11202 = pi19 ? n11201 : n32;
  assign n11203 = pi18 ? n37 : n11202;
  assign n11204 = pi17 ? n37 : n11203;
  assign n11205 = pi16 ? n439 : n11204;
  assign n11206 = pi15 ? n11198 : n11205;
  assign n11207 = pi14 ? n11191 : n11206;
  assign n11208 = pi22 ? n5011 : n685;
  assign n11209 = pi21 ? n11208 : n32;
  assign n11210 = pi20 ? n11209 : n32;
  assign n11211 = pi19 ? n11210 : n32;
  assign n11212 = pi18 ? n37 : n11211;
  assign n11213 = pi17 ? n37 : n11212;
  assign n11214 = pi16 ? n439 : n11213;
  assign n11215 = pi21 ? n2721 : n32;
  assign n11216 = pi20 ? n11215 : n32;
  assign n11217 = pi19 ? n11216 : n32;
  assign n11218 = pi18 ? n37 : n11217;
  assign n11219 = pi17 ? n37 : n11218;
  assign n11220 = pi16 ? n439 : n11219;
  assign n11221 = pi15 ? n11214 : n11220;
  assign n11222 = pi22 ? n3944 : n1475;
  assign n11223 = pi21 ? n11222 : n32;
  assign n11224 = pi20 ? n11223 : n32;
  assign n11225 = pi19 ? n11224 : n32;
  assign n11226 = pi18 ? n37 : n11225;
  assign n11227 = pi17 ? n37 : n11226;
  assign n11228 = pi16 ? n439 : n11227;
  assign n11229 = pi15 ? n11220 : n11228;
  assign n11230 = pi14 ? n11221 : n11229;
  assign n11231 = pi13 ? n11207 : n11230;
  assign n11232 = pi18 ? n9973 : n10321;
  assign n11233 = pi17 ? n99 : n11232;
  assign n11234 = pi16 ? n201 : n11233;
  assign n11235 = pi22 ? n204 : n759;
  assign n11236 = pi21 ? n11235 : n32;
  assign n11237 = pi20 ? n11236 : n32;
  assign n11238 = pi19 ? n11237 : n32;
  assign n11239 = pi18 ? n99 : n11238;
  assign n11240 = pi17 ? n99 : n11239;
  assign n11241 = pi16 ? n744 : n11240;
  assign n11242 = pi15 ? n11234 : n11241;
  assign n11243 = pi21 ? n2200 : n32;
  assign n11244 = pi20 ? n11243 : n32;
  assign n11245 = pi19 ? n11244 : n32;
  assign n11246 = pi18 ? n99 : n11245;
  assign n11247 = pi17 ? n99 : n11246;
  assign n11248 = pi16 ? n744 : n11247;
  assign n11249 = pi18 ? n9985 : n10328;
  assign n11250 = pi17 ? n99 : n11249;
  assign n11251 = pi16 ? n744 : n11250;
  assign n11252 = pi15 ? n11248 : n11251;
  assign n11253 = pi14 ? n11242 : n11252;
  assign n11254 = pi18 ? n5087 : n9458;
  assign n11255 = pi17 ? n99 : n11254;
  assign n11256 = pi16 ? n744 : n11255;
  assign n11257 = pi18 ? n9992 : n9965;
  assign n11258 = pi17 ? n157 : n11257;
  assign n11259 = pi16 ? n7793 : n11258;
  assign n11260 = pi15 ? n11256 : n11259;
  assign n11261 = pi15 ? n11259 : n10831;
  assign n11262 = pi14 ? n11260 : n11261;
  assign n11263 = pi13 ? n11253 : n11262;
  assign n11264 = pi12 ? n11231 : n11263;
  assign n11265 = pi16 ? n744 : n10843;
  assign n11266 = pi15 ? n10841 : n11265;
  assign n11267 = pi19 ? n139 : n7839;
  assign n11268 = pi18 ? n11267 : n10013;
  assign n11269 = pi17 ? n139 : n11268;
  assign n11270 = pi16 ? n915 : n11269;
  assign n11271 = pi16 ? n915 : n10852;
  assign n11272 = pi15 ? n11270 : n11271;
  assign n11273 = pi14 ? n11266 : n11272;
  assign n11274 = pi21 ? n910 : n359;
  assign n11275 = pi20 ? n32 : n11274;
  assign n11276 = pi19 ? n32 : n11275;
  assign n11277 = pi21 ? n139 : n359;
  assign n11278 = pi21 ? n4419 : n349;
  assign n11279 = pi20 ? n350 : n11278;
  assign n11280 = pi19 ? n11277 : n11279;
  assign n11281 = pi18 ? n11276 : n11280;
  assign n11282 = pi17 ? n32 : n11281;
  assign n11283 = pi20 ? n8719 : n1775;
  assign n11284 = pi20 ? n6919 : n5969;
  assign n11285 = pi19 ? n11283 : n11284;
  assign n11286 = pi21 ? n4014 : n4052;
  assign n11287 = pi20 ? n356 : n11286;
  assign n11288 = pi21 ? n3118 : n3617;
  assign n11289 = pi20 ? n11278 : n11288;
  assign n11290 = pi19 ? n11287 : n11289;
  assign n11291 = pi18 ? n11285 : n11290;
  assign n11292 = pi21 ? n1774 : n3617;
  assign n11293 = pi20 ? n8423 : n11292;
  assign n11294 = pi21 ? n1785 : n1027;
  assign n11295 = pi20 ? n8423 : n11294;
  assign n11296 = pi19 ? n11293 : n11295;
  assign n11297 = pi18 ? n11296 : n10013;
  assign n11298 = pi17 ? n11291 : n11297;
  assign n11299 = pi16 ? n11282 : n11298;
  assign n11300 = pi18 ? n9093 : n10880;
  assign n11301 = pi17 ? n32 : n11300;
  assign n11302 = pi16 ? n11301 : n10887;
  assign n11303 = pi15 ? n11299 : n11302;
  assign n11304 = pi14 ? n11303 : n10898;
  assign n11305 = pi13 ? n11273 : n11304;
  assign n11306 = pi22 ? n566 : n139;
  assign n11307 = pi21 ? n910 : n11306;
  assign n11308 = pi20 ? n32 : n11307;
  assign n11309 = pi19 ? n32 : n11308;
  assign n11310 = pi21 ? n139 : n11306;
  assign n11311 = pi21 ? n4990 : n9143;
  assign n11312 = pi20 ? n11311 : n10922;
  assign n11313 = pi19 ? n11310 : n11312;
  assign n11314 = pi18 ? n11309 : n11313;
  assign n11315 = pi17 ? n32 : n11314;
  assign n11316 = pi21 ? n10930 : n9144;
  assign n11317 = pi22 ? n583 : n139;
  assign n11318 = pi21 ? n11317 : n9126;
  assign n11319 = pi20 ? n11316 : n11318;
  assign n11320 = pi19 ? n10929 : n11319;
  assign n11321 = pi21 ? n9126 : n9143;
  assign n11322 = pi20 ? n9126 : n11321;
  assign n11323 = pi21 ? n9144 : n9138;
  assign n11324 = pi20 ? n11323 : n9122;
  assign n11325 = pi19 ? n11322 : n11324;
  assign n11326 = pi18 ? n11320 : n11325;
  assign n11327 = pi22 ? n9123 : n583;
  assign n11328 = pi21 ? n11327 : n9144;
  assign n11329 = pi20 ? n11328 : n9122;
  assign n11330 = pi21 ? n11327 : n9133;
  assign n11331 = pi20 ? n11330 : n10942;
  assign n11332 = pi19 ? n11329 : n11331;
  assign n11333 = pi18 ? n11332 : n2655;
  assign n11334 = pi17 ? n11326 : n11333;
  assign n11335 = pi16 ? n11315 : n11334;
  assign n11336 = pi22 ? n335 : n685;
  assign n11337 = pi21 ? n1079 : n11336;
  assign n11338 = pi20 ? n335 : n11337;
  assign n11339 = pi19 ? n335 : n11338;
  assign n11340 = pi18 ? n11339 : n1824;
  assign n11341 = pi17 ? n335 : n11340;
  assign n11342 = pi16 ? n2035 : n11341;
  assign n11343 = pi15 ? n11335 : n11342;
  assign n11344 = pi14 ? n10917 : n11343;
  assign n11345 = pi18 ? n10963 : n1824;
  assign n11346 = pi17 ? n335 : n11345;
  assign n11347 = pi16 ? n10960 : n11346;
  assign n11348 = pi22 ? n10400 : n2192;
  assign n11349 = pi21 ? n335 : n11348;
  assign n11350 = pi20 ? n335 : n11349;
  assign n11351 = pi19 ? n335 : n11350;
  assign n11352 = pi18 ? n11351 : n32;
  assign n11353 = pi17 ? n335 : n11352;
  assign n11354 = pi16 ? n7943 : n11353;
  assign n11355 = pi15 ? n11347 : n11354;
  assign n11356 = pi14 ? n11355 : n10989;
  assign n11357 = pi13 ? n11344 : n11356;
  assign n11358 = pi12 ? n11305 : n11357;
  assign n11359 = pi11 ? n11264 : n11358;
  assign n11360 = pi10 ? n11177 : n11359;
  assign n11361 = pi09 ? n11003 : n11360;
  assign n11362 = pi08 ? n10995 : n11361;
  assign n11363 = pi07 ? n10431 : n11362;
  assign n11364 = pi06 ? n9606 : n11363;
  assign n11365 = pi20 ? n49 : n32;
  assign n11366 = pi19 ? n11365 : n32;
  assign n11367 = pi18 ? n37 : n11366;
  assign n11368 = pi17 ? n37 : n11367;
  assign n11369 = pi16 ? n83 : n11368;
  assign n11370 = pi15 ? n32 : n11369;
  assign n11371 = pi16 ? n8027 : n11368;
  assign n11372 = pi16 ? n1130 : n11368;
  assign n11373 = pi15 ? n11371 : n11372;
  assign n11374 = pi14 ? n11370 : n11373;
  assign n11375 = pi13 ? n32 : n11374;
  assign n11376 = pi12 ? n32 : n11375;
  assign n11377 = pi11 ? n32 : n11376;
  assign n11378 = pi10 ? n32 : n11377;
  assign n11379 = pi21 ? n37 : n104;
  assign n11380 = pi20 ? n11379 : n32;
  assign n11381 = pi19 ? n11380 : n32;
  assign n11382 = pi18 ? n37 : n11381;
  assign n11383 = pi17 ? n37 : n11382;
  assign n11384 = pi16 ? n9232 : n11383;
  assign n11385 = pi21 ? n37 : n303;
  assign n11386 = pi20 ? n11385 : n32;
  assign n11387 = pi19 ? n11386 : n32;
  assign n11388 = pi18 ? n37 : n11387;
  assign n11389 = pi17 ? n37 : n11388;
  assign n11390 = pi16 ? n2461 : n11389;
  assign n11391 = pi15 ? n11384 : n11390;
  assign n11392 = pi16 ? n10154 : n10458;
  assign n11393 = pi22 ? n335 : n32;
  assign n11394 = pi21 ? n37 : n11393;
  assign n11395 = pi20 ? n11394 : n32;
  assign n11396 = pi19 ? n11395 : n32;
  assign n11397 = pi18 ? n37 : n11396;
  assign n11398 = pi17 ? n37 : n11397;
  assign n11399 = pi16 ? n11011 : n11398;
  assign n11400 = pi15 ? n11392 : n11399;
  assign n11401 = pi14 ? n11391 : n11400;
  assign n11402 = pi22 ? n583 : n32;
  assign n11403 = pi21 ? n37 : n11402;
  assign n11404 = pi20 ? n11403 : n32;
  assign n11405 = pi19 ? n11404 : n32;
  assign n11406 = pi18 ? n37 : n11405;
  assign n11407 = pi17 ? n37 : n11406;
  assign n11408 = pi16 ? n439 : n11407;
  assign n11409 = pi21 ? n180 : n2175;
  assign n11410 = pi20 ? n32 : n11409;
  assign n11411 = pi19 ? n32 : n11410;
  assign n11412 = pi19 ? n2185 : n2963;
  assign n11413 = pi18 ? n11411 : n11412;
  assign n11414 = pi17 ? n32 : n11413;
  assign n11415 = pi21 ? n218 : n2175;
  assign n11416 = pi20 ? n11415 : n2185;
  assign n11417 = pi19 ? n2969 : n11416;
  assign n11418 = pi21 ? n218 : n2160;
  assign n11419 = pi20 ? n2185 : n11418;
  assign n11420 = pi21 ? n181 : n2175;
  assign n11421 = pi20 ? n2185 : n11420;
  assign n11422 = pi19 ? n11419 : n11421;
  assign n11423 = pi18 ? n11417 : n11422;
  assign n11424 = pi21 ? n218 : n2161;
  assign n11425 = pi20 ? n11420 : n11424;
  assign n11426 = pi19 ? n11425 : n2967;
  assign n11427 = pi22 ? n5011 : n32;
  assign n11428 = pi21 ? n2175 : n11427;
  assign n11429 = pi20 ? n11428 : n32;
  assign n11430 = pi19 ? n11429 : n32;
  assign n11431 = pi18 ? n11426 : n11430;
  assign n11432 = pi17 ? n11423 : n11431;
  assign n11433 = pi16 ? n11414 : n11432;
  assign n11434 = pi15 ? n11408 : n11433;
  assign n11435 = pi22 ? n4537 : n32;
  assign n11436 = pi21 ? n99 : n11435;
  assign n11437 = pi20 ? n11436 : n32;
  assign n11438 = pi19 ? n11437 : n32;
  assign n11439 = pi18 ? n99 : n11438;
  assign n11440 = pi17 ? n99 : n11439;
  assign n11441 = pi16 ? n801 : n11440;
  assign n11442 = pi21 ? n796 : n159;
  assign n11443 = pi20 ? n32 : n11442;
  assign n11444 = pi19 ? n32 : n11443;
  assign n11445 = pi20 ? n2238 : n157;
  assign n11446 = pi19 ? n11445 : n157;
  assign n11447 = pi18 ? n11444 : n11446;
  assign n11448 = pi17 ? n32 : n11447;
  assign n11449 = pi21 ? n157 : n11026;
  assign n11450 = pi20 ? n11449 : n32;
  assign n11451 = pi19 ? n11450 : n32;
  assign n11452 = pi18 ? n157 : n11451;
  assign n11453 = pi17 ? n157 : n11452;
  assign n11454 = pi16 ? n11448 : n11453;
  assign n11455 = pi15 ? n11441 : n11454;
  assign n11456 = pi14 ? n11434 : n11455;
  assign n11457 = pi13 ? n11401 : n11456;
  assign n11458 = pi22 ? n7377 : n32;
  assign n11459 = pi21 ? n99 : n11458;
  assign n11460 = pi20 ? n11459 : n32;
  assign n11461 = pi19 ? n11460 : n32;
  assign n11462 = pi18 ? n99 : n11461;
  assign n11463 = pi17 ? n99 : n11462;
  assign n11464 = pi16 ? n744 : n11463;
  assign n11465 = pi22 ? n1682 : n32;
  assign n11466 = pi21 ? n99 : n11465;
  assign n11467 = pi20 ? n11466 : n32;
  assign n11468 = pi19 ? n11467 : n32;
  assign n11469 = pi18 ? n99 : n11468;
  assign n11470 = pi17 ? n99 : n11469;
  assign n11471 = pi16 ? n801 : n11470;
  assign n11472 = pi15 ? n11464 : n11471;
  assign n11473 = pi16 ? n801 : n11043;
  assign n11474 = pi21 ? n796 : n775;
  assign n11475 = pi20 ? n32 : n11474;
  assign n11476 = pi19 ? n32 : n11475;
  assign n11477 = pi18 ? n11476 : n99;
  assign n11478 = pi17 ? n32 : n11477;
  assign n11479 = pi16 ? n11478 : n11053;
  assign n11480 = pi15 ? n11473 : n11479;
  assign n11481 = pi14 ? n11472 : n11480;
  assign n11482 = pi21 ? n796 : n2998;
  assign n11483 = pi20 ? n32 : n11482;
  assign n11484 = pi19 ? n32 : n11483;
  assign n11485 = pi18 ? n11484 : n99;
  assign n11486 = pi17 ? n32 : n11485;
  assign n11487 = pi16 ? n11486 : n11053;
  assign n11488 = pi22 ? n3443 : n32;
  assign n11489 = pi21 ? n99 : n11488;
  assign n11490 = pi20 ? n11489 : n32;
  assign n11491 = pi19 ? n11490 : n32;
  assign n11492 = pi18 ? n99 : n11491;
  assign n11493 = pi17 ? n99 : n11492;
  assign n11494 = pi16 ? n744 : n11493;
  assign n11495 = pi15 ? n11487 : n11494;
  assign n11496 = pi20 ? n5696 : n7571;
  assign n11497 = pi19 ? n11496 : n316;
  assign n11498 = pi18 ? n11497 : n316;
  assign n11499 = pi20 ? n5245 : n32;
  assign n11500 = pi19 ? n11499 : n32;
  assign n11501 = pi18 ? n316 : n11500;
  assign n11502 = pi17 ? n11498 : n11501;
  assign n11503 = pi16 ? n439 : n11502;
  assign n11504 = pi20 ? n37 : n393;
  assign n11505 = pi20 ? n10589 : n3702;
  assign n11506 = pi19 ? n11504 : n11505;
  assign n11507 = pi21 ? n391 : n381;
  assign n11508 = pi20 ? n316 : n11507;
  assign n11509 = pi20 ? n3702 : n316;
  assign n11510 = pi19 ? n11508 : n11509;
  assign n11511 = pi18 ? n11506 : n11510;
  assign n11512 = pi19 ? n316 : n7571;
  assign n11513 = pi18 ? n11512 : n11500;
  assign n11514 = pi17 ? n11511 : n11513;
  assign n11515 = pi16 ? n439 : n11514;
  assign n11516 = pi15 ? n11503 : n11515;
  assign n11517 = pi14 ? n11495 : n11516;
  assign n11518 = pi13 ? n11481 : n11517;
  assign n11519 = pi12 ? n11457 : n11518;
  assign n11520 = pi20 ? n5707 : n11073;
  assign n11521 = pi19 ? n37 : n11520;
  assign n11522 = pi21 ? n139 : n424;
  assign n11523 = pi20 ? n11522 : n37;
  assign n11524 = pi20 ? n382 : n3232;
  assign n11525 = pi19 ? n11523 : n11524;
  assign n11526 = pi18 ? n11521 : n11525;
  assign n11527 = pi21 ? n3617 : n316;
  assign n11528 = pi21 ? n1774 : n3258;
  assign n11529 = pi20 ? n11527 : n11528;
  assign n11530 = pi21 ? n359 : n3258;
  assign n11531 = pi21 ? n424 : n4017;
  assign n11532 = pi20 ? n11530 : n11531;
  assign n11533 = pi19 ? n11529 : n11532;
  assign n11534 = pi22 ? n1784 : n706;
  assign n11535 = pi21 ? n316 : n11534;
  assign n11536 = pi20 ? n11535 : n32;
  assign n11537 = pi19 ? n11536 : n32;
  assign n11538 = pi18 ? n11533 : n11537;
  assign n11539 = pi17 ? n11526 : n11538;
  assign n11540 = pi16 ? n439 : n11539;
  assign n11541 = pi20 ? n4839 : n37;
  assign n11542 = pi20 ? n37 : n5696;
  assign n11543 = pi19 ? n11541 : n11542;
  assign n11544 = pi21 ? n424 : n11083;
  assign n11545 = pi20 ? n11544 : n32;
  assign n11546 = pi19 ? n11545 : n32;
  assign n11547 = pi18 ? n11543 : n11546;
  assign n11548 = pi17 ? n37 : n11547;
  assign n11549 = pi16 ? n439 : n11548;
  assign n11550 = pi15 ? n11540 : n11549;
  assign n11551 = pi19 ? n37 : n3096;
  assign n11552 = pi19 ? n139 : n8765;
  assign n11553 = pi18 ? n11551 : n11552;
  assign n11554 = pi18 ? n139 : n11086;
  assign n11555 = pi17 ? n11553 : n11554;
  assign n11556 = pi16 ? n439 : n11555;
  assign n11557 = pi19 ? n1806 : n8765;
  assign n11558 = pi18 ? n11551 : n11557;
  assign n11559 = pi21 ? n139 : n3156;
  assign n11560 = pi20 ? n11559 : n32;
  assign n11561 = pi19 ? n11560 : n32;
  assign n11562 = pi18 ? n139 : n11561;
  assign n11563 = pi17 ? n11558 : n11562;
  assign n11564 = pi16 ? n439 : n11563;
  assign n11565 = pi15 ? n11556 : n11564;
  assign n11566 = pi14 ? n11550 : n11565;
  assign n11567 = pi19 ? n37 : n139;
  assign n11568 = pi18 ? n37 : n11567;
  assign n11569 = pi22 ? n7513 : n32;
  assign n11570 = pi21 ? n139 : n11569;
  assign n11571 = pi20 ? n11570 : n32;
  assign n11572 = pi19 ? n11571 : n32;
  assign n11573 = pi18 ? n139 : n11572;
  assign n11574 = pi17 ? n11568 : n11573;
  assign n11575 = pi16 ? n439 : n11574;
  assign n11576 = pi20 ? n8209 : n3245;
  assign n11577 = pi19 ? n37 : n11576;
  assign n11578 = pi18 ? n37 : n11577;
  assign n11579 = pi21 ? n1211 : n1529;
  assign n11580 = pi20 ? n11579 : n3557;
  assign n11581 = pi20 ? n1737 : n3913;
  assign n11582 = pi19 ? n11580 : n11581;
  assign n11583 = pi21 ? n295 : n3175;
  assign n11584 = pi20 ? n11583 : n32;
  assign n11585 = pi19 ? n11584 : n32;
  assign n11586 = pi18 ? n11582 : n11585;
  assign n11587 = pi17 ? n11578 : n11586;
  assign n11588 = pi16 ? n439 : n11587;
  assign n11589 = pi21 ? n335 : n3175;
  assign n11590 = pi20 ? n11589 : n32;
  assign n11591 = pi19 ? n11590 : n32;
  assign n11592 = pi18 ? n37 : n11591;
  assign n11593 = pi17 ? n37 : n11592;
  assign n11594 = pi16 ? n439 : n11593;
  assign n11595 = pi15 ? n11588 : n11594;
  assign n11596 = pi14 ? n11575 : n11595;
  assign n11597 = pi13 ? n11566 : n11596;
  assign n11598 = pi19 ? n10957 : n2068;
  assign n11599 = pi18 ? n11598 : n11591;
  assign n11600 = pi17 ? n37 : n11599;
  assign n11601 = pi16 ? n439 : n11600;
  assign n11602 = pi21 ? n569 : n4109;
  assign n11603 = pi20 ? n11602 : n32;
  assign n11604 = pi19 ? n11603 : n32;
  assign n11605 = pi18 ? n37 : n11604;
  assign n11606 = pi17 ? n37 : n11605;
  assign n11607 = pi16 ? n439 : n11606;
  assign n11608 = pi15 ? n11601 : n11607;
  assign n11609 = pi14 ? n11608 : n11607;
  assign n11610 = pi21 ? n569 : n760;
  assign n11611 = pi20 ? n11610 : n32;
  assign n11612 = pi19 ? n11611 : n32;
  assign n11613 = pi18 ? n37 : n11612;
  assign n11614 = pi17 ? n37 : n11613;
  assign n11615 = pi16 ? n439 : n11614;
  assign n11616 = pi22 ? n583 : n2060;
  assign n11617 = pi21 ? n11616 : n2637;
  assign n11618 = pi20 ? n11617 : n32;
  assign n11619 = pi19 ? n11618 : n32;
  assign n11620 = pi18 ? n37 : n11619;
  assign n11621 = pi17 ? n37 : n11620;
  assign n11622 = pi16 ? n439 : n11621;
  assign n11623 = pi15 ? n11615 : n11622;
  assign n11624 = pi21 ? n11616 : n928;
  assign n11625 = pi20 ? n11624 : n32;
  assign n11626 = pi19 ? n11625 : n32;
  assign n11627 = pi18 ? n37 : n11626;
  assign n11628 = pi17 ? n37 : n11627;
  assign n11629 = pi16 ? n439 : n11628;
  assign n11630 = pi21 ? n4975 : n580;
  assign n11631 = pi20 ? n37 : n11630;
  assign n11632 = pi20 ? n37 : n3292;
  assign n11633 = pi19 ? n11631 : n11632;
  assign n11634 = pi18 ? n37 : n11633;
  assign n11635 = pi22 ? n5011 : n233;
  assign n11636 = pi21 ? n11635 : n928;
  assign n11637 = pi20 ? n11636 : n32;
  assign n11638 = pi19 ? n11637 : n32;
  assign n11639 = pi18 ? n37 : n11638;
  assign n11640 = pi17 ? n11634 : n11639;
  assign n11641 = pi16 ? n439 : n11640;
  assign n11642 = pi15 ? n11629 : n11641;
  assign n11643 = pi14 ? n11623 : n11642;
  assign n11644 = pi13 ? n11609 : n11643;
  assign n11645 = pi12 ? n11597 : n11644;
  assign n11646 = pi11 ? n11519 : n11645;
  assign n11647 = pi21 ? n2091 : n1009;
  assign n11648 = pi20 ? n11647 : n32;
  assign n11649 = pi19 ? n11648 : n32;
  assign n11650 = pi18 ? n37 : n11649;
  assign n11651 = pi17 ? n37 : n11650;
  assign n11652 = pi16 ? n439 : n11651;
  assign n11653 = pi20 ? n37 : n561;
  assign n11654 = pi19 ? n37 : n11653;
  assign n11655 = pi18 ? n11654 : n11649;
  assign n11656 = pi17 ? n37 : n11655;
  assign n11657 = pi16 ? n439 : n11656;
  assign n11658 = pi15 ? n11652 : n11657;
  assign n11659 = pi21 ? n2091 : n32;
  assign n11660 = pi20 ? n11659 : n32;
  assign n11661 = pi19 ? n11660 : n32;
  assign n11662 = pi18 ? n37 : n11661;
  assign n11663 = pi17 ? n37 : n11662;
  assign n11664 = pi16 ? n439 : n11663;
  assign n11665 = pi21 ? n2106 : n32;
  assign n11666 = pi20 ? n11665 : n32;
  assign n11667 = pi19 ? n11666 : n32;
  assign n11668 = pi18 ? n37 : n11667;
  assign n11669 = pi17 ? n37 : n11668;
  assign n11670 = pi16 ? n439 : n11669;
  assign n11671 = pi15 ? n11664 : n11670;
  assign n11672 = pi14 ? n11658 : n11671;
  assign n11673 = pi15 ? n11670 : n11220;
  assign n11674 = pi21 ? n685 : n32;
  assign n11675 = pi20 ? n11674 : n32;
  assign n11676 = pi19 ? n11675 : n32;
  assign n11677 = pi18 ? n37 : n11676;
  assign n11678 = pi17 ? n37 : n11677;
  assign n11679 = pi16 ? n439 : n11678;
  assign n11680 = pi23 ? n37 : n7420;
  assign n11681 = pi23 ? n2766 : n316;
  assign n11682 = pi22 ? n11680 : n11681;
  assign n11683 = pi21 ? n11682 : n32;
  assign n11684 = pi20 ? n11683 : n32;
  assign n11685 = pi19 ? n11684 : n32;
  assign n11686 = pi18 ? n37 : n11685;
  assign n11687 = pi17 ? n37 : n11686;
  assign n11688 = pi16 ? n439 : n11687;
  assign n11689 = pi15 ? n11679 : n11688;
  assign n11690 = pi14 ? n11673 : n11689;
  assign n11691 = pi13 ? n11672 : n11690;
  assign n11692 = pi18 ? n99 : n10313;
  assign n11693 = pi17 ? n99 : n11692;
  assign n11694 = pi16 ? n201 : n11693;
  assign n11695 = pi21 ? n2147 : n32;
  assign n11696 = pi20 ? n11695 : n32;
  assign n11697 = pi19 ? n11696 : n32;
  assign n11698 = pi18 ? n99 : n11697;
  assign n11699 = pi17 ? n99 : n11698;
  assign n11700 = pi16 ? n721 : n11699;
  assign n11701 = pi15 ? n11694 : n11700;
  assign n11702 = pi18 ? n5093 : n11245;
  assign n11703 = pi17 ? n99 : n11702;
  assign n11704 = pi16 ? n721 : n11703;
  assign n11705 = pi15 ? n11700 : n11704;
  assign n11706 = pi14 ? n11701 : n11705;
  assign n11707 = pi20 ? n7754 : n685;
  assign n11708 = pi19 ? n99 : n11707;
  assign n11709 = pi18 ? n11708 : n11245;
  assign n11710 = pi17 ? n99 : n11709;
  assign n11711 = pi16 ? n721 : n11710;
  assign n11712 = pi18 ? n9992 : n9458;
  assign n11713 = pi17 ? n157 : n11712;
  assign n11714 = pi16 ? n5910 : n11713;
  assign n11715 = pi15 ? n11711 : n11714;
  assign n11716 = pi18 ? n157 : n5669;
  assign n11717 = pi17 ? n157 : n11716;
  assign n11718 = pi16 ? n5910 : n11717;
  assign n11719 = pi18 ? n1667 : n5669;
  assign n11720 = pi17 ? n99 : n11719;
  assign n11721 = pi16 ? n744 : n11720;
  assign n11722 = pi15 ? n11718 : n11721;
  assign n11723 = pi14 ? n11715 : n11722;
  assign n11724 = pi13 ? n11706 : n11723;
  assign n11725 = pi12 ? n11691 : n11724;
  assign n11726 = pi18 ? n1667 : n4010;
  assign n11727 = pi17 ? n99 : n11726;
  assign n11728 = pi16 ? n744 : n11727;
  assign n11729 = pi21 ? n6472 : n4247;
  assign n11730 = pi20 ? n32 : n11729;
  assign n11731 = pi19 ? n32 : n11730;
  assign n11732 = pi22 ? n812 : n112;
  assign n11733 = pi21 ? n11732 : n4247;
  assign n11734 = pi21 ? n4234 : n4221;
  assign n11735 = pi21 ? n4247 : n4234;
  assign n11736 = pi20 ? n11734 : n11735;
  assign n11737 = pi19 ? n11733 : n11736;
  assign n11738 = pi18 ? n11731 : n11737;
  assign n11739 = pi17 ? n32 : n11738;
  assign n11740 = pi21 ? n99 : n4234;
  assign n11741 = pi22 ? n112 : n139;
  assign n11742 = pi21 ? n4221 : n11741;
  assign n11743 = pi21 ? n4221 : n4247;
  assign n11744 = pi20 ? n11742 : n11743;
  assign n11745 = pi19 ? n11740 : n11744;
  assign n11746 = pi20 ? n4252 : n4247;
  assign n11747 = pi21 ? n4237 : n4221;
  assign n11748 = pi20 ? n11735 : n11747;
  assign n11749 = pi19 ? n11746 : n11748;
  assign n11750 = pi18 ? n11745 : n11749;
  assign n11751 = pi20 ? n11735 : n11734;
  assign n11752 = pi21 ? n248 : n862;
  assign n11753 = pi20 ? n11735 : n11752;
  assign n11754 = pi19 ? n11751 : n11753;
  assign n11755 = pi18 ? n11754 : n4010;
  assign n11756 = pi17 ? n11750 : n11755;
  assign n11757 = pi16 ? n11739 : n11756;
  assign n11758 = pi15 ? n11728 : n11757;
  assign n11759 = pi20 ? n139 : n157;
  assign n11760 = pi19 ? n139 : n11759;
  assign n11761 = pi18 ? n11760 : n3212;
  assign n11762 = pi17 ? n139 : n11761;
  assign n11763 = pi16 ? n915 : n11762;
  assign n11764 = pi20 ? n139 : n5199;
  assign n11765 = pi19 ? n139 : n11764;
  assign n11766 = pi18 ? n11765 : n3212;
  assign n11767 = pi17 ? n139 : n11766;
  assign n11768 = pi16 ? n915 : n11767;
  assign n11769 = pi15 ? n11763 : n11768;
  assign n11770 = pi14 ? n11758 : n11769;
  assign n11771 = pi18 ? n5285 : n316;
  assign n11772 = pi17 ? n32 : n11771;
  assign n11773 = pi18 ? n316 : n3212;
  assign n11774 = pi17 ? n5307 : n11773;
  assign n11775 = pi16 ? n11772 : n11774;
  assign n11776 = pi21 ? n3692 : n316;
  assign n11777 = pi20 ? n32 : n11776;
  assign n11778 = pi19 ? n32 : n11777;
  assign n11779 = pi18 ? n11778 : n316;
  assign n11780 = pi17 ? n32 : n11779;
  assign n11781 = pi17 ? n316 : n11773;
  assign n11782 = pi16 ? n11780 : n11781;
  assign n11783 = pi18 ? n10879 : n316;
  assign n11784 = pi17 ? n32 : n11783;
  assign n11785 = pi21 ? n359 : n316;
  assign n11786 = pi20 ? n11785 : n316;
  assign n11787 = pi19 ? n11786 : n316;
  assign n11788 = pi18 ? n11787 : n316;
  assign n11789 = pi17 ? n11788 : n10886;
  assign n11790 = pi16 ? n11784 : n11789;
  assign n11791 = pi15 ? n11782 : n11790;
  assign n11792 = pi14 ? n11775 : n11791;
  assign n11793 = pi13 ? n11770 : n11792;
  assign n11794 = pi18 ? n9111 : n10013;
  assign n11795 = pi17 ? n139 : n11794;
  assign n11796 = pi16 ? n331 : n11795;
  assign n11797 = pi20 ? n139 : n2353;
  assign n11798 = pi19 ? n139 : n11797;
  assign n11799 = pi18 ? n11798 : n10013;
  assign n11800 = pi17 ? n139 : n11799;
  assign n11801 = pi16 ? n331 : n11800;
  assign n11802 = pi15 ? n11796 : n11801;
  assign n11803 = pi18 ? n6157 : n204;
  assign n11804 = pi17 ? n32 : n11803;
  assign n11805 = pi20 ? n577 : n204;
  assign n11806 = pi19 ? n11805 : n204;
  assign n11807 = pi18 ? n11806 : n204;
  assign n11808 = pi22 ? n204 : n233;
  assign n11809 = pi21 ? n204 : n11808;
  assign n11810 = pi20 ? n204 : n11809;
  assign n11811 = pi19 ? n204 : n11810;
  assign n11812 = pi18 ? n11811 : n2655;
  assign n11813 = pi17 ? n11807 : n11812;
  assign n11814 = pi16 ? n11804 : n11813;
  assign n11815 = pi20 ? n335 : n204;
  assign n11816 = pi19 ? n11815 : n204;
  assign n11817 = pi18 ? n11816 : n204;
  assign n11818 = pi22 ? n335 : n3762;
  assign n11819 = pi21 ? n204 : n11818;
  assign n11820 = pi20 ? n204 : n11819;
  assign n11821 = pi19 ? n204 : n11820;
  assign n11822 = pi18 ? n11821 : n2703;
  assign n11823 = pi17 ? n11817 : n11822;
  assign n11824 = pi16 ? n11804 : n11823;
  assign n11825 = pi15 ? n11814 : n11824;
  assign n11826 = pi14 ? n11802 : n11825;
  assign n11827 = pi20 ? n8857 : n335;
  assign n11828 = pi19 ? n11827 : n335;
  assign n11829 = pi18 ? n11828 : n335;
  assign n11830 = pi22 ? n10400 : n3762;
  assign n11831 = pi21 ? n335 : n11830;
  assign n11832 = pi20 ? n335 : n11831;
  assign n11833 = pi19 ? n335 : n11832;
  assign n11834 = pi18 ? n11833 : n1824;
  assign n11835 = pi17 ? n11829 : n11834;
  assign n11836 = pi16 ? n3351 : n11835;
  assign n11837 = pi22 ? n10400 : n1070;
  assign n11838 = pi21 ? n335 : n11837;
  assign n11839 = pi20 ? n335 : n11838;
  assign n11840 = pi19 ? n335 : n11839;
  assign n11841 = pi18 ? n11840 : n32;
  assign n11842 = pi17 ? n335 : n11841;
  assign n11843 = pi16 ? n2035 : n11842;
  assign n11844 = pi15 ? n11836 : n11843;
  assign n11845 = pi21 ? n716 : n335;
  assign n11846 = pi20 ? n32 : n11845;
  assign n11847 = pi19 ? n32 : n11846;
  assign n11848 = pi18 ? n11847 : n335;
  assign n11849 = pi17 ? n32 : n11848;
  assign n11850 = pi22 ? n3935 : n1070;
  assign n11851 = pi21 ? n335 : n11850;
  assign n11852 = pi20 ? n335 : n11851;
  assign n11853 = pi19 ? n335 : n11852;
  assign n11854 = pi18 ? n11853 : n32;
  assign n11855 = pi17 ? n335 : n11854;
  assign n11856 = pi16 ? n11849 : n11855;
  assign n11857 = pi21 ? n335 : n9430;
  assign n11858 = pi20 ? n335 : n11857;
  assign n11859 = pi19 ? n335 : n11858;
  assign n11860 = pi18 ? n11859 : n32;
  assign n11861 = pi17 ? n335 : n11860;
  assign n11862 = pi16 ? n10118 : n11861;
  assign n11863 = pi15 ? n11856 : n11862;
  assign n11864 = pi14 ? n11844 : n11863;
  assign n11865 = pi13 ? n11826 : n11864;
  assign n11866 = pi12 ? n11793 : n11865;
  assign n11867 = pi11 ? n11725 : n11866;
  assign n11868 = pi10 ? n11646 : n11867;
  assign n11869 = pi09 ? n11378 : n11868;
  assign n11870 = pi15 ? n32 : n11371;
  assign n11871 = pi16 ? n9232 : n11368;
  assign n11872 = pi15 ? n11372 : n11871;
  assign n11873 = pi14 ? n11870 : n11872;
  assign n11874 = pi13 ? n32 : n11873;
  assign n11875 = pi12 ? n32 : n11874;
  assign n11876 = pi11 ? n32 : n11875;
  assign n11877 = pi10 ? n32 : n11876;
  assign n11878 = pi16 ? n2461 : n11383;
  assign n11879 = pi16 ? n10154 : n11389;
  assign n11880 = pi15 ? n11878 : n11879;
  assign n11881 = pi16 ? n11011 : n10458;
  assign n11882 = pi20 ? n32 : n41;
  assign n11883 = pi19 ? n32 : n11882;
  assign n11884 = pi18 ? n11883 : n37;
  assign n11885 = pi17 ? n32 : n11884;
  assign n11886 = pi16 ? n11885 : n11398;
  assign n11887 = pi15 ? n11881 : n11886;
  assign n11888 = pi14 ? n11880 : n11887;
  assign n11889 = pi23 ? n37 : n1342;
  assign n11890 = pi22 ? n11889 : n32;
  assign n11891 = pi21 ? n37 : n11890;
  assign n11892 = pi20 ? n11891 : n32;
  assign n11893 = pi19 ? n11892 : n32;
  assign n11894 = pi18 ? n37 : n11893;
  assign n11895 = pi17 ? n37 : n11894;
  assign n11896 = pi16 ? n439 : n11895;
  assign n11897 = pi20 ? n2165 : n2755;
  assign n11898 = pi19 ? n11897 : n3808;
  assign n11899 = pi18 ? n8057 : n11898;
  assign n11900 = pi17 ? n32 : n11899;
  assign n11901 = pi20 ? n11424 : n2755;
  assign n11902 = pi19 ? n3813 : n11901;
  assign n11903 = pi20 ? n2755 : n11424;
  assign n11904 = pi21 ? n1143 : n2160;
  assign n11905 = pi20 ? n2755 : n11904;
  assign n11906 = pi19 ? n11903 : n11905;
  assign n11907 = pi18 ? n11902 : n11906;
  assign n11908 = pi20 ? n3506 : n11424;
  assign n11909 = pi19 ? n11908 : n3825;
  assign n11910 = pi24 ? n99 : n363;
  assign n11911 = pi23 ? n37 : n11910;
  assign n11912 = pi22 ? n11911 : n32;
  assign n11913 = pi21 ? n2175 : n11912;
  assign n11914 = pi20 ? n11913 : n32;
  assign n11915 = pi19 ? n11914 : n32;
  assign n11916 = pi18 ? n11909 : n11915;
  assign n11917 = pi17 ? n11907 : n11916;
  assign n11918 = pi16 ? n11900 : n11917;
  assign n11919 = pi15 ? n11896 : n11918;
  assign n11920 = pi23 ? n99 : n1432;
  assign n11921 = pi22 ? n11920 : n32;
  assign n11922 = pi21 ? n99 : n11921;
  assign n11923 = pi20 ? n11922 : n32;
  assign n11924 = pi19 ? n11923 : n32;
  assign n11925 = pi18 ? n99 : n11924;
  assign n11926 = pi17 ? n99 : n11925;
  assign n11927 = pi16 ? n801 : n11926;
  assign n11928 = pi22 ? n157 : n2468;
  assign n11929 = pi21 ? n157 : n11928;
  assign n11930 = pi20 ? n11929 : n32;
  assign n11931 = pi19 ? n11930 : n32;
  assign n11932 = pi18 ? n157 : n11931;
  assign n11933 = pi17 ? n157 : n11932;
  assign n11934 = pi16 ? n11448 : n11933;
  assign n11935 = pi15 ? n11927 : n11934;
  assign n11936 = pi14 ? n11919 : n11935;
  assign n11937 = pi13 ? n11888 : n11936;
  assign n11938 = pi22 ? n99 : n2468;
  assign n11939 = pi21 ? n99 : n11938;
  assign n11940 = pi20 ? n11939 : n32;
  assign n11941 = pi19 ? n11940 : n32;
  assign n11942 = pi18 ? n99 : n11941;
  assign n11943 = pi17 ? n99 : n11942;
  assign n11944 = pi16 ? n721 : n11943;
  assign n11945 = pi22 ? n99 : n532;
  assign n11946 = pi21 ? n99 : n11945;
  assign n11947 = pi20 ? n11946 : n32;
  assign n11948 = pi19 ? n11947 : n32;
  assign n11949 = pi18 ? n99 : n11948;
  assign n11950 = pi17 ? n99 : n11949;
  assign n11951 = pi16 ? n801 : n11950;
  assign n11952 = pi15 ? n11944 : n11951;
  assign n11953 = pi22 ? n3492 : n625;
  assign n11954 = pi21 ? n99 : n11953;
  assign n11955 = pi20 ? n11954 : n32;
  assign n11956 = pi19 ? n11955 : n32;
  assign n11957 = pi18 ? n99 : n11956;
  assign n11958 = pi17 ? n99 : n11957;
  assign n11959 = pi16 ? n11478 : n11958;
  assign n11960 = pi15 ? n11951 : n11959;
  assign n11961 = pi14 ? n11952 : n11960;
  assign n11962 = pi24 ? n99 : n335;
  assign n11963 = pi23 ? n99 : n11962;
  assign n11964 = pi22 ? n11963 : n625;
  assign n11965 = pi21 ? n99 : n11964;
  assign n11966 = pi20 ? n11965 : n32;
  assign n11967 = pi19 ? n11966 : n32;
  assign n11968 = pi18 ? n99 : n11967;
  assign n11969 = pi17 ? n99 : n11968;
  assign n11970 = pi16 ? n11486 : n11969;
  assign n11971 = pi22 ? n7377 : n688;
  assign n11972 = pi21 ? n99 : n11971;
  assign n11973 = pi20 ? n11972 : n32;
  assign n11974 = pi19 ? n11973 : n32;
  assign n11975 = pi18 ? n99 : n11974;
  assign n11976 = pi17 ? n99 : n11975;
  assign n11977 = pi16 ? n721 : n11976;
  assign n11978 = pi15 ? n11970 : n11977;
  assign n11979 = pi21 ? n316 : n3494;
  assign n11980 = pi20 ? n11979 : n32;
  assign n11981 = pi19 ? n11980 : n32;
  assign n11982 = pi18 ? n316 : n11981;
  assign n11983 = pi17 ? n11498 : n11982;
  assign n11984 = pi16 ? n439 : n11983;
  assign n11985 = pi20 ? n9544 : n7571;
  assign n11986 = pi19 ? n316 : n11985;
  assign n11987 = pi18 ? n11986 : n11500;
  assign n11988 = pi17 ? n11511 : n11987;
  assign n11989 = pi16 ? n439 : n11988;
  assign n11990 = pi15 ? n11984 : n11989;
  assign n11991 = pi14 ? n11978 : n11990;
  assign n11992 = pi13 ? n11961 : n11991;
  assign n11993 = pi12 ? n11937 : n11992;
  assign n11994 = pi22 ? n8174 : n32;
  assign n11995 = pi21 ? n139 : n11994;
  assign n11996 = pi20 ? n11995 : n32;
  assign n11997 = pi19 ? n11996 : n32;
  assign n11998 = pi18 ? n139 : n11997;
  assign n11999 = pi17 ? n11558 : n11998;
  assign n12000 = pi16 ? n439 : n11999;
  assign n12001 = pi15 ? n11556 : n12000;
  assign n12002 = pi14 ? n11550 : n12001;
  assign n12003 = pi22 ? n8198 : n32;
  assign n12004 = pi21 ? n139 : n12003;
  assign n12005 = pi20 ? n12004 : n32;
  assign n12006 = pi19 ? n12005 : n32;
  assign n12007 = pi18 ? n139 : n12006;
  assign n12008 = pi17 ? n11568 : n12007;
  assign n12009 = pi16 ? n439 : n12008;
  assign n12010 = pi21 ? n1696 : n375;
  assign n12011 = pi20 ? n8209 : n12010;
  assign n12012 = pi19 ? n37 : n12011;
  assign n12013 = pi18 ? n37 : n12012;
  assign n12014 = pi21 ? n1531 : n1696;
  assign n12015 = pi20 ? n11579 : n12014;
  assign n12016 = pi20 ? n12014 : n3579;
  assign n12017 = pi19 ? n12015 : n12016;
  assign n12018 = pi23 ? n204 : n1149;
  assign n12019 = pi22 ? n12018 : n32;
  assign n12020 = pi21 ? n375 : n12019;
  assign n12021 = pi20 ? n12020 : n32;
  assign n12022 = pi19 ? n12021 : n32;
  assign n12023 = pi18 ? n12017 : n12022;
  assign n12024 = pi17 ? n12013 : n12023;
  assign n12025 = pi16 ? n439 : n12024;
  assign n12026 = pi21 ? n335 : n12019;
  assign n12027 = pi20 ? n12026 : n32;
  assign n12028 = pi19 ? n12027 : n32;
  assign n12029 = pi18 ? n37 : n12028;
  assign n12030 = pi17 ? n37 : n12029;
  assign n12031 = pi16 ? n439 : n12030;
  assign n12032 = pi15 ? n12025 : n12031;
  assign n12033 = pi14 ? n12009 : n12032;
  assign n12034 = pi13 ? n12002 : n12033;
  assign n12035 = pi21 ? n569 : n5813;
  assign n12036 = pi20 ? n12035 : n32;
  assign n12037 = pi19 ? n12036 : n32;
  assign n12038 = pi18 ? n37 : n12037;
  assign n12039 = pi17 ? n37 : n12038;
  assign n12040 = pi16 ? n439 : n12039;
  assign n12041 = pi15 ? n11601 : n12040;
  assign n12042 = pi21 ? n569 : n7034;
  assign n12043 = pi20 ? n12042 : n32;
  assign n12044 = pi19 ? n12043 : n32;
  assign n12045 = pi18 ? n37 : n12044;
  assign n12046 = pi17 ? n37 : n12045;
  assign n12047 = pi16 ? n439 : n12046;
  assign n12048 = pi15 ? n11607 : n12047;
  assign n12049 = pi14 ? n12041 : n12048;
  assign n12050 = pi21 ? n2074 : n6416;
  assign n12051 = pi20 ? n12050 : n32;
  assign n12052 = pi19 ? n12051 : n32;
  assign n12053 = pi18 ? n37 : n12052;
  assign n12054 = pi17 ? n37 : n12053;
  assign n12055 = pi16 ? n439 : n12054;
  assign n12056 = pi21 ? n11616 : n760;
  assign n12057 = pi20 ? n12056 : n32;
  assign n12058 = pi19 ? n12057 : n32;
  assign n12059 = pi18 ? n37 : n12058;
  assign n12060 = pi17 ? n37 : n12059;
  assign n12061 = pi16 ? n439 : n12060;
  assign n12062 = pi15 ? n12055 : n12061;
  assign n12063 = pi20 ? n37 : n580;
  assign n12064 = pi19 ? n12063 : n11632;
  assign n12065 = pi18 ? n37 : n12064;
  assign n12066 = pi21 ? n11635 : n882;
  assign n12067 = pi20 ? n12066 : n32;
  assign n12068 = pi19 ? n12067 : n32;
  assign n12069 = pi18 ? n37 : n12068;
  assign n12070 = pi17 ? n12065 : n12069;
  assign n12071 = pi16 ? n439 : n12070;
  assign n12072 = pi15 ? n11622 : n12071;
  assign n12073 = pi14 ? n12062 : n12072;
  assign n12074 = pi13 ? n12049 : n12073;
  assign n12075 = pi12 ? n12034 : n12074;
  assign n12076 = pi11 ? n11993 : n12075;
  assign n12077 = pi21 ? n2091 : n928;
  assign n12078 = pi20 ? n12077 : n32;
  assign n12079 = pi19 ? n12078 : n32;
  assign n12080 = pi18 ? n37 : n12079;
  assign n12081 = pi17 ? n37 : n12080;
  assign n12082 = pi16 ? n439 : n12081;
  assign n12083 = pi18 ? n11654 : n12079;
  assign n12084 = pi17 ? n37 : n12083;
  assign n12085 = pi16 ? n439 : n12084;
  assign n12086 = pi15 ? n12082 : n12085;
  assign n12087 = pi21 ? n2106 : n2678;
  assign n12088 = pi20 ? n12087 : n32;
  assign n12089 = pi19 ? n12088 : n32;
  assign n12090 = pi18 ? n37 : n12089;
  assign n12091 = pi17 ? n37 : n12090;
  assign n12092 = pi16 ? n439 : n12091;
  assign n12093 = pi15 ? n9883 : n12092;
  assign n12094 = pi14 ? n12086 : n12093;
  assign n12095 = pi21 ? n2106 : n2700;
  assign n12096 = pi20 ? n12095 : n32;
  assign n12097 = pi19 ? n12096 : n32;
  assign n12098 = pi18 ? n37 : n12097;
  assign n12099 = pi17 ? n37 : n12098;
  assign n12100 = pi16 ? n439 : n12099;
  assign n12101 = pi21 ? n2721 : n2700;
  assign n12102 = pi20 ? n12101 : n32;
  assign n12103 = pi19 ? n12102 : n32;
  assign n12104 = pi18 ? n37 : n12103;
  assign n12105 = pi17 ? n37 : n12104;
  assign n12106 = pi16 ? n439 : n12105;
  assign n12107 = pi15 ? n12100 : n12106;
  assign n12108 = pi18 ? n37 : n7409;
  assign n12109 = pi17 ? n37 : n12108;
  assign n12110 = pi16 ? n439 : n12109;
  assign n12111 = pi22 ? n295 : n1484;
  assign n12112 = pi21 ? n12111 : n1009;
  assign n12113 = pi20 ? n12112 : n32;
  assign n12114 = pi19 ? n12113 : n32;
  assign n12115 = pi18 ? n37 : n12114;
  assign n12116 = pi17 ? n37 : n12115;
  assign n12117 = pi16 ? n439 : n12116;
  assign n12118 = pi15 ? n12110 : n12117;
  assign n12119 = pi14 ? n12107 : n12118;
  assign n12120 = pi13 ? n12094 : n12119;
  assign n12121 = pi18 ? n99 : n11217;
  assign n12122 = pi17 ? n99 : n12121;
  assign n12123 = pi16 ? n201 : n12122;
  assign n12124 = pi18 ? n99 : n11676;
  assign n12125 = pi17 ? n99 : n12124;
  assign n12126 = pi16 ? n744 : n12125;
  assign n12127 = pi15 ? n12123 : n12126;
  assign n12128 = pi21 ? n5113 : n32;
  assign n12129 = pi20 ? n12128 : n32;
  assign n12130 = pi19 ? n12129 : n32;
  assign n12131 = pi18 ? n99 : n12130;
  assign n12132 = pi17 ? n99 : n12131;
  assign n12133 = pi16 ? n744 : n12132;
  assign n12134 = pi18 ? n5093 : n12130;
  assign n12135 = pi17 ? n99 : n12134;
  assign n12136 = pi16 ? n744 : n12135;
  assign n12137 = pi15 ? n12133 : n12136;
  assign n12138 = pi14 ? n12127 : n12137;
  assign n12139 = pi16 ? n744 : n11710;
  assign n12140 = pi18 ? n9992 : n11245;
  assign n12141 = pi17 ? n157 : n12140;
  assign n12142 = pi16 ? n5910 : n12141;
  assign n12143 = pi15 ? n12139 : n12142;
  assign n12144 = pi16 ? n721 : n11720;
  assign n12145 = pi15 ? n11718 : n12144;
  assign n12146 = pi14 ? n12143 : n12145;
  assign n12147 = pi13 ? n12138 : n12146;
  assign n12148 = pi12 ? n12120 : n12147;
  assign n12149 = pi21 ? n3494 : n32;
  assign n12150 = pi20 ? n12149 : n32;
  assign n12151 = pi19 ? n12150 : n32;
  assign n12152 = pi18 ? n1667 : n12151;
  assign n12153 = pi17 ? n99 : n12152;
  assign n12154 = pi16 ? n721 : n12153;
  assign n12155 = pi23 ? n961 : n99;
  assign n12156 = pi22 ? n12155 : n295;
  assign n12157 = pi21 ? n12156 : n4252;
  assign n12158 = pi20 ? n32 : n12157;
  assign n12159 = pi19 ? n32 : n12158;
  assign n12160 = pi21 ? n4226 : n4252;
  assign n12161 = pi21 ? n4234 : n812;
  assign n12162 = pi20 ? n12161 : n11735;
  assign n12163 = pi19 ? n12160 : n12162;
  assign n12164 = pi18 ? n12159 : n12163;
  assign n12165 = pi17 ? n32 : n12164;
  assign n12166 = pi21 ? n4221 : n4234;
  assign n12167 = pi20 ? n11740 : n12166;
  assign n12168 = pi21 ? n4221 : n1721;
  assign n12169 = pi21 ? n4234 : n4252;
  assign n12170 = pi20 ? n12168 : n12169;
  assign n12171 = pi19 ? n12167 : n12170;
  assign n12172 = pi21 ? n4252 : n4247;
  assign n12173 = pi20 ? n4252 : n12172;
  assign n12174 = pi21 ? n4234 : n4237;
  assign n12175 = pi20 ? n11735 : n12174;
  assign n12176 = pi19 ? n12173 : n12175;
  assign n12177 = pi18 ? n12171 : n12176;
  assign n12178 = pi21 ? n4252 : n139;
  assign n12179 = pi20 ? n12178 : n12174;
  assign n12180 = pi20 ? n12178 : n11752;
  assign n12181 = pi19 ? n12179 : n12180;
  assign n12182 = pi18 ? n12181 : n4010;
  assign n12183 = pi17 ? n12177 : n12182;
  assign n12184 = pi16 ? n12165 : n12183;
  assign n12185 = pi15 ? n12154 : n12184;
  assign n12186 = pi16 ? n2291 : n11762;
  assign n12187 = pi15 ? n12186 : n11768;
  assign n12188 = pi14 ? n12185 : n12187;
  assign n12189 = pi18 ? n9093 : n316;
  assign n12190 = pi17 ? n32 : n12189;
  assign n12191 = pi16 ? n12190 : n11781;
  assign n12192 = pi21 ? n2835 : n32;
  assign n12193 = pi20 ? n12192 : n32;
  assign n12194 = pi19 ? n12193 : n32;
  assign n12195 = pi18 ? n316 : n12194;
  assign n12196 = pi17 ? n11788 : n12195;
  assign n12197 = pi16 ? n12190 : n12196;
  assign n12198 = pi15 ? n12191 : n12197;
  assign n12199 = pi14 ? n11775 : n12198;
  assign n12200 = pi13 ? n12188 : n12199;
  assign n12201 = pi18 ? n11821 : n2655;
  assign n12202 = pi17 ? n11817 : n12201;
  assign n12203 = pi16 ? n11804 : n12202;
  assign n12204 = pi15 ? n11814 : n12203;
  assign n12205 = pi14 ? n11802 : n12204;
  assign n12206 = pi18 ? n11833 : n2655;
  assign n12207 = pi17 ? n11829 : n12206;
  assign n12208 = pi16 ? n3351 : n12207;
  assign n12209 = pi15 ? n12208 : n11843;
  assign n12210 = pi14 ? n12209 : n11863;
  assign n12211 = pi13 ? n12205 : n12210;
  assign n12212 = pi12 ? n12200 : n12211;
  assign n12213 = pi11 ? n12148 : n12212;
  assign n12214 = pi10 ? n12076 : n12213;
  assign n12215 = pi09 ? n11877 : n12214;
  assign n12216 = pi08 ? n11869 : n12215;
  assign n12217 = pi20 ? n86 : n32;
  assign n12218 = pi19 ? n12217 : n32;
  assign n12219 = pi18 ? n37 : n12218;
  assign n12220 = pi17 ? n37 : n12219;
  assign n12221 = pi16 ? n8027 : n12220;
  assign n12222 = pi15 ? n32 : n12221;
  assign n12223 = pi16 ? n1130 : n12220;
  assign n12224 = pi22 ? n37 : n119;
  assign n12225 = pi21 ? n37 : n12224;
  assign n12226 = pi20 ? n12225 : n32;
  assign n12227 = pi19 ? n12226 : n32;
  assign n12228 = pi18 ? n37 : n12227;
  assign n12229 = pi17 ? n37 : n12228;
  assign n12230 = pi16 ? n9232 : n12229;
  assign n12231 = pi15 ? n12223 : n12230;
  assign n12232 = pi14 ? n12222 : n12231;
  assign n12233 = pi13 ? n32 : n12232;
  assign n12234 = pi12 ? n32 : n12233;
  assign n12235 = pi11 ? n32 : n12234;
  assign n12236 = pi10 ? n32 : n12235;
  assign n12237 = pi21 ? n37 : n120;
  assign n12238 = pi20 ? n12237 : n32;
  assign n12239 = pi19 ? n12238 : n32;
  assign n12240 = pi18 ? n37 : n12239;
  assign n12241 = pi17 ? n37 : n12240;
  assign n12242 = pi16 ? n2461 : n12241;
  assign n12243 = pi22 ? n139 : n140;
  assign n12244 = pi21 ? n37 : n12243;
  assign n12245 = pi20 ? n12244 : n32;
  assign n12246 = pi19 ? n12245 : n32;
  assign n12247 = pi18 ? n37 : n12246;
  assign n12248 = pi17 ? n37 : n12247;
  assign n12249 = pi16 ? n10154 : n12248;
  assign n12250 = pi15 ? n12242 : n12249;
  assign n12251 = pi16 ? n11011 : n11389;
  assign n12252 = pi21 ? n37 : n588;
  assign n12253 = pi20 ? n12252 : n32;
  assign n12254 = pi19 ? n12253 : n32;
  assign n12255 = pi18 ? n37 : n12254;
  assign n12256 = pi17 ? n37 : n12255;
  assign n12257 = pi16 ? n11885 : n12256;
  assign n12258 = pi15 ? n12251 : n12257;
  assign n12259 = pi14 ? n12250 : n12258;
  assign n12260 = pi22 ? n37 : n587;
  assign n12261 = pi21 ? n37 : n12260;
  assign n12262 = pi20 ? n12261 : n32;
  assign n12263 = pi19 ? n12262 : n32;
  assign n12264 = pi18 ? n37 : n12263;
  assign n12265 = pi17 ? n37 : n12264;
  assign n12266 = pi16 ? n439 : n12265;
  assign n12267 = pi22 ? n99 : n5631;
  assign n12268 = pi21 ? n99 : n12267;
  assign n12269 = pi20 ? n12268 : n32;
  assign n12270 = pi19 ? n12269 : n32;
  assign n12271 = pi18 ? n99 : n12270;
  assign n12272 = pi17 ? n99 : n12271;
  assign n12273 = pi16 ? n3065 : n12272;
  assign n12274 = pi15 ? n12266 : n12273;
  assign n12275 = pi20 ? n99 : n4619;
  assign n12276 = pi19 ? n12275 : n4624;
  assign n12277 = pi18 ? n742 : n12276;
  assign n12278 = pi17 ? n32 : n12277;
  assign n12279 = pi20 ? n4617 : n3506;
  assign n12280 = pi21 ? n2164 : n2168;
  assign n12281 = pi20 ? n12280 : n11418;
  assign n12282 = pi19 ? n12279 : n12281;
  assign n12283 = pi21 ? n112 : n2168;
  assign n12284 = pi20 ? n11418 : n12283;
  assign n12285 = pi19 ? n12284 : n3882;
  assign n12286 = pi18 ? n12282 : n12285;
  assign n12287 = pi21 ? n218 : n2168;
  assign n12288 = pi20 ? n12287 : n3822;
  assign n12289 = pi21 ? n2162 : n112;
  assign n12290 = pi20 ? n12289 : n2174;
  assign n12291 = pi19 ? n12288 : n12290;
  assign n12292 = pi21 ? n2162 : n12267;
  assign n12293 = pi20 ? n12292 : n32;
  assign n12294 = pi19 ? n12293 : n32;
  assign n12295 = pi18 ? n12291 : n12294;
  assign n12296 = pi17 ? n12286 : n12295;
  assign n12297 = pi16 ? n12278 : n12296;
  assign n12298 = pi21 ? n796 : n777;
  assign n12299 = pi20 ? n32 : n12298;
  assign n12300 = pi19 ? n32 : n12299;
  assign n12301 = pi18 ? n12300 : n11446;
  assign n12302 = pi17 ? n32 : n12301;
  assign n12303 = pi16 ? n12302 : n11933;
  assign n12304 = pi15 ? n12297 : n12303;
  assign n12305 = pi14 ? n12274 : n12304;
  assign n12306 = pi13 ? n12259 : n12305;
  assign n12307 = pi16 ? n801 : n11943;
  assign n12308 = pi15 ? n12307 : n11951;
  assign n12309 = pi22 ? n745 : n625;
  assign n12310 = pi21 ? n99 : n12309;
  assign n12311 = pi20 ? n12310 : n32;
  assign n12312 = pi19 ? n12311 : n32;
  assign n12313 = pi18 ? n99 : n12312;
  assign n12314 = pi17 ? n99 : n12313;
  assign n12315 = pi16 ? n744 : n12314;
  assign n12316 = pi15 ? n11951 : n12315;
  assign n12317 = pi14 ? n12308 : n12316;
  assign n12318 = pi22 ? n1656 : n625;
  assign n12319 = pi21 ? n99 : n12318;
  assign n12320 = pi20 ? n12319 : n32;
  assign n12321 = pi19 ? n12320 : n32;
  assign n12322 = pi18 ? n99 : n12321;
  assign n12323 = pi17 ? n99 : n12322;
  assign n12324 = pi16 ? n744 : n12323;
  assign n12325 = pi22 ? n861 : n688;
  assign n12326 = pi21 ? n139 : n12325;
  assign n12327 = pi20 ? n12326 : n32;
  assign n12328 = pi19 ? n12327 : n32;
  assign n12329 = pi18 ? n139 : n12328;
  assign n12330 = pi17 ? n139 : n12329;
  assign n12331 = pi16 ? n915 : n12330;
  assign n12332 = pi15 ? n12324 : n12331;
  assign n12333 = pi21 ? n3258 : n391;
  assign n12334 = pi20 ? n37 : n12333;
  assign n12335 = pi19 ? n37 : n12334;
  assign n12336 = pi21 ? n316 : n390;
  assign n12337 = pi20 ? n12336 : n8742;
  assign n12338 = pi21 ? n3258 : n3073;
  assign n12339 = pi20 ? n12338 : n12333;
  assign n12340 = pi19 ? n12337 : n12339;
  assign n12341 = pi18 ? n12335 : n12340;
  assign n12342 = pi21 ? n4056 : n4052;
  assign n12343 = pi20 ? n316 : n12342;
  assign n12344 = pi21 ? n381 : n392;
  assign n12345 = pi21 ? n3073 : n392;
  assign n12346 = pi20 ? n12344 : n12345;
  assign n12347 = pi19 ? n12343 : n12346;
  assign n12348 = pi20 ? n5205 : n32;
  assign n12349 = pi19 ? n12348 : n32;
  assign n12350 = pi18 ? n12347 : n12349;
  assign n12351 = pi17 ? n12341 : n12350;
  assign n12352 = pi16 ? n439 : n12351;
  assign n12353 = pi20 ? n6625 : n37;
  assign n12354 = pi19 ? n12353 : n37;
  assign n12355 = pi18 ? n37 : n12354;
  assign n12356 = pi21 ? n3258 : n424;
  assign n12357 = pi21 ? n3118 : n37;
  assign n12358 = pi20 ? n12356 : n12357;
  assign n12359 = pi19 ? n12358 : n11072;
  assign n12360 = pi21 ? n4056 : n5178;
  assign n12361 = pi20 ? n12360 : n32;
  assign n12362 = pi19 ? n12361 : n32;
  assign n12363 = pi18 ? n12359 : n12362;
  assign n12364 = pi17 ? n12355 : n12363;
  assign n12365 = pi16 ? n439 : n12364;
  assign n12366 = pi15 ? n12352 : n12365;
  assign n12367 = pi14 ? n12332 : n12366;
  assign n12368 = pi13 ? n12317 : n12367;
  assign n12369 = pi12 ? n12306 : n12368;
  assign n12370 = pi20 ? n37 : n3083;
  assign n12371 = pi19 ? n37 : n12370;
  assign n12372 = pi18 ? n37 : n12371;
  assign n12373 = pi20 ? n1003 : n385;
  assign n12374 = pi19 ? n12373 : n11072;
  assign n12375 = pi21 ? n37 : n5178;
  assign n12376 = pi20 ? n12375 : n32;
  assign n12377 = pi19 ? n12376 : n32;
  assign n12378 = pi18 ? n12374 : n12377;
  assign n12379 = pi17 ? n12372 : n12378;
  assign n12380 = pi16 ? n439 : n12379;
  assign n12381 = pi22 ? n204 : n317;
  assign n12382 = pi21 ? n37 : n12381;
  assign n12383 = pi20 ? n12382 : n32;
  assign n12384 = pi19 ? n12383 : n32;
  assign n12385 = pi18 ? n37 : n12384;
  assign n12386 = pi17 ? n37 : n12385;
  assign n12387 = pi16 ? n439 : n12386;
  assign n12388 = pi15 ? n12380 : n12387;
  assign n12389 = pi22 ? n1038 : n706;
  assign n12390 = pi21 ? n139 : n12389;
  assign n12391 = pi20 ? n12390 : n32;
  assign n12392 = pi19 ? n12391 : n32;
  assign n12393 = pi18 ? n139 : n12392;
  assign n12394 = pi17 ? n11553 : n12393;
  assign n12395 = pi16 ? n439 : n12394;
  assign n12396 = pi21 ? n139 : n3970;
  assign n12397 = pi20 ? n12396 : n32;
  assign n12398 = pi19 ? n12397 : n32;
  assign n12399 = pi18 ? n139 : n12398;
  assign n12400 = pi17 ? n11558 : n12399;
  assign n12401 = pi16 ? n439 : n12400;
  assign n12402 = pi15 ? n12395 : n12401;
  assign n12403 = pi14 ? n12388 : n12402;
  assign n12404 = pi22 ? n204 : n32;
  assign n12405 = pi21 ? n139 : n12404;
  assign n12406 = pi20 ? n12405 : n32;
  assign n12407 = pi19 ? n12406 : n32;
  assign n12408 = pi18 ? n139 : n12407;
  assign n12409 = pi17 ? n11568 : n12408;
  assign n12410 = pi16 ? n439 : n12409;
  assign n12411 = pi21 ? n37 : n522;
  assign n12412 = pi20 ? n37 : n12411;
  assign n12413 = pi19 ? n37 : n12412;
  assign n12414 = pi18 ? n37 : n12413;
  assign n12415 = pi20 ? n37 : n5733;
  assign n12416 = pi19 ? n12415 : n37;
  assign n12417 = pi21 ? n1056 : n12404;
  assign n12418 = pi20 ? n12417 : n32;
  assign n12419 = pi19 ? n12418 : n32;
  assign n12420 = pi18 ? n12416 : n12419;
  assign n12421 = pi17 ? n12414 : n12420;
  assign n12422 = pi16 ? n439 : n12421;
  assign n12423 = pi21 ? n335 : n12404;
  assign n12424 = pi20 ? n12423 : n32;
  assign n12425 = pi19 ? n12424 : n32;
  assign n12426 = pi18 ? n37 : n12425;
  assign n12427 = pi17 ? n37 : n12426;
  assign n12428 = pi16 ? n439 : n12427;
  assign n12429 = pi15 ? n12422 : n12428;
  assign n12430 = pi14 ? n12410 : n12429;
  assign n12431 = pi13 ? n12403 : n12430;
  assign n12432 = pi21 ? n335 : n7034;
  assign n12433 = pi20 ? n12432 : n32;
  assign n12434 = pi19 ? n12433 : n32;
  assign n12435 = pi18 ? n11598 : n12434;
  assign n12436 = pi17 ? n37 : n12435;
  assign n12437 = pi16 ? n439 : n12436;
  assign n12438 = pi15 ? n12437 : n12047;
  assign n12439 = pi14 ? n12438 : n12047;
  assign n12440 = pi20 ? n37 : n7646;
  assign n12441 = pi19 ? n37 : n12440;
  assign n12442 = pi21 ? n569 : n4101;
  assign n12443 = pi20 ? n12442 : n32;
  assign n12444 = pi19 ? n12443 : n32;
  assign n12445 = pi18 ? n12441 : n12444;
  assign n12446 = pi17 ? n37 : n12445;
  assign n12447 = pi16 ? n439 : n12446;
  assign n12448 = pi21 ? n569 : n6416;
  assign n12449 = pi20 ? n12448 : n32;
  assign n12450 = pi19 ? n12449 : n32;
  assign n12451 = pi18 ? n6374 : n12450;
  assign n12452 = pi17 ? n37 : n12451;
  assign n12453 = pi16 ? n439 : n12452;
  assign n12454 = pi15 ? n12447 : n12453;
  assign n12455 = pi21 ? n2091 : n5829;
  assign n12456 = pi20 ? n12455 : n32;
  assign n12457 = pi19 ? n12456 : n32;
  assign n12458 = pi18 ? n11654 : n12457;
  assign n12459 = pi17 ? n37 : n12458;
  assign n12460 = pi16 ? n439 : n12459;
  assign n12461 = pi18 ? n37 : n12457;
  assign n12462 = pi17 ? n37 : n12461;
  assign n12463 = pi16 ? n439 : n12462;
  assign n12464 = pi15 ? n12460 : n12463;
  assign n12465 = pi14 ? n12454 : n12464;
  assign n12466 = pi13 ? n12439 : n12465;
  assign n12467 = pi12 ? n12431 : n12466;
  assign n12468 = pi11 ? n12369 : n12467;
  assign n12469 = pi21 ? n2091 : n3397;
  assign n12470 = pi20 ? n12469 : n32;
  assign n12471 = pi19 ? n12470 : n32;
  assign n12472 = pi18 ? n37 : n12471;
  assign n12473 = pi17 ? n37 : n12472;
  assign n12474 = pi16 ? n439 : n12473;
  assign n12475 = pi21 ? n1920 : n37;
  assign n12476 = pi20 ? n37 : n12475;
  assign n12477 = pi21 ? n560 : n37;
  assign n12478 = pi20 ? n37 : n12477;
  assign n12479 = pi19 ? n12476 : n12478;
  assign n12480 = pi18 ? n12479 : n12471;
  assign n12481 = pi17 ? n37 : n12480;
  assign n12482 = pi16 ? n439 : n12481;
  assign n12483 = pi15 ? n12474 : n12482;
  assign n12484 = pi15 ? n9883 : n12100;
  assign n12485 = pi14 ? n12483 : n12484;
  assign n12486 = pi21 ? n11208 : n2700;
  assign n12487 = pi20 ? n12486 : n32;
  assign n12488 = pi19 ? n12487 : n32;
  assign n12489 = pi18 ? n37 : n12488;
  assign n12490 = pi17 ? n37 : n12489;
  assign n12491 = pi16 ? n439 : n12490;
  assign n12492 = pi21 ? n2721 : n1009;
  assign n12493 = pi20 ? n12492 : n32;
  assign n12494 = pi19 ? n12493 : n32;
  assign n12495 = pi18 ? n37 : n12494;
  assign n12496 = pi17 ? n37 : n12495;
  assign n12497 = pi16 ? n439 : n12496;
  assign n12498 = pi15 ? n12491 : n12497;
  assign n12499 = pi14 ? n12107 : n12498;
  assign n12500 = pi13 ? n12485 : n12499;
  assign n12501 = pi21 ? n6461 : n32;
  assign n12502 = pi20 ? n12501 : n32;
  assign n12503 = pi19 ? n12502 : n32;
  assign n12504 = pi18 ? n99 : n12503;
  assign n12505 = pi17 ? n99 : n12504;
  assign n12506 = pi16 ? n201 : n12505;
  assign n12507 = pi15 ? n12506 : n12126;
  assign n12508 = pi21 ? n3562 : n32;
  assign n12509 = pi20 ? n12508 : n32;
  assign n12510 = pi19 ? n12509 : n32;
  assign n12511 = pi18 ? n99 : n12510;
  assign n12512 = pi17 ? n99 : n12511;
  assign n12513 = pi16 ? n744 : n12512;
  assign n12514 = pi21 ? n3445 : n32;
  assign n12515 = pi20 ? n12514 : n32;
  assign n12516 = pi19 ? n12515 : n32;
  assign n12517 = pi18 ? n5093 : n12516;
  assign n12518 = pi17 ? n99 : n12517;
  assign n12519 = pi16 ? n744 : n12518;
  assign n12520 = pi15 ? n12513 : n12519;
  assign n12521 = pi14 ? n12507 : n12520;
  assign n12522 = pi18 ? n11708 : n11697;
  assign n12523 = pi17 ? n99 : n12522;
  assign n12524 = pi16 ? n744 : n12523;
  assign n12525 = pi20 ? n157 : n7818;
  assign n12526 = pi19 ? n157 : n12525;
  assign n12527 = pi18 ? n12526 : n11697;
  assign n12528 = pi17 ? n157 : n12527;
  assign n12529 = pi16 ? n7793 : n12528;
  assign n12530 = pi15 ? n12524 : n12529;
  assign n12531 = pi21 ? n7128 : n157;
  assign n12532 = pi20 ? n32 : n12531;
  assign n12533 = pi19 ? n32 : n12532;
  assign n12534 = pi18 ? n12533 : n157;
  assign n12535 = pi17 ? n32 : n12534;
  assign n12536 = pi18 ? n157 : n6937;
  assign n12537 = pi17 ? n157 : n12536;
  assign n12538 = pi16 ? n12535 : n12537;
  assign n12539 = pi18 ? n99 : n6937;
  assign n12540 = pi17 ? n99 : n12539;
  assign n12541 = pi16 ? n744 : n12540;
  assign n12542 = pi15 ? n12538 : n12541;
  assign n12543 = pi14 ? n12530 : n12542;
  assign n12544 = pi13 ? n12521 : n12543;
  assign n12545 = pi12 ? n12500 : n12544;
  assign n12546 = pi18 ? n99 : n5669;
  assign n12547 = pi17 ? n99 : n12546;
  assign n12548 = pi16 ? n744 : n12547;
  assign n12549 = pi18 ? n139 : n5669;
  assign n12550 = pi17 ? n139 : n12549;
  assign n12551 = pi16 ? n915 : n12550;
  assign n12552 = pi15 ? n12548 : n12551;
  assign n12553 = pi18 ? n139 : n4010;
  assign n12554 = pi17 ? n139 : n12553;
  assign n12555 = pi16 ? n915 : n12554;
  assign n12556 = pi19 ? n139 : n1017;
  assign n12557 = pi18 ? n12556 : n4010;
  assign n12558 = pi17 ? n139 : n12557;
  assign n12559 = pi16 ? n915 : n12558;
  assign n12560 = pi15 ? n12555 : n12559;
  assign n12561 = pi14 ? n12552 : n12560;
  assign n12562 = pi21 ? n316 : n4429;
  assign n12563 = pi20 ? n12562 : n316;
  assign n12564 = pi19 ? n12563 : n316;
  assign n12565 = pi18 ? n12564 : n316;
  assign n12566 = pi18 ? n316 : n4010;
  assign n12567 = pi17 ? n12565 : n12566;
  assign n12568 = pi16 ? n7883 : n12567;
  assign n12569 = pi17 ? n316 : n12566;
  assign n12570 = pi16 ? n8445 : n12569;
  assign n12571 = pi22 ? n7145 : n316;
  assign n12572 = pi21 ? n12571 : n316;
  assign n12573 = pi20 ? n32 : n12572;
  assign n12574 = pi19 ? n32 : n12573;
  assign n12575 = pi18 ? n12574 : n316;
  assign n12576 = pi17 ? n32 : n12575;
  assign n12577 = pi21 ? n316 : n1785;
  assign n12578 = pi20 ? n12577 : n316;
  assign n12579 = pi19 ? n12578 : n316;
  assign n12580 = pi18 ? n12579 : n316;
  assign n12581 = pi17 ? n12580 : n11773;
  assign n12582 = pi16 ? n12576 : n12581;
  assign n12583 = pi15 ? n12570 : n12582;
  assign n12584 = pi14 ? n12568 : n12583;
  assign n12585 = pi13 ? n12561 : n12584;
  assign n12586 = pi18 ? n9111 : n3212;
  assign n12587 = pi17 ? n139 : n12586;
  assign n12588 = pi16 ? n1575 : n12587;
  assign n12589 = pi20 ? n139 : n1026;
  assign n12590 = pi19 ? n139 : n12589;
  assign n12591 = pi18 ? n12590 : n3342;
  assign n12592 = pi17 ? n139 : n12591;
  assign n12593 = pi16 ? n1575 : n12592;
  assign n12594 = pi15 ? n12588 : n12593;
  assign n12595 = pi22 ? n7959 : n37;
  assign n12596 = pi21 ? n12595 : n204;
  assign n12597 = pi20 ? n32 : n12596;
  assign n12598 = pi19 ? n32 : n12597;
  assign n12599 = pi18 ? n12598 : n204;
  assign n12600 = pi17 ? n32 : n12599;
  assign n12601 = pi21 ? n1046 : n569;
  assign n12602 = pi20 ? n12601 : n204;
  assign n12603 = pi19 ? n12602 : n204;
  assign n12604 = pi18 ? n12603 : n204;
  assign n12605 = pi18 ? n204 : n2640;
  assign n12606 = pi17 ? n12604 : n12605;
  assign n12607 = pi16 ? n12600 : n12606;
  assign n12608 = pi22 ? n7937 : n37;
  assign n12609 = pi21 ? n12608 : n204;
  assign n12610 = pi20 ? n32 : n12609;
  assign n12611 = pi19 ? n32 : n12610;
  assign n12612 = pi18 ? n12611 : n204;
  assign n12613 = pi17 ? n32 : n12612;
  assign n12614 = pi22 ? n335 : n4079;
  assign n12615 = pi21 ? n204 : n12614;
  assign n12616 = pi20 ? n204 : n12615;
  assign n12617 = pi19 ? n204 : n12616;
  assign n12618 = pi18 ? n12617 : n2640;
  assign n12619 = pi17 ? n11817 : n12618;
  assign n12620 = pi16 ? n12613 : n12619;
  assign n12621 = pi15 ? n12607 : n12620;
  assign n12622 = pi14 ? n12594 : n12621;
  assign n12623 = pi21 ? n12608 : n335;
  assign n12624 = pi20 ? n32 : n12623;
  assign n12625 = pi19 ? n32 : n12624;
  assign n12626 = pi18 ? n12625 : n335;
  assign n12627 = pi17 ? n32 : n12626;
  assign n12628 = pi20 ? n649 : n335;
  assign n12629 = pi19 ? n12628 : n335;
  assign n12630 = pi18 ? n12629 : n335;
  assign n12631 = pi19 ? n335 : n8914;
  assign n12632 = pi18 ? n12631 : n2655;
  assign n12633 = pi17 ? n12630 : n12632;
  assign n12634 = pi16 ? n12627 : n12633;
  assign n12635 = pi22 ? n233 : n6365;
  assign n12636 = pi21 ? n335 : n12635;
  assign n12637 = pi20 ? n335 : n12636;
  assign n12638 = pi19 ? n335 : n12637;
  assign n12639 = pi18 ? n12638 : n1824;
  assign n12640 = pi17 ? n335 : n12639;
  assign n12641 = pi16 ? n7943 : n12640;
  assign n12642 = pi15 ? n12634 : n12641;
  assign n12643 = pi22 ? n5996 : n99;
  assign n12644 = pi21 ? n12643 : n335;
  assign n12645 = pi20 ? n32 : n12644;
  assign n12646 = pi19 ? n32 : n12645;
  assign n12647 = pi18 ? n12646 : n335;
  assign n12648 = pi17 ? n32 : n12647;
  assign n12649 = pi18 ? n12638 : n32;
  assign n12650 = pi17 ? n335 : n12649;
  assign n12651 = pi16 ? n12648 : n12650;
  assign n12652 = pi23 ? n961 : n335;
  assign n12653 = pi22 ? n12652 : n335;
  assign n12654 = pi21 ? n12653 : n335;
  assign n12655 = pi20 ? n32 : n12654;
  assign n12656 = pi19 ? n32 : n12655;
  assign n12657 = pi18 ? n12656 : n335;
  assign n12658 = pi17 ? n32 : n12657;
  assign n12659 = pi22 ? n233 : n1070;
  assign n12660 = pi21 ? n335 : n12659;
  assign n12661 = pi20 ? n335 : n12660;
  assign n12662 = pi19 ? n335 : n12661;
  assign n12663 = pi18 ? n12662 : n32;
  assign n12664 = pi17 ? n335 : n12663;
  assign n12665 = pi16 ? n12658 : n12664;
  assign n12666 = pi15 ? n12651 : n12665;
  assign n12667 = pi14 ? n12642 : n12666;
  assign n12668 = pi13 ? n12622 : n12667;
  assign n12669 = pi12 ? n12585 : n12668;
  assign n12670 = pi11 ? n12545 : n12669;
  assign n12671 = pi10 ? n12468 : n12670;
  assign n12672 = pi09 ? n12236 : n12671;
  assign n12673 = pi15 ? n32 : n12223;
  assign n12674 = pi16 ? n9232 : n12220;
  assign n12675 = pi16 ? n2461 : n12229;
  assign n12676 = pi15 ? n12674 : n12675;
  assign n12677 = pi14 ? n12673 : n12676;
  assign n12678 = pi13 ? n32 : n12677;
  assign n12679 = pi12 ? n32 : n12678;
  assign n12680 = pi11 ? n32 : n12679;
  assign n12681 = pi10 ? n32 : n12680;
  assign n12682 = pi16 ? n10154 : n12241;
  assign n12683 = pi16 ? n11011 : n12248;
  assign n12684 = pi15 ? n12682 : n12683;
  assign n12685 = pi16 ? n11885 : n11389;
  assign n12686 = pi20 ? n32 : n1114;
  assign n12687 = pi19 ? n32 : n12686;
  assign n12688 = pi18 ? n12687 : n37;
  assign n12689 = pi17 ? n32 : n12688;
  assign n12690 = pi16 ? n12689 : n12256;
  assign n12691 = pi15 ? n12685 : n12690;
  assign n12692 = pi14 ? n12684 : n12691;
  assign n12693 = pi21 ? n165 : n5875;
  assign n12694 = pi20 ? n99 : n12693;
  assign n12695 = pi21 ? n168 : n164;
  assign n12696 = pi20 ? n12695 : n10526;
  assign n12697 = pi19 ? n12694 : n12696;
  assign n12698 = pi18 ? n719 : n12697;
  assign n12699 = pi17 ? n32 : n12698;
  assign n12700 = pi21 ? n5875 : n168;
  assign n12701 = pi21 ? n164 : n158;
  assign n12702 = pi20 ? n12700 : n12701;
  assign n12703 = pi22 ? n157 : n893;
  assign n12704 = pi21 ? n165 : n12703;
  assign n12705 = pi22 ? n99 : n889;
  assign n12706 = pi21 ? n12705 : n3013;
  assign n12707 = pi20 ? n12704 : n12706;
  assign n12708 = pi19 ? n12702 : n12707;
  assign n12709 = pi22 ? n158 : n893;
  assign n12710 = pi21 ? n164 : n12709;
  assign n12711 = pi20 ? n12706 : n12710;
  assign n12712 = pi21 ? n12705 : n5875;
  assign n12713 = pi22 ? n158 : n889;
  assign n12714 = pi21 ? n12713 : n5875;
  assign n12715 = pi20 ? n12712 : n12714;
  assign n12716 = pi19 ? n12711 : n12715;
  assign n12717 = pi18 ? n12708 : n12716;
  assign n12718 = pi21 ? n12713 : n12703;
  assign n12719 = pi20 ? n12718 : n3011;
  assign n12720 = pi22 ? n893 : n164;
  assign n12721 = pi21 ? n5875 : n12720;
  assign n12722 = pi20 ? n12721 : n5886;
  assign n12723 = pi19 ? n12719 : n12722;
  assign n12724 = pi22 ? n158 : n1378;
  assign n12725 = pi21 ? n5875 : n12724;
  assign n12726 = pi20 ? n12725 : n32;
  assign n12727 = pi19 ? n12726 : n32;
  assign n12728 = pi18 ? n12723 : n12727;
  assign n12729 = pi17 ? n12717 : n12728;
  assign n12730 = pi16 ? n12699 : n12729;
  assign n12731 = pi22 ? n157 : n1378;
  assign n12732 = pi21 ? n157 : n12731;
  assign n12733 = pi20 ? n12732 : n32;
  assign n12734 = pi19 ? n12733 : n32;
  assign n12735 = pi18 ? n157 : n12734;
  assign n12736 = pi17 ? n157 : n12735;
  assign n12737 = pi16 ? n12302 : n12736;
  assign n12738 = pi15 ? n12730 : n12737;
  assign n12739 = pi14 ? n12274 : n12738;
  assign n12740 = pi13 ? n12692 : n12739;
  assign n12741 = pi21 ? n99 : n5482;
  assign n12742 = pi20 ? n12741 : n32;
  assign n12743 = pi19 ? n12742 : n32;
  assign n12744 = pi18 ? n99 : n12743;
  assign n12745 = pi17 ? n99 : n12744;
  assign n12746 = pi16 ? n801 : n12745;
  assign n12747 = pi22 ? n99 : n2564;
  assign n12748 = pi21 ? n99 : n12747;
  assign n12749 = pi20 ? n12748 : n32;
  assign n12750 = pi19 ? n12749 : n32;
  assign n12751 = pi18 ? n99 : n12750;
  assign n12752 = pi17 ? n99 : n12751;
  assign n12753 = pi16 ? n801 : n12752;
  assign n12754 = pi22 ? n745 : n2564;
  assign n12755 = pi21 ? n99 : n12754;
  assign n12756 = pi20 ? n12755 : n32;
  assign n12757 = pi19 ? n12756 : n32;
  assign n12758 = pi18 ? n99 : n12757;
  assign n12759 = pi17 ? n99 : n12758;
  assign n12760 = pi16 ? n721 : n12759;
  assign n12761 = pi15 ? n12753 : n12760;
  assign n12762 = pi14 ? n12746 : n12761;
  assign n12763 = pi22 ? n1656 : n664;
  assign n12764 = pi21 ? n99 : n12763;
  assign n12765 = pi20 ? n12764 : n32;
  assign n12766 = pi19 ? n12765 : n32;
  assign n12767 = pi18 ? n99 : n12766;
  assign n12768 = pi17 ? n99 : n12767;
  assign n12769 = pi16 ? n721 : n12768;
  assign n12770 = pi22 ? n861 : n664;
  assign n12771 = pi21 ? n139 : n12770;
  assign n12772 = pi20 ? n12771 : n32;
  assign n12773 = pi19 ? n12772 : n32;
  assign n12774 = pi18 ? n139 : n12773;
  assign n12775 = pi17 ? n139 : n12774;
  assign n12776 = pi16 ? n2291 : n12775;
  assign n12777 = pi15 ? n12769 : n12776;
  assign n12778 = pi22 ? n1043 : n390;
  assign n12779 = pi21 ? n3258 : n12778;
  assign n12780 = pi20 ? n9354 : n12779;
  assign n12781 = pi19 ? n37 : n12780;
  assign n12782 = pi22 ? n1043 : n348;
  assign n12783 = pi21 ? n3258 : n12782;
  assign n12784 = pi20 ? n12338 : n12783;
  assign n12785 = pi19 ? n12337 : n12784;
  assign n12786 = pi18 ? n12781 : n12785;
  assign n12787 = pi21 ? n4056 : n4014;
  assign n12788 = pi20 ? n316 : n12787;
  assign n12789 = pi19 ? n12788 : n12346;
  assign n12790 = pi18 ? n12789 : n12349;
  assign n12791 = pi17 ? n12786 : n12790;
  assign n12792 = pi16 ? n439 : n12791;
  assign n12793 = pi15 ? n12792 : n12365;
  assign n12794 = pi14 ? n12777 : n12793;
  assign n12795 = pi13 ? n12762 : n12794;
  assign n12796 = pi12 ? n12740 : n12795;
  assign n12797 = pi21 ? n37 : n5746;
  assign n12798 = pi20 ? n12797 : n32;
  assign n12799 = pi19 ? n12798 : n32;
  assign n12800 = pi18 ? n37 : n12799;
  assign n12801 = pi17 ? n37 : n12800;
  assign n12802 = pi16 ? n439 : n12801;
  assign n12803 = pi15 ? n12380 : n12802;
  assign n12804 = pi14 ? n12803 : n12402;
  assign n12805 = pi20 ? n6947 : n12411;
  assign n12806 = pi19 ? n37 : n12805;
  assign n12807 = pi18 ? n37 : n12806;
  assign n12808 = pi21 ? n506 : n37;
  assign n12809 = pi20 ? n37 : n12808;
  assign n12810 = pi19 ? n12415 : n12809;
  assign n12811 = pi18 ? n12810 : n12419;
  assign n12812 = pi17 ? n12807 : n12811;
  assign n12813 = pi16 ? n439 : n12812;
  assign n12814 = pi15 ? n12813 : n12428;
  assign n12815 = pi14 ? n12410 : n12814;
  assign n12816 = pi13 ? n12804 : n12815;
  assign n12817 = pi21 ? n569 : n650;
  assign n12818 = pi20 ? n12817 : n32;
  assign n12819 = pi19 ? n12818 : n32;
  assign n12820 = pi18 ? n37 : n12819;
  assign n12821 = pi17 ? n37 : n12820;
  assign n12822 = pi16 ? n439 : n12821;
  assign n12823 = pi15 ? n12047 : n12822;
  assign n12824 = pi14 ? n12438 : n12823;
  assign n12825 = pi22 ? n2121 : n32;
  assign n12826 = pi21 ? n569 : n12825;
  assign n12827 = pi20 ? n12826 : n32;
  assign n12828 = pi19 ? n12827 : n32;
  assign n12829 = pi18 ? n12441 : n12828;
  assign n12830 = pi17 ? n37 : n12829;
  assign n12831 = pi16 ? n439 : n12830;
  assign n12832 = pi21 ? n569 : n7041;
  assign n12833 = pi20 ? n12832 : n32;
  assign n12834 = pi19 ? n12833 : n32;
  assign n12835 = pi18 ? n6374 : n12834;
  assign n12836 = pi17 ? n37 : n12835;
  assign n12837 = pi16 ? n439 : n12836;
  assign n12838 = pi15 ? n12831 : n12837;
  assign n12839 = pi21 ? n2091 : n760;
  assign n12840 = pi20 ? n12839 : n32;
  assign n12841 = pi19 ? n12840 : n32;
  assign n12842 = pi18 ? n11654 : n12841;
  assign n12843 = pi17 ? n37 : n12842;
  assign n12844 = pi16 ? n439 : n12843;
  assign n12845 = pi21 ? n2091 : n7048;
  assign n12846 = pi20 ? n12845 : n32;
  assign n12847 = pi19 ? n12846 : n32;
  assign n12848 = pi18 ? n37 : n12847;
  assign n12849 = pi17 ? n37 : n12848;
  assign n12850 = pi16 ? n439 : n12849;
  assign n12851 = pi15 ? n12844 : n12850;
  assign n12852 = pi14 ? n12838 : n12851;
  assign n12853 = pi13 ? n12824 : n12852;
  assign n12854 = pi12 ? n12816 : n12853;
  assign n12855 = pi11 ? n12796 : n12854;
  assign n12856 = pi21 ? n2091 : n3339;
  assign n12857 = pi20 ? n12856 : n32;
  assign n12858 = pi19 ? n12857 : n32;
  assign n12859 = pi18 ? n37 : n12858;
  assign n12860 = pi17 ? n37 : n12859;
  assign n12861 = pi16 ? n439 : n12860;
  assign n12862 = pi18 ? n12479 : n12858;
  assign n12863 = pi17 ? n37 : n12862;
  assign n12864 = pi16 ? n439 : n12863;
  assign n12865 = pi15 ? n12861 : n12864;
  assign n12866 = pi21 ? n2091 : n2578;
  assign n12867 = pi20 ? n12866 : n32;
  assign n12868 = pi19 ? n12867 : n32;
  assign n12869 = pi18 ? n37 : n12868;
  assign n12870 = pi17 ? n37 : n12869;
  assign n12871 = pi16 ? n439 : n12870;
  assign n12872 = pi21 ? n2106 : n2637;
  assign n12873 = pi20 ? n12872 : n32;
  assign n12874 = pi19 ? n12873 : n32;
  assign n12875 = pi18 ? n37 : n12874;
  assign n12876 = pi17 ? n37 : n12875;
  assign n12877 = pi16 ? n439 : n12876;
  assign n12878 = pi15 ? n12871 : n12877;
  assign n12879 = pi14 ? n12865 : n12878;
  assign n12880 = pi22 ? n7024 : n685;
  assign n12881 = pi21 ? n12880 : n2637;
  assign n12882 = pi20 ? n12881 : n32;
  assign n12883 = pi19 ? n12882 : n32;
  assign n12884 = pi18 ? n37 : n12883;
  assign n12885 = pi17 ? n37 : n12884;
  assign n12886 = pi16 ? n439 : n12885;
  assign n12887 = pi21 ? n2721 : n2637;
  assign n12888 = pi20 ? n12887 : n32;
  assign n12889 = pi19 ? n12888 : n32;
  assign n12890 = pi18 ? n37 : n12889;
  assign n12891 = pi17 ? n37 : n12890;
  assign n12892 = pi16 ? n439 : n12891;
  assign n12893 = pi15 ? n12886 : n12892;
  assign n12894 = pi21 ? n11208 : n2637;
  assign n12895 = pi20 ? n12894 : n32;
  assign n12896 = pi19 ? n12895 : n32;
  assign n12897 = pi18 ? n37 : n12896;
  assign n12898 = pi17 ? n37 : n12897;
  assign n12899 = pi16 ? n439 : n12898;
  assign n12900 = pi21 ? n2721 : n928;
  assign n12901 = pi20 ? n12900 : n32;
  assign n12902 = pi19 ? n12901 : n32;
  assign n12903 = pi18 ? n37 : n12902;
  assign n12904 = pi17 ? n37 : n12903;
  assign n12905 = pi16 ? n439 : n12904;
  assign n12906 = pi15 ? n12899 : n12905;
  assign n12907 = pi14 ? n12893 : n12906;
  assign n12908 = pi13 ? n12879 : n12907;
  assign n12909 = pi21 ? n6461 : n2700;
  assign n12910 = pi20 ? n12909 : n32;
  assign n12911 = pi19 ? n12910 : n32;
  assign n12912 = pi18 ? n99 : n12911;
  assign n12913 = pi17 ? n99 : n12912;
  assign n12914 = pi16 ? n201 : n12913;
  assign n12915 = pi18 ? n99 : n7409;
  assign n12916 = pi17 ? n99 : n12915;
  assign n12917 = pi16 ? n721 : n12916;
  assign n12918 = pi15 ? n12914 : n12917;
  assign n12919 = pi21 ? n3562 : n1009;
  assign n12920 = pi20 ? n12919 : n32;
  assign n12921 = pi19 ? n12920 : n32;
  assign n12922 = pi18 ? n99 : n12921;
  assign n12923 = pi17 ? n99 : n12922;
  assign n12924 = pi16 ? n721 : n12923;
  assign n12925 = pi21 ? n3445 : n1009;
  assign n12926 = pi20 ? n12925 : n32;
  assign n12927 = pi19 ? n12926 : n32;
  assign n12928 = pi18 ? n5093 : n12927;
  assign n12929 = pi17 ? n99 : n12928;
  assign n12930 = pi16 ? n721 : n12929;
  assign n12931 = pi15 ? n12924 : n12930;
  assign n12932 = pi14 ? n12918 : n12931;
  assign n12933 = pi18 ? n11708 : n12130;
  assign n12934 = pi17 ? n99 : n12933;
  assign n12935 = pi16 ? n721 : n12934;
  assign n12936 = pi18 ? n12526 : n12130;
  assign n12937 = pi17 ? n157 : n12936;
  assign n12938 = pi16 ? n5910 : n12937;
  assign n12939 = pi15 ? n12935 : n12938;
  assign n12940 = pi16 ? n721 : n12540;
  assign n12941 = pi15 ? n12538 : n12940;
  assign n12942 = pi14 ? n12939 : n12941;
  assign n12943 = pi13 ? n12932 : n12942;
  assign n12944 = pi12 ? n12908 : n12943;
  assign n12945 = pi16 ? n721 : n12547;
  assign n12946 = pi16 ? n2291 : n12550;
  assign n12947 = pi15 ? n12945 : n12946;
  assign n12948 = pi16 ? n2291 : n12554;
  assign n12949 = pi16 ? n2291 : n12558;
  assign n12950 = pi15 ? n12948 : n12949;
  assign n12951 = pi14 ? n12947 : n12950;
  assign n12952 = pi16 ? n7883 : n12569;
  assign n12953 = pi16 ? n11772 : n12581;
  assign n12954 = pi15 ? n12952 : n12953;
  assign n12955 = pi14 ? n12568 : n12954;
  assign n12956 = pi13 ? n12951 : n12955;
  assign n12957 = pi16 ? n331 : n12587;
  assign n12958 = pi21 ? n7244 : n32;
  assign n12959 = pi20 ? n12958 : n32;
  assign n12960 = pi19 ? n12959 : n32;
  assign n12961 = pi18 ? n12590 : n12960;
  assign n12962 = pi17 ? n139 : n12961;
  assign n12963 = pi16 ? n331 : n12962;
  assign n12964 = pi15 ? n12957 : n12963;
  assign n12965 = pi22 ? n2390 : n37;
  assign n12966 = pi21 ? n12965 : n204;
  assign n12967 = pi20 ? n32 : n12966;
  assign n12968 = pi19 ? n32 : n12967;
  assign n12969 = pi18 ? n12968 : n204;
  assign n12970 = pi17 ? n32 : n12969;
  assign n12971 = pi18 ? n204 : n5832;
  assign n12972 = pi17 ? n12604 : n12971;
  assign n12973 = pi16 ? n12970 : n12972;
  assign n12974 = pi22 ? n335 : n4883;
  assign n12975 = pi21 ? n204 : n12974;
  assign n12976 = pi20 ? n204 : n12975;
  assign n12977 = pi19 ? n204 : n12976;
  assign n12978 = pi18 ? n12977 : n5832;
  assign n12979 = pi17 ? n11817 : n12978;
  assign n12980 = pi16 ? n12613 : n12979;
  assign n12981 = pi15 ? n12973 : n12980;
  assign n12982 = pi14 ? n12964 : n12981;
  assign n12983 = pi22 ? n233 : n4925;
  assign n12984 = pi21 ? n335 : n12983;
  assign n12985 = pi20 ? n335 : n12984;
  assign n12986 = pi19 ? n335 : n12985;
  assign n12987 = pi18 ? n12986 : n1824;
  assign n12988 = pi17 ? n335 : n12987;
  assign n12989 = pi16 ? n10980 : n12988;
  assign n12990 = pi15 ? n12634 : n12989;
  assign n12991 = pi18 ? n12986 : n32;
  assign n12992 = pi17 ? n335 : n12991;
  assign n12993 = pi16 ? n12648 : n12992;
  assign n12994 = pi22 ? n233 : n2121;
  assign n12995 = pi21 ? n335 : n12994;
  assign n12996 = pi20 ? n335 : n12995;
  assign n12997 = pi19 ? n335 : n12996;
  assign n12998 = pi18 ? n12997 : n32;
  assign n12999 = pi17 ? n335 : n12998;
  assign n13000 = pi16 ? n12658 : n12999;
  assign n13001 = pi15 ? n12993 : n13000;
  assign n13002 = pi14 ? n12990 : n13001;
  assign n13003 = pi13 ? n12982 : n13002;
  assign n13004 = pi12 ? n12956 : n13003;
  assign n13005 = pi11 ? n12944 : n13004;
  assign n13006 = pi10 ? n12855 : n13005;
  assign n13007 = pi09 ? n12681 : n13006;
  assign n13008 = pi08 ? n12672 : n13007;
  assign n13009 = pi07 ? n12216 : n13008;
  assign n13010 = pi20 ? n1619 : n32;
  assign n13011 = pi19 ? n13010 : n32;
  assign n13012 = pi18 ? n37 : n13011;
  assign n13013 = pi17 ? n37 : n13012;
  assign n13014 = pi16 ? n1130 : n13013;
  assign n13015 = pi15 ? n32 : n13014;
  assign n13016 = pi16 ? n9232 : n13013;
  assign n13017 = pi16 ? n2461 : n13013;
  assign n13018 = pi15 ? n13016 : n13017;
  assign n13019 = pi14 ? n13015 : n13018;
  assign n13020 = pi13 ? n32 : n13019;
  assign n13021 = pi12 ? n32 : n13020;
  assign n13022 = pi11 ? n32 : n13021;
  assign n13023 = pi10 ? n32 : n13022;
  assign n13024 = pi22 ? n37 : n3831;
  assign n13025 = pi21 ? n37 : n13024;
  assign n13026 = pi20 ? n13025 : n32;
  assign n13027 = pi19 ? n13026 : n32;
  assign n13028 = pi18 ? n37 : n13027;
  assign n13029 = pi17 ? n37 : n13028;
  assign n13030 = pi16 ? n10154 : n13029;
  assign n13031 = pi22 ? n37 : n9628;
  assign n13032 = pi21 ? n37 : n13031;
  assign n13033 = pi20 ? n13032 : n32;
  assign n13034 = pi19 ? n13033 : n32;
  assign n13035 = pi18 ? n37 : n13034;
  assign n13036 = pi17 ? n37 : n13035;
  assign n13037 = pi16 ? n11011 : n13036;
  assign n13038 = pi15 ? n13030 : n13037;
  assign n13039 = pi22 ? n37 : n140;
  assign n13040 = pi21 ? n37 : n13039;
  assign n13041 = pi20 ? n13040 : n32;
  assign n13042 = pi19 ? n13041 : n32;
  assign n13043 = pi18 ? n37 : n13042;
  assign n13044 = pi17 ? n37 : n13043;
  assign n13045 = pi16 ? n11885 : n13044;
  assign n13046 = pi16 ? n12689 : n13044;
  assign n13047 = pi15 ? n13045 : n13046;
  assign n13048 = pi14 ? n13038 : n13047;
  assign n13049 = pi22 ? n37 : n1344;
  assign n13050 = pi21 ? n37 : n13049;
  assign n13051 = pi20 ? n13050 : n32;
  assign n13052 = pi19 ? n13051 : n32;
  assign n13053 = pi18 ? n37 : n13052;
  assign n13054 = pi17 ? n37 : n13053;
  assign n13055 = pi16 ? n439 : n13054;
  assign n13056 = pi21 ? n99 : n5444;
  assign n13057 = pi20 ? n13056 : n32;
  assign n13058 = pi19 ? n13057 : n32;
  assign n13059 = pi18 ? n99 : n13058;
  assign n13060 = pi17 ? n99 : n13059;
  assign n13061 = pi16 ? n3065 : n13060;
  assign n13062 = pi15 ? n13055 : n13061;
  assign n13063 = pi21 ? n3060 : n777;
  assign n13064 = pi20 ? n32 : n13063;
  assign n13065 = pi19 ? n32 : n13064;
  assign n13066 = pi18 ? n13065 : n157;
  assign n13067 = pi17 ? n32 : n13066;
  assign n13068 = pi16 ? n13067 : n12736;
  assign n13069 = pi20 ? n2243 : n6523;
  assign n13070 = pi20 ? n6508 : n7818;
  assign n13071 = pi19 ? n13069 : n13070;
  assign n13072 = pi18 ? n12300 : n13071;
  assign n13073 = pi17 ? n32 : n13072;
  assign n13074 = pi19 ? n6531 : n157;
  assign n13075 = pi18 ? n13074 : n157;
  assign n13076 = pi17 ? n13075 : n12735;
  assign n13077 = pi16 ? n13073 : n13076;
  assign n13078 = pi15 ? n13068 : n13077;
  assign n13079 = pi14 ? n13062 : n13078;
  assign n13080 = pi13 ? n13048 : n13079;
  assign n13081 = pi16 ? n744 : n12745;
  assign n13082 = pi15 ? n12746 : n13081;
  assign n13083 = pi16 ? n744 : n12752;
  assign n13084 = pi15 ? n12753 : n13083;
  assign n13085 = pi14 ? n13082 : n13084;
  assign n13086 = pi22 ? n99 : n664;
  assign n13087 = pi21 ? n99 : n13086;
  assign n13088 = pi20 ? n13087 : n32;
  assign n13089 = pi19 ? n13088 : n32;
  assign n13090 = pi18 ? n99 : n13089;
  assign n13091 = pi17 ? n99 : n13090;
  assign n13092 = pi16 ? n721 : n13091;
  assign n13093 = pi20 ? n941 : n139;
  assign n13094 = pi20 ? n941 : n37;
  assign n13095 = pi19 ? n13093 : n13094;
  assign n13096 = pi18 ? n2364 : n13095;
  assign n13097 = pi17 ? n32 : n13096;
  assign n13098 = pi19 ? n13094 : n37;
  assign n13099 = pi18 ? n37 : n13098;
  assign n13100 = pi20 ? n139 : n941;
  assign n13101 = pi19 ? n13100 : n13094;
  assign n13102 = pi22 ? n139 : n664;
  assign n13103 = pi21 ? n139 : n13102;
  assign n13104 = pi20 ? n13103 : n32;
  assign n13105 = pi19 ? n13104 : n32;
  assign n13106 = pi18 ? n13101 : n13105;
  assign n13107 = pi17 ? n13099 : n13106;
  assign n13108 = pi16 ? n13097 : n13107;
  assign n13109 = pi15 ? n13092 : n13108;
  assign n13110 = pi19 ? n37 : n8743;
  assign n13111 = pi20 ? n398 : n32;
  assign n13112 = pi19 ? n13111 : n32;
  assign n13113 = pi18 ? n13110 : n13112;
  assign n13114 = pi17 ? n37 : n13113;
  assign n13115 = pi16 ? n439 : n13114;
  assign n13116 = pi21 ? n1696 : n3668;
  assign n13117 = pi19 ? n9824 : n13116;
  assign n13118 = pi21 ? n37 : n1531;
  assign n13119 = pi21 ? n1696 : n1211;
  assign n13120 = pi20 ? n13118 : n13119;
  assign n13121 = pi21 ? n37 : n1211;
  assign n13122 = pi19 ? n13120 : n13121;
  assign n13123 = pi18 ? n13117 : n13122;
  assign n13124 = pi20 ? n37 : n376;
  assign n13125 = pi20 ? n37 : n1003;
  assign n13126 = pi19 ? n13124 : n13125;
  assign n13127 = pi22 ? n1784 : n396;
  assign n13128 = pi21 ? n820 : n13127;
  assign n13129 = pi20 ? n13128 : n32;
  assign n13130 = pi19 ? n13129 : n32;
  assign n13131 = pi18 ? n13126 : n13130;
  assign n13132 = pi17 ? n13123 : n13131;
  assign n13133 = pi16 ? n439 : n13132;
  assign n13134 = pi15 ? n13115 : n13133;
  assign n13135 = pi14 ? n13109 : n13134;
  assign n13136 = pi13 ? n13085 : n13135;
  assign n13137 = pi12 ? n13080 : n13136;
  assign n13138 = pi21 ? n375 : n3668;
  assign n13139 = pi21 ? n820 : n3668;
  assign n13140 = pi20 ? n13138 : n13139;
  assign n13141 = pi19 ? n37 : n13140;
  assign n13142 = pi20 ? n13121 : n1694;
  assign n13143 = pi21 ? n37 : n1043;
  assign n13144 = pi20 ? n13143 : n13121;
  assign n13145 = pi19 ? n13142 : n13144;
  assign n13146 = pi18 ? n13141 : n13145;
  assign n13147 = pi21 ? n1696 : n37;
  assign n13148 = pi20 ? n37 : n13147;
  assign n13149 = pi19 ? n12370 : n13148;
  assign n13150 = pi21 ? n297 : n13127;
  assign n13151 = pi20 ? n13150 : n32;
  assign n13152 = pi19 ? n13151 : n32;
  assign n13153 = pi18 ? n13149 : n13152;
  assign n13154 = pi17 ? n13146 : n13153;
  assign n13155 = pi16 ? n439 : n13154;
  assign n13156 = pi20 ? n1003 : n3104;
  assign n13157 = pi20 ? n3104 : n3086;
  assign n13158 = pi19 ? n13156 : n13157;
  assign n13159 = pi22 ? n1038 : n317;
  assign n13160 = pi21 ? n37 : n13159;
  assign n13161 = pi20 ? n13160 : n32;
  assign n13162 = pi19 ? n13161 : n32;
  assign n13163 = pi18 ? n13158 : n13162;
  assign n13164 = pi17 ? n12372 : n13163;
  assign n13165 = pi16 ? n439 : n13164;
  assign n13166 = pi15 ? n13155 : n13165;
  assign n13167 = pi19 ? n37 : n3086;
  assign n13168 = pi20 ? n3086 : n3083;
  assign n13169 = pi19 ? n3086 : n13168;
  assign n13170 = pi18 ? n13167 : n13169;
  assign n13171 = pi20 ? n3104 : n297;
  assign n13172 = pi19 ? n13156 : n13171;
  assign n13173 = pi21 ? n297 : n318;
  assign n13174 = pi20 ? n13173 : n32;
  assign n13175 = pi19 ? n13174 : n32;
  assign n13176 = pi18 ? n13172 : n13175;
  assign n13177 = pi17 ? n13170 : n13176;
  assign n13178 = pi16 ? n439 : n13177;
  assign n13179 = pi21 ? n3668 : n37;
  assign n13180 = pi20 ? n13179 : n37;
  assign n13181 = pi19 ? n13180 : n1806;
  assign n13182 = pi18 ? n37 : n13181;
  assign n13183 = pi19 ? n3578 : n139;
  assign n13184 = pi21 ? n139 : n4736;
  assign n13185 = pi20 ? n13184 : n32;
  assign n13186 = pi19 ? n13185 : n32;
  assign n13187 = pi18 ? n13183 : n13186;
  assign n13188 = pi17 ? n13182 : n13187;
  assign n13189 = pi16 ? n439 : n13188;
  assign n13190 = pi15 ? n13178 : n13189;
  assign n13191 = pi14 ? n13166 : n13190;
  assign n13192 = pi20 ? n3086 : n139;
  assign n13193 = pi19 ? n37 : n13192;
  assign n13194 = pi18 ? n37 : n13193;
  assign n13195 = pi21 ? n139 : n4748;
  assign n13196 = pi20 ? n13195 : n32;
  assign n13197 = pi19 ? n13196 : n32;
  assign n13198 = pi18 ? n139 : n13197;
  assign n13199 = pi17 ? n13194 : n13198;
  assign n13200 = pi16 ? n439 : n13199;
  assign n13201 = pi20 ? n3074 : n3625;
  assign n13202 = pi19 ? n37 : n13201;
  assign n13203 = pi18 ? n37 : n13202;
  assign n13204 = pi20 ? n2512 : n3656;
  assign n13205 = pi19 ? n139 : n13204;
  assign n13206 = pi21 ? n1531 : n4748;
  assign n13207 = pi20 ? n13206 : n32;
  assign n13208 = pi19 ? n13207 : n32;
  assign n13209 = pi18 ? n13205 : n13208;
  assign n13210 = pi17 ? n13203 : n13209;
  assign n13211 = pi16 ? n439 : n13210;
  assign n13212 = pi15 ? n13200 : n13211;
  assign n13213 = pi21 ? n1313 : n1056;
  assign n13214 = pi21 ? n485 : n37;
  assign n13215 = pi20 ? n13213 : n13214;
  assign n13216 = pi21 ? n499 : n1046;
  assign n13217 = pi21 ? n499 : n522;
  assign n13218 = pi20 ? n13216 : n13217;
  assign n13219 = pi19 ? n13215 : n13218;
  assign n13220 = pi21 ? n1056 : n4748;
  assign n13221 = pi20 ? n13220 : n32;
  assign n13222 = pi19 ? n13221 : n32;
  assign n13223 = pi18 ? n13219 : n13222;
  assign n13224 = pi17 ? n37 : n13223;
  assign n13225 = pi16 ? n439 : n13224;
  assign n13226 = pi21 ? n583 : n567;
  assign n13227 = pi20 ? n4971 : n13226;
  assign n13228 = pi19 ? n37 : n13227;
  assign n13229 = pi18 ? n37 : n13228;
  assign n13230 = pi22 ? n583 : n448;
  assign n13231 = pi21 ? n13230 : n476;
  assign n13232 = pi21 ? n1278 : n1943;
  assign n13233 = pi20 ? n13231 : n13232;
  assign n13234 = pi21 ? n567 : n8833;
  assign n13235 = pi20 ? n1983 : n13234;
  assign n13236 = pi19 ? n13233 : n13235;
  assign n13237 = pi21 ? n1943 : n650;
  assign n13238 = pi20 ? n13237 : n32;
  assign n13239 = pi19 ? n13238 : n32;
  assign n13240 = pi18 ? n13236 : n13239;
  assign n13241 = pi17 ? n13229 : n13240;
  assign n13242 = pi16 ? n439 : n13241;
  assign n13243 = pi15 ? n13225 : n13242;
  assign n13244 = pi14 ? n13212 : n13243;
  assign n13245 = pi13 ? n13191 : n13244;
  assign n13246 = pi21 ? n1943 : n335;
  assign n13247 = pi20 ? n37 : n13246;
  assign n13248 = pi19 ? n37 : n13247;
  assign n13249 = pi18 ? n37 : n13248;
  assign n13250 = pi21 ? n2061 : n4902;
  assign n13251 = pi21 ? n4908 : n335;
  assign n13252 = pi20 ? n13250 : n13251;
  assign n13253 = pi22 ? n335 : n559;
  assign n13254 = pi21 ? n335 : n13253;
  assign n13255 = pi20 ? n13251 : n13254;
  assign n13256 = pi19 ? n13252 : n13255;
  assign n13257 = pi21 ? n335 : n650;
  assign n13258 = pi20 ? n13257 : n32;
  assign n13259 = pi19 ? n13258 : n32;
  assign n13260 = pi18 ? n13256 : n13259;
  assign n13261 = pi17 ? n13249 : n13260;
  assign n13262 = pi16 ? n439 : n13261;
  assign n13263 = pi21 ? n569 : n696;
  assign n13264 = pi20 ? n13263 : n32;
  assign n13265 = pi19 ? n13264 : n32;
  assign n13266 = pi18 ? n37 : n13265;
  assign n13267 = pi17 ? n37 : n13266;
  assign n13268 = pi16 ? n439 : n13267;
  assign n13269 = pi15 ? n13262 : n13268;
  assign n13270 = pi18 ? n6374 : n12819;
  assign n13271 = pi17 ? n37 : n13270;
  assign n13272 = pi16 ? n439 : n13271;
  assign n13273 = pi21 ? n37 : n1943;
  assign n13274 = pi20 ? n37 : n13273;
  assign n13275 = pi21 ? n569 : n2007;
  assign n13276 = pi20 ? n37 : n13275;
  assign n13277 = pi19 ? n13274 : n13276;
  assign n13278 = pi23 ? n1342 : n335;
  assign n13279 = pi22 ? n37 : n13278;
  assign n13280 = pi22 ? n233 : n688;
  assign n13281 = pi21 ? n13279 : n13280;
  assign n13282 = pi20 ? n13281 : n32;
  assign n13283 = pi19 ? n13282 : n32;
  assign n13284 = pi18 ? n13277 : n13283;
  assign n13285 = pi17 ? n37 : n13284;
  assign n13286 = pi16 ? n439 : n13285;
  assign n13287 = pi15 ? n13272 : n13286;
  assign n13288 = pi14 ? n13269 : n13287;
  assign n13289 = pi21 ? n2007 : n570;
  assign n13290 = pi20 ? n37 : n13289;
  assign n13291 = pi19 ? n13274 : n13290;
  assign n13292 = pi21 ? n569 : n4926;
  assign n13293 = pi20 ? n13292 : n32;
  assign n13294 = pi19 ? n13293 : n32;
  assign n13295 = pi18 ? n13291 : n13294;
  assign n13296 = pi17 ? n37 : n13295;
  assign n13297 = pi16 ? n439 : n13296;
  assign n13298 = pi21 ? n584 : n567;
  assign n13299 = pi20 ? n37 : n13298;
  assign n13300 = pi21 ? n2007 : n1943;
  assign n13301 = pi20 ? n2008 : n13300;
  assign n13302 = pi19 ? n13299 : n13301;
  assign n13303 = pi21 ? n569 : n7723;
  assign n13304 = pi20 ? n13303 : n32;
  assign n13305 = pi19 ? n13304 : n32;
  assign n13306 = pi18 ? n13302 : n13305;
  assign n13307 = pi17 ? n37 : n13306;
  assign n13308 = pi16 ? n439 : n13307;
  assign n13309 = pi15 ? n13297 : n13308;
  assign n13310 = pi21 ? n37 : n7334;
  assign n13311 = pi21 ? n5012 : n5015;
  assign n13312 = pi20 ? n13310 : n13311;
  assign n13313 = pi19 ? n8569 : n13312;
  assign n13314 = pi23 ? n233 : n2766;
  assign n13315 = pi22 ? n13314 : n32;
  assign n13316 = pi21 ? n3392 : n13315;
  assign n13317 = pi20 ? n13316 : n32;
  assign n13318 = pi19 ? n13317 : n32;
  assign n13319 = pi18 ? n13313 : n13318;
  assign n13320 = pi17 ? n37 : n13319;
  assign n13321 = pi16 ? n439 : n13320;
  assign n13322 = pi21 ? n2091 : n6416;
  assign n13323 = pi20 ? n13322 : n32;
  assign n13324 = pi19 ? n13323 : n32;
  assign n13325 = pi18 ? n6356 : n13324;
  assign n13326 = pi17 ? n37 : n13325;
  assign n13327 = pi16 ? n439 : n13326;
  assign n13328 = pi15 ? n13321 : n13327;
  assign n13329 = pi14 ? n13309 : n13328;
  assign n13330 = pi13 ? n13288 : n13329;
  assign n13331 = pi12 ? n13245 : n13330;
  assign n13332 = pi11 ? n13137 : n13331;
  assign n13333 = pi19 ? n2095 : n6355;
  assign n13334 = pi18 ? n13333 : n12858;
  assign n13335 = pi17 ? n37 : n13334;
  assign n13336 = pi16 ? n439 : n13335;
  assign n13337 = pi20 ? n37 : n233;
  assign n13338 = pi19 ? n2095 : n13337;
  assign n13339 = pi21 ? n233 : n2578;
  assign n13340 = pi20 ? n13339 : n32;
  assign n13341 = pi19 ? n13340 : n32;
  assign n13342 = pi18 ? n13338 : n13341;
  assign n13343 = pi17 ? n37 : n13342;
  assign n13344 = pi16 ? n439 : n13343;
  assign n13345 = pi15 ? n13336 : n13344;
  assign n13346 = pi21 ? n37 : n2117;
  assign n13347 = pi20 ? n37 : n13346;
  assign n13348 = pi21 ? n4891 : n2117;
  assign n13349 = pi22 ? n559 : n2116;
  assign n13350 = pi21 ? n13349 : n2048;
  assign n13351 = pi20 ? n13348 : n13350;
  assign n13352 = pi19 ? n13347 : n13351;
  assign n13353 = pi21 ? n3409 : n2637;
  assign n13354 = pi20 ? n13353 : n32;
  assign n13355 = pi19 ? n13354 : n32;
  assign n13356 = pi18 ? n13352 : n13355;
  assign n13357 = pi17 ? n37 : n13356;
  assign n13358 = pi16 ? n439 : n13357;
  assign n13359 = pi15 ? n13358 : n12877;
  assign n13360 = pi14 ? n13345 : n13359;
  assign n13361 = pi21 ? n2759 : n928;
  assign n13362 = pi20 ? n13361 : n32;
  assign n13363 = pi19 ? n13362 : n32;
  assign n13364 = pi18 ? n37 : n13363;
  assign n13365 = pi17 ? n37 : n13364;
  assign n13366 = pi16 ? n439 : n13365;
  assign n13367 = pi15 ? n12877 : n13366;
  assign n13368 = pi14 ? n12877 : n13367;
  assign n13369 = pi13 ? n13360 : n13368;
  assign n13370 = pi16 ? n744 : n12913;
  assign n13371 = pi20 ? n99 : n777;
  assign n13372 = pi19 ? n99 : n13371;
  assign n13373 = pi18 ? n13372 : n12911;
  assign n13374 = pi17 ? n99 : n13373;
  assign n13375 = pi16 ? n744 : n13374;
  assign n13376 = pi15 ? n13370 : n13375;
  assign n13377 = pi19 ? n99 : n6091;
  assign n13378 = pi21 ? n6461 : n1009;
  assign n13379 = pi20 ? n13378 : n32;
  assign n13380 = pi19 ? n13379 : n32;
  assign n13381 = pi18 ? n13377 : n13380;
  assign n13382 = pi17 ? n99 : n13381;
  assign n13383 = pi16 ? n744 : n13382;
  assign n13384 = pi21 ? n777 : n767;
  assign n13385 = pi20 ? n99 : n13384;
  assign n13386 = pi19 ? n13385 : n99;
  assign n13387 = pi18 ? n99 : n13386;
  assign n13388 = pi20 ? n5085 : n685;
  assign n13389 = pi19 ? n99 : n13388;
  assign n13390 = pi18 ? n13389 : n11676;
  assign n13391 = pi17 ? n13387 : n13390;
  assign n13392 = pi16 ? n744 : n13391;
  assign n13393 = pi15 ? n13383 : n13392;
  assign n13394 = pi14 ? n13376 : n13393;
  assign n13395 = pi18 ? n157 : n11676;
  assign n13396 = pi17 ? n157 : n13395;
  assign n13397 = pi16 ? n7793 : n13396;
  assign n13398 = pi21 ? n316 : n32;
  assign n13399 = pi20 ? n13398 : n32;
  assign n13400 = pi19 ? n13399 : n32;
  assign n13401 = pi18 ? n157 : n13400;
  assign n13402 = pi17 ? n157 : n13401;
  assign n13403 = pi16 ? n7793 : n13402;
  assign n13404 = pi15 ? n13397 : n13403;
  assign n13405 = pi18 ? n99 : n13400;
  assign n13406 = pi17 ? n99 : n13405;
  assign n13407 = pi16 ? n744 : n13406;
  assign n13408 = pi22 ? n1484 : n396;
  assign n13409 = pi21 ? n13408 : n32;
  assign n13410 = pi20 ? n13409 : n32;
  assign n13411 = pi19 ? n13410 : n32;
  assign n13412 = pi18 ? n99 : n13411;
  assign n13413 = pi17 ? n99 : n13412;
  assign n13414 = pi16 ? n744 : n13413;
  assign n13415 = pi15 ? n13407 : n13414;
  assign n13416 = pi14 ? n13404 : n13415;
  assign n13417 = pi13 ? n13394 : n13416;
  assign n13418 = pi12 ? n13369 : n13417;
  assign n13419 = pi21 ? n139 : n4252;
  assign n13420 = pi20 ? n139 : n13419;
  assign n13421 = pi19 ? n139 : n13420;
  assign n13422 = pi18 ? n13421 : n6937;
  assign n13423 = pi17 ? n139 : n13422;
  assign n13424 = pi16 ? n915 : n13423;
  assign n13425 = pi18 ? n1821 : n6937;
  assign n13426 = pi17 ? n139 : n13425;
  assign n13427 = pi16 ? n915 : n13426;
  assign n13428 = pi15 ? n13424 : n13427;
  assign n13429 = pi21 ? n12381 : n32;
  assign n13430 = pi20 ? n13429 : n32;
  assign n13431 = pi19 ? n13430 : n32;
  assign n13432 = pi18 ? n12590 : n13431;
  assign n13433 = pi17 ? n139 : n13432;
  assign n13434 = pi16 ? n915 : n13433;
  assign n13435 = pi15 ? n12551 : n13434;
  assign n13436 = pi14 ? n13428 : n13435;
  assign n13437 = pi19 ? n9068 : n316;
  assign n13438 = pi18 ? n13437 : n316;
  assign n13439 = pi17 ? n13438 : n6225;
  assign n13440 = pi16 ? n7883 : n13439;
  assign n13441 = pi22 ? n4338 : n204;
  assign n13442 = pi21 ? n13441 : n316;
  assign n13443 = pi20 ? n32 : n13442;
  assign n13444 = pi19 ? n32 : n13443;
  assign n13445 = pi18 ? n13444 : n316;
  assign n13446 = pi17 ? n32 : n13445;
  assign n13447 = pi21 ? n316 : n4712;
  assign n13448 = pi21 ? n916 : n316;
  assign n13449 = pi20 ? n13447 : n13448;
  assign n13450 = pi19 ? n13449 : n316;
  assign n13451 = pi18 ? n13450 : n316;
  assign n13452 = pi17 ? n13451 : n12566;
  assign n13453 = pi16 ? n13446 : n13452;
  assign n13454 = pi15 ? n12570 : n13453;
  assign n13455 = pi14 ? n13440 : n13454;
  assign n13456 = pi13 ? n13436 : n13455;
  assign n13457 = pi21 ? n1549 : n204;
  assign n13458 = pi20 ? n32 : n13457;
  assign n13459 = pi19 ? n32 : n13458;
  assign n13460 = pi18 ? n13459 : n204;
  assign n13461 = pi17 ? n32 : n13460;
  assign n13462 = pi20 ? n2318 : n139;
  assign n13463 = pi19 ? n13462 : n204;
  assign n13464 = pi18 ? n13463 : n204;
  assign n13465 = pi22 ? n2299 : n706;
  assign n13466 = pi21 ? n13465 : n32;
  assign n13467 = pi20 ? n13466 : n32;
  assign n13468 = pi19 ? n13467 : n32;
  assign n13469 = pi18 ? n204 : n13468;
  assign n13470 = pi17 ? n13464 : n13469;
  assign n13471 = pi16 ? n13461 : n13470;
  assign n13472 = pi22 ? n4375 : n204;
  assign n13473 = pi21 ? n13472 : n204;
  assign n13474 = pi20 ? n32 : n13473;
  assign n13475 = pi19 ? n32 : n13474;
  assign n13476 = pi18 ? n13475 : n204;
  assign n13477 = pi17 ? n32 : n13476;
  assign n13478 = pi20 ? n1063 : n1057;
  assign n13479 = pi19 ? n13478 : n204;
  assign n13480 = pi18 ? n13479 : n204;
  assign n13481 = pi25 ? n315 : n32;
  assign n13482 = pi24 ? n685 : n13481;
  assign n13483 = pi23 ? n204 : n13482;
  assign n13484 = pi22 ? n13483 : n32;
  assign n13485 = pi21 ? n13484 : n32;
  assign n13486 = pi20 ? n13485 : n32;
  assign n13487 = pi19 ? n13486 : n32;
  assign n13488 = pi18 ? n204 : n13487;
  assign n13489 = pi17 ? n13480 : n13488;
  assign n13490 = pi16 ? n13477 : n13489;
  assign n13491 = pi15 ? n13471 : n13490;
  assign n13492 = pi18 ? n2394 : n204;
  assign n13493 = pi17 ? n32 : n13492;
  assign n13494 = pi20 ? n1063 : n4878;
  assign n13495 = pi19 ? n13494 : n204;
  assign n13496 = pi18 ? n13495 : n204;
  assign n13497 = pi18 ? n204 : n6419;
  assign n13498 = pi17 ? n13496 : n13497;
  assign n13499 = pi16 ? n13493 : n13498;
  assign n13500 = pi19 ? n335 : n7944;
  assign n13501 = pi18 ? n13500 : n5832;
  assign n13502 = pi17 ? n335 : n13501;
  assign n13503 = pi16 ? n7943 : n13502;
  assign n13504 = pi15 ? n13499 : n13503;
  assign n13505 = pi14 ? n13491 : n13504;
  assign n13506 = pi20 ? n610 : n4939;
  assign n13507 = pi19 ? n13506 : n335;
  assign n13508 = pi18 ? n13507 : n335;
  assign n13509 = pi22 ? n335 : n673;
  assign n13510 = pi21 ? n335 : n13509;
  assign n13511 = pi20 ? n335 : n13510;
  assign n13512 = pi19 ? n335 : n13511;
  assign n13513 = pi18 ? n13512 : n2655;
  assign n13514 = pi17 ? n13508 : n13513;
  assign n13515 = pi16 ? n7943 : n13514;
  assign n13516 = pi22 ? n335 : n1457;
  assign n13517 = pi21 ? n335 : n13516;
  assign n13518 = pi20 ? n335 : n13517;
  assign n13519 = pi19 ? n335 : n13518;
  assign n13520 = pi18 ? n13519 : n2703;
  assign n13521 = pi17 ? n335 : n13520;
  assign n13522 = pi16 ? n10980 : n13521;
  assign n13523 = pi15 ? n13515 : n13522;
  assign n13524 = pi18 ? n12631 : n2703;
  assign n13525 = pi17 ? n335 : n13524;
  assign n13526 = pi16 ? n10980 : n13525;
  assign n13527 = pi21 ? n335 : n233;
  assign n13528 = pi20 ? n335 : n13527;
  assign n13529 = pi19 ? n335 : n13528;
  assign n13530 = pi18 ? n12656 : n13529;
  assign n13531 = pi17 ? n32 : n13530;
  assign n13532 = pi20 ? n335 : n233;
  assign n13533 = pi19 ? n13532 : n233;
  assign n13534 = pi18 ? n335 : n13533;
  assign n13535 = pi20 ? n13527 : n233;
  assign n13536 = pi19 ? n7985 : n13535;
  assign n13537 = pi18 ? n13536 : n1824;
  assign n13538 = pi17 ? n13534 : n13537;
  assign n13539 = pi16 ? n13531 : n13538;
  assign n13540 = pi15 ? n13526 : n13539;
  assign n13541 = pi14 ? n13523 : n13540;
  assign n13542 = pi13 ? n13505 : n13541;
  assign n13543 = pi12 ? n13456 : n13542;
  assign n13544 = pi11 ? n13418 : n13543;
  assign n13545 = pi10 ? n13332 : n13544;
  assign n13546 = pi09 ? n13023 : n13545;
  assign n13547 = pi15 ? n32 : n13016;
  assign n13548 = pi16 ? n10154 : n13013;
  assign n13549 = pi15 ? n13017 : n13548;
  assign n13550 = pi14 ? n13547 : n13549;
  assign n13551 = pi13 ? n32 : n13550;
  assign n13552 = pi12 ? n32 : n13551;
  assign n13553 = pi11 ? n32 : n13552;
  assign n13554 = pi10 ? n32 : n13553;
  assign n13555 = pi16 ? n11011 : n13029;
  assign n13556 = pi16 ? n11885 : n13036;
  assign n13557 = pi15 ? n13555 : n13556;
  assign n13558 = pi20 ? n32 : n57;
  assign n13559 = pi19 ? n32 : n13558;
  assign n13560 = pi18 ? n13559 : n37;
  assign n13561 = pi17 ? n32 : n13560;
  assign n13562 = pi16 ? n13561 : n13044;
  assign n13563 = pi15 ? n13046 : n13562;
  assign n13564 = pi14 ? n13557 : n13563;
  assign n13565 = pi21 ? n157 : n6115;
  assign n13566 = pi20 ? n13565 : n32;
  assign n13567 = pi19 ? n13566 : n32;
  assign n13568 = pi18 ? n157 : n13567;
  assign n13569 = pi17 ? n157 : n13568;
  assign n13570 = pi16 ? n13067 : n13569;
  assign n13571 = pi17 ? n13075 : n13568;
  assign n13572 = pi16 ? n13073 : n13571;
  assign n13573 = pi15 ? n13570 : n13572;
  assign n13574 = pi14 ? n13062 : n13573;
  assign n13575 = pi13 ? n13564 : n13574;
  assign n13576 = pi22 ? n99 : n6114;
  assign n13577 = pi21 ? n99 : n13576;
  assign n13578 = pi20 ? n13577 : n32;
  assign n13579 = pi19 ? n13578 : n32;
  assign n13580 = pi18 ? n99 : n13579;
  assign n13581 = pi17 ? n99 : n13580;
  assign n13582 = pi16 ? n801 : n13581;
  assign n13583 = pi16 ? n721 : n13581;
  assign n13584 = pi15 ? n13582 : n13583;
  assign n13585 = pi22 ? n99 : n3174;
  assign n13586 = pi21 ? n99 : n13585;
  assign n13587 = pi20 ? n13586 : n32;
  assign n13588 = pi19 ? n13587 : n32;
  assign n13589 = pi18 ? n99 : n13588;
  assign n13590 = pi17 ? n99 : n13589;
  assign n13591 = pi16 ? n801 : n13590;
  assign n13592 = pi16 ? n744 : n13590;
  assign n13593 = pi15 ? n13591 : n13592;
  assign n13594 = pi14 ? n13584 : n13593;
  assign n13595 = pi22 ? n99 : n1388;
  assign n13596 = pi21 ? n99 : n13595;
  assign n13597 = pi20 ? n13596 : n32;
  assign n13598 = pi19 ? n13597 : n32;
  assign n13599 = pi18 ? n99 : n13598;
  assign n13600 = pi17 ? n99 : n13599;
  assign n13601 = pi16 ? n721 : n13600;
  assign n13602 = pi22 ? n139 : n1388;
  assign n13603 = pi21 ? n139 : n13602;
  assign n13604 = pi20 ? n13603 : n32;
  assign n13605 = pi19 ? n13604 : n32;
  assign n13606 = pi18 ? n13101 : n13605;
  assign n13607 = pi17 ? n13099 : n13606;
  assign n13608 = pi16 ? n13097 : n13607;
  assign n13609 = pi15 ? n13601 : n13608;
  assign n13610 = pi19 ? n13180 : n37;
  assign n13611 = pi18 ? n37 : n13610;
  assign n13612 = pi21 ? n3073 : n1696;
  assign n13613 = pi21 ? n375 : n37;
  assign n13614 = pi20 ? n13612 : n13613;
  assign n13615 = pi20 ? n13613 : n8742;
  assign n13616 = pi19 ? n13614 : n13615;
  assign n13617 = pi18 ? n13616 : n13112;
  assign n13618 = pi17 ? n13611 : n13617;
  assign n13619 = pi16 ? n439 : n13618;
  assign n13620 = pi15 ? n13619 : n13133;
  assign n13621 = pi14 ? n13609 : n13620;
  assign n13622 = pi13 ? n13594 : n13621;
  assign n13623 = pi12 ? n13575 : n13622;
  assign n13624 = pi23 ? n37 : n5612;
  assign n13625 = pi22 ? n37 : n13624;
  assign n13626 = pi23 ? n7420 : n32;
  assign n13627 = pi22 ? n139 : n13626;
  assign n13628 = pi21 ? n13625 : n13627;
  assign n13629 = pi20 ? n13628 : n32;
  assign n13630 = pi19 ? n13629 : n32;
  assign n13631 = pi18 ? n13158 : n13630;
  assign n13632 = pi17 ? n12372 : n13631;
  assign n13633 = pi16 ? n439 : n13632;
  assign n13634 = pi15 ? n13155 : n13633;
  assign n13635 = pi21 ? n139 : n4669;
  assign n13636 = pi20 ? n13635 : n32;
  assign n13637 = pi19 ? n13636 : n32;
  assign n13638 = pi18 ? n13183 : n13637;
  assign n13639 = pi17 ? n13182 : n13638;
  assign n13640 = pi16 ? n439 : n13639;
  assign n13641 = pi15 ? n13178 : n13640;
  assign n13642 = pi14 ? n13634 : n13641;
  assign n13643 = pi20 ? n3086 : n3245;
  assign n13644 = pi19 ? n37 : n13643;
  assign n13645 = pi18 ? n37 : n13644;
  assign n13646 = pi20 ? n11579 : n1737;
  assign n13647 = pi20 ? n1737 : n3656;
  assign n13648 = pi19 ? n13646 : n13647;
  assign n13649 = pi21 ? n375 : n5632;
  assign n13650 = pi20 ? n13649 : n32;
  assign n13651 = pi19 ? n13650 : n32;
  assign n13652 = pi18 ? n13648 : n13651;
  assign n13653 = pi17 ? n13645 : n13652;
  assign n13654 = pi16 ? n439 : n13653;
  assign n13655 = pi15 ? n13200 : n13654;
  assign n13656 = pi21 ? n506 : n499;
  assign n13657 = pi20 ? n37 : n13656;
  assign n13658 = pi19 ? n37 : n13657;
  assign n13659 = pi18 ? n37 : n13658;
  assign n13660 = pi21 ? n457 : n1056;
  assign n13661 = pi21 ? n485 : n506;
  assign n13662 = pi20 ? n13660 : n13661;
  assign n13663 = pi21 ? n499 : n2395;
  assign n13664 = pi21 ? n499 : n204;
  assign n13665 = pi20 ? n13663 : n13664;
  assign n13666 = pi19 ? n13662 : n13665;
  assign n13667 = pi18 ? n13666 : n13222;
  assign n13668 = pi17 ? n13659 : n13667;
  assign n13669 = pi16 ? n439 : n13668;
  assign n13670 = pi21 ? n567 : n1936;
  assign n13671 = pi20 ? n1983 : n13670;
  assign n13672 = pi19 ? n13233 : n13671;
  assign n13673 = pi21 ? n1943 : n8937;
  assign n13674 = pi20 ? n13673 : n32;
  assign n13675 = pi19 ? n13674 : n32;
  assign n13676 = pi18 ? n13672 : n13675;
  assign n13677 = pi17 ? n13229 : n13676;
  assign n13678 = pi16 ? n439 : n13677;
  assign n13679 = pi15 ? n13669 : n13678;
  assign n13680 = pi14 ? n13655 : n13679;
  assign n13681 = pi13 ? n13642 : n13680;
  assign n13682 = pi20 ? n13251 : n6377;
  assign n13683 = pi19 ? n13252 : n13682;
  assign n13684 = pi18 ? n13683 : n13259;
  assign n13685 = pi17 ? n13249 : n13684;
  assign n13686 = pi16 ? n439 : n13685;
  assign n13687 = pi22 ? n685 : n532;
  assign n13688 = pi21 ? n569 : n13687;
  assign n13689 = pi20 ? n13688 : n32;
  assign n13690 = pi19 ? n13689 : n32;
  assign n13691 = pi18 ? n37 : n13690;
  assign n13692 = pi17 ? n37 : n13691;
  assign n13693 = pi16 ? n439 : n13692;
  assign n13694 = pi15 ? n13686 : n13693;
  assign n13695 = pi21 ? n2074 : n650;
  assign n13696 = pi20 ? n13695 : n32;
  assign n13697 = pi19 ? n13696 : n32;
  assign n13698 = pi18 ? n6374 : n13697;
  assign n13699 = pi17 ? n37 : n13698;
  assign n13700 = pi16 ? n439 : n13699;
  assign n13701 = pi21 ? n584 : n650;
  assign n13702 = pi20 ? n13701 : n32;
  assign n13703 = pi19 ? n13702 : n32;
  assign n13704 = pi18 ? n13277 : n13703;
  assign n13705 = pi17 ? n37 : n13704;
  assign n13706 = pi16 ? n439 : n13705;
  assign n13707 = pi15 ? n13700 : n13706;
  assign n13708 = pi14 ? n13694 : n13707;
  assign n13709 = pi21 ? n569 : n5758;
  assign n13710 = pi20 ? n13709 : n32;
  assign n13711 = pi19 ? n13710 : n32;
  assign n13712 = pi18 ? n13291 : n13711;
  assign n13713 = pi17 ? n37 : n13712;
  assign n13714 = pi16 ? n439 : n13713;
  assign n13715 = pi15 ? n13714 : n13308;
  assign n13716 = pi21 ? n6401 : n9666;
  assign n13717 = pi20 ? n37 : n13716;
  assign n13718 = pi21 ? n5012 : n7326;
  assign n13719 = pi21 ? n5012 : n9657;
  assign n13720 = pi20 ? n13718 : n13719;
  assign n13721 = pi19 ? n13717 : n13720;
  assign n13722 = pi22 ? n4925 : n32;
  assign n13723 = pi21 ? n3392 : n13722;
  assign n13724 = pi20 ? n13723 : n32;
  assign n13725 = pi19 ? n13724 : n32;
  assign n13726 = pi18 ? n13721 : n13725;
  assign n13727 = pi17 ? n37 : n13726;
  assign n13728 = pi16 ? n439 : n13727;
  assign n13729 = pi21 ? n2091 : n12825;
  assign n13730 = pi20 ? n13729 : n32;
  assign n13731 = pi19 ? n13730 : n32;
  assign n13732 = pi18 ? n6356 : n13731;
  assign n13733 = pi17 ? n37 : n13732;
  assign n13734 = pi16 ? n439 : n13733;
  assign n13735 = pi15 ? n13728 : n13734;
  assign n13736 = pi14 ? n13715 : n13735;
  assign n13737 = pi13 ? n13708 : n13736;
  assign n13738 = pi12 ? n13681 : n13737;
  assign n13739 = pi11 ? n13623 : n13738;
  assign n13740 = pi18 ? n13333 : n13731;
  assign n13741 = pi17 ? n37 : n13740;
  assign n13742 = pi16 ? n439 : n13741;
  assign n13743 = pi21 ? n233 : n4109;
  assign n13744 = pi20 ? n13743 : n32;
  assign n13745 = pi19 ? n13744 : n32;
  assign n13746 = pi18 ? n13338 : n13745;
  assign n13747 = pi17 ? n37 : n13746;
  assign n13748 = pi16 ? n439 : n13747;
  assign n13749 = pi15 ? n13742 : n13748;
  assign n13750 = pi21 ? n4891 : n1920;
  assign n13751 = pi21 ? n4891 : n560;
  assign n13752 = pi20 ? n13750 : n13751;
  assign n13753 = pi19 ? n13347 : n13752;
  assign n13754 = pi21 ? n2117 : n760;
  assign n13755 = pi20 ? n13754 : n32;
  assign n13756 = pi19 ? n13755 : n32;
  assign n13757 = pi18 ? n13753 : n13756;
  assign n13758 = pi17 ? n37 : n13757;
  assign n13759 = pi16 ? n439 : n13758;
  assign n13760 = pi21 ? n2106 : n760;
  assign n13761 = pi20 ? n13760 : n32;
  assign n13762 = pi19 ? n13761 : n32;
  assign n13763 = pi18 ? n37 : n13762;
  assign n13764 = pi17 ? n37 : n13763;
  assign n13765 = pi16 ? n439 : n13764;
  assign n13766 = pi15 ? n13759 : n13765;
  assign n13767 = pi14 ? n13749 : n13766;
  assign n13768 = pi21 ? n2759 : n882;
  assign n13769 = pi20 ? n13768 : n32;
  assign n13770 = pi19 ? n13769 : n32;
  assign n13771 = pi18 ? n37 : n13770;
  assign n13772 = pi17 ? n37 : n13771;
  assign n13773 = pi16 ? n439 : n13772;
  assign n13774 = pi15 ? n13765 : n13773;
  assign n13775 = pi14 ? n13765 : n13774;
  assign n13776 = pi13 ? n13767 : n13775;
  assign n13777 = pi21 ? n6461 : n2637;
  assign n13778 = pi20 ? n13777 : n32;
  assign n13779 = pi19 ? n13778 : n32;
  assign n13780 = pi18 ? n99 : n13779;
  assign n13781 = pi17 ? n99 : n13780;
  assign n13782 = pi16 ? n721 : n13781;
  assign n13783 = pi21 ? n6461 : n928;
  assign n13784 = pi20 ? n13783 : n32;
  assign n13785 = pi19 ? n13784 : n32;
  assign n13786 = pi18 ? n13372 : n13785;
  assign n13787 = pi17 ? n99 : n13786;
  assign n13788 = pi16 ? n721 : n13787;
  assign n13789 = pi15 ? n13782 : n13788;
  assign n13790 = pi18 ? n13377 : n13785;
  assign n13791 = pi17 ? n99 : n13790;
  assign n13792 = pi16 ? n721 : n13791;
  assign n13793 = pi21 ? n685 : n1009;
  assign n13794 = pi20 ? n13793 : n32;
  assign n13795 = pi19 ? n13794 : n32;
  assign n13796 = pi18 ? n13389 : n13795;
  assign n13797 = pi17 ? n13387 : n13796;
  assign n13798 = pi16 ? n721 : n13797;
  assign n13799 = pi15 ? n13792 : n13798;
  assign n13800 = pi14 ? n13789 : n13799;
  assign n13801 = pi18 ? n157 : n13795;
  assign n13802 = pi17 ? n157 : n13801;
  assign n13803 = pi16 ? n5910 : n13802;
  assign n13804 = pi16 ? n5910 : n13402;
  assign n13805 = pi15 ? n13803 : n13804;
  assign n13806 = pi16 ? n721 : n13413;
  assign n13807 = pi15 ? n13407 : n13806;
  assign n13808 = pi14 ? n13805 : n13807;
  assign n13809 = pi13 ? n13800 : n13808;
  assign n13810 = pi12 ? n13776 : n13809;
  assign n13811 = pi19 ? n139 : n6592;
  assign n13812 = pi18 ? n13811 : n6937;
  assign n13813 = pi17 ? n139 : n13812;
  assign n13814 = pi16 ? n2291 : n13813;
  assign n13815 = pi16 ? n2291 : n13426;
  assign n13816 = pi15 ? n13814 : n13815;
  assign n13817 = pi16 ? n2291 : n13433;
  assign n13818 = pi15 ? n12946 : n13817;
  assign n13819 = pi14 ? n13816 : n13818;
  assign n13820 = pi21 ? n5186 : n316;
  assign n13821 = pi20 ? n32 : n13820;
  assign n13822 = pi19 ? n32 : n13821;
  assign n13823 = pi18 ? n13822 : n316;
  assign n13824 = pi17 ? n32 : n13823;
  assign n13825 = pi16 ? n13824 : n13452;
  assign n13826 = pi15 ? n12952 : n13825;
  assign n13827 = pi14 ? n13440 : n13826;
  assign n13828 = pi13 ? n13819 : n13827;
  assign n13829 = pi21 ? n326 : n204;
  assign n13830 = pi20 ? n32 : n13829;
  assign n13831 = pi19 ? n32 : n13830;
  assign n13832 = pi18 ? n13831 : n204;
  assign n13833 = pi17 ? n32 : n13832;
  assign n13834 = pi23 ? n204 : n8133;
  assign n13835 = pi22 ? n13834 : n706;
  assign n13836 = pi21 ? n13835 : n32;
  assign n13837 = pi20 ? n13836 : n32;
  assign n13838 = pi19 ? n13837 : n32;
  assign n13839 = pi18 ? n204 : n13838;
  assign n13840 = pi17 ? n13464 : n13839;
  assign n13841 = pi16 ? n13833 : n13840;
  assign n13842 = pi21 ? n1037 : n204;
  assign n13843 = pi20 ? n32 : n13842;
  assign n13844 = pi19 ? n32 : n13843;
  assign n13845 = pi18 ? n13844 : n204;
  assign n13846 = pi17 ? n32 : n13845;
  assign n13847 = pi18 ? n204 : n4097;
  assign n13848 = pi17 ? n13480 : n13847;
  assign n13849 = pi16 ? n13846 : n13848;
  assign n13850 = pi15 ? n13841 : n13849;
  assign n13851 = pi18 ? n204 : n4104;
  assign n13852 = pi17 ? n13496 : n13851;
  assign n13853 = pi16 ? n13493 : n13852;
  assign n13854 = pi18 ? n13500 : n4118;
  assign n13855 = pi17 ? n335 : n13854;
  assign n13856 = pi16 ? n7943 : n13855;
  assign n13857 = pi15 ? n13853 : n13856;
  assign n13858 = pi14 ? n13850 : n13857;
  assign n13859 = pi18 ? n13512 : n10013;
  assign n13860 = pi17 ? n13508 : n13859;
  assign n13861 = pi16 ? n7943 : n13860;
  assign n13862 = pi18 ? n13519 : n2640;
  assign n13863 = pi17 ? n335 : n13862;
  assign n13864 = pi16 ? n10980 : n13863;
  assign n13865 = pi15 ? n13861 : n13864;
  assign n13866 = pi18 ? n12631 : n2640;
  assign n13867 = pi17 ? n335 : n13866;
  assign n13868 = pi16 ? n10980 : n13867;
  assign n13869 = pi18 ? n13536 : n2655;
  assign n13870 = pi17 ? n13534 : n13869;
  assign n13871 = pi16 ? n13531 : n13870;
  assign n13872 = pi15 ? n13868 : n13871;
  assign n13873 = pi14 ? n13865 : n13872;
  assign n13874 = pi13 ? n13858 : n13873;
  assign n13875 = pi12 ? n13828 : n13874;
  assign n13876 = pi11 ? n13810 : n13875;
  assign n13877 = pi10 ? n13739 : n13876;
  assign n13878 = pi09 ? n13554 : n13877;
  assign n13879 = pi08 ? n13546 : n13878;
  assign n13880 = pi20 ? n37 : n32;
  assign n13881 = pi19 ? n13880 : n32;
  assign n13882 = pi18 ? n37 : n13881;
  assign n13883 = pi17 ? n37 : n13882;
  assign n13884 = pi16 ? n9232 : n13883;
  assign n13885 = pi15 ? n32 : n13884;
  assign n13886 = pi16 ? n2461 : n13883;
  assign n13887 = pi16 ? n10154 : n13883;
  assign n13888 = pi15 ? n13886 : n13887;
  assign n13889 = pi14 ? n13885 : n13888;
  assign n13890 = pi13 ? n32 : n13889;
  assign n13891 = pi12 ? n32 : n13890;
  assign n13892 = pi11 ? n32 : n13891;
  assign n13893 = pi10 ? n32 : n13892;
  assign n13894 = pi20 ? n5077 : n32;
  assign n13895 = pi19 ? n13894 : n32;
  assign n13896 = pi18 ? n37 : n13895;
  assign n13897 = pi17 ? n37 : n13896;
  assign n13898 = pi16 ? n11011 : n13897;
  assign n13899 = pi20 ? n3086 : n32;
  assign n13900 = pi19 ? n13899 : n32;
  assign n13901 = pi18 ? n37 : n13900;
  assign n13902 = pi17 ? n37 : n13901;
  assign n13903 = pi16 ? n11885 : n13902;
  assign n13904 = pi15 ? n13898 : n13903;
  assign n13905 = pi20 ? n649 : n32;
  assign n13906 = pi19 ? n13905 : n32;
  assign n13907 = pi18 ? n37 : n13906;
  assign n13908 = pi17 ? n37 : n13907;
  assign n13909 = pi16 ? n12689 : n13908;
  assign n13910 = pi21 ? n37 : n6789;
  assign n13911 = pi20 ? n13910 : n32;
  assign n13912 = pi19 ? n13911 : n32;
  assign n13913 = pi18 ? n37 : n13912;
  assign n13914 = pi17 ? n37 : n13913;
  assign n13915 = pi16 ? n13561 : n13914;
  assign n13916 = pi15 ? n13909 : n13915;
  assign n13917 = pi14 ? n13904 : n13916;
  assign n13918 = pi23 ? n99 : n586;
  assign n13919 = pi22 ? n99 : n13918;
  assign n13920 = pi21 ? n99 : n13919;
  assign n13921 = pi20 ? n13920 : n32;
  assign n13922 = pi19 ? n13921 : n32;
  assign n13923 = pi18 ? n99 : n13922;
  assign n13924 = pi17 ? n99 : n13923;
  assign n13925 = pi16 ? n3065 : n13924;
  assign n13926 = pi16 ? n801 : n13924;
  assign n13927 = pi15 ? n13925 : n13926;
  assign n13928 = pi21 ? n3060 : n5899;
  assign n13929 = pi20 ? n32 : n13928;
  assign n13930 = pi19 ? n32 : n13929;
  assign n13931 = pi18 ? n13930 : n157;
  assign n13932 = pi17 ? n32 : n13931;
  assign n13933 = pi23 ? n157 : n5630;
  assign n13934 = pi22 ? n157 : n13933;
  assign n13935 = pi21 ? n157 : n13934;
  assign n13936 = pi20 ? n13935 : n32;
  assign n13937 = pi19 ? n13936 : n32;
  assign n13938 = pi18 ? n157 : n13937;
  assign n13939 = pi17 ? n157 : n13938;
  assign n13940 = pi16 ? n13932 : n13939;
  assign n13941 = pi21 ? n739 : n168;
  assign n13942 = pi20 ? n32 : n13941;
  assign n13943 = pi19 ? n32 : n13942;
  assign n13944 = pi20 ? n776 : n2238;
  assign n13945 = pi19 ? n13944 : n9715;
  assign n13946 = pi18 ? n13943 : n13945;
  assign n13947 = pi17 ? n32 : n13946;
  assign n13948 = pi21 ? n777 : n99;
  assign n13949 = pi20 ? n13948 : n776;
  assign n13950 = pi20 ? n7818 : n9015;
  assign n13951 = pi19 ? n13949 : n13950;
  assign n13952 = pi21 ? n12703 : n775;
  assign n13953 = pi20 ? n9015 : n13952;
  assign n13954 = pi21 ? n164 : n157;
  assign n13955 = pi20 ? n13954 : n7823;
  assign n13956 = pi19 ? n13953 : n13955;
  assign n13957 = pi18 ? n13951 : n13956;
  assign n13958 = pi19 ? n157 : n787;
  assign n13959 = pi22 ? n157 : n10510;
  assign n13960 = pi21 ? n157 : n13959;
  assign n13961 = pi20 ? n13960 : n32;
  assign n13962 = pi19 ? n13961 : n32;
  assign n13963 = pi18 ? n13958 : n13962;
  assign n13964 = pi17 ? n13957 : n13963;
  assign n13965 = pi16 ? n13947 : n13964;
  assign n13966 = pi15 ? n13940 : n13965;
  assign n13967 = pi14 ? n13927 : n13966;
  assign n13968 = pi13 ? n13917 : n13967;
  assign n13969 = pi23 ? n37 : n1149;
  assign n13970 = pi22 ? n99 : n13969;
  assign n13971 = pi21 ? n99 : n13970;
  assign n13972 = pi20 ? n13971 : n32;
  assign n13973 = pi19 ? n13972 : n32;
  assign n13974 = pi18 ? n99 : n13973;
  assign n13975 = pi17 ? n99 : n13974;
  assign n13976 = pi16 ? n801 : n13975;
  assign n13977 = pi16 ? n744 : n13975;
  assign n13978 = pi15 ? n13976 : n13977;
  assign n13979 = pi20 ? n1187 : n32;
  assign n13980 = pi19 ? n13979 : n32;
  assign n13981 = pi18 ? n99 : n13980;
  assign n13982 = pi17 ? n99 : n13981;
  assign n13983 = pi16 ? n744 : n13982;
  assign n13984 = pi23 ? n3491 : n531;
  assign n13985 = pi22 ? n99 : n13984;
  assign n13986 = pi21 ? n99 : n13985;
  assign n13987 = pi20 ? n13986 : n32;
  assign n13988 = pi19 ? n13987 : n32;
  assign n13989 = pi18 ? n99 : n13988;
  assign n13990 = pi17 ? n99 : n13989;
  assign n13991 = pi16 ? n801 : n13990;
  assign n13992 = pi15 ? n13983 : n13991;
  assign n13993 = pi14 ? n13978 : n13992;
  assign n13994 = pi21 ? n739 : n2164;
  assign n13995 = pi20 ? n32 : n13994;
  assign n13996 = pi19 ? n32 : n13995;
  assign n13997 = pi20 ? n4616 : n2189;
  assign n13998 = pi20 ? n3506 : n3805;
  assign n13999 = pi19 ? n13997 : n13998;
  assign n14000 = pi18 ? n13996 : n13999;
  assign n14001 = pi17 ? n32 : n14000;
  assign n14002 = pi19 ? n6045 : n3807;
  assign n14003 = pi20 ? n2752 : n3807;
  assign n14004 = pi19 ? n14003 : n2962;
  assign n14005 = pi18 ? n14002 : n14004;
  assign n14006 = pi20 ? n2163 : n4619;
  assign n14007 = pi19 ? n14006 : n2755;
  assign n14008 = pi23 ? n11962 : n624;
  assign n14009 = pi22 ? n99 : n14008;
  assign n14010 = pi21 ? n2162 : n14009;
  assign n14011 = pi20 ? n14010 : n32;
  assign n14012 = pi19 ? n14011 : n32;
  assign n14013 = pi18 ? n14007 : n14012;
  assign n14014 = pi17 ? n14005 : n14013;
  assign n14015 = pi16 ? n14001 : n14014;
  assign n14016 = pi18 ? n990 : n13095;
  assign n14017 = pi17 ? n32 : n14016;
  assign n14018 = pi23 ? n3134 : n687;
  assign n14019 = pi22 ? n139 : n14018;
  assign n14020 = pi21 ? n139 : n14019;
  assign n14021 = pi20 ? n14020 : n32;
  assign n14022 = pi19 ? n14021 : n32;
  assign n14023 = pi18 ? n13101 : n14022;
  assign n14024 = pi17 ? n13099 : n14023;
  assign n14025 = pi16 ? n14017 : n14024;
  assign n14026 = pi15 ? n14015 : n14025;
  assign n14027 = pi21 ? n37 : n346;
  assign n14028 = pi20 ? n14027 : n32;
  assign n14029 = pi19 ? n14028 : n32;
  assign n14030 = pi18 ? n37 : n14029;
  assign n14031 = pi17 ? n37 : n14030;
  assign n14032 = pi16 ? n439 : n14031;
  assign n14033 = pi20 ? n37 : n8707;
  assign n14034 = pi21 ? n3668 : n1696;
  assign n14035 = pi20 ? n8707 : n14034;
  assign n14036 = pi19 ? n14033 : n14035;
  assign n14037 = pi20 ? n5257 : n37;
  assign n14038 = pi21 ? n1211 : n37;
  assign n14039 = pi21 ? n1211 : n1696;
  assign n14040 = pi20 ? n14038 : n14039;
  assign n14041 = pi19 ? n14037 : n14040;
  assign n14042 = pi18 ? n14036 : n14041;
  assign n14043 = pi21 ? n1529 : n297;
  assign n14044 = pi20 ? n1715 : n14043;
  assign n14045 = pi20 ? n1707 : n1693;
  assign n14046 = pi19 ? n14044 : n14045;
  assign n14047 = pi21 ? n1711 : n346;
  assign n14048 = pi20 ? n14047 : n32;
  assign n14049 = pi19 ? n14048 : n32;
  assign n14050 = pi18 ? n14046 : n14049;
  assign n14051 = pi17 ? n14042 : n14050;
  assign n14052 = pi16 ? n439 : n14051;
  assign n14053 = pi15 ? n14032 : n14052;
  assign n14054 = pi14 ? n14026 : n14053;
  assign n14055 = pi13 ? n13993 : n14054;
  assign n14056 = pi12 ? n13968 : n14055;
  assign n14057 = pi21 ? n3668 : n820;
  assign n14058 = pi20 ? n3083 : n14057;
  assign n14059 = pi19 ? n37 : n14058;
  assign n14060 = pi20 ? n14038 : n37;
  assign n14061 = pi21 ? n1043 : n37;
  assign n14062 = pi21 ? n1043 : n820;
  assign n14063 = pi20 ? n14061 : n14062;
  assign n14064 = pi19 ? n14060 : n14063;
  assign n14065 = pi18 ? n14059 : n14064;
  assign n14066 = pi21 ? n820 : n1696;
  assign n14067 = pi20 ? n14039 : n14066;
  assign n14068 = pi21 ? n820 : n1043;
  assign n14069 = pi20 ? n14068 : n1757;
  assign n14070 = pi19 ? n14067 : n14069;
  assign n14071 = pi20 ? n8782 : n32;
  assign n14072 = pi19 ? n14071 : n32;
  assign n14073 = pi18 ? n14070 : n14072;
  assign n14074 = pi17 ? n14065 : n14073;
  assign n14075 = pi16 ? n439 : n14074;
  assign n14076 = pi21 ? n375 : n1698;
  assign n14077 = pi21 ? n1529 : n1698;
  assign n14078 = pi20 ? n14076 : n14077;
  assign n14079 = pi19 ? n8743 : n14078;
  assign n14080 = pi20 ? n5269 : n2543;
  assign n14081 = pi19 ? n14080 : n2528;
  assign n14082 = pi18 ? n14079 : n14081;
  assign n14083 = pi20 ? n2510 : n139;
  assign n14084 = pi19 ? n13646 : n14083;
  assign n14085 = pi22 ? n139 : n430;
  assign n14086 = pi21 ? n139 : n14085;
  assign n14087 = pi20 ? n14086 : n32;
  assign n14088 = pi19 ? n14087 : n32;
  assign n14089 = pi18 ? n14084 : n14088;
  assign n14090 = pi17 ? n14082 : n14089;
  assign n14091 = pi16 ? n439 : n14090;
  assign n14092 = pi15 ? n14075 : n14091;
  assign n14093 = pi19 ? n37 : n13121;
  assign n14094 = pi20 ? n3086 : n1707;
  assign n14095 = pi20 ? n1707 : n3245;
  assign n14096 = pi19 ? n14094 : n14095;
  assign n14097 = pi18 ? n14093 : n14096;
  assign n14098 = pi21 ? n295 : n14085;
  assign n14099 = pi20 ? n14098 : n32;
  assign n14100 = pi19 ? n14099 : n32;
  assign n14101 = pi18 ? n13648 : n14100;
  assign n14102 = pi17 ? n14097 : n14101;
  assign n14103 = pi16 ? n439 : n14102;
  assign n14104 = pi20 ? n37 : n13143;
  assign n14105 = pi19 ? n14104 : n6596;
  assign n14106 = pi18 ? n37 : n14105;
  assign n14107 = pi21 ? n139 : n6184;
  assign n14108 = pi20 ? n14107 : n32;
  assign n14109 = pi19 ? n14108 : n32;
  assign n14110 = pi18 ? n13183 : n14109;
  assign n14111 = pi17 ? n14106 : n14110;
  assign n14112 = pi16 ? n439 : n14111;
  assign n14113 = pi15 ? n14103 : n14112;
  assign n14114 = pi14 ? n14092 : n14113;
  assign n14115 = pi19 ? n37 : n9795;
  assign n14116 = pi18 ? n37 : n14115;
  assign n14117 = pi21 ? n139 : n6194;
  assign n14118 = pi20 ? n14117 : n32;
  assign n14119 = pi19 ? n14118 : n32;
  assign n14120 = pi18 ? n139 : n14119;
  assign n14121 = pi17 ? n14116 : n14120;
  assign n14122 = pi16 ? n439 : n14121;
  assign n14123 = pi22 ? n566 : n204;
  assign n14124 = pi22 ? n456 : n566;
  assign n14125 = pi21 ? n14123 : n14124;
  assign n14126 = pi21 ? n522 : n14124;
  assign n14127 = pi20 ? n14125 : n14126;
  assign n14128 = pi21 ? n522 : n580;
  assign n14129 = pi21 ? n522 : n569;
  assign n14130 = pi20 ? n14128 : n14129;
  assign n14131 = pi19 ? n14127 : n14130;
  assign n14132 = pi21 ? n1046 : n6194;
  assign n14133 = pi20 ? n14132 : n32;
  assign n14134 = pi19 ? n14133 : n32;
  assign n14135 = pi18 ? n14131 : n14134;
  assign n14136 = pi17 ? n12414 : n14135;
  assign n14137 = pi16 ? n439 : n14136;
  assign n14138 = pi15 ? n14122 : n14137;
  assign n14139 = pi21 ? n1079 : n485;
  assign n14140 = pi21 ? n1083 : n485;
  assign n14141 = pi20 ? n14139 : n14140;
  assign n14142 = pi19 ? n14141 : n14129;
  assign n14143 = pi21 ? n1046 : n6270;
  assign n14144 = pi20 ? n14143 : n32;
  assign n14145 = pi19 ? n14144 : n32;
  assign n14146 = pi18 ? n14142 : n14145;
  assign n14147 = pi17 ? n12414 : n14146;
  assign n14148 = pi16 ? n439 : n14147;
  assign n14149 = pi19 ? n37 : n8802;
  assign n14150 = pi18 ? n37 : n14149;
  assign n14151 = pi21 ? n570 : n2007;
  assign n14152 = pi20 ? n13275 : n14151;
  assign n14153 = pi20 ? n2014 : n4980;
  assign n14154 = pi19 ? n14152 : n14153;
  assign n14155 = pi22 ? n233 : n2564;
  assign n14156 = pi21 ? n583 : n14155;
  assign n14157 = pi20 ? n14156 : n32;
  assign n14158 = pi19 ? n14157 : n32;
  assign n14159 = pi18 ? n14154 : n14158;
  assign n14160 = pi17 ? n14150 : n14159;
  assign n14161 = pi16 ? n439 : n14160;
  assign n14162 = pi15 ? n14148 : n14161;
  assign n14163 = pi14 ? n14138 : n14162;
  assign n14164 = pi13 ? n14114 : n14163;
  assign n14165 = pi18 ? n37 : n7686;
  assign n14166 = pi20 ? n604 : n335;
  assign n14167 = pi19 ? n14166 : n335;
  assign n14168 = pi22 ? n233 : n1407;
  assign n14169 = pi21 ? n335 : n14168;
  assign n14170 = pi20 ? n14169 : n32;
  assign n14171 = pi19 ? n14170 : n32;
  assign n14172 = pi18 ? n14167 : n14171;
  assign n14173 = pi17 ? n14165 : n14172;
  assign n14174 = pi16 ? n439 : n14173;
  assign n14175 = pi22 ? n685 : n664;
  assign n14176 = pi21 ? n569 : n14175;
  assign n14177 = pi20 ? n14176 : n32;
  assign n14178 = pi19 ? n14177 : n32;
  assign n14179 = pi18 ? n37 : n14178;
  assign n14180 = pi17 ? n37 : n14179;
  assign n14181 = pi16 ? n439 : n14180;
  assign n14182 = pi15 ? n14174 : n14181;
  assign n14183 = pi21 ? n569 : n8916;
  assign n14184 = pi20 ? n14183 : n32;
  assign n14185 = pi19 ? n14184 : n32;
  assign n14186 = pi18 ? n13291 : n14185;
  assign n14187 = pi17 ? n37 : n14186;
  assign n14188 = pi16 ? n439 : n14187;
  assign n14189 = pi19 ? n6373 : n11632;
  assign n14190 = pi21 ? n569 : n14168;
  assign n14191 = pi20 ? n14190 : n32;
  assign n14192 = pi19 ? n14191 : n32;
  assign n14193 = pi18 ? n14189 : n14192;
  assign n14194 = pi17 ? n37 : n14193;
  assign n14195 = pi16 ? n439 : n14194;
  assign n14196 = pi15 ? n14188 : n14195;
  assign n14197 = pi14 ? n14182 : n14196;
  assign n14198 = pi20 ? n37 : n3289;
  assign n14199 = pi19 ? n14198 : n13290;
  assign n14200 = pi18 ? n14199 : n14185;
  assign n14201 = pi17 ? n37 : n14200;
  assign n14202 = pi16 ? n439 : n14201;
  assign n14203 = pi21 ? n335 : n4902;
  assign n14204 = pi20 ? n605 : n14203;
  assign n14205 = pi19 ? n8867 : n14204;
  assign n14206 = pi21 ? n335 : n8486;
  assign n14207 = pi20 ? n14206 : n32;
  assign n14208 = pi19 ? n14207 : n32;
  assign n14209 = pi18 ? n14205 : n14208;
  assign n14210 = pi17 ? n37 : n14209;
  assign n14211 = pi16 ? n439 : n14210;
  assign n14212 = pi15 ? n14202 : n14211;
  assign n14213 = pi22 ? n363 : n2116;
  assign n14214 = pi21 ? n37 : n14213;
  assign n14215 = pi20 ? n37 : n14214;
  assign n14216 = pi19 ? n37 : n14215;
  assign n14217 = pi21 ? n3392 : n8486;
  assign n14218 = pi20 ? n14217 : n32;
  assign n14219 = pi19 ? n14218 : n32;
  assign n14220 = pi18 ? n14216 : n14219;
  assign n14221 = pi17 ? n37 : n14220;
  assign n14222 = pi16 ? n439 : n14221;
  assign n14223 = pi21 ? n233 : n2048;
  assign n14224 = pi20 ? n7705 : n14223;
  assign n14225 = pi19 ? n8928 : n14224;
  assign n14226 = pi21 ? n233 : n2320;
  assign n14227 = pi20 ? n14226 : n32;
  assign n14228 = pi19 ? n14227 : n32;
  assign n14229 = pi18 ? n14225 : n14228;
  assign n14230 = pi17 ? n37 : n14229;
  assign n14231 = pi16 ? n439 : n14230;
  assign n14232 = pi15 ? n14222 : n14231;
  assign n14233 = pi14 ? n14212 : n14232;
  assign n14234 = pi13 ? n14197 : n14233;
  assign n14235 = pi12 ? n14164 : n14234;
  assign n14236 = pi11 ? n14056 : n14235;
  assign n14237 = pi20 ? n37 : n6360;
  assign n14238 = pi21 ? n560 : n2048;
  assign n14239 = pi20 ? n37 : n14238;
  assign n14240 = pi19 ? n14237 : n14239;
  assign n14241 = pi18 ? n14240 : n13731;
  assign n14242 = pi17 ? n37 : n14241;
  assign n14243 = pi16 ? n439 : n14242;
  assign n14244 = pi15 ? n14243 : n13748;
  assign n14245 = pi23 ? n37 : n685;
  assign n14246 = pi22 ? n14245 : n37;
  assign n14247 = pi21 ? n14246 : n5015;
  assign n14248 = pi20 ? n37 : n14247;
  assign n14249 = pi19 ? n37 : n14248;
  assign n14250 = pi18 ? n14249 : n13762;
  assign n14251 = pi17 ? n37 : n14250;
  assign n14252 = pi16 ? n439 : n14251;
  assign n14253 = pi15 ? n14252 : n13765;
  assign n14254 = pi14 ? n14244 : n14253;
  assign n14255 = pi22 ? n363 : n686;
  assign n14256 = pi21 ? n14255 : n760;
  assign n14257 = pi20 ? n14256 : n32;
  assign n14258 = pi19 ? n14257 : n32;
  assign n14259 = pi18 ? n37 : n14258;
  assign n14260 = pi17 ? n37 : n14259;
  assign n14261 = pi16 ? n439 : n14260;
  assign n14262 = pi21 ? n685 : n5829;
  assign n14263 = pi20 ? n14262 : n32;
  assign n14264 = pi19 ? n14263 : n32;
  assign n14265 = pi18 ? n37 : n14264;
  assign n14266 = pi17 ? n37 : n14265;
  assign n14267 = pi16 ? n439 : n14266;
  assign n14268 = pi15 ? n14261 : n14267;
  assign n14269 = pi14 ? n13765 : n14268;
  assign n14270 = pi13 ? n14254 : n14269;
  assign n14271 = pi21 ? n6089 : n775;
  assign n14272 = pi20 ? n99 : n14271;
  assign n14273 = pi19 ? n99 : n14272;
  assign n14274 = pi18 ? n14273 : n13779;
  assign n14275 = pi17 ? n99 : n14274;
  assign n14276 = pi16 ? n744 : n14275;
  assign n14277 = pi22 ? n685 : n157;
  assign n14278 = pi21 ? n14277 : n157;
  assign n14279 = pi20 ? n1665 : n14278;
  assign n14280 = pi19 ? n99 : n14279;
  assign n14281 = pi18 ? n14280 : n13785;
  assign n14282 = pi17 ? n99 : n14281;
  assign n14283 = pi16 ? n744 : n14282;
  assign n14284 = pi15 ? n14276 : n14283;
  assign n14285 = pi20 ? n802 : n99;
  assign n14286 = pi19 ? n2255 : n14285;
  assign n14287 = pi18 ? n99 : n14286;
  assign n14288 = pi20 ? n99 : n6089;
  assign n14289 = pi19 ? n99 : n14288;
  assign n14290 = pi18 ? n14289 : n13785;
  assign n14291 = pi17 ? n14287 : n14290;
  assign n14292 = pi16 ? n744 : n14291;
  assign n14293 = pi21 ? n777 : n6461;
  assign n14294 = pi20 ? n99 : n14293;
  assign n14295 = pi21 ? n6089 : n99;
  assign n14296 = pi20 ? n14295 : n13948;
  assign n14297 = pi19 ? n14294 : n14296;
  assign n14298 = pi18 ? n99 : n14297;
  assign n14299 = pi18 ? n13389 : n7409;
  assign n14300 = pi17 ? n14298 : n14299;
  assign n14301 = pi16 ? n744 : n14300;
  assign n14302 = pi15 ? n14292 : n14301;
  assign n14303 = pi14 ? n14284 : n14302;
  assign n14304 = pi16 ? n7793 : n13802;
  assign n14305 = pi20 ? n1010 : n32;
  assign n14306 = pi19 ? n14305 : n32;
  assign n14307 = pi18 ? n157 : n14306;
  assign n14308 = pi17 ? n157 : n14307;
  assign n14309 = pi16 ? n7793 : n14308;
  assign n14310 = pi15 ? n14304 : n14309;
  assign n14311 = pi15 ? n13407 : n12513;
  assign n14312 = pi14 ? n14310 : n14311;
  assign n14313 = pi13 ? n14303 : n14312;
  assign n14314 = pi12 ? n14270 : n14313;
  assign n14315 = pi18 ? n139 : n13400;
  assign n14316 = pi17 ? n139 : n14315;
  assign n14317 = pi16 ? n915 : n14316;
  assign n14318 = pi20 ? n139 : n1008;
  assign n14319 = pi19 ? n14318 : n139;
  assign n14320 = pi18 ? n139 : n14319;
  assign n14321 = pi21 ? n7890 : n32;
  assign n14322 = pi20 ? n14321 : n32;
  assign n14323 = pi19 ? n14322 : n32;
  assign n14324 = pi18 ? n139 : n14323;
  assign n14325 = pi17 ? n14320 : n14324;
  assign n14326 = pi16 ? n915 : n14325;
  assign n14327 = pi21 ? n491 : n32;
  assign n14328 = pi20 ? n14327 : n32;
  assign n14329 = pi19 ? n14328 : n32;
  assign n14330 = pi18 ? n12590 : n14329;
  assign n14331 = pi17 ? n14320 : n14330;
  assign n14332 = pi16 ? n915 : n14331;
  assign n14333 = pi15 ? n14326 : n14332;
  assign n14334 = pi14 ? n14317 : n14333;
  assign n14335 = pi21 ? n4020 : n2319;
  assign n14336 = pi20 ? n316 : n14335;
  assign n14337 = pi19 ? n14336 : n316;
  assign n14338 = pi18 ? n14337 : n316;
  assign n14339 = pi17 ? n14338 : n6938;
  assign n14340 = pi16 ? n11772 : n14339;
  assign n14341 = pi16 ? n7883 : n6226;
  assign n14342 = pi21 ? n1044 : n316;
  assign n14343 = pi20 ? n3731 : n14342;
  assign n14344 = pi19 ? n14343 : n316;
  assign n14345 = pi18 ? n14344 : n316;
  assign n14346 = pi17 ? n14345 : n6225;
  assign n14347 = pi16 ? n13824 : n14346;
  assign n14348 = pi15 ? n14341 : n14347;
  assign n14349 = pi14 ? n14340 : n14348;
  assign n14350 = pi13 ? n14334 : n14349;
  assign n14351 = pi22 ? n204 : n706;
  assign n14352 = pi21 ? n14351 : n32;
  assign n14353 = pi20 ? n14352 : n32;
  assign n14354 = pi19 ? n14353 : n32;
  assign n14355 = pi18 ? n204 : n14354;
  assign n14356 = pi17 ? n13464 : n14355;
  assign n14357 = pi16 ? n13833 : n14356;
  assign n14358 = pi21 ? n37 : n1578;
  assign n14359 = pi20 ? n204 : n14358;
  assign n14360 = pi19 ? n14359 : n204;
  assign n14361 = pi18 ? n14360 : n204;
  assign n14362 = pi24 ? n13481 : n32;
  assign n14363 = pi23 ? n14362 : n32;
  assign n14364 = pi22 ? n204 : n14363;
  assign n14365 = pi21 ? n14364 : n32;
  assign n14366 = pi20 ? n14365 : n32;
  assign n14367 = pi19 ? n14366 : n32;
  assign n14368 = pi18 ? n204 : n14367;
  assign n14369 = pi17 ? n14361 : n14368;
  assign n14370 = pi16 ? n13846 : n14369;
  assign n14371 = pi15 ? n14357 : n14370;
  assign n14372 = pi21 ? n37 : n516;
  assign n14373 = pi20 ? n204 : n14372;
  assign n14374 = pi19 ? n14373 : n204;
  assign n14375 = pi18 ? n14374 : n204;
  assign n14376 = pi22 ? n4883 : n32;
  assign n14377 = pi21 ? n14376 : n32;
  assign n14378 = pi20 ? n14377 : n32;
  assign n14379 = pi19 ? n14378 : n32;
  assign n14380 = pi18 ? n204 : n14379;
  assign n14381 = pi17 ? n14375 : n14380;
  assign n14382 = pi16 ? n13846 : n14381;
  assign n14383 = pi21 ? n335 : n10684;
  assign n14384 = pi20 ? n335 : n14383;
  assign n14385 = pi19 ? n335 : n14384;
  assign n14386 = pi21 ? n13722 : n32;
  assign n14387 = pi20 ? n14386 : n32;
  assign n14388 = pi19 ? n14387 : n32;
  assign n14389 = pi18 ? n14385 : n14388;
  assign n14390 = pi17 ? n335 : n14389;
  assign n14391 = pi16 ? n2035 : n14390;
  assign n14392 = pi15 ? n14382 : n14391;
  assign n14393 = pi14 ? n14371 : n14392;
  assign n14394 = pi20 ? n335 : n577;
  assign n14395 = pi19 ? n14394 : n335;
  assign n14396 = pi18 ? n14395 : n335;
  assign n14397 = pi21 ? n12825 : n32;
  assign n14398 = pi20 ? n14397 : n32;
  assign n14399 = pi19 ? n14398 : n32;
  assign n14400 = pi18 ? n14385 : n14399;
  assign n14401 = pi17 ? n14396 : n14400;
  assign n14402 = pi16 ? n2035 : n14401;
  assign n14403 = pi22 ? n335 : n3935;
  assign n14404 = pi21 ? n335 : n14403;
  assign n14405 = pi20 ? n335 : n14404;
  assign n14406 = pi19 ? n335 : n14405;
  assign n14407 = pi18 ? n14406 : n6419;
  assign n14408 = pi17 ? n335 : n14407;
  assign n14409 = pi16 ? n10980 : n14408;
  assign n14410 = pi15 ? n14402 : n14409;
  assign n14411 = pi19 ? n8914 : n335;
  assign n14412 = pi18 ? n335 : n14411;
  assign n14413 = pi22 ? n335 : n3944;
  assign n14414 = pi21 ? n335 : n14413;
  assign n14415 = pi20 ? n335 : n14414;
  assign n14416 = pi19 ? n335 : n14415;
  assign n14417 = pi18 ? n14416 : n3342;
  assign n14418 = pi17 ? n14412 : n14417;
  assign n14419 = pi16 ? n10118 : n14418;
  assign n14420 = pi18 ? n13536 : n3342;
  assign n14421 = pi17 ? n13534 : n14420;
  assign n14422 = pi16 ? n13531 : n14421;
  assign n14423 = pi15 ? n14419 : n14422;
  assign n14424 = pi14 ? n14410 : n14423;
  assign n14425 = pi13 ? n14393 : n14424;
  assign n14426 = pi12 ? n14350 : n14425;
  assign n14427 = pi11 ? n14314 : n14426;
  assign n14428 = pi10 ? n14236 : n14427;
  assign n14429 = pi09 ? n13893 : n14428;
  assign n14430 = pi15 ? n32 : n13886;
  assign n14431 = pi16 ? n11011 : n13883;
  assign n14432 = pi15 ? n13887 : n14431;
  assign n14433 = pi14 ? n14430 : n14432;
  assign n14434 = pi13 ? n32 : n14433;
  assign n14435 = pi12 ? n32 : n14434;
  assign n14436 = pi11 ? n32 : n14435;
  assign n14437 = pi10 ? n32 : n14436;
  assign n14438 = pi16 ? n11885 : n13897;
  assign n14439 = pi16 ? n12689 : n13902;
  assign n14440 = pi15 ? n14438 : n14439;
  assign n14441 = pi16 ? n13561 : n13908;
  assign n14442 = pi20 ? n32 : n2443;
  assign n14443 = pi19 ? n32 : n14442;
  assign n14444 = pi18 ? n14443 : n37;
  assign n14445 = pi17 ? n32 : n14444;
  assign n14446 = pi16 ? n14445 : n13914;
  assign n14447 = pi15 ? n14441 : n14446;
  assign n14448 = pi14 ? n14440 : n14447;
  assign n14449 = pi20 ? n157 : n32;
  assign n14450 = pi19 ? n14449 : n32;
  assign n14451 = pi18 ? n157 : n14450;
  assign n14452 = pi17 ? n157 : n14451;
  assign n14453 = pi16 ? n13932 : n14452;
  assign n14454 = pi21 ? n716 : n168;
  assign n14455 = pi20 ? n32 : n14454;
  assign n14456 = pi19 ? n32 : n14455;
  assign n14457 = pi18 ? n14456 : n13945;
  assign n14458 = pi17 ? n32 : n14457;
  assign n14459 = pi20 ? n7818 : n787;
  assign n14460 = pi19 ? n13949 : n14459;
  assign n14461 = pi22 ? n157 : n112;
  assign n14462 = pi21 ? n14461 : n775;
  assign n14463 = pi20 ? n787 : n14462;
  assign n14464 = pi21 ? n165 : n157;
  assign n14465 = pi20 ? n14464 : n7823;
  assign n14466 = pi19 ? n14463 : n14465;
  assign n14467 = pi18 ? n14460 : n14466;
  assign n14468 = pi21 ? n157 : n3013;
  assign n14469 = pi20 ? n14468 : n32;
  assign n14470 = pi19 ? n14469 : n32;
  assign n14471 = pi18 ? n13958 : n14470;
  assign n14472 = pi17 ? n14467 : n14471;
  assign n14473 = pi16 ? n14458 : n14472;
  assign n14474 = pi15 ? n14453 : n14473;
  assign n14475 = pi14 ? n13927 : n14474;
  assign n14476 = pi13 ? n14448 : n14475;
  assign n14477 = pi22 ? n99 : n893;
  assign n14478 = pi21 ? n99 : n14477;
  assign n14479 = pi20 ? n14478 : n32;
  assign n14480 = pi19 ? n14479 : n32;
  assign n14481 = pi18 ? n99 : n14480;
  assign n14482 = pi17 ? n99 : n14481;
  assign n14483 = pi16 ? n801 : n14482;
  assign n14484 = pi23 ? n37 : n170;
  assign n14485 = pi22 ? n99 : n14484;
  assign n14486 = pi21 ? n99 : n14485;
  assign n14487 = pi20 ? n14486 : n32;
  assign n14488 = pi19 ? n14487 : n32;
  assign n14489 = pi18 ? n99 : n14488;
  assign n14490 = pi17 ? n99 : n14489;
  assign n14491 = pi16 ? n744 : n14490;
  assign n14492 = pi15 ? n14483 : n14491;
  assign n14493 = pi20 ? n1684 : n32;
  assign n14494 = pi19 ? n14493 : n32;
  assign n14495 = pi18 ? n99 : n14494;
  assign n14496 = pi17 ? n99 : n14495;
  assign n14497 = pi16 ? n721 : n14496;
  assign n14498 = pi21 ? n99 : n7395;
  assign n14499 = pi20 ? n14498 : n32;
  assign n14500 = pi19 ? n14499 : n32;
  assign n14501 = pi18 ? n99 : n14500;
  assign n14502 = pi17 ? n99 : n14501;
  assign n14503 = pi16 ? n801 : n14502;
  assign n14504 = pi15 ? n14497 : n14503;
  assign n14505 = pi14 ? n14492 : n14504;
  assign n14506 = pi22 ? n55 : n2160;
  assign n14507 = pi21 ? n14506 : n112;
  assign n14508 = pi20 ? n32 : n14507;
  assign n14509 = pi19 ? n32 : n14508;
  assign n14510 = pi21 ? n2175 : n2957;
  assign n14511 = pi20 ? n14510 : n5496;
  assign n14512 = pi21 ? n2156 : n2981;
  assign n14513 = pi21 ? n2156 : n2175;
  assign n14514 = pi20 ? n14512 : n14513;
  assign n14515 = pi19 ? n14511 : n14514;
  assign n14516 = pi18 ? n14509 : n14515;
  assign n14517 = pi17 ? n32 : n14516;
  assign n14518 = pi21 ? n2981 : n2156;
  assign n14519 = pi20 ? n2970 : n14518;
  assign n14520 = pi21 ? n2160 : n2156;
  assign n14521 = pi21 ? n2175 : n2156;
  assign n14522 = pi20 ? n14520 : n14521;
  assign n14523 = pi19 ? n14519 : n14522;
  assign n14524 = pi21 ? n37 : n2156;
  assign n14525 = pi20 ? n14524 : n5501;
  assign n14526 = pi21 ? n2175 : n112;
  assign n14527 = pi20 ? n14526 : n14521;
  assign n14528 = pi19 ? n14525 : n14527;
  assign n14529 = pi18 ? n14523 : n14528;
  assign n14530 = pi21 ? n2981 : n37;
  assign n14531 = pi20 ? n14530 : n2974;
  assign n14532 = pi20 ? n2974 : n2958;
  assign n14533 = pi19 ? n14531 : n14532;
  assign n14534 = pi22 ? n99 : n10720;
  assign n14535 = pi21 ? n2156 : n14534;
  assign n14536 = pi20 ? n14535 : n32;
  assign n14537 = pi19 ? n14536 : n32;
  assign n14538 = pi18 ? n14533 : n14537;
  assign n14539 = pi17 ? n14529 : n14538;
  assign n14540 = pi16 ? n14517 : n14539;
  assign n14541 = pi22 ? n139 : n3472;
  assign n14542 = pi21 ? n139 : n14541;
  assign n14543 = pi20 ? n14542 : n32;
  assign n14544 = pi19 ? n14543 : n32;
  assign n14545 = pi18 ? n13101 : n14544;
  assign n14546 = pi17 ? n13099 : n14545;
  assign n14547 = pi16 ? n14017 : n14546;
  assign n14548 = pi15 ? n14540 : n14547;
  assign n14549 = pi21 ? n37 : n1785;
  assign n14550 = pi20 ? n14549 : n32;
  assign n14551 = pi19 ? n14550 : n32;
  assign n14552 = pi18 ? n37 : n14551;
  assign n14553 = pi17 ? n37 : n14552;
  assign n14554 = pi16 ? n439 : n14553;
  assign n14555 = pi21 ? n1711 : n1785;
  assign n14556 = pi20 ? n14555 : n32;
  assign n14557 = pi19 ? n14556 : n32;
  assign n14558 = pi18 ? n14046 : n14557;
  assign n14559 = pi17 ? n14042 : n14558;
  assign n14560 = pi16 ? n439 : n14559;
  assign n14561 = pi15 ? n14554 : n14560;
  assign n14562 = pi14 ? n14548 : n14561;
  assign n14563 = pi13 ? n14505 : n14562;
  assign n14564 = pi12 ? n14476 : n14563;
  assign n14565 = pi21 ? n1696 : n1785;
  assign n14566 = pi20 ? n14565 : n32;
  assign n14567 = pi19 ? n14566 : n32;
  assign n14568 = pi18 ? n14070 : n14567;
  assign n14569 = pi17 ? n14065 : n14568;
  assign n14570 = pi16 ? n439 : n14569;
  assign n14571 = pi20 ? n8209 : n1705;
  assign n14572 = pi19 ? n8743 : n14571;
  assign n14573 = pi21 ? n1696 : n295;
  assign n14574 = pi20 ? n14573 : n5269;
  assign n14575 = pi19 ? n14574 : n1743;
  assign n14576 = pi18 ? n14572 : n14575;
  assign n14577 = pi21 ? n1531 : n1043;
  assign n14578 = pi20 ? n14577 : n1715;
  assign n14579 = pi19 ? n13646 : n14578;
  assign n14580 = pi21 ? n1711 : n14085;
  assign n14581 = pi20 ? n14580 : n32;
  assign n14582 = pi19 ? n14581 : n32;
  assign n14583 = pi18 ? n14579 : n14582;
  assign n14584 = pi17 ? n14576 : n14583;
  assign n14585 = pi16 ? n439 : n14584;
  assign n14586 = pi15 ? n14570 : n14585;
  assign n14587 = pi14 ? n14586 : n14113;
  assign n14588 = pi20 ? n37 : n13217;
  assign n14589 = pi19 ? n37 : n14588;
  assign n14590 = pi18 ? n37 : n14589;
  assign n14591 = pi21 ? n204 : n485;
  assign n14592 = pi20 ? n14126 : n14591;
  assign n14593 = pi19 ? n14127 : n14592;
  assign n14594 = pi21 ? n522 : n6194;
  assign n14595 = pi20 ? n14594 : n32;
  assign n14596 = pi19 ? n14595 : n32;
  assign n14597 = pi18 ? n14593 : n14596;
  assign n14598 = pi17 ? n14590 : n14597;
  assign n14599 = pi16 ? n439 : n14598;
  assign n14600 = pi15 ? n14122 : n14599;
  assign n14601 = pi21 ? n522 : n485;
  assign n14602 = pi20 ? n14601 : n14591;
  assign n14603 = pi19 ? n14141 : n14602;
  assign n14604 = pi21 ? n522 : n6270;
  assign n14605 = pi20 ? n14604 : n32;
  assign n14606 = pi19 ? n14605 : n32;
  assign n14607 = pi18 ? n14603 : n14606;
  assign n14608 = pi17 ? n12414 : n14607;
  assign n14609 = pi16 ? n439 : n14608;
  assign n14610 = pi18 ? n37 : n8868;
  assign n14611 = pi21 ? n4938 : n1943;
  assign n14612 = pi21 ? n4990 : n1943;
  assign n14613 = pi20 ? n14611 : n14612;
  assign n14614 = pi21 ? n335 : n583;
  assign n14615 = pi20 ? n14614 : n4980;
  assign n14616 = pi19 ? n14613 : n14615;
  assign n14617 = pi21 ? n1943 : n14155;
  assign n14618 = pi20 ? n14617 : n32;
  assign n14619 = pi19 ? n14618 : n32;
  assign n14620 = pi18 ? n14616 : n14619;
  assign n14621 = pi17 ? n14610 : n14620;
  assign n14622 = pi16 ? n439 : n14621;
  assign n14623 = pi15 ? n14609 : n14622;
  assign n14624 = pi14 ? n14600 : n14623;
  assign n14625 = pi13 ? n14587 : n14624;
  assign n14626 = pi25 ? n232 : n32;
  assign n14627 = pi24 ? n233 : n14626;
  assign n14628 = pi23 ? n14627 : n32;
  assign n14629 = pi22 ? n233 : n14628;
  assign n14630 = pi21 ? n569 : n14629;
  assign n14631 = pi20 ? n14630 : n32;
  assign n14632 = pi19 ? n14631 : n32;
  assign n14633 = pi18 ? n14189 : n14632;
  assign n14634 = pi17 ? n37 : n14633;
  assign n14635 = pi16 ? n439 : n14634;
  assign n14636 = pi15 ? n14188 : n14635;
  assign n14637 = pi14 ? n14182 : n14636;
  assign n14638 = pi21 ? n569 : n8272;
  assign n14639 = pi20 ? n14638 : n32;
  assign n14640 = pi19 ? n14639 : n32;
  assign n14641 = pi18 ? n14199 : n14640;
  assign n14642 = pi17 ? n37 : n14641;
  assign n14643 = pi16 ? n439 : n14642;
  assign n14644 = pi21 ? n335 : n696;
  assign n14645 = pi20 ? n14644 : n32;
  assign n14646 = pi19 ? n14645 : n32;
  assign n14647 = pi18 ? n14205 : n14646;
  assign n14648 = pi17 ? n37 : n14647;
  assign n14649 = pi16 ? n439 : n14648;
  assign n14650 = pi15 ? n14643 : n14649;
  assign n14651 = pi21 ? n3392 : n696;
  assign n14652 = pi20 ? n14651 : n32;
  assign n14653 = pi19 ? n14652 : n32;
  assign n14654 = pi18 ? n14216 : n14653;
  assign n14655 = pi17 ? n37 : n14654;
  assign n14656 = pi16 ? n439 : n14655;
  assign n14657 = pi21 ? n233 : n3523;
  assign n14658 = pi20 ? n14657 : n32;
  assign n14659 = pi19 ? n14658 : n32;
  assign n14660 = pi18 ? n14225 : n14659;
  assign n14661 = pi17 ? n37 : n14660;
  assign n14662 = pi16 ? n439 : n14661;
  assign n14663 = pi15 ? n14656 : n14662;
  assign n14664 = pi14 ? n14650 : n14663;
  assign n14665 = pi13 ? n14637 : n14664;
  assign n14666 = pi12 ? n14625 : n14665;
  assign n14667 = pi11 ? n14564 : n14666;
  assign n14668 = pi21 ? n2091 : n5758;
  assign n14669 = pi20 ? n14668 : n32;
  assign n14670 = pi19 ? n14669 : n32;
  assign n14671 = pi18 ? n14240 : n14670;
  assign n14672 = pi17 ? n37 : n14671;
  assign n14673 = pi16 ? n439 : n14672;
  assign n14674 = pi21 ? n233 : n7034;
  assign n14675 = pi20 ? n14674 : n32;
  assign n14676 = pi19 ? n14675 : n32;
  assign n14677 = pi18 ? n13338 : n14676;
  assign n14678 = pi17 ? n37 : n14677;
  assign n14679 = pi16 ? n439 : n14678;
  assign n14680 = pi15 ? n14673 : n14679;
  assign n14681 = pi21 ? n2106 : n7723;
  assign n14682 = pi20 ? n14681 : n32;
  assign n14683 = pi19 ? n14682 : n32;
  assign n14684 = pi18 ? n14249 : n14683;
  assign n14685 = pi17 ? n37 : n14684;
  assign n14686 = pi16 ? n439 : n14685;
  assign n14687 = pi18 ? n37 : n14683;
  assign n14688 = pi17 ? n37 : n14687;
  assign n14689 = pi16 ? n439 : n14688;
  assign n14690 = pi15 ? n14686 : n14689;
  assign n14691 = pi14 ? n14680 : n14690;
  assign n14692 = pi21 ? n363 : n7723;
  assign n14693 = pi20 ? n14692 : n32;
  assign n14694 = pi19 ? n14693 : n32;
  assign n14695 = pi18 ? n37 : n14694;
  assign n14696 = pi17 ? n37 : n14695;
  assign n14697 = pi16 ? n439 : n14696;
  assign n14698 = pi21 ? n685 : n7048;
  assign n14699 = pi20 ? n14698 : n32;
  assign n14700 = pi19 ? n14699 : n32;
  assign n14701 = pi18 ? n37 : n14700;
  assign n14702 = pi17 ? n37 : n14701;
  assign n14703 = pi16 ? n439 : n14702;
  assign n14704 = pi15 ? n14697 : n14703;
  assign n14705 = pi14 ? n14689 : n14704;
  assign n14706 = pi13 ? n14691 : n14705;
  assign n14707 = pi21 ? n6461 : n760;
  assign n14708 = pi20 ? n14707 : n32;
  assign n14709 = pi19 ? n14708 : n32;
  assign n14710 = pi18 ? n14273 : n14709;
  assign n14711 = pi17 ? n99 : n14710;
  assign n14712 = pi16 ? n721 : n14711;
  assign n14713 = pi21 ? n6461 : n882;
  assign n14714 = pi20 ? n14713 : n32;
  assign n14715 = pi19 ? n14714 : n32;
  assign n14716 = pi18 ? n14280 : n14715;
  assign n14717 = pi17 ? n99 : n14716;
  assign n14718 = pi16 ? n721 : n14717;
  assign n14719 = pi15 ? n14712 : n14718;
  assign n14720 = pi18 ? n14289 : n14715;
  assign n14721 = pi17 ? n14287 : n14720;
  assign n14722 = pi16 ? n721 : n14721;
  assign n14723 = pi21 ? n685 : n928;
  assign n14724 = pi20 ? n14723 : n32;
  assign n14725 = pi19 ? n14724 : n32;
  assign n14726 = pi18 ? n13389 : n14725;
  assign n14727 = pi17 ? n14298 : n14726;
  assign n14728 = pi16 ? n721 : n14727;
  assign n14729 = pi15 ? n14722 : n14728;
  assign n14730 = pi14 ? n14719 : n14729;
  assign n14731 = pi18 ? n157 : n14725;
  assign n14732 = pi17 ? n157 : n14731;
  assign n14733 = pi16 ? n5910 : n14732;
  assign n14734 = pi16 ? n5910 : n14308;
  assign n14735 = pi15 ? n14733 : n14734;
  assign n14736 = pi18 ? n99 : n14306;
  assign n14737 = pi17 ? n99 : n14736;
  assign n14738 = pi16 ? n744 : n14737;
  assign n14739 = pi16 ? n744 : n12923;
  assign n14740 = pi15 ? n14738 : n14739;
  assign n14741 = pi14 ? n14735 : n14740;
  assign n14742 = pi13 ? n14730 : n14741;
  assign n14743 = pi12 ? n14706 : n14742;
  assign n14744 = pi18 ? n139 : n14306;
  assign n14745 = pi17 ? n139 : n14744;
  assign n14746 = pi16 ? n915 : n14745;
  assign n14747 = pi22 ? n316 : n1070;
  assign n14748 = pi21 ? n14747 : n32;
  assign n14749 = pi20 ? n14748 : n32;
  assign n14750 = pi19 ? n14749 : n32;
  assign n14751 = pi18 ? n139 : n14750;
  assign n14752 = pi17 ? n14320 : n14751;
  assign n14753 = pi16 ? n915 : n14752;
  assign n14754 = pi20 ? n1101 : n32;
  assign n14755 = pi19 ? n14754 : n32;
  assign n14756 = pi18 ? n12590 : n14755;
  assign n14757 = pi17 ? n14320 : n14756;
  assign n14758 = pi16 ? n2291 : n14757;
  assign n14759 = pi15 ? n14753 : n14758;
  assign n14760 = pi14 ? n14746 : n14759;
  assign n14761 = pi22 ? n962 : n316;
  assign n14762 = pi21 ? n14761 : n316;
  assign n14763 = pi20 ? n32 : n14762;
  assign n14764 = pi19 ? n32 : n14763;
  assign n14765 = pi18 ? n14764 : n316;
  assign n14766 = pi17 ? n32 : n14765;
  assign n14767 = pi18 ? n316 : n13400;
  assign n14768 = pi17 ? n14338 : n14767;
  assign n14769 = pi16 ? n14766 : n14768;
  assign n14770 = pi16 ? n7883 : n6939;
  assign n14771 = pi21 ? n2395 : n316;
  assign n14772 = pi20 ? n3731 : n14771;
  assign n14773 = pi19 ? n14772 : n316;
  assign n14774 = pi18 ? n14773 : n316;
  assign n14775 = pi17 ? n14774 : n6938;
  assign n14776 = pi16 ? n13824 : n14775;
  assign n14777 = pi15 ? n14770 : n14776;
  assign n14778 = pi14 ? n14769 : n14777;
  assign n14779 = pi13 ? n14760 : n14778;
  assign n14780 = pi18 ? n204 : n13431;
  assign n14781 = pi17 ? n13464 : n14780;
  assign n14782 = pi16 ? n13833 : n14781;
  assign n14783 = pi17 ? n14361 : n14355;
  assign n14784 = pi16 ? n13846 : n14783;
  assign n14785 = pi15 ? n14782 : n14784;
  assign n14786 = pi20 ? n204 : n1912;
  assign n14787 = pi19 ? n14786 : n204;
  assign n14788 = pi18 ? n14787 : n204;
  assign n14789 = pi22 ? n4079 : n706;
  assign n14790 = pi21 ? n14789 : n32;
  assign n14791 = pi20 ? n14790 : n32;
  assign n14792 = pi19 ? n14791 : n32;
  assign n14793 = pi18 ? n204 : n14792;
  assign n14794 = pi17 ? n14788 : n14793;
  assign n14795 = pi16 ? n13846 : n14794;
  assign n14796 = pi18 ? n14385 : n7044;
  assign n14797 = pi17 ? n335 : n14796;
  assign n14798 = pi16 ? n2035 : n14797;
  assign n14799 = pi15 ? n14795 : n14798;
  assign n14800 = pi14 ? n14785 : n14799;
  assign n14801 = pi18 ? n14385 : n4104;
  assign n14802 = pi17 ? n14396 : n14801;
  assign n14803 = pi16 ? n2035 : n14802;
  assign n14804 = pi15 ? n14803 : n14409;
  assign n14805 = pi14 ? n14804 : n14423;
  assign n14806 = pi13 ? n14800 : n14805;
  assign n14807 = pi12 ? n14779 : n14806;
  assign n14808 = pi11 ? n14743 : n14807;
  assign n14809 = pi10 ? n14667 : n14808;
  assign n14810 = pi09 ? n14437 : n14809;
  assign n14811 = pi08 ? n14429 : n14810;
  assign n14812 = pi07 ? n13879 : n14811;
  assign n14813 = pi06 ? n13009 : n14812;
  assign n14814 = pi05 ? n11364 : n14813;
  assign n14815 = pi20 ? n37 : n2934;
  assign n14816 = pi19 ? n14815 : n32;
  assign n14817 = pi18 ? n37 : n14816;
  assign n14818 = pi17 ? n37 : n14817;
  assign n14819 = pi16 ? n2461 : n14818;
  assign n14820 = pi15 ? n32 : n14819;
  assign n14821 = pi16 ? n10154 : n14818;
  assign n14822 = pi16 ? n11011 : n14818;
  assign n14823 = pi15 ? n14821 : n14822;
  assign n14824 = pi14 ? n14820 : n14823;
  assign n14825 = pi13 ? n32 : n14824;
  assign n14826 = pi12 ? n32 : n14825;
  assign n14827 = pi11 ? n32 : n14826;
  assign n14828 = pi10 ? n32 : n14827;
  assign n14829 = pi21 ? n8008 : n32;
  assign n14830 = pi20 ? n99 : n14829;
  assign n14831 = pi19 ? n14830 : n32;
  assign n14832 = pi18 ? n37 : n14831;
  assign n14833 = pi17 ? n37 : n14832;
  assign n14834 = pi16 ? n11885 : n14833;
  assign n14835 = pi21 ? n8015 : n32;
  assign n14836 = pi20 ? n99 : n14835;
  assign n14837 = pi19 ? n14836 : n32;
  assign n14838 = pi18 ? n37 : n14837;
  assign n14839 = pi17 ? n37 : n14838;
  assign n14840 = pi16 ? n12689 : n14839;
  assign n14841 = pi15 ? n14834 : n14840;
  assign n14842 = pi19 ? n37 : n99;
  assign n14843 = pi18 ? n14842 : n99;
  assign n14844 = pi21 ? n37 : n99;
  assign n14845 = pi19 ? n99 : n14844;
  assign n14846 = pi21 ? n99 : n139;
  assign n14847 = pi21 ? n8557 : n32;
  assign n14848 = pi20 ? n14846 : n14847;
  assign n14849 = pi19 ? n14848 : n32;
  assign n14850 = pi18 ? n14845 : n14849;
  assign n14851 = pi17 ? n14843 : n14850;
  assign n14852 = pi16 ? n13561 : n14851;
  assign n14853 = pi21 ? n92 : n99;
  assign n14854 = pi20 ? n32 : n14853;
  assign n14855 = pi19 ? n32 : n14854;
  assign n14856 = pi18 ? n14855 : n99;
  assign n14857 = pi17 ? n32 : n14856;
  assign n14858 = pi20 ? n14846 : n32;
  assign n14859 = pi19 ? n14858 : n32;
  assign n14860 = pi18 ? n99 : n14859;
  assign n14861 = pi17 ? n99 : n14860;
  assign n14862 = pi16 ? n14857 : n14861;
  assign n14863 = pi15 ? n14852 : n14862;
  assign n14864 = pi14 ? n14841 : n14863;
  assign n14865 = pi22 ? n99 : n335;
  assign n14866 = pi21 ? n99 : n14865;
  assign n14867 = pi20 ? n14866 : n32;
  assign n14868 = pi19 ? n14867 : n32;
  assign n14869 = pi18 ? n99 : n14868;
  assign n14870 = pi17 ? n99 : n14869;
  assign n14871 = pi16 ? n3065 : n14870;
  assign n14872 = pi20 ? n1658 : n32;
  assign n14873 = pi19 ? n14872 : n32;
  assign n14874 = pi18 ? n99 : n14873;
  assign n14875 = pi17 ? n99 : n14874;
  assign n14876 = pi16 ? n801 : n14875;
  assign n14877 = pi15 ? n14871 : n14876;
  assign n14878 = pi21 ? n3060 : n37;
  assign n14879 = pi20 ? n32 : n14878;
  assign n14880 = pi19 ? n32 : n14879;
  assign n14881 = pi18 ? n14880 : n37;
  assign n14882 = pi17 ? n32 : n14881;
  assign n14883 = pi19 ? n37 : n2970;
  assign n14884 = pi22 ? n37 : n164;
  assign n14885 = pi21 ? n14884 : n2175;
  assign n14886 = pi20 ? n14885 : n2970;
  assign n14887 = pi21 ? n218 : n37;
  assign n14888 = pi19 ? n14886 : n14887;
  assign n14889 = pi18 ? n14883 : n14888;
  assign n14890 = pi21 ? n157 : n2981;
  assign n14891 = pi20 ? n5878 : n14890;
  assign n14892 = pi21 ? n6433 : n218;
  assign n14893 = pi20 ? n14892 : n3039;
  assign n14894 = pi19 ? n14891 : n14893;
  assign n14895 = pi20 ? n6508 : n32;
  assign n14896 = pi19 ? n14895 : n32;
  assign n14897 = pi18 ? n14894 : n14896;
  assign n14898 = pi17 ? n14889 : n14897;
  assign n14899 = pi16 ? n14882 : n14898;
  assign n14900 = pi21 ? n12705 : n99;
  assign n14901 = pi20 ? n14900 : n99;
  assign n14902 = pi19 ? n14901 : n99;
  assign n14903 = pi18 ? n99 : n14902;
  assign n14904 = pi21 ? n12705 : n5877;
  assign n14905 = pi20 ? n14904 : n99;
  assign n14906 = pi21 ? n14477 : n99;
  assign n14907 = pi20 ? n14906 : n99;
  assign n14908 = pi19 ? n14905 : n14907;
  assign n14909 = pi21 ? n2998 : n14477;
  assign n14910 = pi20 ? n14909 : n32;
  assign n14911 = pi19 ? n14910 : n32;
  assign n14912 = pi18 ? n14908 : n14911;
  assign n14913 = pi17 ? n14903 : n14912;
  assign n14914 = pi16 ? n744 : n14913;
  assign n14915 = pi15 ? n14899 : n14914;
  assign n14916 = pi14 ? n14877 : n14915;
  assign n14917 = pi13 ? n14864 : n14916;
  assign n14918 = pi21 ? n99 : n214;
  assign n14919 = pi20 ? n14918 : n32;
  assign n14920 = pi19 ? n14919 : n32;
  assign n14921 = pi18 ? n99 : n14920;
  assign n14922 = pi17 ? n99 : n14921;
  assign n14923 = pi16 ? n744 : n14922;
  assign n14924 = pi15 ? n14923 : n14483;
  assign n14925 = pi18 ? n742 : n4584;
  assign n14926 = pi17 ? n32 : n14925;
  assign n14927 = pi21 ? n99 : n6823;
  assign n14928 = pi20 ? n14927 : n32;
  assign n14929 = pi19 ? n14928 : n32;
  assign n14930 = pi18 ? n99 : n14929;
  assign n14931 = pi17 ? n99 : n14930;
  assign n14932 = pi16 ? n14926 : n14931;
  assign n14933 = pi19 ? n5134 : n99;
  assign n14934 = pi18 ? n719 : n14933;
  assign n14935 = pi17 ? n32 : n14934;
  assign n14936 = pi22 ? n99 : n11047;
  assign n14937 = pi21 ? n99 : n14936;
  assign n14938 = pi20 ? n14937 : n32;
  assign n14939 = pi19 ? n14938 : n32;
  assign n14940 = pi18 ? n99 : n14939;
  assign n14941 = pi17 ? n99 : n14940;
  assign n14942 = pi16 ? n14935 : n14941;
  assign n14943 = pi15 ? n14932 : n14942;
  assign n14944 = pi14 ? n14924 : n14943;
  assign n14945 = pi21 ? n1564 : n37;
  assign n14946 = pi20 ? n32 : n14945;
  assign n14947 = pi19 ? n32 : n14946;
  assign n14948 = pi20 ? n5269 : n1747;
  assign n14949 = pi19 ? n37 : n14948;
  assign n14950 = pi18 ? n14947 : n14949;
  assign n14951 = pi17 ? n32 : n14950;
  assign n14952 = pi22 ? n139 : n6833;
  assign n14953 = pi21 ? n139 : n14952;
  assign n14954 = pi20 ? n14953 : n32;
  assign n14955 = pi19 ? n14954 : n32;
  assign n14956 = pi18 ? n139 : n14955;
  assign n14957 = pi17 ? n139 : n14956;
  assign n14958 = pi16 ? n14951 : n14957;
  assign n14959 = pi21 ? n8143 : n37;
  assign n14960 = pi20 ? n32 : n14959;
  assign n14961 = pi19 ? n32 : n14960;
  assign n14962 = pi20 ? n947 : n139;
  assign n14963 = pi19 ? n37 : n14962;
  assign n14964 = pi18 ? n14961 : n14963;
  assign n14965 = pi17 ? n32 : n14964;
  assign n14966 = pi18 ? n139 : n14544;
  assign n14967 = pi17 ? n139 : n14966;
  assign n14968 = pi16 ? n14965 : n14967;
  assign n14969 = pi15 ? n14958 : n14968;
  assign n14970 = pi20 ? n5269 : n2513;
  assign n14971 = pi19 ? n8743 : n14970;
  assign n14972 = pi20 ? n1738 : n2513;
  assign n14973 = pi20 ? n2513 : n5273;
  assign n14974 = pi19 ? n14972 : n14973;
  assign n14975 = pi18 ? n14971 : n14974;
  assign n14976 = pi20 ? n2521 : n1715;
  assign n14977 = pi19 ? n139 : n14976;
  assign n14978 = pi22 ? n139 : n6380;
  assign n14979 = pi21 ? n1711 : n14978;
  assign n14980 = pi20 ? n14979 : n1822;
  assign n14981 = pi19 ? n14980 : n32;
  assign n14982 = pi18 ? n14977 : n14981;
  assign n14983 = pi17 ? n14975 : n14982;
  assign n14984 = pi16 ? n439 : n14983;
  assign n14985 = pi21 ? n297 : n1211;
  assign n14986 = pi20 ? n13121 : n14985;
  assign n14987 = pi19 ? n37 : n14986;
  assign n14988 = pi21 ? n297 : n1531;
  assign n14989 = pi20 ? n14988 : n942;
  assign n14990 = pi19 ? n14989 : n139;
  assign n14991 = pi18 ? n14987 : n14990;
  assign n14992 = pi21 ? n139 : n14978;
  assign n14993 = pi20 ? n14992 : n1822;
  assign n14994 = pi19 ? n14993 : n32;
  assign n14995 = pi18 ? n139 : n14994;
  assign n14996 = pi17 ? n14991 : n14995;
  assign n14997 = pi16 ? n439 : n14996;
  assign n14998 = pi15 ? n14984 : n14997;
  assign n14999 = pi14 ? n14969 : n14998;
  assign n15000 = pi13 ? n14944 : n14999;
  assign n15001 = pi12 ? n14917 : n15000;
  assign n15002 = pi20 ? n37 : n3104;
  assign n15003 = pi19 ? n37 : n15002;
  assign n15004 = pi20 ? n37 : n3645;
  assign n15005 = pi19 ? n15004 : n139;
  assign n15006 = pi18 ? n15003 : n15005;
  assign n15007 = pi22 ? n139 : n705;
  assign n15008 = pi21 ? n139 : n15007;
  assign n15009 = pi20 ? n15008 : n1822;
  assign n15010 = pi19 ? n15009 : n32;
  assign n15011 = pi18 ? n139 : n15010;
  assign n15012 = pi17 ? n15006 : n15011;
  assign n15013 = pi16 ? n439 : n15012;
  assign n15014 = pi19 ? n3083 : n3104;
  assign n15015 = pi18 ? n374 : n15014;
  assign n15016 = pi17 ? n32 : n15015;
  assign n15017 = pi20 ? n3104 : n820;
  assign n15018 = pi20 ? n297 : n3090;
  assign n15019 = pi19 ? n15017 : n15018;
  assign n15020 = pi20 ? n3104 : n947;
  assign n15021 = pi19 ? n15020 : n9769;
  assign n15022 = pi18 ? n15019 : n15021;
  assign n15023 = pi20 ? n1786 : n32;
  assign n15024 = pi19 ? n15023 : n32;
  assign n15025 = pi18 ? n139 : n15024;
  assign n15026 = pi17 ? n15022 : n15025;
  assign n15027 = pi16 ? n15016 : n15026;
  assign n15028 = pi15 ? n15013 : n15027;
  assign n15029 = pi19 ? n37 : n8765;
  assign n15030 = pi18 ? n37 : n15029;
  assign n15031 = pi17 ? n15030 : n15025;
  assign n15032 = pi16 ? n439 : n15031;
  assign n15033 = pi20 ? n1003 : n297;
  assign n15034 = pi19 ? n15033 : n3086;
  assign n15035 = pi18 ? n374 : n15034;
  assign n15036 = pi17 ? n32 : n15035;
  assign n15037 = pi20 ? n997 : n820;
  assign n15038 = pi19 ? n13168 : n15037;
  assign n15039 = pi20 ? n3104 : n941;
  assign n15040 = pi19 ? n15039 : n1806;
  assign n15041 = pi18 ? n15038 : n15040;
  assign n15042 = pi21 ? n139 : n8175;
  assign n15043 = pi20 ? n15042 : n32;
  assign n15044 = pi19 ? n15043 : n32;
  assign n15045 = pi18 ? n139 : n15044;
  assign n15046 = pi17 ? n15041 : n15045;
  assign n15047 = pi16 ? n15036 : n15046;
  assign n15048 = pi15 ? n15032 : n15047;
  assign n15049 = pi14 ? n15028 : n15048;
  assign n15050 = pi22 ? n37 : n9827;
  assign n15051 = pi21 ? n3073 : n15050;
  assign n15052 = pi20 ? n37 : n15051;
  assign n15053 = pi19 ? n37 : n15052;
  assign n15054 = pi18 ? n37 : n15053;
  assign n15055 = pi22 ? n9827 : n295;
  assign n15056 = pi21 ? n6676 : n15055;
  assign n15057 = pi22 ? n204 : n9827;
  assign n15058 = pi21 ? n15057 : n15055;
  assign n15059 = pi20 ? n15056 : n15058;
  assign n15060 = pi22 ? n9827 : n204;
  assign n15061 = pi21 ? n9126 : n15060;
  assign n15062 = pi20 ? n15058 : n15061;
  assign n15063 = pi19 ? n15059 : n15062;
  assign n15064 = pi21 ? n9827 : n7621;
  assign n15065 = pi20 ? n15064 : n32;
  assign n15066 = pi19 ? n15065 : n32;
  assign n15067 = pi18 ? n15063 : n15066;
  assign n15068 = pi17 ? n15054 : n15067;
  assign n15069 = pi16 ? n439 : n15068;
  assign n15070 = pi18 ? n37 : n7677;
  assign n15071 = pi20 ? n335 : n1084;
  assign n15072 = pi20 ? n1084 : n3311;
  assign n15073 = pi19 ? n15071 : n15072;
  assign n15074 = pi22 ? n204 : n8198;
  assign n15075 = pi21 ? n335 : n15074;
  assign n15076 = pi20 ? n15075 : n32;
  assign n15077 = pi19 ? n15076 : n32;
  assign n15078 = pi18 ? n15073 : n15077;
  assign n15079 = pi17 ? n15070 : n15078;
  assign n15080 = pi16 ? n439 : n15079;
  assign n15081 = pi15 ? n15069 : n15080;
  assign n15082 = pi19 ? n10681 : n335;
  assign n15083 = pi21 ? n335 : n7597;
  assign n15084 = pi20 ? n15083 : n32;
  assign n15085 = pi19 ? n15084 : n32;
  assign n15086 = pi18 ? n15082 : n15085;
  assign n15087 = pi17 ? n37 : n15086;
  assign n15088 = pi16 ? n439 : n15087;
  assign n15089 = pi22 ? n335 : n1159;
  assign n15090 = pi21 ? n335 : n15089;
  assign n15091 = pi20 ? n15090 : n32;
  assign n15092 = pi19 ? n15091 : n32;
  assign n15093 = pi18 ? n12629 : n15092;
  assign n15094 = pi17 ? n37 : n15093;
  assign n15095 = pi16 ? n439 : n15094;
  assign n15096 = pi15 ? n15088 : n15095;
  assign n15097 = pi14 ? n15081 : n15096;
  assign n15098 = pi13 ? n15049 : n15097;
  assign n15099 = pi19 ? n7685 : n335;
  assign n15100 = pi22 ? n335 : n1388;
  assign n15101 = pi21 ? n335 : n15100;
  assign n15102 = pi20 ? n15101 : n32;
  assign n15103 = pi19 ? n15102 : n32;
  assign n15104 = pi18 ? n15099 : n15103;
  assign n15105 = pi17 ? n37 : n15104;
  assign n15106 = pi16 ? n439 : n15105;
  assign n15107 = pi23 ? n37 : n6960;
  assign n15108 = pi22 ? n15107 : n1388;
  assign n15109 = pi21 ? n37 : n15108;
  assign n15110 = pi20 ? n15109 : n32;
  assign n15111 = pi19 ? n15110 : n32;
  assign n15112 = pi18 ? n9381 : n15111;
  assign n15113 = pi17 ? n37 : n15112;
  assign n15114 = pi16 ? n439 : n15113;
  assign n15115 = pi15 ? n15106 : n15114;
  assign n15116 = pi21 ? n569 : n4975;
  assign n15117 = pi20 ? n568 : n15116;
  assign n15118 = pi19 ? n37 : n15117;
  assign n15119 = pi22 ? n10730 : n759;
  assign n15120 = pi21 ? n570 : n15119;
  assign n15121 = pi20 ? n15120 : n32;
  assign n15122 = pi19 ? n15121 : n32;
  assign n15123 = pi18 ? n15118 : n15122;
  assign n15124 = pi17 ? n37 : n15123;
  assign n15125 = pi16 ? n439 : n15124;
  assign n15126 = pi15 ? n15114 : n15125;
  assign n15127 = pi14 ? n15115 : n15126;
  assign n15128 = pi19 ? n37 : n3285;
  assign n15129 = pi18 ? n37 : n15128;
  assign n15130 = pi19 ? n8802 : n639;
  assign n15131 = pi21 ? n1920 : n7668;
  assign n15132 = pi20 ? n15131 : n32;
  assign n15133 = pi19 ? n15132 : n32;
  assign n15134 = pi18 ? n15130 : n15133;
  assign n15135 = pi17 ? n15129 : n15134;
  assign n15136 = pi16 ? n439 : n15135;
  assign n15137 = pi20 ? n3289 : n37;
  assign n15138 = pi19 ? n37 : n15137;
  assign n15139 = pi18 ? n37 : n15138;
  assign n15140 = pi21 ? n580 : n4973;
  assign n15141 = pi20 ? n15140 : n2019;
  assign n15142 = pi19 ? n8802 : n15141;
  assign n15143 = pi22 ? n566 : n559;
  assign n15144 = pi21 ? n15143 : n8916;
  assign n15145 = pi20 ? n15144 : n32;
  assign n15146 = pi19 ? n15145 : n32;
  assign n15147 = pi18 ? n15142 : n15146;
  assign n15148 = pi17 ? n15139 : n15147;
  assign n15149 = pi16 ? n439 : n15148;
  assign n15150 = pi15 ? n15136 : n15149;
  assign n15151 = pi21 ? n2091 : n2707;
  assign n15152 = pi20 ? n37 : n15151;
  assign n15153 = pi19 ? n37 : n15152;
  assign n15154 = pi21 ? n2091 : n8916;
  assign n15155 = pi20 ? n15154 : n32;
  assign n15156 = pi19 ? n15155 : n32;
  assign n15157 = pi18 ? n15153 : n15156;
  assign n15158 = pi17 ? n37 : n15157;
  assign n15159 = pi16 ? n439 : n15158;
  assign n15160 = pi20 ? n2049 : n233;
  assign n15161 = pi19 ? n37 : n15160;
  assign n15162 = pi21 ? n233 : n5758;
  assign n15163 = pi20 ? n15162 : n32;
  assign n15164 = pi19 ? n15163 : n32;
  assign n15165 = pi18 ? n15161 : n15164;
  assign n15166 = pi17 ? n37 : n15165;
  assign n15167 = pi16 ? n439 : n15166;
  assign n15168 = pi15 ? n15159 : n15167;
  assign n15169 = pi14 ? n15150 : n15168;
  assign n15170 = pi13 ? n15127 : n15169;
  assign n15171 = pi12 ? n15098 : n15170;
  assign n15172 = pi11 ? n15001 : n15171;
  assign n15173 = pi21 ? n3392 : n37;
  assign n15174 = pi20 ? n15173 : n37;
  assign n15175 = pi19 ? n37 : n15174;
  assign n15176 = pi18 ? n37 : n15175;
  assign n15177 = pi21 ? n2707 : n233;
  assign n15178 = pi20 ? n8927 : n15177;
  assign n15179 = pi19 ? n37 : n15178;
  assign n15180 = pi21 ? n5014 : n5758;
  assign n15181 = pi20 ? n15180 : n32;
  assign n15182 = pi19 ? n15181 : n32;
  assign n15183 = pi18 ? n15179 : n15182;
  assign n15184 = pi17 ? n15176 : n15183;
  assign n15185 = pi16 ? n439 : n15184;
  assign n15186 = pi23 ? n685 : n363;
  assign n15187 = pi22 ? n686 : n15186;
  assign n15188 = pi21 ? n363 : n15187;
  assign n15189 = pi20 ? n3393 : n15188;
  assign n15190 = pi19 ? n37 : n15189;
  assign n15191 = pi18 ? n15190 : n14694;
  assign n15192 = pi17 ? n15176 : n15191;
  assign n15193 = pi16 ? n439 : n15192;
  assign n15194 = pi15 ? n15185 : n15193;
  assign n15195 = pi20 ? n2107 : n685;
  assign n15196 = pi19 ? n37 : n15195;
  assign n15197 = pi21 ? n685 : n7723;
  assign n15198 = pi20 ? n15197 : n32;
  assign n15199 = pi19 ? n15198 : n32;
  assign n15200 = pi18 ? n15196 : n15199;
  assign n15201 = pi17 ? n37 : n15200;
  assign n15202 = pi16 ? n439 : n15201;
  assign n15203 = pi15 ? n15202 : n14689;
  assign n15204 = pi14 ? n15194 : n15203;
  assign n15205 = pi19 ? n99 : n7746;
  assign n15206 = pi18 ? n15205 : n14683;
  assign n15207 = pi17 ? n99 : n15206;
  assign n15208 = pi16 ? n201 : n15207;
  assign n15209 = pi21 ? n767 : n7048;
  assign n15210 = pi20 ? n15209 : n32;
  assign n15211 = pi19 ? n15210 : n32;
  assign n15212 = pi18 ? n99 : n15211;
  assign n15213 = pi17 ? n99 : n15212;
  assign n15214 = pi16 ? n744 : n15213;
  assign n15215 = pi15 ? n15208 : n15214;
  assign n15216 = pi14 ? n14689 : n15215;
  assign n15217 = pi13 ? n15204 : n15216;
  assign n15218 = pi20 ? n775 : n99;
  assign n15219 = pi19 ? n2242 : n15218;
  assign n15220 = pi18 ? n99 : n15219;
  assign n15221 = pi21 ? n777 : n6089;
  assign n15222 = pi20 ? n99 : n15221;
  assign n15223 = pi19 ? n99 : n15222;
  assign n15224 = pi18 ? n15223 : n14709;
  assign n15225 = pi17 ? n15220 : n15224;
  assign n15226 = pi16 ? n744 : n15225;
  assign n15227 = pi21 ? n6461 : n775;
  assign n15228 = pi20 ? n15227 : n787;
  assign n15229 = pi19 ? n7845 : n15228;
  assign n15230 = pi18 ? n99 : n15229;
  assign n15231 = pi20 ? n99 : n775;
  assign n15232 = pi21 ? n777 : n14277;
  assign n15233 = pi20 ? n99 : n15232;
  assign n15234 = pi19 ? n15231 : n15233;
  assign n15235 = pi21 ? n6461 : n5829;
  assign n15236 = pi20 ? n15235 : n32;
  assign n15237 = pi19 ? n15236 : n32;
  assign n15238 = pi18 ? n15234 : n15237;
  assign n15239 = pi17 ? n15230 : n15238;
  assign n15240 = pi16 ? n744 : n15239;
  assign n15241 = pi15 ? n15226 : n15240;
  assign n15242 = pi19 ? n14285 : n99;
  assign n15243 = pi18 ? n742 : n15242;
  assign n15244 = pi17 ? n32 : n15243;
  assign n15245 = pi20 ? n776 : n99;
  assign n15246 = pi19 ? n14285 : n15245;
  assign n15247 = pi20 ? n99 : n6523;
  assign n15248 = pi19 ? n15247 : n157;
  assign n15249 = pi18 ? n15246 : n15248;
  assign n15250 = pi20 ? n787 : n7818;
  assign n15251 = pi21 ? n775 : n6089;
  assign n15252 = pi20 ? n787 : n15251;
  assign n15253 = pi19 ? n15250 : n15252;
  assign n15254 = pi21 ? n157 : n5829;
  assign n15255 = pi20 ? n15254 : n32;
  assign n15256 = pi19 ? n15255 : n32;
  assign n15257 = pi18 ? n15253 : n15256;
  assign n15258 = pi17 ? n15249 : n15257;
  assign n15259 = pi16 ? n15244 : n15258;
  assign n15260 = pi21 ? n7128 : n777;
  assign n15261 = pi20 ? n32 : n15260;
  assign n15262 = pi19 ? n32 : n15261;
  assign n15263 = pi21 ? n157 : n99;
  assign n15264 = pi20 ? n15263 : n6508;
  assign n15265 = pi19 ? n15263 : n15264;
  assign n15266 = pi18 ? n15262 : n15265;
  assign n15267 = pi17 ? n32 : n15266;
  assign n15268 = pi21 ? n157 : n2998;
  assign n15269 = pi20 ? n6523 : n15268;
  assign n15270 = pi19 ? n15269 : n14459;
  assign n15271 = pi20 ? n787 : n157;
  assign n15272 = pi21 ? n685 : n157;
  assign n15273 = pi20 ? n15272 : n157;
  assign n15274 = pi19 ? n15271 : n15273;
  assign n15275 = pi18 ? n15270 : n15274;
  assign n15276 = pi21 ? n685 : n6089;
  assign n15277 = pi20 ? n9021 : n15276;
  assign n15278 = pi19 ? n157 : n15277;
  assign n15279 = pi21 ? n14277 : n2637;
  assign n15280 = pi20 ? n15279 : n32;
  assign n15281 = pi19 ? n15280 : n32;
  assign n15282 = pi18 ? n15278 : n15281;
  assign n15283 = pi17 ? n15275 : n15282;
  assign n15284 = pi16 ? n15267 : n15283;
  assign n15285 = pi15 ? n15259 : n15284;
  assign n15286 = pi14 ? n15241 : n15285;
  assign n15287 = pi21 ? n157 : n928;
  assign n15288 = pi20 ? n15287 : n32;
  assign n15289 = pi19 ? n15288 : n32;
  assign n15290 = pi18 ? n157 : n15289;
  assign n15291 = pi17 ? n157 : n15290;
  assign n15292 = pi16 ? n7793 : n15291;
  assign n15293 = pi24 ? n157 : n204;
  assign n15294 = pi23 ? n157 : n15293;
  assign n15295 = pi22 ? n99 : n15294;
  assign n15296 = pi21 ? n15295 : n928;
  assign n15297 = pi20 ? n15296 : n32;
  assign n15298 = pi19 ? n15297 : n32;
  assign n15299 = pi18 ? n99 : n15298;
  assign n15300 = pi17 ? n99 : n15299;
  assign n15301 = pi16 ? n1510 : n15300;
  assign n15302 = pi21 ? n14506 : n3520;
  assign n15303 = pi20 ? n32 : n15302;
  assign n15304 = pi19 ? n32 : n15303;
  assign n15305 = pi22 ? n112 : n157;
  assign n15306 = pi21 ? n4221 : n15305;
  assign n15307 = pi18 ? n15304 : n15306;
  assign n15308 = pi17 ? n32 : n15307;
  assign n15309 = pi21 ? n11732 : n775;
  assign n15310 = pi21 ? n3520 : n181;
  assign n15311 = pi20 ? n15309 : n15310;
  assign n15312 = pi22 ? n2160 : n812;
  assign n15313 = pi21 ? n3520 : n15312;
  assign n15314 = pi21 ? n15305 : n4221;
  assign n15315 = pi20 ? n15313 : n15314;
  assign n15316 = pi19 ? n15311 : n15315;
  assign n15317 = pi21 ? n775 : n3520;
  assign n15318 = pi22 ? n157 : n812;
  assign n15319 = pi21 ? n4221 : n15318;
  assign n15320 = pi20 ? n15317 : n15319;
  assign n15321 = pi22 ? n316 : n812;
  assign n15322 = pi21 ? n15321 : n15318;
  assign n15323 = pi21 ? n775 : n4247;
  assign n15324 = pi20 ? n15322 : n15323;
  assign n15325 = pi19 ? n15320 : n15324;
  assign n15326 = pi18 ? n15316 : n15325;
  assign n15327 = pi20 ? n3520 : n11747;
  assign n15328 = pi20 ? n15317 : n11747;
  assign n15329 = pi19 ? n15327 : n15328;
  assign n15330 = pi20 ? n980 : n32;
  assign n15331 = pi19 ? n15330 : n32;
  assign n15332 = pi18 ? n15329 : n15331;
  assign n15333 = pi17 ? n15326 : n15332;
  assign n15334 = pi16 ? n15308 : n15333;
  assign n15335 = pi15 ? n15301 : n15334;
  assign n15336 = pi14 ? n15292 : n15335;
  assign n15337 = pi13 ? n15286 : n15336;
  assign n15338 = pi12 ? n15217 : n15337;
  assign n15339 = pi20 ? n9773 : n139;
  assign n15340 = pi19 ? n139 : n15339;
  assign n15341 = pi18 ? n139 : n15340;
  assign n15342 = pi20 ? n929 : n32;
  assign n15343 = pi19 ? n15342 : n32;
  assign n15344 = pi18 ? n139 : n15343;
  assign n15345 = pi17 ? n15341 : n15344;
  assign n15346 = pi16 ? n915 : n15345;
  assign n15347 = pi20 ? n5317 : n975;
  assign n15348 = pi19 ? n1820 : n15347;
  assign n15349 = pi18 ? n139 : n15348;
  assign n15350 = pi21 ? n1785 : n356;
  assign n15351 = pi20 ? n139 : n15350;
  assign n15352 = pi19 ? n139 : n15351;
  assign n15353 = pi18 ? n15352 : n15331;
  assign n15354 = pi17 ? n15349 : n15353;
  assign n15355 = pi16 ? n915 : n15354;
  assign n15356 = pi15 ? n15346 : n15355;
  assign n15357 = pi20 ? n350 : n139;
  assign n15358 = pi19 ? n15357 : n139;
  assign n15359 = pi19 ? n2352 : n316;
  assign n15360 = pi18 ? n15358 : n15359;
  assign n15361 = pi20 ? n2353 : n5317;
  assign n15362 = pi19 ? n15361 : n9071;
  assign n15363 = pi18 ? n15362 : n14306;
  assign n15364 = pi17 ? n15360 : n15363;
  assign n15365 = pi16 ? n915 : n15364;
  assign n15366 = pi19 ? n15339 : n139;
  assign n15367 = pi18 ? n15366 : n15359;
  assign n15368 = pi20 ? n975 : n927;
  assign n15369 = pi19 ? n316 : n15368;
  assign n15370 = pi21 ? n3990 : n1009;
  assign n15371 = pi20 ? n15370 : n32;
  assign n15372 = pi19 ? n15371 : n32;
  assign n15373 = pi18 ? n15369 : n15372;
  assign n15374 = pi17 ? n15367 : n15373;
  assign n15375 = pi16 ? n915 : n15374;
  assign n15376 = pi15 ? n15365 : n15375;
  assign n15377 = pi14 ? n15356 : n15376;
  assign n15378 = pi19 ? n10892 : n316;
  assign n15379 = pi18 ? n15378 : n316;
  assign n15380 = pi18 ? n316 : n14306;
  assign n15381 = pi17 ? n15379 : n15380;
  assign n15382 = pi16 ? n11772 : n15381;
  assign n15383 = pi20 ? n1030 : n32;
  assign n15384 = pi19 ? n15383 : n32;
  assign n15385 = pi18 ? n316 : n15384;
  assign n15386 = pi17 ? n15379 : n15385;
  assign n15387 = pi16 ? n11772 : n15386;
  assign n15388 = pi15 ? n15382 : n15387;
  assign n15389 = pi18 ? n10060 : n316;
  assign n15390 = pi17 ? n32 : n15389;
  assign n15391 = pi18 ? n15378 : n10893;
  assign n15392 = pi18 ? n10893 : n13400;
  assign n15393 = pi17 ? n15391 : n15392;
  assign n15394 = pi16 ? n15390 : n15393;
  assign n15395 = pi21 ? n910 : n204;
  assign n15396 = pi20 ? n32 : n15395;
  assign n15397 = pi19 ? n32 : n15396;
  assign n15398 = pi20 ? n2318 : n204;
  assign n15399 = pi19 ? n2318 : n15398;
  assign n15400 = pi18 ? n15397 : n15399;
  assign n15401 = pi17 ? n32 : n15400;
  assign n15402 = pi20 ? n1016 : n2318;
  assign n15403 = pi19 ? n15402 : n15398;
  assign n15404 = pi18 ? n15403 : n204;
  assign n15405 = pi20 ? n204 : n2318;
  assign n15406 = pi19 ? n204 : n15405;
  assign n15407 = pi21 ? n10417 : n32;
  assign n15408 = pi20 ? n15407 : n32;
  assign n15409 = pi19 ? n15408 : n32;
  assign n15410 = pi18 ? n15406 : n15409;
  assign n15411 = pi17 ? n15404 : n15410;
  assign n15412 = pi16 ? n15401 : n15411;
  assign n15413 = pi15 ? n15394 : n15412;
  assign n15414 = pi14 ? n15388 : n15413;
  assign n15415 = pi13 ? n15377 : n15414;
  assign n15416 = pi21 ? n555 : n204;
  assign n15417 = pi20 ? n32 : n15416;
  assign n15418 = pi19 ? n32 : n15417;
  assign n15419 = pi18 ? n15418 : n204;
  assign n15420 = pi17 ? n32 : n15419;
  assign n15421 = pi21 ? n204 : n37;
  assign n15422 = pi20 ? n204 : n15421;
  assign n15423 = pi19 ? n15422 : n204;
  assign n15424 = pi18 ? n15423 : n204;
  assign n15425 = pi18 ? n204 : n15409;
  assign n15426 = pi17 ? n15424 : n15425;
  assign n15427 = pi16 ? n15420 : n15426;
  assign n15428 = pi20 ? n204 : n9180;
  assign n15429 = pi19 ? n15428 : n6749;
  assign n15430 = pi18 ? n15429 : n204;
  assign n15431 = pi17 ? n15430 : n14780;
  assign n15432 = pi16 ? n15420 : n15431;
  assign n15433 = pi15 ? n15427 : n15432;
  assign n15434 = pi21 ? n1929 : n335;
  assign n15435 = pi20 ? n15434 : n335;
  assign n15436 = pi19 ? n335 : n15435;
  assign n15437 = pi18 ? n335 : n15436;
  assign n15438 = pi19 ? n335 : n13532;
  assign n15439 = pi22 ? n4079 : n317;
  assign n15440 = pi21 ? n15439 : n32;
  assign n15441 = pi20 ? n15440 : n32;
  assign n15442 = pi19 ? n15441 : n32;
  assign n15443 = pi18 ? n15438 : n15442;
  assign n15444 = pi17 ? n15437 : n15443;
  assign n15445 = pi16 ? n2035 : n15444;
  assign n15446 = pi21 ? n13280 : n32;
  assign n15447 = pi20 ? n15446 : n32;
  assign n15448 = pi19 ? n15447 : n32;
  assign n15449 = pi18 ? n335 : n15448;
  assign n15450 = pi17 ? n335 : n15449;
  assign n15451 = pi16 ? n2035 : n15450;
  assign n15452 = pi15 ? n15445 : n15451;
  assign n15453 = pi14 ? n15433 : n15452;
  assign n15454 = pi18 ? n14385 : n6369;
  assign n15455 = pi17 ? n335 : n15454;
  assign n15456 = pi16 ? n2035 : n15455;
  assign n15457 = pi21 ? n6376 : n335;
  assign n15458 = pi20 ? n15457 : n335;
  assign n15459 = pi19 ? n335 : n15458;
  assign n15460 = pi18 ? n335 : n15459;
  assign n15461 = pi18 ? n12631 : n7044;
  assign n15462 = pi17 ? n15460 : n15461;
  assign n15463 = pi16 ? n10118 : n15462;
  assign n15464 = pi15 ? n15456 : n15463;
  assign n15465 = pi21 ? n233 : n6361;
  assign n15466 = pi20 ? n15465 : n335;
  assign n15467 = pi19 ? n8914 : n15466;
  assign n15468 = pi18 ? n335 : n15467;
  assign n15469 = pi21 ? n6361 : n335;
  assign n15470 = pi20 ? n15469 : n335;
  assign n15471 = pi19 ? n15470 : n8914;
  assign n15472 = pi18 ? n15471 : n3979;
  assign n15473 = pi17 ? n15468 : n15472;
  assign n15474 = pi16 ? n11849 : n15473;
  assign n15475 = pi22 ? n962 : n233;
  assign n15476 = pi21 ? n15475 : n335;
  assign n15477 = pi20 ? n32 : n15476;
  assign n15478 = pi19 ? n32 : n15477;
  assign n15479 = pi21 ? n6376 : n9122;
  assign n15480 = pi21 ? n335 : n9122;
  assign n15481 = pi20 ? n15479 : n15480;
  assign n15482 = pi20 ? n15480 : n335;
  assign n15483 = pi19 ? n15481 : n15482;
  assign n15484 = pi18 ? n15478 : n15483;
  assign n15485 = pi17 ? n32 : n15484;
  assign n15486 = pi21 ? n335 : n9143;
  assign n15487 = pi20 ? n233 : n15486;
  assign n15488 = pi20 ? n13527 : n335;
  assign n15489 = pi19 ? n15487 : n15488;
  assign n15490 = pi18 ? n15489 : n13533;
  assign n15491 = pi18 ? n233 : n4104;
  assign n15492 = pi17 ? n15490 : n15491;
  assign n15493 = pi16 ? n15485 : n15492;
  assign n15494 = pi15 ? n15474 : n15493;
  assign n15495 = pi14 ? n15464 : n15494;
  assign n15496 = pi13 ? n15453 : n15495;
  assign n15497 = pi12 ? n15415 : n15496;
  assign n15498 = pi11 ? n15338 : n15497;
  assign n15499 = pi10 ? n15172 : n15498;
  assign n15500 = pi09 ? n14828 : n15499;
  assign n15501 = pi15 ? n32 : n14821;
  assign n15502 = pi16 ? n11885 : n14818;
  assign n15503 = pi15 ? n14822 : n15502;
  assign n15504 = pi14 ? n15501 : n15503;
  assign n15505 = pi13 ? n32 : n15504;
  assign n15506 = pi12 ? n32 : n15505;
  assign n15507 = pi11 ? n32 : n15506;
  assign n15508 = pi10 ? n32 : n15507;
  assign n15509 = pi16 ? n12689 : n14833;
  assign n15510 = pi16 ? n13561 : n14839;
  assign n15511 = pi15 ? n15509 : n15510;
  assign n15512 = pi16 ? n14445 : n14851;
  assign n15513 = pi21 ? n3779 : n99;
  assign n15514 = pi20 ? n32 : n15513;
  assign n15515 = pi19 ? n32 : n15514;
  assign n15516 = pi18 ? n15515 : n99;
  assign n15517 = pi17 ? n32 : n15516;
  assign n15518 = pi16 ? n15517 : n14861;
  assign n15519 = pi15 ? n15512 : n15518;
  assign n15520 = pi14 ? n15511 : n15519;
  assign n15521 = pi16 ? n801 : n14870;
  assign n15522 = pi16 ? n721 : n14875;
  assign n15523 = pi15 ? n15521 : n15522;
  assign n15524 = pi21 ? n796 : n112;
  assign n15525 = pi20 ? n32 : n15524;
  assign n15526 = pi19 ? n32 : n15525;
  assign n15527 = pi20 ? n5501 : n2962;
  assign n15528 = pi19 ? n15527 : n6039;
  assign n15529 = pi18 ? n15526 : n15528;
  assign n15530 = pi17 ? n32 : n15529;
  assign n15531 = pi19 ? n14003 : n4616;
  assign n15532 = pi18 ? n14002 : n15531;
  assign n15533 = pi21 ? n157 : n2746;
  assign n15534 = pi20 ? n2191 : n15533;
  assign n15535 = pi19 ? n15534 : n4619;
  assign n15536 = pi20 ? n6508 : n2470;
  assign n15537 = pi19 ? n15536 : n32;
  assign n15538 = pi18 ? n15535 : n15537;
  assign n15539 = pi17 ? n15532 : n15538;
  assign n15540 = pi16 ? n15530 : n15539;
  assign n15541 = pi19 ? n3050 : n99;
  assign n15542 = pi18 ? n99 : n15541;
  assign n15543 = pi20 ? n3046 : n99;
  assign n15544 = pi19 ? n15543 : n3050;
  assign n15545 = pi21 ? n2998 : n2164;
  assign n15546 = pi20 ? n15545 : n2470;
  assign n15547 = pi19 ? n15546 : n32;
  assign n15548 = pi18 ? n15544 : n15547;
  assign n15549 = pi17 ? n15542 : n15548;
  assign n15550 = pi16 ? n744 : n15549;
  assign n15551 = pi15 ? n15540 : n15550;
  assign n15552 = pi14 ? n15523 : n15551;
  assign n15553 = pi13 ? n15520 : n15552;
  assign n15554 = pi20 ? n220 : n2470;
  assign n15555 = pi19 ? n15554 : n32;
  assign n15556 = pi18 ? n99 : n15555;
  assign n15557 = pi17 ? n99 : n15556;
  assign n15558 = pi16 ? n721 : n15557;
  assign n15559 = pi20 ? n14478 : n2554;
  assign n15560 = pi19 ? n15559 : n32;
  assign n15561 = pi18 ? n99 : n15560;
  assign n15562 = pi17 ? n99 : n15561;
  assign n15563 = pi16 ? n801 : n15562;
  assign n15564 = pi15 ? n15558 : n15563;
  assign n15565 = pi20 ? n14927 : n2554;
  assign n15566 = pi19 ? n15565 : n32;
  assign n15567 = pi18 ? n99 : n15566;
  assign n15568 = pi17 ? n99 : n15567;
  assign n15569 = pi16 ? n14926 : n15568;
  assign n15570 = pi20 ? n14937 : n2679;
  assign n15571 = pi19 ? n15570 : n32;
  assign n15572 = pi18 ? n99 : n15571;
  assign n15573 = pi17 ? n99 : n15572;
  assign n15574 = pi16 ? n721 : n15573;
  assign n15575 = pi15 ? n15569 : n15574;
  assign n15576 = pi14 ? n15564 : n15575;
  assign n15577 = pi20 ? n5269 : n1761;
  assign n15578 = pi19 ? n37 : n15577;
  assign n15579 = pi18 ? n374 : n15578;
  assign n15580 = pi17 ? n32 : n15579;
  assign n15581 = pi20 ? n14953 : n2679;
  assign n15582 = pi19 ? n15581 : n32;
  assign n15583 = pi18 ? n139 : n15582;
  assign n15584 = pi17 ? n139 : n15583;
  assign n15585 = pi16 ? n15580 : n15584;
  assign n15586 = pi18 ? n374 : n14963;
  assign n15587 = pi17 ? n32 : n15586;
  assign n15588 = pi20 ? n14542 : n2701;
  assign n15589 = pi19 ? n15588 : n32;
  assign n15590 = pi18 ? n139 : n15589;
  assign n15591 = pi17 ? n139 : n15590;
  assign n15592 = pi16 ? n15587 : n15591;
  assign n15593 = pi15 ? n15585 : n15592;
  assign n15594 = pi21 ? n1211 : n375;
  assign n15595 = pi20 ? n12010 : n15594;
  assign n15596 = pi19 ? n37 : n15595;
  assign n15597 = pi20 ? n1699 : n1738;
  assign n15598 = pi20 ? n1738 : n11579;
  assign n15599 = pi19 ? n15597 : n15598;
  assign n15600 = pi18 ? n15596 : n15599;
  assign n15601 = pi20 ? n1715 : n1707;
  assign n15602 = pi20 ? n1707 : n1714;
  assign n15603 = pi19 ? n15601 : n15602;
  assign n15604 = pi20 ? n14979 : n2701;
  assign n15605 = pi19 ? n15604 : n32;
  assign n15606 = pi18 ? n15603 : n15605;
  assign n15607 = pi17 ? n15600 : n15606;
  assign n15608 = pi16 ? n439 : n15607;
  assign n15609 = pi15 ? n15608 : n14997;
  assign n15610 = pi14 ? n15593 : n15609;
  assign n15611 = pi13 ? n15576 : n15610;
  assign n15612 = pi12 ? n15553 : n15611;
  assign n15613 = pi23 ? n139 : n8133;
  assign n15614 = pi22 ? n139 : n15613;
  assign n15615 = pi21 ? n139 : n15614;
  assign n15616 = pi20 ? n15615 : n32;
  assign n15617 = pi19 ? n15616 : n32;
  assign n15618 = pi18 ? n139 : n15617;
  assign n15619 = pi17 ? n15030 : n15618;
  assign n15620 = pi16 ? n439 : n15619;
  assign n15621 = pi20 ? n1219 : n32;
  assign n15622 = pi19 ? n15621 : n32;
  assign n15623 = pi18 ? n139 : n15622;
  assign n15624 = pi17 ? n15041 : n15623;
  assign n15625 = pi16 ? n15036 : n15624;
  assign n15626 = pi15 ? n15620 : n15625;
  assign n15627 = pi14 ? n15028 : n15626;
  assign n15628 = pi22 ? n583 : n295;
  assign n15629 = pi21 ? n15057 : n15628;
  assign n15630 = pi20 ? n15629 : n13670;
  assign n15631 = pi19 ? n15059 : n15630;
  assign n15632 = pi22 ? n9827 : n583;
  assign n15633 = pi21 ? n15632 : n7621;
  assign n15634 = pi20 ? n15633 : n32;
  assign n15635 = pi19 ? n15634 : n32;
  assign n15636 = pi18 ? n15631 : n15635;
  assign n15637 = pi17 ? n15054 : n15636;
  assign n15638 = pi16 ? n439 : n15637;
  assign n15639 = pi22 ? n204 : n7513;
  assign n15640 = pi21 ? n335 : n15639;
  assign n15641 = pi20 ? n15640 : n32;
  assign n15642 = pi19 ? n15641 : n32;
  assign n15643 = pi18 ? n15073 : n15642;
  assign n15644 = pi17 ? n15070 : n15643;
  assign n15645 = pi16 ? n439 : n15644;
  assign n15646 = pi15 ? n15638 : n15645;
  assign n15647 = pi22 ? n335 : n6405;
  assign n15648 = pi21 ? n335 : n15647;
  assign n15649 = pi20 ? n15648 : n32;
  assign n15650 = pi19 ? n15649 : n32;
  assign n15651 = pi18 ? n12629 : n15650;
  assign n15652 = pi17 ? n37 : n15651;
  assign n15653 = pi16 ? n439 : n15652;
  assign n15654 = pi15 ? n15088 : n15653;
  assign n15655 = pi14 ? n15646 : n15654;
  assign n15656 = pi13 ? n15627 : n15655;
  assign n15657 = pi22 ? n583 : n1388;
  assign n15658 = pi21 ? n37 : n15657;
  assign n15659 = pi20 ? n15658 : n32;
  assign n15660 = pi19 ? n15659 : n32;
  assign n15661 = pi18 ? n9381 : n15660;
  assign n15662 = pi17 ? n37 : n15661;
  assign n15663 = pi16 ? n439 : n15662;
  assign n15664 = pi15 ? n15106 : n15663;
  assign n15665 = pi21 ? n37 : n11199;
  assign n15666 = pi20 ? n15665 : n32;
  assign n15667 = pi19 ? n15666 : n32;
  assign n15668 = pi18 ? n9381 : n15667;
  assign n15669 = pi17 ? n37 : n15668;
  assign n15670 = pi16 ? n439 : n15669;
  assign n15671 = pi21 ? n570 : n9413;
  assign n15672 = pi20 ? n15671 : n32;
  assign n15673 = pi19 ? n15672 : n32;
  assign n15674 = pi18 ? n15118 : n15673;
  assign n15675 = pi17 ? n37 : n15674;
  assign n15676 = pi16 ? n439 : n15675;
  assign n15677 = pi15 ? n15670 : n15676;
  assign n15678 = pi14 ? n15664 : n15677;
  assign n15679 = pi21 ? n1920 : n9413;
  assign n15680 = pi20 ? n15679 : n32;
  assign n15681 = pi19 ? n15680 : n32;
  assign n15682 = pi18 ? n15130 : n15681;
  assign n15683 = pi17 ? n15129 : n15682;
  assign n15684 = pi16 ? n439 : n15683;
  assign n15685 = pi21 ? n580 : n584;
  assign n15686 = pi21 ? n580 : n2007;
  assign n15687 = pi20 ? n15685 : n15686;
  assign n15688 = pi19 ? n8802 : n15687;
  assign n15689 = pi22 ? n233 : n4146;
  assign n15690 = pi21 ? n15143 : n15689;
  assign n15691 = pi20 ? n15690 : n32;
  assign n15692 = pi19 ? n15691 : n32;
  assign n15693 = pi18 ? n15688 : n15692;
  assign n15694 = pi17 ? n15139 : n15693;
  assign n15695 = pi16 ? n439 : n15694;
  assign n15696 = pi15 ? n15684 : n15695;
  assign n15697 = pi23 ? n2120 : n395;
  assign n15698 = pi22 ? n233 : n15697;
  assign n15699 = pi21 ? n2091 : n15698;
  assign n15700 = pi20 ? n15699 : n32;
  assign n15701 = pi19 ? n15700 : n32;
  assign n15702 = pi18 ? n15153 : n15701;
  assign n15703 = pi17 ? n37 : n15702;
  assign n15704 = pi16 ? n439 : n15703;
  assign n15705 = pi21 ? n233 : n8272;
  assign n15706 = pi20 ? n15705 : n32;
  assign n15707 = pi19 ? n15706 : n32;
  assign n15708 = pi18 ? n15161 : n15707;
  assign n15709 = pi17 ? n37 : n15708;
  assign n15710 = pi16 ? n439 : n15709;
  assign n15711 = pi15 ? n15704 : n15710;
  assign n15712 = pi14 ? n15696 : n15711;
  assign n15713 = pi13 ? n15678 : n15712;
  assign n15714 = pi12 ? n15656 : n15713;
  assign n15715 = pi11 ? n15612 : n15714;
  assign n15716 = pi21 ? n5014 : n650;
  assign n15717 = pi20 ? n15716 : n32;
  assign n15718 = pi19 ? n15717 : n32;
  assign n15719 = pi18 ? n15179 : n15718;
  assign n15720 = pi17 ? n15176 : n15719;
  assign n15721 = pi16 ? n439 : n15720;
  assign n15722 = pi21 ? n363 : n696;
  assign n15723 = pi20 ? n15722 : n32;
  assign n15724 = pi19 ? n15723 : n32;
  assign n15725 = pi18 ? n15190 : n15724;
  assign n15726 = pi17 ? n15176 : n15725;
  assign n15727 = pi16 ? n439 : n15726;
  assign n15728 = pi15 ? n15721 : n15727;
  assign n15729 = pi21 ? n685 : n696;
  assign n15730 = pi20 ? n15729 : n32;
  assign n15731 = pi19 ? n15730 : n32;
  assign n15732 = pi18 ? n15196 : n15731;
  assign n15733 = pi17 ? n37 : n15732;
  assign n15734 = pi16 ? n439 : n15733;
  assign n15735 = pi21 ? n2106 : n696;
  assign n15736 = pi20 ? n15735 : n32;
  assign n15737 = pi19 ? n15736 : n32;
  assign n15738 = pi18 ? n37 : n15737;
  assign n15739 = pi17 ? n37 : n15738;
  assign n15740 = pi16 ? n439 : n15739;
  assign n15741 = pi15 ? n15734 : n15740;
  assign n15742 = pi14 ? n15728 : n15741;
  assign n15743 = pi18 ? n15205 : n15737;
  assign n15744 = pi17 ? n99 : n15743;
  assign n15745 = pi16 ? n201 : n15744;
  assign n15746 = pi20 ? n1477 : n32;
  assign n15747 = pi19 ? n15746 : n32;
  assign n15748 = pi18 ? n99 : n15747;
  assign n15749 = pi17 ? n99 : n15748;
  assign n15750 = pi16 ? n721 : n15749;
  assign n15751 = pi15 ? n15745 : n15750;
  assign n15752 = pi14 ? n15740 : n15751;
  assign n15753 = pi13 ? n15742 : n15752;
  assign n15754 = pi21 ? n6461 : n7723;
  assign n15755 = pi20 ? n15754 : n32;
  assign n15756 = pi19 ? n15755 : n32;
  assign n15757 = pi18 ? n15223 : n15756;
  assign n15758 = pi17 ? n15220 : n15757;
  assign n15759 = pi16 ? n721 : n15758;
  assign n15760 = pi21 ? n6461 : n7048;
  assign n15761 = pi20 ? n15760 : n32;
  assign n15762 = pi19 ? n15761 : n32;
  assign n15763 = pi18 ? n15234 : n15762;
  assign n15764 = pi17 ? n15230 : n15763;
  assign n15765 = pi16 ? n721 : n15764;
  assign n15766 = pi15 ? n15759 : n15765;
  assign n15767 = pi18 ? n719 : n15242;
  assign n15768 = pi17 ? n32 : n15767;
  assign n15769 = pi21 ? n157 : n7048;
  assign n15770 = pi20 ? n15769 : n32;
  assign n15771 = pi19 ? n15770 : n32;
  assign n15772 = pi18 ? n15253 : n15771;
  assign n15773 = pi17 ? n15249 : n15772;
  assign n15774 = pi16 ? n15768 : n15773;
  assign n15775 = pi21 ? n6519 : n777;
  assign n15776 = pi20 ? n32 : n15775;
  assign n15777 = pi19 ? n32 : n15776;
  assign n15778 = pi18 ? n15777 : n15265;
  assign n15779 = pi17 ? n32 : n15778;
  assign n15780 = pi21 ? n14277 : n5829;
  assign n15781 = pi20 ? n15780 : n32;
  assign n15782 = pi19 ? n15781 : n32;
  assign n15783 = pi18 ? n15278 : n15782;
  assign n15784 = pi17 ? n15275 : n15783;
  assign n15785 = pi16 ? n15779 : n15784;
  assign n15786 = pi15 ? n15774 : n15785;
  assign n15787 = pi14 ? n15766 : n15786;
  assign n15788 = pi20 ? n883 : n32;
  assign n15789 = pi19 ? n15788 : n32;
  assign n15790 = pi18 ? n157 : n15789;
  assign n15791 = pi17 ? n157 : n15790;
  assign n15792 = pi16 ? n5910 : n15791;
  assign n15793 = pi16 ? n5910 : n15291;
  assign n15794 = pi15 ? n15792 : n15793;
  assign n15795 = pi21 ? n777 : n928;
  assign n15796 = pi20 ? n15795 : n32;
  assign n15797 = pi19 ? n15796 : n32;
  assign n15798 = pi18 ? n99 : n15797;
  assign n15799 = pi17 ? n99 : n15798;
  assign n15800 = pi16 ? n801 : n15799;
  assign n15801 = pi21 ? n8143 : n3520;
  assign n15802 = pi20 ? n32 : n15801;
  assign n15803 = pi19 ? n32 : n15802;
  assign n15804 = pi21 ? n4221 : n1526;
  assign n15805 = pi18 ? n15803 : n15804;
  assign n15806 = pi17 ? n32 : n15805;
  assign n15807 = pi21 ? n4226 : n15318;
  assign n15808 = pi22 ? n1043 : n99;
  assign n15809 = pi21 ? n248 : n15808;
  assign n15810 = pi20 ? n15807 : n15809;
  assign n15811 = pi22 ? n1043 : n812;
  assign n15812 = pi21 ? n248 : n15811;
  assign n15813 = pi21 ? n1526 : n4234;
  assign n15814 = pi20 ? n15812 : n15813;
  assign n15815 = pi19 ? n15810 : n15814;
  assign n15816 = pi21 ? n4221 : n5540;
  assign n15817 = pi20 ? n15317 : n15816;
  assign n15818 = pi21 ? n356 : n15318;
  assign n15819 = pi21 ? n15318 : n4252;
  assign n15820 = pi20 ? n15818 : n15819;
  assign n15821 = pi19 ? n15817 : n15820;
  assign n15822 = pi18 ? n15815 : n15821;
  assign n15823 = pi21 ? n248 : n3520;
  assign n15824 = pi20 ? n15823 : n11734;
  assign n15825 = pi21 ? n775 : n248;
  assign n15826 = pi20 ? n15825 : n11734;
  assign n15827 = pi19 ? n15824 : n15826;
  assign n15828 = pi18 ? n15827 : n15331;
  assign n15829 = pi17 ? n15822 : n15828;
  assign n15830 = pi16 ? n15806 : n15829;
  assign n15831 = pi15 ? n15800 : n15830;
  assign n15832 = pi14 ? n15794 : n15831;
  assign n15833 = pi13 ? n15787 : n15832;
  assign n15834 = pi12 ? n15753 : n15833;
  assign n15835 = pi16 ? n12576 : n15381;
  assign n15836 = pi16 ? n12576 : n15386;
  assign n15837 = pi15 ? n15835 : n15836;
  assign n15838 = pi22 ? n8447 : n139;
  assign n15839 = pi21 ? n15838 : n316;
  assign n15840 = pi20 ? n32 : n15839;
  assign n15841 = pi19 ? n32 : n15840;
  assign n15842 = pi18 ? n15841 : n316;
  assign n15843 = pi17 ? n32 : n15842;
  assign n15844 = pi16 ? n15843 : n15393;
  assign n15845 = pi21 ? n963 : n204;
  assign n15846 = pi20 ? n32 : n15845;
  assign n15847 = pi19 ? n32 : n15846;
  assign n15848 = pi18 ? n15847 : n15399;
  assign n15849 = pi17 ? n32 : n15848;
  assign n15850 = pi20 ? n1601 : n32;
  assign n15851 = pi19 ? n15850 : n32;
  assign n15852 = pi18 ? n15406 : n15851;
  assign n15853 = pi17 ? n15404 : n15852;
  assign n15854 = pi16 ? n15849 : n15853;
  assign n15855 = pi15 ? n15844 : n15854;
  assign n15856 = pi14 ? n15837 : n15855;
  assign n15857 = pi13 ? n15377 : n15856;
  assign n15858 = pi20 ? n1072 : n32;
  assign n15859 = pi19 ? n15858 : n32;
  assign n15860 = pi18 ? n204 : n15859;
  assign n15861 = pi17 ? n15424 : n15860;
  assign n15862 = pi16 ? n15420 : n15861;
  assign n15863 = pi23 ? n8133 : n32;
  assign n15864 = pi22 ? n204 : n15863;
  assign n15865 = pi21 ? n15864 : n32;
  assign n15866 = pi20 ? n15865 : n32;
  assign n15867 = pi19 ? n15866 : n32;
  assign n15868 = pi18 ? n204 : n15867;
  assign n15869 = pi17 ? n15430 : n15868;
  assign n15870 = pi16 ? n15420 : n15869;
  assign n15871 = pi15 ? n15862 : n15870;
  assign n15872 = pi19 ? n335 : n4940;
  assign n15873 = pi18 ? n335 : n15872;
  assign n15874 = pi22 ? n4079 : n1407;
  assign n15875 = pi21 ? n15874 : n32;
  assign n15876 = pi20 ? n15875 : n32;
  assign n15877 = pi19 ? n15876 : n32;
  assign n15878 = pi18 ? n15438 : n15877;
  assign n15879 = pi17 ? n15873 : n15878;
  assign n15880 = pi16 ? n2035 : n15879;
  assign n15881 = pi21 ? n10119 : n32;
  assign n15882 = pi20 ? n15881 : n32;
  assign n15883 = pi19 ? n15882 : n32;
  assign n15884 = pi18 ? n335 : n15883;
  assign n15885 = pi17 ? n335 : n15884;
  assign n15886 = pi16 ? n2035 : n15885;
  assign n15887 = pi15 ? n15880 : n15886;
  assign n15888 = pi14 ? n15871 : n15887;
  assign n15889 = pi22 ? n6365 : n317;
  assign n15890 = pi21 ? n15889 : n32;
  assign n15891 = pi20 ? n15890 : n32;
  assign n15892 = pi19 ? n15891 : n32;
  assign n15893 = pi18 ? n14385 : n15892;
  assign n15894 = pi17 ? n335 : n15893;
  assign n15895 = pi16 ? n2035 : n15894;
  assign n15896 = pi15 ? n15895 : n15463;
  assign n15897 = pi18 ? n233 : n14399;
  assign n15898 = pi17 ? n15490 : n15897;
  assign n15899 = pi16 ? n15485 : n15898;
  assign n15900 = pi15 ? n15474 : n15899;
  assign n15901 = pi14 ? n15896 : n15900;
  assign n15902 = pi13 ? n15888 : n15901;
  assign n15903 = pi12 ? n15857 : n15902;
  assign n15904 = pi11 ? n15834 : n15903;
  assign n15905 = pi10 ? n15715 : n15904;
  assign n15906 = pi09 ? n15508 : n15905;
  assign n15907 = pi08 ? n15500 : n15906;
  assign n15908 = pi20 ? n37 : n2947;
  assign n15909 = pi19 ? n15908 : n32;
  assign n15910 = pi18 ? n37 : n15909;
  assign n15911 = pi17 ? n37 : n15910;
  assign n15912 = pi16 ? n10154 : n15911;
  assign n15913 = pi15 ? n32 : n15912;
  assign n15914 = pi16 ? n11011 : n15911;
  assign n15915 = pi16 ? n11885 : n15911;
  assign n15916 = pi15 ? n15914 : n15915;
  assign n15917 = pi14 ? n15913 : n15916;
  assign n15918 = pi13 ? n32 : n15917;
  assign n15919 = pi12 ? n32 : n15918;
  assign n15920 = pi11 ? n32 : n15919;
  assign n15921 = pi10 ? n32 : n15920;
  assign n15922 = pi20 ? n99 : n2990;
  assign n15923 = pi19 ? n15922 : n32;
  assign n15924 = pi18 ? n37 : n15923;
  assign n15925 = pi17 ? n37 : n15924;
  assign n15926 = pi16 ? n12689 : n15925;
  assign n15927 = pi20 ? n99 : n3023;
  assign n15928 = pi19 ? n15927 : n32;
  assign n15929 = pi18 ? n37 : n15928;
  assign n15930 = pi17 ? n37 : n15929;
  assign n15931 = pi16 ? n13561 : n15930;
  assign n15932 = pi15 ? n15926 : n15931;
  assign n15933 = pi20 ? n14846 : n3067;
  assign n15934 = pi19 ? n15933 : n32;
  assign n15935 = pi18 ? n14845 : n15934;
  assign n15936 = pi17 ? n14843 : n15935;
  assign n15937 = pi16 ? n14445 : n15936;
  assign n15938 = pi22 ? n39 : n99;
  assign n15939 = pi21 ? n15938 : n99;
  assign n15940 = pi20 ? n32 : n15939;
  assign n15941 = pi19 ? n32 : n15940;
  assign n15942 = pi18 ? n15941 : n99;
  assign n15943 = pi17 ? n32 : n15942;
  assign n15944 = pi20 ? n14846 : n14835;
  assign n15945 = pi19 ? n15944 : n32;
  assign n15946 = pi18 ? n99 : n15945;
  assign n15947 = pi17 ? n99 : n15946;
  assign n15948 = pi16 ? n15943 : n15947;
  assign n15949 = pi15 ? n15937 : n15948;
  assign n15950 = pi14 ? n15932 : n15949;
  assign n15951 = pi20 ? n3039 : n37;
  assign n15952 = pi19 ? n15951 : n37;
  assign n15953 = pi18 ? n14880 : n15952;
  assign n15954 = pi17 ? n32 : n15953;
  assign n15955 = pi21 ? n2957 : n2156;
  assign n15956 = pi20 ? n3870 : n15955;
  assign n15957 = pi19 ? n37 : n15956;
  assign n15958 = pi21 ? n2957 : n2162;
  assign n15959 = pi20 ? n15958 : n3870;
  assign n15960 = pi21 ? n2981 : n218;
  assign n15961 = pi19 ? n15959 : n15960;
  assign n15962 = pi18 ? n15957 : n15961;
  assign n15963 = pi20 ? n2959 : n2755;
  assign n15964 = pi21 ? n37 : n2160;
  assign n15965 = pi19 ? n15963 : n15964;
  assign n15966 = pi20 ? n4616 : n14847;
  assign n15967 = pi19 ? n15966 : n32;
  assign n15968 = pi18 ? n15965 : n15967;
  assign n15969 = pi17 ? n15962 : n15968;
  assign n15970 = pi16 ? n15954 : n15969;
  assign n15971 = pi20 ? n99 : n14847;
  assign n15972 = pi19 ? n15971 : n32;
  assign n15973 = pi18 ? n99 : n15972;
  assign n15974 = pi17 ? n99 : n15973;
  assign n15975 = pi16 ? n744 : n15974;
  assign n15976 = pi15 ? n15970 : n15975;
  assign n15977 = pi19 ? n9710 : n99;
  assign n15978 = pi21 ? n8044 : n32;
  assign n15979 = pi20 ? n3014 : n15978;
  assign n15980 = pi19 ? n15979 : n32;
  assign n15981 = pi18 ? n15977 : n15980;
  assign n15982 = pi17 ? n99 : n15981;
  assign n15983 = pi16 ? n721 : n15982;
  assign n15984 = pi20 ? n221 : n2470;
  assign n15985 = pi19 ? n15984 : n32;
  assign n15986 = pi18 ? n99 : n15985;
  assign n15987 = pi17 ? n99 : n15986;
  assign n15988 = pi16 ? n801 : n15987;
  assign n15989 = pi15 ? n15983 : n15988;
  assign n15990 = pi14 ? n15976 : n15989;
  assign n15991 = pi13 ? n15950 : n15990;
  assign n15992 = pi16 ? n744 : n15557;
  assign n15993 = pi20 ? n99 : n2554;
  assign n15994 = pi19 ? n15993 : n32;
  assign n15995 = pi18 ? n99 : n15994;
  assign n15996 = pi17 ? n99 : n15995;
  assign n15997 = pi16 ? n721 : n15996;
  assign n15998 = pi15 ? n15992 : n15997;
  assign n15999 = pi20 ? n2191 : n3825;
  assign n16000 = pi19 ? n15999 : n99;
  assign n16001 = pi18 ? n799 : n16000;
  assign n16002 = pi17 ? n32 : n16001;
  assign n16003 = pi16 ? n16002 : n15996;
  assign n16004 = pi22 ? n738 : n2160;
  assign n16005 = pi21 ? n16004 : n2168;
  assign n16006 = pi20 ? n32 : n16005;
  assign n16007 = pi19 ? n32 : n16006;
  assign n16008 = pi21 ? n2156 : n37;
  assign n16009 = pi20 ? n16008 : n15964;
  assign n16010 = pi19 ? n16009 : n3508;
  assign n16011 = pi18 ? n16007 : n16010;
  assign n16012 = pi17 ? n32 : n16011;
  assign n16013 = pi19 ? n3889 : n99;
  assign n16014 = pi18 ? n16013 : n99;
  assign n16015 = pi20 ? n10836 : n2679;
  assign n16016 = pi19 ? n16015 : n32;
  assign n16017 = pi18 ? n99 : n16016;
  assign n16018 = pi17 ? n16014 : n16017;
  assign n16019 = pi16 ? n16012 : n16018;
  assign n16020 = pi15 ? n16003 : n16019;
  assign n16021 = pi14 ? n15998 : n16020;
  assign n16022 = pi20 ? n3083 : n1747;
  assign n16023 = pi20 ? n5273 : n139;
  assign n16024 = pi19 ? n16022 : n16023;
  assign n16025 = pi18 ? n16024 : n139;
  assign n16026 = pi21 ? n139 : n9828;
  assign n16027 = pi20 ? n16026 : n2679;
  assign n16028 = pi19 ? n16027 : n32;
  assign n16029 = pi18 ? n139 : n16028;
  assign n16030 = pi17 ? n16025 : n16029;
  assign n16031 = pi16 ? n439 : n16030;
  assign n16032 = pi20 ? n1761 : n139;
  assign n16033 = pi19 ? n37 : n16032;
  assign n16034 = pi18 ? n16033 : n139;
  assign n16035 = pi23 ? n139 : n3134;
  assign n16036 = pi22 ? n139 : n16035;
  assign n16037 = pi21 ? n139 : n16036;
  assign n16038 = pi20 ? n16037 : n2701;
  assign n16039 = pi19 ? n16038 : n32;
  assign n16040 = pi18 ? n139 : n16039;
  assign n16041 = pi17 ? n16034 : n16040;
  assign n16042 = pi16 ? n439 : n16041;
  assign n16043 = pi15 ? n16031 : n16042;
  assign n16044 = pi20 ? n13121 : n942;
  assign n16045 = pi19 ? n9824 : n16044;
  assign n16046 = pi18 ? n37 : n16045;
  assign n16047 = pi21 ? n820 : n1721;
  assign n16048 = pi20 ? n139 : n16047;
  assign n16049 = pi19 ? n16048 : n939;
  assign n16050 = pi21 ? n820 : n1785;
  assign n16051 = pi20 ? n16050 : n2653;
  assign n16052 = pi19 ? n16051 : n32;
  assign n16053 = pi18 ? n16049 : n16052;
  assign n16054 = pi17 ? n16046 : n16053;
  assign n16055 = pi16 ? n439 : n16054;
  assign n16056 = pi19 ? n37 : n13125;
  assign n16057 = pi20 ? n37 : n3078;
  assign n16058 = pi21 ? n297 : n375;
  assign n16059 = pi20 ? n3078 : n16058;
  assign n16060 = pi19 ? n16057 : n16059;
  assign n16061 = pi18 ? n16056 : n16060;
  assign n16062 = pi20 ? n3092 : n3084;
  assign n16063 = pi20 ? n1693 : n1714;
  assign n16064 = pi19 ? n16062 : n16063;
  assign n16065 = pi21 ? n1696 : n1793;
  assign n16066 = pi20 ? n16065 : n2653;
  assign n16067 = pi19 ? n16066 : n32;
  assign n16068 = pi18 ? n16064 : n16067;
  assign n16069 = pi17 ? n16061 : n16068;
  assign n16070 = pi16 ? n439 : n16069;
  assign n16071 = pi15 ? n16055 : n16070;
  assign n16072 = pi14 ? n16043 : n16071;
  assign n16073 = pi13 ? n16021 : n16072;
  assign n16074 = pi12 ? n15991 : n16073;
  assign n16075 = pi20 ? n3083 : n13118;
  assign n16076 = pi19 ? n12370 : n16075;
  assign n16077 = pi18 ? n37 : n16076;
  assign n16078 = pi21 ? n1531 : n375;
  assign n16079 = pi20 ? n16058 : n16078;
  assign n16080 = pi20 ? n5257 : n3092;
  assign n16081 = pi19 ? n16079 : n16080;
  assign n16082 = pi20 ? n3645 : n2653;
  assign n16083 = pi19 ? n16082 : n32;
  assign n16084 = pi18 ? n16081 : n16083;
  assign n16085 = pi17 ? n16077 : n16084;
  assign n16086 = pi16 ? n439 : n16085;
  assign n16087 = pi20 ? n139 : n1822;
  assign n16088 = pi19 ? n16087 : n32;
  assign n16089 = pi18 ? n139 : n16088;
  assign n16090 = pi17 ? n15030 : n16089;
  assign n16091 = pi16 ? n439 : n16090;
  assign n16092 = pi15 ? n16086 : n16091;
  assign n16093 = pi19 ? n37 : n9814;
  assign n16094 = pi18 ? n37 : n16093;
  assign n16095 = pi20 ? n1026 : n1822;
  assign n16096 = pi19 ? n16095 : n32;
  assign n16097 = pi18 ? n139 : n16096;
  assign n16098 = pi17 ? n16094 : n16097;
  assign n16099 = pi16 ? n439 : n16098;
  assign n16100 = pi20 ? n1794 : n32;
  assign n16101 = pi19 ? n16100 : n32;
  assign n16102 = pi18 ? n139 : n16101;
  assign n16103 = pi17 ? n16094 : n16102;
  assign n16104 = pi16 ? n439 : n16103;
  assign n16105 = pi15 ? n16099 : n16104;
  assign n16106 = pi14 ? n16092 : n16105;
  assign n16107 = pi21 ? n1056 : n506;
  assign n16108 = pi21 ? n1046 : n506;
  assign n16109 = pi20 ? n16107 : n16108;
  assign n16110 = pi21 ? n1046 : n455;
  assign n16111 = pi21 ? n1046 : n516;
  assign n16112 = pi20 ? n16110 : n16111;
  assign n16113 = pi19 ? n16109 : n16112;
  assign n16114 = pi21 ? n506 : n204;
  assign n16115 = pi20 ? n16114 : n32;
  assign n16116 = pi19 ? n16115 : n32;
  assign n16117 = pi18 ? n16113 : n16116;
  assign n16118 = pi17 ? n37 : n16117;
  assign n16119 = pi16 ? n439 : n16118;
  assign n16120 = pi21 ? n1083 : n10663;
  assign n16121 = pi20 ? n6947 : n16120;
  assign n16122 = pi21 ? n1083 : n455;
  assign n16123 = pi20 ? n16122 : n4870;
  assign n16124 = pi19 ? n16121 : n16123;
  assign n16125 = pi21 ? n10663 : n204;
  assign n16126 = pi20 ? n16125 : n32;
  assign n16127 = pi19 ? n16126 : n32;
  assign n16128 = pi18 ? n16124 : n16127;
  assign n16129 = pi17 ? n37 : n16128;
  assign n16130 = pi16 ? n439 : n16129;
  assign n16131 = pi15 ? n16119 : n16130;
  assign n16132 = pi19 ? n13247 : n335;
  assign n16133 = pi20 ? n6377 : n32;
  assign n16134 = pi19 ? n16133 : n32;
  assign n16135 = pi18 ? n16132 : n16134;
  assign n16136 = pi17 ? n37 : n16135;
  assign n16137 = pi16 ? n439 : n16136;
  assign n16138 = pi19 ? n7676 : n335;
  assign n16139 = pi20 ? n2062 : n32;
  assign n16140 = pi19 ? n16139 : n32;
  assign n16141 = pi18 ? n16138 : n16140;
  assign n16142 = pi17 ? n37 : n16141;
  assign n16143 = pi16 ? n439 : n16142;
  assign n16144 = pi15 ? n16137 : n16143;
  assign n16145 = pi14 ? n16131 : n16144;
  assign n16146 = pi13 ? n16106 : n16145;
  assign n16147 = pi19 ? n6373 : n335;
  assign n16148 = pi20 ? n13510 : n32;
  assign n16149 = pi19 ? n16148 : n32;
  assign n16150 = pi18 ? n16147 : n16149;
  assign n16151 = pi17 ? n37 : n16150;
  assign n16152 = pi16 ? n439 : n16151;
  assign n16153 = pi20 ? n2016 : n15116;
  assign n16154 = pi19 ? n8802 : n16153;
  assign n16155 = pi21 ? n1943 : n13516;
  assign n16156 = pi20 ? n16155 : n32;
  assign n16157 = pi19 ? n16156 : n32;
  assign n16158 = pi18 ? n16154 : n16157;
  assign n16159 = pi17 ? n37 : n16158;
  assign n16160 = pi16 ? n439 : n16159;
  assign n16161 = pi15 ? n16152 : n16160;
  assign n16162 = pi19 ? n37 : n16153;
  assign n16163 = pi21 ? n1943 : n6376;
  assign n16164 = pi20 ? n16163 : n32;
  assign n16165 = pi19 ? n16164 : n32;
  assign n16166 = pi18 ? n16162 : n16165;
  assign n16167 = pi17 ? n37 : n16166;
  assign n16168 = pi16 ? n439 : n16167;
  assign n16169 = pi21 ? n569 : n11199;
  assign n16170 = pi20 ? n2016 : n16169;
  assign n16171 = pi19 ? n37 : n16170;
  assign n16172 = pi21 ? n1943 : n8860;
  assign n16173 = pi20 ? n16172 : n32;
  assign n16174 = pi19 ? n16173 : n32;
  assign n16175 = pi18 ? n16171 : n16174;
  assign n16176 = pi17 ? n37 : n16175;
  assign n16177 = pi16 ? n439 : n16176;
  assign n16178 = pi15 ? n16168 : n16177;
  assign n16179 = pi14 ? n16161 : n16178;
  assign n16180 = pi20 ? n603 : n6377;
  assign n16181 = pi19 ? n37 : n16180;
  assign n16182 = pi21 ? n335 : n8869;
  assign n16183 = pi20 ? n16182 : n32;
  assign n16184 = pi19 ? n16183 : n32;
  assign n16185 = pi18 ? n16181 : n16184;
  assign n16186 = pi17 ? n37 : n16185;
  assign n16187 = pi16 ? n439 : n16186;
  assign n16188 = pi21 ? n37 : n9657;
  assign n16189 = pi21 ? n11635 : n2707;
  assign n16190 = pi20 ? n16188 : n16189;
  assign n16191 = pi19 ? n37 : n16190;
  assign n16192 = pi21 ? n9666 : n9430;
  assign n16193 = pi20 ? n16192 : n32;
  assign n16194 = pi19 ? n16193 : n32;
  assign n16195 = pi18 ? n16191 : n16194;
  assign n16196 = pi17 ? n37 : n16195;
  assign n16197 = pi16 ? n439 : n16196;
  assign n16198 = pi15 ? n16187 : n16197;
  assign n16199 = pi21 ? n5012 : n2707;
  assign n16200 = pi20 ? n37 : n16199;
  assign n16201 = pi19 ? n37 : n16200;
  assign n16202 = pi22 ? n5011 : n3338;
  assign n16203 = pi21 ? n3392 : n16202;
  assign n16204 = pi20 ? n16203 : n32;
  assign n16205 = pi19 ? n16204 : n32;
  assign n16206 = pi18 ? n16201 : n16205;
  assign n16207 = pi17 ? n37 : n16206;
  assign n16208 = pi16 ? n439 : n16207;
  assign n16209 = pi19 ? n37 : n13337;
  assign n16210 = pi22 ? n559 : n664;
  assign n16211 = pi21 ? n233 : n16210;
  assign n16212 = pi20 ? n16211 : n32;
  assign n16213 = pi19 ? n16212 : n32;
  assign n16214 = pi18 ? n16209 : n16213;
  assign n16215 = pi17 ? n37 : n16214;
  assign n16216 = pi16 ? n439 : n16215;
  assign n16217 = pi15 ? n16208 : n16216;
  assign n16218 = pi14 ? n16198 : n16217;
  assign n16219 = pi13 ? n16179 : n16218;
  assign n16220 = pi12 ? n16146 : n16219;
  assign n16221 = pi11 ? n16074 : n16220;
  assign n16222 = pi20 ? n37 : n10496;
  assign n16223 = pi19 ? n37 : n16222;
  assign n16224 = pi21 ? n363 : n16210;
  assign n16225 = pi20 ? n16224 : n32;
  assign n16226 = pi19 ? n16225 : n32;
  assign n16227 = pi18 ? n16223 : n16226;
  assign n16228 = pi17 ? n37 : n16227;
  assign n16229 = pi16 ? n439 : n16228;
  assign n16230 = pi22 ? n14245 : n1407;
  assign n16231 = pi21 ? n363 : n16230;
  assign n16232 = pi20 ? n16231 : n32;
  assign n16233 = pi19 ? n16232 : n32;
  assign n16234 = pi18 ? n16223 : n16233;
  assign n16235 = pi17 ? n15176 : n16234;
  assign n16236 = pi16 ? n439 : n16235;
  assign n16237 = pi15 ? n16229 : n16236;
  assign n16238 = pi20 ? n37 : n685;
  assign n16239 = pi19 ? n37 : n16238;
  assign n16240 = pi20 ? n2214 : n32;
  assign n16241 = pi19 ? n16240 : n32;
  assign n16242 = pi18 ? n16239 : n16241;
  assign n16243 = pi17 ? n37 : n16242;
  assign n16244 = pi16 ? n439 : n16243;
  assign n16245 = pi21 ? n2106 : n1423;
  assign n16246 = pi20 ? n16245 : n32;
  assign n16247 = pi19 ? n16246 : n32;
  assign n16248 = pi18 ? n37 : n16247;
  assign n16249 = pi17 ? n37 : n16248;
  assign n16250 = pi16 ? n439 : n16249;
  assign n16251 = pi15 ? n16244 : n16250;
  assign n16252 = pi14 ? n16237 : n16251;
  assign n16253 = pi21 ? n2106 : n1416;
  assign n16254 = pi20 ? n16253 : n32;
  assign n16255 = pi19 ? n16254 : n32;
  assign n16256 = pi18 ? n37 : n16255;
  assign n16257 = pi17 ? n37 : n16256;
  assign n16258 = pi16 ? n439 : n16257;
  assign n16259 = pi15 ? n16250 : n16258;
  assign n16260 = pi18 ? n15205 : n16247;
  assign n16261 = pi17 ? n99 : n16260;
  assign n16262 = pi16 ? n201 : n16261;
  assign n16263 = pi21 ? n99 : n5464;
  assign n16264 = pi20 ? n99 : n16263;
  assign n16265 = pi19 ? n99 : n16264;
  assign n16266 = pi22 ? n2244 : n317;
  assign n16267 = pi21 ? n767 : n16266;
  assign n16268 = pi20 ? n16267 : n32;
  assign n16269 = pi19 ? n16268 : n32;
  assign n16270 = pi18 ? n16265 : n16269;
  assign n16271 = pi17 ? n99 : n16270;
  assign n16272 = pi16 ? n744 : n16271;
  assign n16273 = pi15 ? n16262 : n16272;
  assign n16274 = pi14 ? n16259 : n16273;
  assign n16275 = pi13 ? n16252 : n16274;
  assign n16276 = pi20 ? n157 : n99;
  assign n16277 = pi19 ? n99 : n16276;
  assign n16278 = pi18 ? n99 : n16277;
  assign n16279 = pi21 ? n157 : n14277;
  assign n16280 = pi20 ? n99 : n16279;
  assign n16281 = pi19 ? n14285 : n16280;
  assign n16282 = pi20 ? n4297 : n32;
  assign n16283 = pi19 ? n16282 : n32;
  assign n16284 = pi18 ? n16281 : n16283;
  assign n16285 = pi17 ? n16278 : n16284;
  assign n16286 = pi16 ? n744 : n16285;
  assign n16287 = pi21 ? n777 : n2998;
  assign n16288 = pi20 ? n16287 : n99;
  assign n16289 = pi19 ? n16288 : n99;
  assign n16290 = pi19 ? n7845 : n6532;
  assign n16291 = pi18 ? n16289 : n16290;
  assign n16292 = pi20 ? n6503 : n157;
  assign n16293 = pi21 ? n99 : n14277;
  assign n16294 = pi20 ? n99 : n16293;
  assign n16295 = pi19 ? n16292 : n16294;
  assign n16296 = pi22 ? n158 : n7377;
  assign n16297 = pi21 ? n16296 : n2245;
  assign n16298 = pi20 ? n16297 : n32;
  assign n16299 = pi19 ? n16298 : n32;
  assign n16300 = pi18 ? n16295 : n16299;
  assign n16301 = pi17 ? n16291 : n16300;
  assign n16302 = pi16 ? n744 : n16301;
  assign n16303 = pi15 ? n16286 : n16302;
  assign n16304 = pi21 ? n5168 : n99;
  assign n16305 = pi20 ? n32 : n16304;
  assign n16306 = pi19 ? n32 : n16305;
  assign n16307 = pi20 ? n157 : n2243;
  assign n16308 = pi19 ? n16307 : n2243;
  assign n16309 = pi18 ? n16306 : n16308;
  assign n16310 = pi17 ? n32 : n16309;
  assign n16311 = pi20 ? n15263 : n157;
  assign n16312 = pi20 ? n3484 : n2238;
  assign n16313 = pi19 ? n16311 : n16312;
  assign n16314 = pi18 ? n16313 : n6510;
  assign n16315 = pi20 ? n157 : n15251;
  assign n16316 = pi19 ? n157 : n16315;
  assign n16317 = pi22 ? n1484 : n706;
  assign n16318 = pi21 ? n157 : n16317;
  assign n16319 = pi20 ? n16318 : n32;
  assign n16320 = pi19 ? n16319 : n32;
  assign n16321 = pi18 ? n16316 : n16320;
  assign n16322 = pi17 ? n16314 : n16321;
  assign n16323 = pi16 ? n16310 : n16322;
  assign n16324 = pi19 ? n157 : n16307;
  assign n16325 = pi20 ? n2283 : n32;
  assign n16326 = pi19 ? n16325 : n32;
  assign n16327 = pi18 ? n16324 : n16326;
  assign n16328 = pi17 ? n157 : n16327;
  assign n16329 = pi16 ? n5910 : n16328;
  assign n16330 = pi15 ? n16323 : n16329;
  assign n16331 = pi14 ? n16303 : n16330;
  assign n16332 = pi23 ? n4262 : n99;
  assign n16333 = pi22 ? n16332 : n157;
  assign n16334 = pi21 ? n16333 : n157;
  assign n16335 = pi20 ? n32 : n16334;
  assign n16336 = pi19 ? n32 : n16335;
  assign n16337 = pi18 ? n16336 : n157;
  assign n16338 = pi17 ? n32 : n16337;
  assign n16339 = pi21 ? n157 : n2320;
  assign n16340 = pi20 ? n16339 : n32;
  assign n16341 = pi19 ? n16340 : n32;
  assign n16342 = pi18 ? n157 : n16341;
  assign n16343 = pi17 ? n157 : n16342;
  assign n16344 = pi16 ? n16338 : n16343;
  assign n16345 = pi21 ? n6519 : n157;
  assign n16346 = pi20 ? n32 : n16345;
  assign n16347 = pi19 ? n32 : n16346;
  assign n16348 = pi18 ? n16347 : n157;
  assign n16349 = pi17 ? n32 : n16348;
  assign n16350 = pi22 ? n6146 : n32;
  assign n16351 = pi21 ? n777 : n16350;
  assign n16352 = pi20 ? n16351 : n32;
  assign n16353 = pi19 ? n16352 : n32;
  assign n16354 = pi18 ? n157 : n16353;
  assign n16355 = pi17 ? n157 : n16354;
  assign n16356 = pi16 ? n16349 : n16355;
  assign n16357 = pi15 ? n16344 : n16356;
  assign n16358 = pi22 ? n430 : n32;
  assign n16359 = pi21 ? n777 : n16358;
  assign n16360 = pi20 ? n16359 : n32;
  assign n16361 = pi19 ? n16360 : n32;
  assign n16362 = pi18 ? n99 : n16361;
  assign n16363 = pi17 ? n99 : n16362;
  assign n16364 = pi16 ? n721 : n16363;
  assign n16365 = pi21 ? n963 : n248;
  assign n16366 = pi20 ? n32 : n16365;
  assign n16367 = pi19 ? n32 : n16366;
  assign n16368 = pi18 ? n16367 : n2281;
  assign n16369 = pi17 ? n32 : n16368;
  assign n16370 = pi20 ? n876 : n875;
  assign n16371 = pi21 ? n244 : n139;
  assign n16372 = pi20 ? n16371 : n875;
  assign n16373 = pi19 ? n16370 : n16372;
  assign n16374 = pi21 ? n258 : n248;
  assign n16375 = pi20 ? n16374 : n876;
  assign n16376 = pi20 ? n1001 : n2292;
  assign n16377 = pi19 ? n16375 : n16376;
  assign n16378 = pi18 ? n16373 : n16377;
  assign n16379 = pi20 ? n248 : n139;
  assign n16380 = pi20 ? n16374 : n1008;
  assign n16381 = pi19 ? n16379 : n16380;
  assign n16382 = pi21 ? n316 : n3339;
  assign n16383 = pi20 ? n16382 : n32;
  assign n16384 = pi19 ? n16383 : n32;
  assign n16385 = pi18 ? n16381 : n16384;
  assign n16386 = pi17 ? n16378 : n16385;
  assign n16387 = pi16 ? n16369 : n16386;
  assign n16388 = pi15 ? n16364 : n16387;
  assign n16389 = pi14 ? n16357 : n16388;
  assign n16390 = pi13 ? n16331 : n16389;
  assign n16391 = pi12 ? n16275 : n16390;
  assign n16392 = pi20 ? n976 : n139;
  assign n16393 = pi19 ? n139 : n16392;
  assign n16394 = pi18 ? n139 : n16393;
  assign n16395 = pi21 ? n2319 : n882;
  assign n16396 = pi20 ? n16395 : n32;
  assign n16397 = pi19 ? n16396 : n32;
  assign n16398 = pi18 ? n139 : n16397;
  assign n16399 = pi17 ? n16394 : n16398;
  assign n16400 = pi16 ? n2291 : n16399;
  assign n16401 = pi20 ? n316 : n975;
  assign n16402 = pi19 ? n139 : n16401;
  assign n16403 = pi18 ? n139 : n16402;
  assign n16404 = pi19 ? n5312 : n14318;
  assign n16405 = pi18 ? n16404 : n9757;
  assign n16406 = pi17 ? n16403 : n16405;
  assign n16407 = pi16 ? n2291 : n16406;
  assign n16408 = pi15 ? n16400 : n16407;
  assign n16409 = pi20 ? n15350 : n139;
  assign n16410 = pi19 ? n16409 : n139;
  assign n16411 = pi18 ? n16410 : n15359;
  assign n16412 = pi20 ? n4437 : n11785;
  assign n16413 = pi19 ? n316 : n16412;
  assign n16414 = pi18 ? n16413 : n15331;
  assign n16415 = pi17 ? n16411 : n16414;
  assign n16416 = pi16 ? n2291 : n16415;
  assign n16417 = pi20 ? n1001 : n139;
  assign n16418 = pi19 ? n16417 : n139;
  assign n16419 = pi18 ? n16418 : n15359;
  assign n16420 = pi21 ? n3990 : n928;
  assign n16421 = pi20 ? n16420 : n32;
  assign n16422 = pi19 ? n16421 : n32;
  assign n16423 = pi18 ? n15369 : n16422;
  assign n16424 = pi17 ? n16419 : n16423;
  assign n16425 = pi16 ? n915 : n16424;
  assign n16426 = pi15 ? n16416 : n16425;
  assign n16427 = pi14 ? n16408 : n16426;
  assign n16428 = pi21 ? n4429 : n316;
  assign n16429 = pi20 ? n16428 : n316;
  assign n16430 = pi19 ? n316 : n16429;
  assign n16431 = pi18 ? n16430 : n316;
  assign n16432 = pi18 ? n316 : n15331;
  assign n16433 = pi17 ? n16431 : n16432;
  assign n16434 = pi16 ? n11772 : n16433;
  assign n16435 = pi20 ? n9082 : n316;
  assign n16436 = pi19 ? n10892 : n16435;
  assign n16437 = pi18 ? n16436 : n316;
  assign n16438 = pi22 ? n204 : n2299;
  assign n16439 = pi21 ? n16438 : n928;
  assign n16440 = pi20 ? n16439 : n32;
  assign n16441 = pi19 ? n16440 : n32;
  assign n16442 = pi18 ? n316 : n16441;
  assign n16443 = pi17 ? n16437 : n16442;
  assign n16444 = pi16 ? n11772 : n16443;
  assign n16445 = pi15 ? n16434 : n16444;
  assign n16446 = pi21 ? n10057 : n139;
  assign n16447 = pi20 ? n32 : n16446;
  assign n16448 = pi19 ? n32 : n16447;
  assign n16449 = pi21 ? n3617 : n359;
  assign n16450 = pi20 ? n16449 : n11277;
  assign n16451 = pi19 ? n16450 : n11277;
  assign n16452 = pi18 ? n16448 : n16451;
  assign n16453 = pi17 ? n32 : n16452;
  assign n16454 = pi21 ? n4429 : n349;
  assign n16455 = pi20 ? n350 : n16454;
  assign n16456 = pi20 ? n8719 : n3172;
  assign n16457 = pi19 ? n16455 : n16456;
  assign n16458 = pi20 ? n6919 : n4433;
  assign n16459 = pi21 ? n4429 : n1785;
  assign n16460 = pi20 ? n11277 : n16459;
  assign n16461 = pi19 ? n16458 : n16460;
  assign n16462 = pi18 ? n16457 : n16461;
  assign n16463 = pi20 ? n8719 : n3617;
  assign n16464 = pi20 ? n16454 : n5961;
  assign n16465 = pi19 ? n16463 : n16464;
  assign n16466 = pi22 ? n1038 : n2299;
  assign n16467 = pi21 ? n16466 : n1009;
  assign n16468 = pi20 ? n16467 : n32;
  assign n16469 = pi19 ? n16468 : n32;
  assign n16470 = pi18 ? n16465 : n16469;
  assign n16471 = pi17 ? n16462 : n16470;
  assign n16472 = pi16 ? n16453 : n16471;
  assign n16473 = pi20 ? n139 : n204;
  assign n16474 = pi19 ? n15402 : n16473;
  assign n16475 = pi18 ? n16474 : n204;
  assign n16476 = pi21 ? n16438 : n32;
  assign n16477 = pi20 ? n16476 : n32;
  assign n16478 = pi19 ? n16477 : n32;
  assign n16479 = pi18 ? n15406 : n16478;
  assign n16480 = pi17 ? n16475 : n16479;
  assign n16481 = pi16 ? n15401 : n16480;
  assign n16482 = pi15 ? n16472 : n16481;
  assign n16483 = pi14 ? n16445 : n16482;
  assign n16484 = pi13 ? n16427 : n16483;
  assign n16485 = pi22 ? n2390 : n335;
  assign n16486 = pi21 ? n16485 : n204;
  assign n16487 = pi20 ? n32 : n16486;
  assign n16488 = pi19 ? n32 : n16487;
  assign n16489 = pi18 ? n16488 : n204;
  assign n16490 = pi17 ? n32 : n16489;
  assign n16491 = pi21 ? n204 : n570;
  assign n16492 = pi20 ? n204 : n16491;
  assign n16493 = pi21 ? n1313 : n204;
  assign n16494 = pi20 ? n16493 : n204;
  assign n16495 = pi19 ? n16492 : n16494;
  assign n16496 = pi18 ? n16495 : n204;
  assign n16497 = pi18 ? n204 : n16478;
  assign n16498 = pi17 ? n16496 : n16497;
  assign n16499 = pi16 ? n16490 : n16498;
  assign n16500 = pi21 ? n7938 : n204;
  assign n16501 = pi20 ? n32 : n16500;
  assign n16502 = pi19 ? n32 : n16501;
  assign n16503 = pi18 ? n16502 : n204;
  assign n16504 = pi17 ? n32 : n16503;
  assign n16505 = pi22 ? n204 : n430;
  assign n16506 = pi21 ? n16505 : n32;
  assign n16507 = pi20 ? n16506 : n32;
  assign n16508 = pi19 ? n16507 : n32;
  assign n16509 = pi18 ? n204 : n16508;
  assign n16510 = pi17 ? n15430 : n16509;
  assign n16511 = pi16 ? n16504 : n16510;
  assign n16512 = pi15 ? n16499 : n16511;
  assign n16513 = pi18 ? n15438 : n9443;
  assign n16514 = pi17 ? n335 : n16513;
  assign n16515 = pi16 ? n7943 : n16514;
  assign n16516 = pi20 ? n603 : n335;
  assign n16517 = pi19 ? n335 : n16516;
  assign n16518 = pi18 ? n16517 : n335;
  assign n16519 = pi21 ? n14168 : n32;
  assign n16520 = pi20 ? n16519 : n32;
  assign n16521 = pi19 ? n16520 : n32;
  assign n16522 = pi18 ? n335 : n16521;
  assign n16523 = pi17 ? n16518 : n16522;
  assign n16524 = pi16 ? n10399 : n16523;
  assign n16525 = pi15 ? n16515 : n16524;
  assign n16526 = pi14 ? n16512 : n16525;
  assign n16527 = pi18 ? n335 : n8919;
  assign n16528 = pi17 ? n16518 : n16527;
  assign n16529 = pi16 ? n10399 : n16528;
  assign n16530 = pi21 ? n6376 : n6361;
  assign n16531 = pi20 ? n16530 : n335;
  assign n16532 = pi19 ? n335 : n16531;
  assign n16533 = pi18 ? n335 : n16532;
  assign n16534 = pi18 ? n12631 : n15448;
  assign n16535 = pi17 ? n16533 : n16534;
  assign n16536 = pi16 ? n2425 : n16535;
  assign n16537 = pi15 ? n16529 : n16536;
  assign n16538 = pi22 ? n2419 : n99;
  assign n16539 = pi21 ? n16538 : n335;
  assign n16540 = pi20 ? n32 : n16539;
  assign n16541 = pi19 ? n32 : n16540;
  assign n16542 = pi18 ? n16541 : n335;
  assign n16543 = pi17 ? n32 : n16542;
  assign n16544 = pi21 ? n6376 : n233;
  assign n16545 = pi20 ? n16544 : n15469;
  assign n16546 = pi19 ? n335 : n16545;
  assign n16547 = pi18 ? n335 : n16546;
  assign n16548 = pi20 ? n7980 : n335;
  assign n16549 = pi19 ? n16548 : n8914;
  assign n16550 = pi18 ? n16549 : n5761;
  assign n16551 = pi17 ? n16547 : n16550;
  assign n16552 = pi16 ? n16543 : n16551;
  assign n16553 = pi22 ? n2419 : n233;
  assign n16554 = pi21 ? n16553 : n335;
  assign n16555 = pi20 ? n32 : n16554;
  assign n16556 = pi19 ? n32 : n16555;
  assign n16557 = pi21 ? n6376 : n4902;
  assign n16558 = pi20 ? n16557 : n14203;
  assign n16559 = pi19 ? n16558 : n14203;
  assign n16560 = pi18 ? n16556 : n16559;
  assign n16561 = pi17 ? n32 : n16560;
  assign n16562 = pi22 ? n4899 : n335;
  assign n16563 = pi21 ? n4908 : n16562;
  assign n16564 = pi20 ? n233 : n16563;
  assign n16565 = pi20 ? n13527 : n2062;
  assign n16566 = pi19 ? n16564 : n16565;
  assign n16567 = pi21 ? n4902 : n335;
  assign n16568 = pi20 ? n16567 : n233;
  assign n16569 = pi19 ? n16568 : n233;
  assign n16570 = pi18 ? n16566 : n16569;
  assign n16571 = pi18 ? n233 : n5761;
  assign n16572 = pi17 ? n16570 : n16571;
  assign n16573 = pi16 ? n16561 : n16572;
  assign n16574 = pi15 ? n16552 : n16573;
  assign n16575 = pi14 ? n16537 : n16574;
  assign n16576 = pi13 ? n16526 : n16575;
  assign n16577 = pi12 ? n16484 : n16576;
  assign n16578 = pi11 ? n16391 : n16577;
  assign n16579 = pi10 ? n16221 : n16578;
  assign n16580 = pi09 ? n15921 : n16579;
  assign n16581 = pi15 ? n32 : n15914;
  assign n16582 = pi16 ? n12689 : n15911;
  assign n16583 = pi15 ? n15915 : n16582;
  assign n16584 = pi14 ? n16581 : n16583;
  assign n16585 = pi13 ? n32 : n16584;
  assign n16586 = pi12 ? n32 : n16585;
  assign n16587 = pi11 ? n32 : n16586;
  assign n16588 = pi10 ? n32 : n16587;
  assign n16589 = pi16 ? n13561 : n15925;
  assign n16590 = pi16 ? n14445 : n15930;
  assign n16591 = pi15 ? n16589 : n16590;
  assign n16592 = pi20 ? n32 : n3780;
  assign n16593 = pi19 ? n32 : n16592;
  assign n16594 = pi18 ? n16593 : n37;
  assign n16595 = pi17 ? n32 : n16594;
  assign n16596 = pi16 ? n16595 : n15936;
  assign n16597 = pi21 ? n127 : n99;
  assign n16598 = pi20 ? n32 : n16597;
  assign n16599 = pi19 ? n32 : n16598;
  assign n16600 = pi18 ? n16599 : n99;
  assign n16601 = pi17 ? n32 : n16600;
  assign n16602 = pi16 ? n16601 : n15947;
  assign n16603 = pi15 ? n16596 : n16602;
  assign n16604 = pi14 ? n16591 : n16603;
  assign n16605 = pi18 ? n374 : n15952;
  assign n16606 = pi17 ? n32 : n16605;
  assign n16607 = pi20 ? n14518 : n14524;
  assign n16608 = pi19 ? n37 : n16607;
  assign n16609 = pi20 ? n14524 : n14518;
  assign n16610 = pi19 ? n16609 : n3039;
  assign n16611 = pi18 ? n16608 : n16610;
  assign n16612 = pi20 ? n14530 : n2959;
  assign n16613 = pi19 ? n16612 : n2974;
  assign n16614 = pi21 ? n218 : n2164;
  assign n16615 = pi20 ? n16614 : n14847;
  assign n16616 = pi19 ? n16615 : n32;
  assign n16617 = pi18 ? n16613 : n16616;
  assign n16618 = pi17 ? n16611 : n16617;
  assign n16619 = pi16 ? n16606 : n16618;
  assign n16620 = pi15 ? n16619 : n15975;
  assign n16621 = pi21 ? n9246 : n32;
  assign n16622 = pi20 ? n3014 : n16621;
  assign n16623 = pi19 ? n16622 : n32;
  assign n16624 = pi18 ? n15977 : n16623;
  assign n16625 = pi17 ? n99 : n16624;
  assign n16626 = pi16 ? n744 : n16625;
  assign n16627 = pi20 ? n221 : n16621;
  assign n16628 = pi19 ? n16627 : n32;
  assign n16629 = pi18 ? n99 : n16628;
  assign n16630 = pi17 ? n99 : n16629;
  assign n16631 = pi16 ? n801 : n16630;
  assign n16632 = pi15 ? n16626 : n16631;
  assign n16633 = pi14 ? n16620 : n16632;
  assign n16634 = pi13 ? n16604 : n16633;
  assign n16635 = pi20 ? n220 : n16621;
  assign n16636 = pi19 ? n16635 : n32;
  assign n16637 = pi18 ? n99 : n16636;
  assign n16638 = pi17 ? n99 : n16637;
  assign n16639 = pi16 ? n744 : n16638;
  assign n16640 = pi20 ? n99 : n2566;
  assign n16641 = pi19 ? n16640 : n32;
  assign n16642 = pi18 ? n99 : n16641;
  assign n16643 = pi17 ? n99 : n16642;
  assign n16644 = pi16 ? n744 : n16643;
  assign n16645 = pi15 ? n16639 : n16644;
  assign n16646 = pi20 ? n220 : n14844;
  assign n16647 = pi19 ? n16646 : n99;
  assign n16648 = pi18 ? n799 : n16647;
  assign n16649 = pi17 ? n32 : n16648;
  assign n16650 = pi16 ? n16649 : n16643;
  assign n16651 = pi20 ? n37 : n14513;
  assign n16652 = pi19 ? n37 : n16651;
  assign n16653 = pi18 ? n374 : n16652;
  assign n16654 = pi17 ? n32 : n16653;
  assign n16655 = pi20 ? n3814 : n8060;
  assign n16656 = pi19 ? n16655 : n99;
  assign n16657 = pi18 ? n16656 : n99;
  assign n16658 = pi21 ? n837 : n4237;
  assign n16659 = pi20 ? n16658 : n2579;
  assign n16660 = pi19 ? n16659 : n32;
  assign n16661 = pi18 ? n99 : n16660;
  assign n16662 = pi17 ? n16657 : n16661;
  assign n16663 = pi16 ? n16654 : n16662;
  assign n16664 = pi15 ? n16650 : n16663;
  assign n16665 = pi14 ? n16645 : n16664;
  assign n16666 = pi20 ? n3083 : n1761;
  assign n16667 = pi19 ? n16666 : n9769;
  assign n16668 = pi18 ? n16667 : n139;
  assign n16669 = pi20 ? n16026 : n2579;
  assign n16670 = pi19 ? n16669 : n32;
  assign n16671 = pi18 ? n139 : n16670;
  assign n16672 = pi17 ? n16668 : n16671;
  assign n16673 = pi16 ? n439 : n16672;
  assign n16674 = pi20 ? n13119 : n139;
  assign n16675 = pi19 ? n37 : n16674;
  assign n16676 = pi18 ? n16675 : n139;
  assign n16677 = pi20 ? n139 : n2653;
  assign n16678 = pi19 ? n16677 : n32;
  assign n16679 = pi18 ? n139 : n16678;
  assign n16680 = pi17 ? n16676 : n16679;
  assign n16681 = pi16 ? n439 : n16680;
  assign n16682 = pi15 ? n16673 : n16681;
  assign n16683 = pi20 ? n947 : n2653;
  assign n16684 = pi19 ? n16683 : n32;
  assign n16685 = pi18 ? n16049 : n16684;
  assign n16686 = pi17 ? n16046 : n16685;
  assign n16687 = pi16 ? n439 : n16686;
  assign n16688 = pi20 ? n3916 : n14988;
  assign n16689 = pi19 ? n16057 : n16688;
  assign n16690 = pi18 ? n16056 : n16689;
  assign n16691 = pi20 ? n2512 : n3654;
  assign n16692 = pi19 ? n16691 : n1715;
  assign n16693 = pi20 ? n2543 : n2653;
  assign n16694 = pi19 ? n16693 : n32;
  assign n16695 = pi18 ? n16692 : n16694;
  assign n16696 = pi17 ? n16690 : n16695;
  assign n16697 = pi16 ? n439 : n16696;
  assign n16698 = pi15 ? n16687 : n16697;
  assign n16699 = pi14 ? n16682 : n16698;
  assign n16700 = pi13 ? n16665 : n16699;
  assign n16701 = pi12 ? n16634 : n16700;
  assign n16702 = pi21 ? n37 : n1711;
  assign n16703 = pi21 ? n375 : n1531;
  assign n16704 = pi20 ? n16702 : n16703;
  assign n16705 = pi19 ? n12370 : n16704;
  assign n16706 = pi18 ? n37 : n16705;
  assign n16707 = pi20 ? n16078 : n2512;
  assign n16708 = pi19 ? n16079 : n16707;
  assign n16709 = pi20 ? n1708 : n2653;
  assign n16710 = pi19 ? n16709 : n32;
  assign n16711 = pi18 ? n16708 : n16710;
  assign n16712 = pi17 ? n16706 : n16711;
  assign n16713 = pi16 ? n439 : n16712;
  assign n16714 = pi15 ? n16713 : n16091;
  assign n16715 = pi14 ? n16714 : n16105;
  assign n16716 = pi13 ? n16715 : n16145;
  assign n16717 = pi23 ? n6960 : n233;
  assign n16718 = pi22 ? n335 : n16717;
  assign n16719 = pi21 ? n335 : n16718;
  assign n16720 = pi20 ? n16719 : n32;
  assign n16721 = pi19 ? n16720 : n32;
  assign n16722 = pi18 ? n16147 : n16721;
  assign n16723 = pi17 ? n37 : n16722;
  assign n16724 = pi16 ? n439 : n16723;
  assign n16725 = pi21 ? n1943 : n16718;
  assign n16726 = pi20 ? n16725 : n32;
  assign n16727 = pi19 ? n16726 : n32;
  assign n16728 = pi18 ? n16154 : n16727;
  assign n16729 = pi17 ? n37 : n16728;
  assign n16730 = pi16 ? n439 : n16729;
  assign n16731 = pi15 ? n16724 : n16730;
  assign n16732 = pi20 ? n16725 : n2679;
  assign n16733 = pi19 ? n16732 : n32;
  assign n16734 = pi18 ? n16162 : n16733;
  assign n16735 = pi17 ? n37 : n16734;
  assign n16736 = pi16 ? n439 : n16735;
  assign n16737 = pi15 ? n16736 : n16177;
  assign n16738 = pi14 ? n16731 : n16737;
  assign n16739 = pi21 ? n335 : n8860;
  assign n16740 = pi20 ? n16739 : n32;
  assign n16741 = pi19 ? n16740 : n32;
  assign n16742 = pi18 ? n16181 : n16741;
  assign n16743 = pi17 ? n37 : n16742;
  assign n16744 = pi16 ? n439 : n16743;
  assign n16745 = pi21 ? n9666 : n1389;
  assign n16746 = pi20 ? n16745 : n32;
  assign n16747 = pi19 ? n16746 : n32;
  assign n16748 = pi18 ? n16191 : n16747;
  assign n16749 = pi17 ? n37 : n16748;
  assign n16750 = pi16 ? n439 : n16749;
  assign n16751 = pi15 ? n16744 : n16750;
  assign n16752 = pi22 ? n5011 : n1070;
  assign n16753 = pi21 ? n3392 : n16752;
  assign n16754 = pi20 ? n16753 : n32;
  assign n16755 = pi19 ? n16754 : n32;
  assign n16756 = pi18 ? n16201 : n16755;
  assign n16757 = pi17 ? n37 : n16756;
  assign n16758 = pi16 ? n439 : n16757;
  assign n16759 = pi22 ? n559 : n1388;
  assign n16760 = pi21 ? n233 : n16759;
  assign n16761 = pi20 ? n16760 : n32;
  assign n16762 = pi19 ? n16761 : n32;
  assign n16763 = pi18 ? n16209 : n16762;
  assign n16764 = pi17 ? n37 : n16763;
  assign n16765 = pi16 ? n439 : n16764;
  assign n16766 = pi15 ? n16758 : n16765;
  assign n16767 = pi14 ? n16751 : n16766;
  assign n16768 = pi13 ? n16738 : n16767;
  assign n16769 = pi12 ? n16716 : n16768;
  assign n16770 = pi11 ? n16701 : n16769;
  assign n16771 = pi23 ? n363 : n687;
  assign n16772 = pi22 ? n559 : n16771;
  assign n16773 = pi21 ? n363 : n16772;
  assign n16774 = pi20 ? n16773 : n32;
  assign n16775 = pi19 ? n16774 : n32;
  assign n16776 = pi18 ? n16223 : n16775;
  assign n16777 = pi17 ? n37 : n16776;
  assign n16778 = pi16 ? n439 : n16777;
  assign n16779 = pi22 ? n14245 : n759;
  assign n16780 = pi21 ? n363 : n16779;
  assign n16781 = pi20 ? n16780 : n32;
  assign n16782 = pi19 ? n16781 : n32;
  assign n16783 = pi18 ? n16223 : n16782;
  assign n16784 = pi17 ? n15176 : n16783;
  assign n16785 = pi16 ? n439 : n16784;
  assign n16786 = pi15 ? n16778 : n16785;
  assign n16787 = pi21 ? n685 : n2147;
  assign n16788 = pi20 ? n16787 : n32;
  assign n16789 = pi19 ? n16788 : n32;
  assign n16790 = pi18 ? n16239 : n16789;
  assign n16791 = pi17 ? n37 : n16790;
  assign n16792 = pi16 ? n439 : n16791;
  assign n16793 = pi21 ? n2106 : n2147;
  assign n16794 = pi20 ? n16793 : n32;
  assign n16795 = pi19 ? n16794 : n32;
  assign n16796 = pi18 ? n37 : n16795;
  assign n16797 = pi17 ? n37 : n16796;
  assign n16798 = pi16 ? n439 : n16797;
  assign n16799 = pi15 ? n16792 : n16798;
  assign n16800 = pi14 ? n16786 : n16799;
  assign n16801 = pi22 ? n686 : n759;
  assign n16802 = pi21 ? n2106 : n16801;
  assign n16803 = pi20 ? n16802 : n32;
  assign n16804 = pi19 ? n16803 : n32;
  assign n16805 = pi18 ? n37 : n16804;
  assign n16806 = pi17 ? n37 : n16805;
  assign n16807 = pi16 ? n439 : n16806;
  assign n16808 = pi15 ? n16798 : n16807;
  assign n16809 = pi18 ? n15205 : n16795;
  assign n16810 = pi17 ? n99 : n16809;
  assign n16811 = pi16 ? n201 : n16810;
  assign n16812 = pi22 ? n2244 : n396;
  assign n16813 = pi21 ? n767 : n16812;
  assign n16814 = pi20 ? n16813 : n32;
  assign n16815 = pi19 ? n16814 : n32;
  assign n16816 = pi18 ? n16265 : n16815;
  assign n16817 = pi17 ? n99 : n16816;
  assign n16818 = pi16 ? n721 : n16817;
  assign n16819 = pi15 ? n16811 : n16818;
  assign n16820 = pi14 ? n16808 : n16819;
  assign n16821 = pi13 ? n16800 : n16820;
  assign n16822 = pi22 ? n2244 : n1407;
  assign n16823 = pi21 ? n157 : n16822;
  assign n16824 = pi20 ? n16823 : n32;
  assign n16825 = pi19 ? n16824 : n32;
  assign n16826 = pi18 ? n16281 : n16825;
  assign n16827 = pi17 ? n16278 : n16826;
  assign n16828 = pi16 ? n721 : n16827;
  assign n16829 = pi21 ? n168 : n16266;
  assign n16830 = pi20 ? n16829 : n32;
  assign n16831 = pi19 ? n16830 : n32;
  assign n16832 = pi18 ? n16295 : n16831;
  assign n16833 = pi17 ? n16291 : n16832;
  assign n16834 = pi16 ? n721 : n16833;
  assign n16835 = pi15 ? n16828 : n16834;
  assign n16836 = pi21 ? n7414 : n99;
  assign n16837 = pi20 ? n32 : n16836;
  assign n16838 = pi19 ? n32 : n16837;
  assign n16839 = pi18 ? n16838 : n16308;
  assign n16840 = pi17 ? n32 : n16839;
  assign n16841 = pi22 ? n1484 : n317;
  assign n16842 = pi21 ? n157 : n16841;
  assign n16843 = pi20 ? n16842 : n32;
  assign n16844 = pi19 ? n16843 : n32;
  assign n16845 = pi18 ? n16316 : n16844;
  assign n16846 = pi17 ? n16314 : n16845;
  assign n16847 = pi16 ? n16840 : n16846;
  assign n16848 = pi16 ? n7419 : n16328;
  assign n16849 = pi15 ? n16847 : n16848;
  assign n16850 = pi14 ? n16835 : n16849;
  assign n16851 = pi16 ? n12535 : n16343;
  assign n16852 = pi20 ? n1486 : n32;
  assign n16853 = pi19 ? n16852 : n32;
  assign n16854 = pi18 ? n157 : n16853;
  assign n16855 = pi17 ? n157 : n16854;
  assign n16856 = pi16 ? n12535 : n16855;
  assign n16857 = pi15 ? n16851 : n16856;
  assign n16858 = pi21 ? n777 : n2300;
  assign n16859 = pi20 ? n16858 : n32;
  assign n16860 = pi19 ? n16859 : n32;
  assign n16861 = pi18 ? n99 : n16860;
  assign n16862 = pi17 ? n99 : n16861;
  assign n16863 = pi16 ? n744 : n16862;
  assign n16864 = pi21 ? n910 : n248;
  assign n16865 = pi20 ? n32 : n16864;
  assign n16866 = pi19 ? n32 : n16865;
  assign n16867 = pi18 ? n16866 : n2281;
  assign n16868 = pi17 ? n32 : n16867;
  assign n16869 = pi21 ? n316 : n4109;
  assign n16870 = pi20 ? n16869 : n32;
  assign n16871 = pi19 ? n16870 : n32;
  assign n16872 = pi18 ? n16381 : n16871;
  assign n16873 = pi17 ? n16378 : n16872;
  assign n16874 = pi16 ? n16868 : n16873;
  assign n16875 = pi15 ? n16863 : n16874;
  assign n16876 = pi14 ? n16857 : n16875;
  assign n16877 = pi13 ? n16850 : n16876;
  assign n16878 = pi12 ? n16821 : n16877;
  assign n16879 = pi21 ? n2319 : n2835;
  assign n16880 = pi20 ? n16879 : n32;
  assign n16881 = pi19 ? n16880 : n32;
  assign n16882 = pi18 ? n139 : n16881;
  assign n16883 = pi17 ? n16394 : n16882;
  assign n16884 = pi16 ? n915 : n16883;
  assign n16885 = pi16 ? n915 : n16406;
  assign n16886 = pi15 ? n16884 : n16885;
  assign n16887 = pi16 ? n915 : n16415;
  assign n16888 = pi15 ? n16887 : n16425;
  assign n16889 = pi14 ? n16886 : n16888;
  assign n16890 = pi24 ? n139 : n204;
  assign n16891 = pi23 ? n16890 : n316;
  assign n16892 = pi22 ? n204 : n16891;
  assign n16893 = pi21 ? n16892 : n928;
  assign n16894 = pi20 ? n16893 : n32;
  assign n16895 = pi19 ? n16894 : n32;
  assign n16896 = pi18 ? n316 : n16895;
  assign n16897 = pi17 ? n16437 : n16896;
  assign n16898 = pi16 ? n11772 : n16897;
  assign n16899 = pi15 ? n16434 : n16898;
  assign n16900 = pi20 ? n3656 : n2512;
  assign n16901 = pi19 ? n16900 : n2512;
  assign n16902 = pi18 ? n1573 : n16901;
  assign n16903 = pi17 ? n32 : n16902;
  assign n16904 = pi21 ? n3617 : n1531;
  assign n16905 = pi20 ? n16904 : n11579;
  assign n16906 = pi22 ? n348 : n1043;
  assign n16907 = pi21 ? n16906 : n1785;
  assign n16908 = pi20 ? n11277 : n16907;
  assign n16909 = pi19 ? n16905 : n16908;
  assign n16910 = pi18 ? n16457 : n16909;
  assign n16911 = pi21 ? n1211 : n3617;
  assign n16912 = pi20 ? n8719 : n16911;
  assign n16913 = pi20 ? n3245 : n5961;
  assign n16914 = pi19 ? n16912 : n16913;
  assign n16915 = pi22 ? n1038 : n3762;
  assign n16916 = pi21 ? n16915 : n1009;
  assign n16917 = pi20 ? n16916 : n32;
  assign n16918 = pi19 ? n16917 : n32;
  assign n16919 = pi18 ? n16914 : n16918;
  assign n16920 = pi17 ? n16910 : n16919;
  assign n16921 = pi16 ? n16903 : n16920;
  assign n16922 = pi23 ? n204 : n2120;
  assign n16923 = pi22 ? n204 : n16922;
  assign n16924 = pi21 ? n16923 : n1009;
  assign n16925 = pi20 ? n16924 : n32;
  assign n16926 = pi19 ? n16925 : n32;
  assign n16927 = pi18 ? n15406 : n16926;
  assign n16928 = pi17 ? n16475 : n16927;
  assign n16929 = pi16 ? n15849 : n16928;
  assign n16930 = pi15 ? n16921 : n16929;
  assign n16931 = pi14 ? n16899 : n16930;
  assign n16932 = pi13 ? n16889 : n16931;
  assign n16933 = pi22 ? n204 : n3318;
  assign n16934 = pi21 ? n16933 : n32;
  assign n16935 = pi20 ? n16934 : n32;
  assign n16936 = pi19 ? n16935 : n32;
  assign n16937 = pi18 ? n204 : n16936;
  assign n16938 = pi17 ? n15430 : n16937;
  assign n16939 = pi16 ? n16504 : n16938;
  assign n16940 = pi15 ? n16499 : n16939;
  assign n16941 = pi18 ? n15438 : n9433;
  assign n16942 = pi17 ? n335 : n16941;
  assign n16943 = pi16 ? n7943 : n16942;
  assign n16944 = pi21 ? n10981 : n32;
  assign n16945 = pi20 ? n16944 : n32;
  assign n16946 = pi19 ? n16945 : n32;
  assign n16947 = pi18 ? n335 : n16946;
  assign n16948 = pi17 ? n16518 : n16947;
  assign n16949 = pi16 ? n2035 : n16948;
  assign n16950 = pi15 ? n16943 : n16949;
  assign n16951 = pi14 ? n16940 : n16950;
  assign n16952 = pi16 ? n2035 : n16528;
  assign n16953 = pi16 ? n10980 : n16535;
  assign n16954 = pi15 ? n16952 : n16953;
  assign n16955 = pi16 ? n12648 : n16551;
  assign n16956 = pi22 ? n12652 : n233;
  assign n16957 = pi21 ? n16956 : n335;
  assign n16958 = pi20 ? n32 : n16957;
  assign n16959 = pi19 ? n32 : n16958;
  assign n16960 = pi18 ? n16959 : n16559;
  assign n16961 = pi17 ? n32 : n16960;
  assign n16962 = pi16 ? n16961 : n16572;
  assign n16963 = pi15 ? n16955 : n16962;
  assign n16964 = pi14 ? n16954 : n16963;
  assign n16965 = pi13 ? n16951 : n16964;
  assign n16966 = pi12 ? n16932 : n16965;
  assign n16967 = pi11 ? n16878 : n16966;
  assign n16968 = pi10 ? n16770 : n16967;
  assign n16969 = pi09 ? n16588 : n16968;
  assign n16970 = pi08 ? n16580 : n16969;
  assign n16971 = pi07 ? n15907 : n16970;
  assign n16972 = pi20 ? n37 : n3792;
  assign n16973 = pi19 ? n16972 : n32;
  assign n16974 = pi18 ? n37 : n16973;
  assign n16975 = pi17 ? n37 : n16974;
  assign n16976 = pi16 ? n11011 : n16975;
  assign n16977 = pi15 ? n32 : n16976;
  assign n16978 = pi16 ? n11885 : n16975;
  assign n16979 = pi16 ? n12689 : n16975;
  assign n16980 = pi15 ? n16978 : n16979;
  assign n16981 = pi14 ? n16977 : n16980;
  assign n16982 = pi13 ? n32 : n16981;
  assign n16983 = pi12 ? n32 : n16982;
  assign n16984 = pi11 ? n32 : n16983;
  assign n16985 = pi10 ? n32 : n16984;
  assign n16986 = pi20 ? n99 : n3833;
  assign n16987 = pi19 ? n16986 : n32;
  assign n16988 = pi18 ? n37 : n16987;
  assign n16989 = pi17 ? n37 : n16988;
  assign n16990 = pi16 ? n13561 : n16989;
  assign n16991 = pi21 ? n9629 : n32;
  assign n16992 = pi20 ? n99 : n16991;
  assign n16993 = pi19 ? n16992 : n32;
  assign n16994 = pi18 ? n37 : n16993;
  assign n16995 = pi17 ? n37 : n16994;
  assign n16996 = pi16 ? n14445 : n16995;
  assign n16997 = pi15 ? n16990 : n16996;
  assign n16998 = pi18 ? n37 : n15952;
  assign n16999 = pi20 ? n37 : n2973;
  assign n17000 = pi19 ? n16999 : n37;
  assign n17001 = pi21 ? n11994 : n32;
  assign n17002 = pi20 ? n181 : n17001;
  assign n17003 = pi19 ? n17002 : n32;
  assign n17004 = pi18 ? n17000 : n17003;
  assign n17005 = pi17 ? n16998 : n17004;
  assign n17006 = pi16 ? n16595 : n17005;
  assign n17007 = pi20 ? n32 : n66;
  assign n17008 = pi19 ? n32 : n17007;
  assign n17009 = pi18 ? n17008 : n37;
  assign n17010 = pi17 ? n32 : n17009;
  assign n17011 = pi19 ? n37 : n5077;
  assign n17012 = pi20 ? n7747 : n37;
  assign n17013 = pi20 ? n37 : n5077;
  assign n17014 = pi19 ? n17012 : n17013;
  assign n17015 = pi18 ? n17011 : n17014;
  assign n17016 = pi20 ? n221 : n7745;
  assign n17017 = pi20 ? n11420 : n5077;
  assign n17018 = pi19 ? n17016 : n17017;
  assign n17019 = pi18 ? n17018 : n15928;
  assign n17020 = pi17 ? n17015 : n17019;
  assign n17021 = pi16 ? n17010 : n17020;
  assign n17022 = pi15 ? n17006 : n17021;
  assign n17023 = pi14 ? n16997 : n17022;
  assign n17024 = pi21 ? n2168 : n37;
  assign n17025 = pi20 ? n37 : n17024;
  assign n17026 = pi19 ? n17025 : n37;
  assign n17027 = pi20 ? n2970 : n3067;
  assign n17028 = pi19 ? n17027 : n32;
  assign n17029 = pi18 ? n17026 : n17028;
  assign n17030 = pi17 ? n37 : n17029;
  assign n17031 = pi16 ? n439 : n17030;
  assign n17032 = pi21 ? n9238 : n32;
  assign n17033 = pi20 ? n37 : n17032;
  assign n17034 = pi19 ? n17033 : n32;
  assign n17035 = pi18 ? n37 : n17034;
  assign n17036 = pi17 ? n37 : n17035;
  assign n17037 = pi16 ? n439 : n17036;
  assign n17038 = pi15 ? n17031 : n17037;
  assign n17039 = pi20 ? n7745 : n16621;
  assign n17040 = pi19 ? n17039 : n32;
  assign n17041 = pi18 ? n37 : n17040;
  assign n17042 = pi17 ? n37 : n17041;
  assign n17043 = pi16 ? n439 : n17042;
  assign n17044 = pi22 ? n171 : n32;
  assign n17045 = pi21 ? n17044 : n32;
  assign n17046 = pi20 ? n7745 : n17045;
  assign n17047 = pi19 ? n17046 : n32;
  assign n17048 = pi18 ? n37 : n17047;
  assign n17049 = pi17 ? n37 : n17048;
  assign n17050 = pi16 ? n439 : n17049;
  assign n17051 = pi15 ? n17043 : n17050;
  assign n17052 = pi14 ? n17038 : n17051;
  assign n17053 = pi13 ? n17023 : n17052;
  assign n17054 = pi20 ? n99 : n17045;
  assign n17055 = pi19 ? n17054 : n32;
  assign n17056 = pi18 ? n99 : n17055;
  assign n17057 = pi17 ? n99 : n17056;
  assign n17058 = pi16 ? n201 : n17057;
  assign n17059 = pi16 ? n801 : n16643;
  assign n17060 = pi15 ? n17058 : n17059;
  assign n17061 = pi19 ? n37 : n9824;
  assign n17062 = pi18 ? n374 : n17061;
  assign n17063 = pi17 ? n32 : n17062;
  assign n17064 = pi20 ? n139 : n2579;
  assign n17065 = pi19 ? n17064 : n32;
  assign n17066 = pi18 ? n139 : n17065;
  assign n17067 = pi17 ? n139 : n17066;
  assign n17068 = pi16 ? n17063 : n17067;
  assign n17069 = pi15 ? n16644 : n17068;
  assign n17070 = pi14 ? n17060 : n17069;
  assign n17071 = pi20 ? n37 : n16047;
  assign n17072 = pi19 ? n17071 : n139;
  assign n17073 = pi18 ? n17072 : n139;
  assign n17074 = pi17 ? n17073 : n17066;
  assign n17075 = pi16 ? n439 : n17074;
  assign n17076 = pi20 ? n376 : n942;
  assign n17077 = pi19 ? n37 : n17076;
  assign n17078 = pi21 ? n3668 : n1721;
  assign n17079 = pi20 ? n17078 : n139;
  assign n17080 = pi19 ? n17079 : n139;
  assign n17081 = pi18 ? n17077 : n17080;
  assign n17082 = pi20 ? n139 : n10011;
  assign n17083 = pi19 ? n17082 : n32;
  assign n17084 = pi18 ? n139 : n17083;
  assign n17085 = pi17 ? n17081 : n17084;
  assign n17086 = pi16 ? n439 : n17085;
  assign n17087 = pi15 ? n17075 : n17086;
  assign n17088 = pi19 ? n8743 : n16059;
  assign n17089 = pi18 ? n37 : n17088;
  assign n17090 = pi20 ? n3090 : n3086;
  assign n17091 = pi20 ? n3086 : n3074;
  assign n17092 = pi19 ? n17090 : n17091;
  assign n17093 = pi20 ? n3096 : n10011;
  assign n17094 = pi19 ? n17093 : n32;
  assign n17095 = pi18 ? n17092 : n17094;
  assign n17096 = pi17 ? n17089 : n17095;
  assign n17097 = pi16 ? n439 : n17096;
  assign n17098 = pi20 ? n8742 : n37;
  assign n17099 = pi19 ? n37 : n17098;
  assign n17100 = pi18 ? n37 : n17099;
  assign n17101 = pi20 ? n37 : n3074;
  assign n17102 = pi19 ? n37 : n17101;
  assign n17103 = pi18 ? n17102 : n17094;
  assign n17104 = pi17 ? n17100 : n17103;
  assign n17105 = pi16 ? n439 : n17104;
  assign n17106 = pi15 ? n17097 : n17105;
  assign n17107 = pi14 ? n17087 : n17106;
  assign n17108 = pi13 ? n17070 : n17107;
  assign n17109 = pi12 ? n17053 : n17108;
  assign n17110 = pi20 ? n37 : n13118;
  assign n17111 = pi19 ? n37 : n17110;
  assign n17112 = pi18 ? n37 : n17111;
  assign n17113 = pi23 ? n8160 : n395;
  assign n17114 = pi22 ? n17113 : n32;
  assign n17115 = pi21 ? n17114 : n32;
  assign n17116 = pi20 ? n3645 : n17115;
  assign n17117 = pi19 ? n17116 : n32;
  assign n17118 = pi18 ? n16081 : n17117;
  assign n17119 = pi17 ? n17112 : n17118;
  assign n17120 = pi16 ? n439 : n17119;
  assign n17121 = pi23 ? n8160 : n32;
  assign n17122 = pi22 ? n17121 : n32;
  assign n17123 = pi21 ? n17122 : n32;
  assign n17124 = pi20 ? n139 : n17123;
  assign n17125 = pi19 ? n17124 : n32;
  assign n17126 = pi18 ? n139 : n17125;
  assign n17127 = pi17 ? n16094 : n17126;
  assign n17128 = pi16 ? n439 : n17127;
  assign n17129 = pi15 ? n17120 : n17128;
  assign n17130 = pi21 ? n139 : n1313;
  assign n17131 = pi20 ? n17130 : n14847;
  assign n17132 = pi19 ? n17131 : n32;
  assign n17133 = pi18 ? n9770 : n17132;
  assign n17134 = pi17 ? n37 : n17133;
  assign n17135 = pi16 ? n439 : n17134;
  assign n17136 = pi21 ? n1696 : n1529;
  assign n17137 = pi20 ? n17136 : n12014;
  assign n17138 = pi19 ? n17137 : n14578;
  assign n17139 = pi21 ? n1529 : n2585;
  assign n17140 = pi20 ? n17139 : n2554;
  assign n17141 = pi19 ? n17140 : n32;
  assign n17142 = pi18 ? n17138 : n17141;
  assign n17143 = pi17 ? n37 : n17142;
  assign n17144 = pi16 ? n439 : n17143;
  assign n17145 = pi15 ? n17135 : n17144;
  assign n17146 = pi14 ? n17129 : n17145;
  assign n17147 = pi21 ? n522 : n520;
  assign n17148 = pi20 ? n5733 : n17147;
  assign n17149 = pi22 ? n448 : n455;
  assign n17150 = pi21 ? n522 : n17149;
  assign n17151 = pi22 ? n448 : n204;
  assign n17152 = pi21 ? n204 : n17151;
  assign n17153 = pi20 ? n17150 : n17152;
  assign n17154 = pi19 ? n17148 : n17153;
  assign n17155 = pi21 ? n464 : n204;
  assign n17156 = pi20 ? n17155 : n15978;
  assign n17157 = pi19 ? n17156 : n32;
  assign n17158 = pi18 ? n17154 : n17157;
  assign n17159 = pi17 ? n37 : n17158;
  assign n17160 = pi16 ? n439 : n17159;
  assign n17161 = pi21 ? n457 : n485;
  assign n17162 = pi20 ? n37 : n17161;
  assign n17163 = pi21 ? n522 : n1940;
  assign n17164 = pi21 ? n204 : n1940;
  assign n17165 = pi20 ? n17163 : n17164;
  assign n17166 = pi19 ? n17162 : n17165;
  assign n17167 = pi21 ? n464 : n8842;
  assign n17168 = pi20 ? n17167 : n2554;
  assign n17169 = pi19 ? n17168 : n32;
  assign n17170 = pi18 ? n17166 : n17169;
  assign n17171 = pi17 ? n37 : n17170;
  assign n17172 = pi16 ? n439 : n17171;
  assign n17173 = pi15 ? n17160 : n17172;
  assign n17174 = pi21 ? n1920 : n4893;
  assign n17175 = pi20 ? n37 : n17174;
  assign n17176 = pi21 ? n3411 : n4893;
  assign n17177 = pi21 ? n233 : n4893;
  assign n17178 = pi20 ? n17176 : n17177;
  assign n17179 = pi19 ? n17175 : n17178;
  assign n17180 = pi21 ? n559 : n4912;
  assign n17181 = pi20 ? n17180 : n2470;
  assign n17182 = pi19 ? n17181 : n32;
  assign n17183 = pi18 ? n17179 : n17182;
  assign n17184 = pi17 ? n37 : n17183;
  assign n17185 = pi16 ? n439 : n17184;
  assign n17186 = pi21 ? n4900 : n4908;
  assign n17187 = pi21 ? n4903 : n4908;
  assign n17188 = pi20 ? n17186 : n17187;
  assign n17189 = pi19 ? n11653 : n17188;
  assign n17190 = pi21 ? n2060 : n4899;
  assign n17191 = pi20 ? n17190 : n2679;
  assign n17192 = pi19 ? n17191 : n32;
  assign n17193 = pi18 ? n17189 : n17192;
  assign n17194 = pi17 ? n37 : n17193;
  assign n17195 = pi16 ? n439 : n17194;
  assign n17196 = pi15 ? n17185 : n17195;
  assign n17197 = pi14 ? n17173 : n17196;
  assign n17198 = pi13 ? n17146 : n17197;
  assign n17199 = pi20 ? n13527 : n2554;
  assign n17200 = pi19 ? n17199 : n32;
  assign n17201 = pi18 ? n9856 : n17200;
  assign n17202 = pi17 ? n37 : n17201;
  assign n17203 = pi16 ? n439 : n17202;
  assign n17204 = pi20 ? n37 : n335;
  assign n17205 = pi19 ? n37 : n17204;
  assign n17206 = pi23 ? n6960 : n316;
  assign n17207 = pi22 ? n37 : n17206;
  assign n17208 = pi21 ? n335 : n17207;
  assign n17209 = pi20 ? n17208 : n2679;
  assign n17210 = pi19 ? n17209 : n32;
  assign n17211 = pi18 ? n17205 : n17210;
  assign n17212 = pi17 ? n37 : n17211;
  assign n17213 = pi16 ? n439 : n17212;
  assign n17214 = pi15 ? n17203 : n17213;
  assign n17215 = pi20 ? n37 : n605;
  assign n17216 = pi19 ? n37 : n17215;
  assign n17217 = pi22 ? n37 : n16717;
  assign n17218 = pi21 ? n569 : n17217;
  assign n17219 = pi20 ? n17218 : n2679;
  assign n17220 = pi19 ? n17219 : n32;
  assign n17221 = pi18 ? n17216 : n17220;
  assign n17222 = pi17 ? n37 : n17221;
  assign n17223 = pi16 ? n439 : n17222;
  assign n17224 = pi20 ? n37 : n569;
  assign n17225 = pi19 ? n37 : n17224;
  assign n17226 = pi23 ? n10729 : n685;
  assign n17227 = pi22 ? n37 : n17226;
  assign n17228 = pi21 ? n569 : n17227;
  assign n17229 = pi20 ? n17228 : n2701;
  assign n17230 = pi19 ? n17229 : n32;
  assign n17231 = pi18 ? n17225 : n17230;
  assign n17232 = pi17 ? n37 : n17231;
  assign n17233 = pi16 ? n439 : n17232;
  assign n17234 = pi15 ? n17223 : n17233;
  assign n17235 = pi14 ? n17214 : n17234;
  assign n17236 = pi21 ? n2007 : n3392;
  assign n17237 = pi20 ? n37 : n17236;
  assign n17238 = pi19 ? n37 : n17237;
  assign n17239 = pi23 ? n1991 : n685;
  assign n17240 = pi22 ? n583 : n17239;
  assign n17241 = pi21 ? n569 : n17240;
  assign n17242 = pi20 ? n17241 : n1822;
  assign n17243 = pi19 ? n17242 : n32;
  assign n17244 = pi18 ? n17238 : n17243;
  assign n17245 = pi17 ? n37 : n17244;
  assign n17246 = pi16 ? n439 : n17245;
  assign n17247 = pi21 ? n37 : n10282;
  assign n17248 = pi20 ? n17247 : n32;
  assign n17249 = pi19 ? n17248 : n32;
  assign n17250 = pi18 ? n37 : n17249;
  assign n17251 = pi17 ? n37 : n17250;
  assign n17252 = pi16 ? n439 : n17251;
  assign n17253 = pi15 ? n17246 : n17252;
  assign n17254 = pi20 ? n37 : n2092;
  assign n17255 = pi19 ? n37 : n17254;
  assign n17256 = pi22 ? n7024 : n2121;
  assign n17257 = pi21 ? n1920 : n17256;
  assign n17258 = pi20 ? n17257 : n32;
  assign n17259 = pi19 ? n17258 : n32;
  assign n17260 = pi18 ? n17255 : n17259;
  assign n17261 = pi17 ? n37 : n17260;
  assign n17262 = pi16 ? n439 : n17261;
  assign n17263 = pi21 ? n2091 : n1389;
  assign n17264 = pi20 ? n17263 : n32;
  assign n17265 = pi19 ? n17264 : n32;
  assign n17266 = pi18 ? n17255 : n17265;
  assign n17267 = pi17 ? n37 : n17266;
  assign n17268 = pi16 ? n439 : n17267;
  assign n17269 = pi15 ? n17262 : n17268;
  assign n17270 = pi14 ? n17253 : n17269;
  assign n17271 = pi13 ? n17235 : n17270;
  assign n17272 = pi12 ? n17198 : n17271;
  assign n17273 = pi11 ? n17109 : n17272;
  assign n17274 = pi21 ? n2106 : n37;
  assign n17275 = pi20 ? n37 : n17274;
  assign n17276 = pi19 ? n37 : n17275;
  assign n17277 = pi22 ? n685 : n14245;
  assign n17278 = pi21 ? n17277 : n2139;
  assign n17279 = pi20 ? n17278 : n32;
  assign n17280 = pi19 ? n17279 : n32;
  assign n17281 = pi18 ? n17276 : n17280;
  assign n17282 = pi17 ? n37 : n17281;
  assign n17283 = pi16 ? n439 : n17282;
  assign n17284 = pi22 ? n5011 : n759;
  assign n17285 = pi21 ? n2106 : n17284;
  assign n17286 = pi20 ? n17285 : n32;
  assign n17287 = pi19 ? n17286 : n32;
  assign n17288 = pi18 ? n37 : n17287;
  assign n17289 = pi17 ? n37 : n17288;
  assign n17290 = pi16 ? n439 : n17289;
  assign n17291 = pi15 ? n17283 : n17290;
  assign n17292 = pi21 ? n2106 : n16779;
  assign n17293 = pi20 ? n17292 : n32;
  assign n17294 = pi19 ? n17293 : n32;
  assign n17295 = pi18 ? n37 : n17294;
  assign n17296 = pi17 ? n37 : n17295;
  assign n17297 = pi16 ? n439 : n17296;
  assign n17298 = pi21 ? n37 : n16779;
  assign n17299 = pi20 ? n17298 : n32;
  assign n17300 = pi19 ? n17299 : n32;
  assign n17301 = pi18 ? n37 : n17300;
  assign n17302 = pi17 ? n37 : n17301;
  assign n17303 = pi16 ? n439 : n17302;
  assign n17304 = pi15 ? n17297 : n17303;
  assign n17305 = pi14 ? n17291 : n17304;
  assign n17306 = pi19 ? n99 : n4583;
  assign n17307 = pi21 ? n2175 : n16779;
  assign n17308 = pi20 ? n17307 : n32;
  assign n17309 = pi19 ? n17308 : n32;
  assign n17310 = pi18 ? n17306 : n17309;
  assign n17311 = pi17 ? n99 : n17310;
  assign n17312 = pi16 ? n744 : n17311;
  assign n17313 = pi21 ? n3444 : n685;
  assign n17314 = pi20 ? n99 : n17313;
  assign n17315 = pi19 ? n99 : n17314;
  assign n17316 = pi22 ? n3443 : n2192;
  assign n17317 = pi21 ? n685 : n17316;
  assign n17318 = pi20 ? n17317 : n32;
  assign n17319 = pi19 ? n17318 : n32;
  assign n17320 = pi18 ? n17315 : n17319;
  assign n17321 = pi17 ? n99 : n17320;
  assign n17322 = pi16 ? n744 : n17321;
  assign n17323 = pi15 ? n17312 : n17322;
  assign n17324 = pi14 ? n17303 : n17323;
  assign n17325 = pi13 ? n17305 : n17324;
  assign n17326 = pi19 ? n99 : n15271;
  assign n17327 = pi18 ? n99 : n17326;
  assign n17328 = pi20 ? n7818 : n2243;
  assign n17329 = pi20 ? n15263 : n776;
  assign n17330 = pi19 ? n17328 : n17329;
  assign n17331 = pi21 ? n6089 : n1423;
  assign n17332 = pi20 ? n17331 : n32;
  assign n17333 = pi19 ? n17332 : n32;
  assign n17334 = pi18 ? n17330 : n17333;
  assign n17335 = pi17 ? n17327 : n17334;
  assign n17336 = pi16 ? n744 : n17335;
  assign n17337 = pi21 ? n99 : n5899;
  assign n17338 = pi20 ? n17337 : n99;
  assign n17339 = pi19 ? n17338 : n99;
  assign n17340 = pi19 ? n99 : n157;
  assign n17341 = pi18 ? n17339 : n17340;
  assign n17342 = pi20 ? n157 : n776;
  assign n17343 = pi19 ? n157 : n17342;
  assign n17344 = pi20 ? n2231 : n32;
  assign n17345 = pi19 ? n17344 : n32;
  assign n17346 = pi18 ? n17343 : n17345;
  assign n17347 = pi17 ? n17341 : n17346;
  assign n17348 = pi16 ? n744 : n17347;
  assign n17349 = pi15 ? n17336 : n17348;
  assign n17350 = pi21 ? n7815 : n777;
  assign n17351 = pi20 ? n17350 : n157;
  assign n17352 = pi19 ? n157 : n17351;
  assign n17353 = pi18 ? n17352 : n157;
  assign n17354 = pi20 ? n157 : n5085;
  assign n17355 = pi19 ? n157 : n17354;
  assign n17356 = pi18 ? n17355 : n17345;
  assign n17357 = pi17 ? n17353 : n17356;
  assign n17358 = pi16 ? n9291 : n17357;
  assign n17359 = pi20 ? n157 : n802;
  assign n17360 = pi19 ? n157 : n17359;
  assign n17361 = pi18 ? n17360 : n16320;
  assign n17362 = pi17 ? n157 : n17361;
  assign n17363 = pi16 ? n5910 : n17362;
  assign n17364 = pi15 ? n17358 : n17363;
  assign n17365 = pi14 ? n17349 : n17364;
  assign n17366 = pi21 ? n157 : n7429;
  assign n17367 = pi20 ? n157 : n17366;
  assign n17368 = pi19 ? n157 : n17367;
  assign n17369 = pi21 ? n3562 : n2320;
  assign n17370 = pi20 ? n17369 : n32;
  assign n17371 = pi19 ? n17370 : n32;
  assign n17372 = pi18 ? n17368 : n17371;
  assign n17373 = pi17 ? n157 : n17372;
  assign n17374 = pi16 ? n5910 : n17373;
  assign n17375 = pi22 ? n316 : n99;
  assign n17376 = pi21 ? n165 : n17375;
  assign n17377 = pi20 ? n157 : n17376;
  assign n17378 = pi19 ? n157 : n17377;
  assign n17379 = pi18 ? n17378 : n10596;
  assign n17380 = pi17 ? n157 : n17379;
  assign n17381 = pi16 ? n9291 : n17380;
  assign n17382 = pi15 ? n17374 : n17381;
  assign n17383 = pi21 ? n7128 : n204;
  assign n17384 = pi20 ? n32 : n17383;
  assign n17385 = pi19 ? n32 : n17384;
  assign n17386 = pi18 ? n17385 : n204;
  assign n17387 = pi17 ? n32 : n17386;
  assign n17388 = pi20 ? n157 : n204;
  assign n17389 = pi19 ? n204 : n17388;
  assign n17390 = pi21 ? n316 : n157;
  assign n17391 = pi20 ? n7909 : n17390;
  assign n17392 = pi19 ? n204 : n17391;
  assign n17393 = pi18 ? n17389 : n17392;
  assign n17394 = pi21 ? n204 : n157;
  assign n17395 = pi21 ? n157 : n204;
  assign n17396 = pi20 ? n17394 : n17395;
  assign n17397 = pi21 ? n775 : n7429;
  assign n17398 = pi20 ? n204 : n17397;
  assign n17399 = pi19 ? n17396 : n17398;
  assign n17400 = pi18 ? n17399 : n10596;
  assign n17401 = pi17 ? n17393 : n17400;
  assign n17402 = pi16 ? n17387 : n17401;
  assign n17403 = pi20 ? n16047 : n204;
  assign n17404 = pi19 ? n204 : n17403;
  assign n17405 = pi20 ? n7909 : n316;
  assign n17406 = pi19 ? n204 : n17405;
  assign n17407 = pi18 ? n17404 : n17406;
  assign n17408 = pi20 ? n7909 : n1016;
  assign n17409 = pi20 ? n204 : n2353;
  assign n17410 = pi19 ? n17408 : n17409;
  assign n17411 = pi18 ? n17410 : n10596;
  assign n17412 = pi17 ? n17407 : n17411;
  assign n17413 = pi16 ? n13833 : n17412;
  assign n17414 = pi15 ? n17402 : n17413;
  assign n17415 = pi14 ? n17382 : n17414;
  assign n17416 = pi13 ? n17365 : n17415;
  assign n17417 = pi12 ? n17325 : n17416;
  assign n17418 = pi19 ? n139 : n999;
  assign n17419 = pi18 ? n139 : n17418;
  assign n17420 = pi20 ? n5317 : n139;
  assign n17421 = pi20 ? n1022 : n1008;
  assign n17422 = pi19 ? n17420 : n17421;
  assign n17423 = pi18 ? n17422 : n10596;
  assign n17424 = pi17 ? n17419 : n17423;
  assign n17425 = pi16 ? n1575 : n17424;
  assign n17426 = pi20 ? n347 : n360;
  assign n17427 = pi19 ? n17426 : n139;
  assign n17428 = pi18 ? n17427 : n17418;
  assign n17429 = pi19 ? n316 : n16401;
  assign n17430 = pi18 ? n17429 : n10596;
  assign n17431 = pi17 ? n17428 : n17430;
  assign n17432 = pi16 ? n1575 : n17431;
  assign n17433 = pi15 ? n17425 : n17432;
  assign n17434 = pi21 ? n316 : n428;
  assign n17435 = pi20 ? n17434 : n316;
  assign n17436 = pi19 ? n316 : n17435;
  assign n17437 = pi18 ? n17436 : n316;
  assign n17438 = pi18 ? n17429 : n9757;
  assign n17439 = pi17 ? n17437 : n17438;
  assign n17440 = pi16 ? n6235 : n17439;
  assign n17441 = pi18 ? n10068 : n316;
  assign n17442 = pi17 ? n32 : n17441;
  assign n17443 = pi19 ? n316 : n9066;
  assign n17444 = pi18 ? n17443 : n316;
  assign n17445 = pi17 ? n17444 : n9758;
  assign n17446 = pi16 ? n17442 : n17445;
  assign n17447 = pi15 ? n17440 : n17446;
  assign n17448 = pi14 ? n17433 : n17447;
  assign n17449 = pi19 ? n139 : n6655;
  assign n17450 = pi20 ? n2354 : n32;
  assign n17451 = pi19 ? n17450 : n32;
  assign n17452 = pi18 ? n17449 : n17451;
  assign n17453 = pi17 ? n139 : n17452;
  assign n17454 = pi16 ? n1773 : n17453;
  assign n17455 = pi15 ? n17446 : n17454;
  assign n17456 = pi22 ? n139 : n3762;
  assign n17457 = pi21 ? n17456 : n2700;
  assign n17458 = pi20 ? n17457 : n32;
  assign n17459 = pi19 ? n17458 : n32;
  assign n17460 = pi18 ? n139 : n17459;
  assign n17461 = pi17 ? n139 : n17460;
  assign n17462 = pi16 ? n915 : n17461;
  assign n17463 = pi22 ? n204 : n13834;
  assign n17464 = pi21 ? n17463 : n1009;
  assign n17465 = pi20 ? n17464 : n32;
  assign n17466 = pi19 ? n17465 : n32;
  assign n17467 = pi18 ? n204 : n17466;
  assign n17468 = pi17 ? n204 : n17467;
  assign n17469 = pi16 ? n11804 : n17468;
  assign n17470 = pi15 ? n17462 : n17469;
  assign n17471 = pi14 ? n17455 : n17470;
  assign n17472 = pi13 ? n17448 : n17471;
  assign n17473 = pi18 ? n374 : n14149;
  assign n17474 = pi17 ? n32 : n17473;
  assign n17475 = pi19 ? n10957 : n37;
  assign n17476 = pi19 ? n17204 : n335;
  assign n17477 = pi18 ? n17475 : n17476;
  assign n17478 = pi20 ? n335 : n9180;
  assign n17479 = pi19 ? n335 : n17478;
  assign n17480 = pi18 ? n17479 : n17466;
  assign n17481 = pi17 ? n17477 : n17480;
  assign n17482 = pi16 ? n17474 : n17481;
  assign n17483 = pi20 ? n577 : n37;
  assign n17484 = pi19 ? n17483 : n37;
  assign n17485 = pi18 ? n17484 : n15099;
  assign n17486 = pi20 ? n335 : n15457;
  assign n17487 = pi19 ? n335 : n17486;
  assign n17488 = pi18 ? n17487 : n10299;
  assign n17489 = pi17 ? n17485 : n17488;
  assign n17490 = pi16 ? n439 : n17489;
  assign n17491 = pi15 ? n17482 : n17490;
  assign n17492 = pi20 ? n603 : n7980;
  assign n17493 = pi19 ? n37 : n17492;
  assign n17494 = pi18 ? n37 : n17493;
  assign n17495 = pi20 ? n577 : n649;
  assign n17496 = pi19 ? n2068 : n17495;
  assign n17497 = pi18 ? n17496 : n10299;
  assign n17498 = pi17 ? n17494 : n17497;
  assign n17499 = pi16 ? n439 : n17498;
  assign n17500 = pi20 ? n335 : n649;
  assign n17501 = pi20 ? n649 : n577;
  assign n17502 = pi19 ? n17500 : n17501;
  assign n17503 = pi18 ? n558 : n17502;
  assign n17504 = pi17 ? n32 : n17503;
  assign n17505 = pi21 ? n570 : n4938;
  assign n17506 = pi20 ? n17505 : n335;
  assign n17507 = pi19 ? n335 : n17506;
  assign n17508 = pi18 ? n17507 : n335;
  assign n17509 = pi22 ? n233 : n6415;
  assign n17510 = pi21 ? n17509 : n32;
  assign n17511 = pi20 ? n17510 : n32;
  assign n17512 = pi19 ? n17511 : n32;
  assign n17513 = pi18 ? n335 : n17512;
  assign n17514 = pi17 ? n17508 : n17513;
  assign n17515 = pi16 ? n17504 : n17514;
  assign n17516 = pi15 ? n17499 : n17515;
  assign n17517 = pi14 ? n17491 : n17516;
  assign n17518 = pi20 ? n6969 : n649;
  assign n17519 = pi19 ? n17518 : n649;
  assign n17520 = pi18 ? n3284 : n17519;
  assign n17521 = pi17 ? n32 : n17520;
  assign n17522 = pi20 ? n7646 : n335;
  assign n17523 = pi19 ? n335 : n17522;
  assign n17524 = pi18 ? n17523 : n335;
  assign n17525 = pi18 ? n17487 : n16946;
  assign n17526 = pi17 ? n17524 : n17525;
  assign n17527 = pi16 ? n17521 : n17526;
  assign n17528 = pi21 ? n1592 : n335;
  assign n17529 = pi20 ? n32 : n17528;
  assign n17530 = pi19 ? n32 : n17529;
  assign n17531 = pi18 ? n17530 : n335;
  assign n17532 = pi17 ? n32 : n17531;
  assign n17533 = pi20 ? n13527 : n7980;
  assign n17534 = pi19 ? n335 : n17533;
  assign n17535 = pi18 ? n335 : n17534;
  assign n17536 = pi18 ? n17487 : n16521;
  assign n17537 = pi17 ? n17535 : n17536;
  assign n17538 = pi16 ? n17532 : n17537;
  assign n17539 = pi15 ? n17527 : n17538;
  assign n17540 = pi19 ? n335 : n13535;
  assign n17541 = pi18 ? n335 : n17540;
  assign n17542 = pi20 ? n233 : n335;
  assign n17543 = pi20 ? n7980 : n15457;
  assign n17544 = pi19 ? n17542 : n17543;
  assign n17545 = pi18 ? n17544 : n8275;
  assign n17546 = pi17 ? n17541 : n17545;
  assign n17547 = pi16 ? n10118 : n17546;
  assign n17548 = pi22 ? n363 : n335;
  assign n17549 = pi21 ? n17548 : n335;
  assign n17550 = pi20 ? n335 : n17549;
  assign n17551 = pi19 ? n15488 : n17550;
  assign n17552 = pi19 ? n13528 : n233;
  assign n17553 = pi18 ? n17551 : n17552;
  assign n17554 = pi18 ? n233 : n8919;
  assign n17555 = pi17 ? n17553 : n17554;
  assign n17556 = pi16 ? n2425 : n17555;
  assign n17557 = pi15 ? n17547 : n17556;
  assign n17558 = pi14 ? n17539 : n17557;
  assign n17559 = pi13 ? n17517 : n17558;
  assign n17560 = pi12 ? n17472 : n17559;
  assign n17561 = pi11 ? n17417 : n17560;
  assign n17562 = pi10 ? n17273 : n17561;
  assign n17563 = pi09 ? n16985 : n17562;
  assign n17564 = pi23 ? n5612 : n586;
  assign n17565 = pi22 ? n17564 : n32;
  assign n17566 = pi21 ? n17565 : n32;
  assign n17567 = pi20 ? n181 : n17566;
  assign n17568 = pi19 ? n17567 : n32;
  assign n17569 = pi18 ? n17000 : n17568;
  assign n17570 = pi17 ? n16998 : n17569;
  assign n17571 = pi16 ? n16595 : n17570;
  assign n17572 = pi15 ? n17571 : n17021;
  assign n17573 = pi14 ? n16997 : n17572;
  assign n17574 = pi23 ? n11962 : n32;
  assign n17575 = pi22 ? n17574 : n32;
  assign n17576 = pi21 ? n17575 : n32;
  assign n17577 = pi20 ? n2970 : n17576;
  assign n17578 = pi19 ? n17577 : n32;
  assign n17579 = pi18 ? n37 : n17578;
  assign n17580 = pi17 ? n37 : n17579;
  assign n17581 = pi16 ? n439 : n17580;
  assign n17582 = pi23 ? n1432 : n32;
  assign n17583 = pi22 ? n17582 : n32;
  assign n17584 = pi21 ? n17583 : n32;
  assign n17585 = pi20 ? n37 : n17584;
  assign n17586 = pi19 ? n17585 : n32;
  assign n17587 = pi18 ? n37 : n17586;
  assign n17588 = pi17 ? n37 : n17587;
  assign n17589 = pi16 ? n439 : n17588;
  assign n17590 = pi15 ? n17581 : n17589;
  assign n17591 = pi21 ? n10174 : n32;
  assign n17592 = pi20 ? n7745 : n17591;
  assign n17593 = pi19 ? n17592 : n32;
  assign n17594 = pi18 ? n37 : n17593;
  assign n17595 = pi17 ? n37 : n17594;
  assign n17596 = pi16 ? n439 : n17595;
  assign n17597 = pi20 ? n7745 : n3849;
  assign n17598 = pi19 ? n17597 : n32;
  assign n17599 = pi18 ? n37 : n17598;
  assign n17600 = pi17 ? n37 : n17599;
  assign n17601 = pi16 ? n439 : n17600;
  assign n17602 = pi15 ? n17596 : n17601;
  assign n17603 = pi14 ? n17590 : n17602;
  assign n17604 = pi13 ? n17573 : n17603;
  assign n17605 = pi20 ? n99 : n3849;
  assign n17606 = pi19 ? n17605 : n32;
  assign n17607 = pi18 ? n99 : n17606;
  assign n17608 = pi17 ? n99 : n17607;
  assign n17609 = pi16 ? n201 : n17608;
  assign n17610 = pi21 ? n10188 : n32;
  assign n17611 = pi20 ? n99 : n17610;
  assign n17612 = pi19 ? n17611 : n32;
  assign n17613 = pi18 ? n99 : n17612;
  assign n17614 = pi17 ? n99 : n17613;
  assign n17615 = pi16 ? n1510 : n17614;
  assign n17616 = pi15 ? n17609 : n17615;
  assign n17617 = pi16 ? n721 : n17614;
  assign n17618 = pi22 ? n6069 : n32;
  assign n17619 = pi21 ? n17618 : n32;
  assign n17620 = pi20 ? n139 : n17619;
  assign n17621 = pi19 ? n17620 : n32;
  assign n17622 = pi18 ? n139 : n17621;
  assign n17623 = pi17 ? n139 : n17622;
  assign n17624 = pi16 ? n17063 : n17623;
  assign n17625 = pi15 ? n17617 : n17624;
  assign n17626 = pi14 ? n17616 : n17625;
  assign n17627 = pi20 ? n37 : n8731;
  assign n17628 = pi19 ? n17627 : n139;
  assign n17629 = pi18 ? n17628 : n139;
  assign n17630 = pi22 ? n6077 : n32;
  assign n17631 = pi21 ? n17630 : n32;
  assign n17632 = pi20 ? n139 : n17631;
  assign n17633 = pi19 ? n17632 : n32;
  assign n17634 = pi18 ? n139 : n17633;
  assign n17635 = pi17 ? n17629 : n17634;
  assign n17636 = pi16 ? n439 : n17635;
  assign n17637 = pi20 ? n13118 : n942;
  assign n17638 = pi19 ? n37 : n17637;
  assign n17639 = pi20 ? n1722 : n139;
  assign n17640 = pi19 ? n17639 : n139;
  assign n17641 = pi18 ? n17638 : n17640;
  assign n17642 = pi17 ? n17641 : n17084;
  assign n17643 = pi16 ? n439 : n17642;
  assign n17644 = pi15 ? n17636 : n17643;
  assign n17645 = pi19 ? n8743 : n16688;
  assign n17646 = pi18 ? n37 : n17645;
  assign n17647 = pi20 ? n8731 : n3913;
  assign n17648 = pi19 ? n17647 : n3579;
  assign n17649 = pi20 ? n3645 : n10011;
  assign n17650 = pi19 ? n17649 : n32;
  assign n17651 = pi18 ? n17648 : n17650;
  assign n17652 = pi17 ? n17646 : n17651;
  assign n17653 = pi16 ? n439 : n17652;
  assign n17654 = pi20 ? n8742 : n8209;
  assign n17655 = pi19 ? n37 : n17654;
  assign n17656 = pi18 ? n37 : n17655;
  assign n17657 = pi19 ? n13124 : n17101;
  assign n17658 = pi18 ? n17657 : n17094;
  assign n17659 = pi17 ? n17656 : n17658;
  assign n17660 = pi16 ? n439 : n17659;
  assign n17661 = pi15 ? n17653 : n17660;
  assign n17662 = pi14 ? n17644 : n17661;
  assign n17663 = pi13 ? n17626 : n17662;
  assign n17664 = pi12 ? n17604 : n17663;
  assign n17665 = pi20 ? n1708 : n10011;
  assign n17666 = pi19 ? n17665 : n32;
  assign n17667 = pi18 ? n16708 : n17666;
  assign n17668 = pi17 ? n17112 : n17667;
  assign n17669 = pi16 ? n439 : n17668;
  assign n17670 = pi20 ? n139 : n2566;
  assign n17671 = pi19 ? n17670 : n32;
  assign n17672 = pi18 ? n139 : n17671;
  assign n17673 = pi17 ? n16094 : n17672;
  assign n17674 = pi16 ? n439 : n17673;
  assign n17675 = pi15 ? n17669 : n17674;
  assign n17676 = pi20 ? n17130 : n2566;
  assign n17677 = pi19 ? n17676 : n32;
  assign n17678 = pi18 ? n9770 : n17677;
  assign n17679 = pi17 ? n37 : n17678;
  assign n17680 = pi16 ? n439 : n17679;
  assign n17681 = pi21 ? n375 : n1696;
  assign n17682 = pi20 ? n8707 : n17681;
  assign n17683 = pi20 ? n1694 : n1693;
  assign n17684 = pi19 ? n17682 : n17683;
  assign n17685 = pi21 ? n1696 : n2585;
  assign n17686 = pi20 ? n17685 : n2566;
  assign n17687 = pi19 ? n17686 : n32;
  assign n17688 = pi18 ? n17684 : n17687;
  assign n17689 = pi17 ? n37 : n17688;
  assign n17690 = pi16 ? n439 : n17689;
  assign n17691 = pi15 ? n17680 : n17690;
  assign n17692 = pi14 ? n17675 : n17691;
  assign n17693 = pi21 ? n522 : n8834;
  assign n17694 = pi21 ? n522 : n14123;
  assign n17695 = pi20 ? n17693 : n17694;
  assign n17696 = pi19 ? n17148 : n17695;
  assign n17697 = pi21 ? n14124 : n522;
  assign n17698 = pi20 ? n17697 : n2566;
  assign n17699 = pi19 ? n17698 : n32;
  assign n17700 = pi18 ? n17696 : n17699;
  assign n17701 = pi17 ? n37 : n17700;
  assign n17702 = pi16 ? n439 : n17701;
  assign n17703 = pi21 ? n522 : n567;
  assign n17704 = pi19 ? n17162 : n17703;
  assign n17705 = pi22 ? n204 : n11047;
  assign n17706 = pi21 ? n14124 : n17705;
  assign n17707 = pi20 ? n17706 : n2579;
  assign n17708 = pi19 ? n17707 : n32;
  assign n17709 = pi18 ? n17704 : n17708;
  assign n17710 = pi17 ? n37 : n17709;
  assign n17711 = pi16 ? n439 : n17710;
  assign n17712 = pi15 ? n17702 : n17711;
  assign n17713 = pi21 ? n3411 : n569;
  assign n17714 = pi19 ? n17175 : n17713;
  assign n17715 = pi21 ? n560 : n6361;
  assign n17716 = pi20 ? n17715 : n2579;
  assign n17717 = pi19 ? n17716 : n32;
  assign n17718 = pi18 ? n17714 : n17717;
  assign n17719 = pi17 ? n37 : n17718;
  assign n17720 = pi16 ? n439 : n17719;
  assign n17721 = pi21 ? n4900 : n567;
  assign n17722 = pi22 ? n4899 : n559;
  assign n17723 = pi21 ? n17722 : n567;
  assign n17724 = pi20 ? n17721 : n17723;
  assign n17725 = pi19 ? n11653 : n17724;
  assign n17726 = pi22 ? n2060 : n566;
  assign n17727 = pi21 ? n17726 : n16562;
  assign n17728 = pi20 ? n17727 : n2579;
  assign n17729 = pi19 ? n17728 : n32;
  assign n17730 = pi18 ? n17725 : n17729;
  assign n17731 = pi17 ? n37 : n17730;
  assign n17732 = pi16 ? n439 : n17731;
  assign n17733 = pi15 ? n17720 : n17732;
  assign n17734 = pi14 ? n17712 : n17733;
  assign n17735 = pi13 ? n17692 : n17734;
  assign n17736 = pi20 ? n13527 : n2579;
  assign n17737 = pi19 ? n17736 : n32;
  assign n17738 = pi18 ? n9856 : n17737;
  assign n17739 = pi17 ? n37 : n17738;
  assign n17740 = pi16 ? n439 : n17739;
  assign n17741 = pi22 ? n37 : n6380;
  assign n17742 = pi21 ? n335 : n17741;
  assign n17743 = pi20 ? n17742 : n2579;
  assign n17744 = pi19 ? n17743 : n32;
  assign n17745 = pi18 ? n17205 : n17744;
  assign n17746 = pi17 ? n37 : n17745;
  assign n17747 = pi16 ? n439 : n17746;
  assign n17748 = pi15 ? n17740 : n17747;
  assign n17749 = pi21 ? n569 : n2074;
  assign n17750 = pi20 ? n17749 : n2579;
  assign n17751 = pi19 ? n17750 : n32;
  assign n17752 = pi18 ? n17216 : n17751;
  assign n17753 = pi17 ? n37 : n17752;
  assign n17754 = pi16 ? n439 : n17753;
  assign n17755 = pi22 ? n37 : n5782;
  assign n17756 = pi21 ? n569 : n17755;
  assign n17757 = pi20 ? n17756 : n2638;
  assign n17758 = pi19 ? n17757 : n32;
  assign n17759 = pi18 ? n17225 : n17758;
  assign n17760 = pi17 ? n37 : n17759;
  assign n17761 = pi16 ? n439 : n17760;
  assign n17762 = pi15 ? n17754 : n17761;
  assign n17763 = pi14 ? n17748 : n17762;
  assign n17764 = pi22 ? n37 : n686;
  assign n17765 = pi21 ? n584 : n17764;
  assign n17766 = pi20 ? n17765 : n2653;
  assign n17767 = pi19 ? n17766 : n32;
  assign n17768 = pi18 ? n5030 : n17767;
  assign n17769 = pi17 ? n37 : n17768;
  assign n17770 = pi16 ? n439 : n17769;
  assign n17771 = pi20 ? n17247 : n1822;
  assign n17772 = pi19 ? n17771 : n32;
  assign n17773 = pi18 ? n37 : n17772;
  assign n17774 = pi17 ? n37 : n17773;
  assign n17775 = pi16 ? n439 : n17774;
  assign n17776 = pi15 ? n17770 : n17775;
  assign n17777 = pi21 ? n1920 : n2091;
  assign n17778 = pi20 ? n17777 : n1822;
  assign n17779 = pi19 ? n17778 : n32;
  assign n17780 = pi18 ? n17255 : n17779;
  assign n17781 = pi17 ? n37 : n17780;
  assign n17782 = pi16 ? n439 : n17781;
  assign n17783 = pi20 ? n7705 : n32;
  assign n17784 = pi19 ? n17783 : n32;
  assign n17785 = pi18 ? n17255 : n17784;
  assign n17786 = pi17 ? n37 : n17785;
  assign n17787 = pi16 ? n439 : n17786;
  assign n17788 = pi15 ? n17782 : n17787;
  assign n17789 = pi14 ? n17776 : n17788;
  assign n17790 = pi13 ? n17763 : n17789;
  assign n17791 = pi12 ? n17735 : n17790;
  assign n17792 = pi11 ? n17664 : n17791;
  assign n17793 = pi21 ? n17277 : n2721;
  assign n17794 = pi20 ? n17793 : n32;
  assign n17795 = pi19 ? n17794 : n32;
  assign n17796 = pi18 ? n17276 : n17795;
  assign n17797 = pi17 ? n37 : n17796;
  assign n17798 = pi16 ? n439 : n17797;
  assign n17799 = pi21 ? n2106 : n11208;
  assign n17800 = pi20 ? n17799 : n32;
  assign n17801 = pi19 ? n17800 : n32;
  assign n17802 = pi18 ? n37 : n17801;
  assign n17803 = pi17 ? n37 : n17802;
  assign n17804 = pi16 ? n439 : n17803;
  assign n17805 = pi15 ? n17798 : n17804;
  assign n17806 = pi22 ? n14245 : n685;
  assign n17807 = pi21 ? n2106 : n17806;
  assign n17808 = pi20 ? n17807 : n32;
  assign n17809 = pi19 ? n17808 : n32;
  assign n17810 = pi18 ? n37 : n17809;
  assign n17811 = pi17 ? n37 : n17810;
  assign n17812 = pi16 ? n439 : n17811;
  assign n17813 = pi21 ? n37 : n17806;
  assign n17814 = pi20 ? n17813 : n32;
  assign n17815 = pi19 ? n17814 : n32;
  assign n17816 = pi18 ? n37 : n17815;
  assign n17817 = pi17 ? n37 : n17816;
  assign n17818 = pi16 ? n439 : n17817;
  assign n17819 = pi15 ? n17812 : n17818;
  assign n17820 = pi14 ? n17805 : n17819;
  assign n17821 = pi21 ? n2161 : n17806;
  assign n17822 = pi20 ? n17821 : n32;
  assign n17823 = pi19 ? n17822 : n32;
  assign n17824 = pi18 ? n17306 : n17823;
  assign n17825 = pi17 ? n99 : n17824;
  assign n17826 = pi16 ? n744 : n17825;
  assign n17827 = pi21 ? n685 : n4193;
  assign n17828 = pi20 ? n17827 : n32;
  assign n17829 = pi19 ? n17828 : n32;
  assign n17830 = pi18 ? n17315 : n17829;
  assign n17831 = pi17 ? n99 : n17830;
  assign n17832 = pi16 ? n744 : n17831;
  assign n17833 = pi15 ? n17826 : n17832;
  assign n17834 = pi14 ? n17818 : n17833;
  assign n17835 = pi13 ? n17820 : n17834;
  assign n17836 = pi21 ? n6089 : n2200;
  assign n17837 = pi20 ? n17836 : n32;
  assign n17838 = pi19 ? n17837 : n32;
  assign n17839 = pi18 ? n17330 : n17838;
  assign n17840 = pi17 ? n17327 : n17839;
  assign n17841 = pi16 ? n744 : n17840;
  assign n17842 = pi21 ? n99 : n10325;
  assign n17843 = pi20 ? n17842 : n32;
  assign n17844 = pi19 ? n17843 : n32;
  assign n17845 = pi18 ? n17343 : n17844;
  assign n17846 = pi17 ? n17341 : n17845;
  assign n17847 = pi16 ? n744 : n17846;
  assign n17848 = pi15 ? n17841 : n17847;
  assign n17849 = pi16 ? n7793 : n17362;
  assign n17850 = pi15 ? n17358 : n17849;
  assign n17851 = pi14 ? n17848 : n17850;
  assign n17852 = pi20 ? n3563 : n32;
  assign n17853 = pi19 ? n17852 : n32;
  assign n17854 = pi18 ? n17368 : n17853;
  assign n17855 = pi17 ? n157 : n17854;
  assign n17856 = pi16 ? n7419 : n17855;
  assign n17857 = pi18 ? n17378 : n11500;
  assign n17858 = pi17 ? n157 : n17857;
  assign n17859 = pi16 ? n8620 : n17858;
  assign n17860 = pi15 ? n17856 : n17859;
  assign n17861 = pi14 ? n17860 : n17414;
  assign n17862 = pi13 ? n17851 : n17861;
  assign n17863 = pi12 ? n17835 : n17862;
  assign n17864 = pi16 ? n331 : n17424;
  assign n17865 = pi16 ? n331 : n17431;
  assign n17866 = pi15 ? n17864 : n17865;
  assign n17867 = pi20 ? n2836 : n32;
  assign n17868 = pi19 ? n17867 : n32;
  assign n17869 = pi18 ? n17429 : n17868;
  assign n17870 = pi17 ? n17437 : n17869;
  assign n17871 = pi16 ? n6235 : n17870;
  assign n17872 = pi18 ? n316 : n17868;
  assign n17873 = pi17 ? n17444 : n17872;
  assign n17874 = pi16 ? n17442 : n17873;
  assign n17875 = pi15 ? n17871 : n17874;
  assign n17876 = pi14 ? n17866 : n17875;
  assign n17877 = pi21 ? n17456 : n928;
  assign n17878 = pi20 ? n17877 : n32;
  assign n17879 = pi19 ? n17878 : n32;
  assign n17880 = pi18 ? n139 : n17879;
  assign n17881 = pi17 ? n139 : n17880;
  assign n17882 = pi16 ? n915 : n17881;
  assign n17883 = pi21 ? n8842 : n928;
  assign n17884 = pi20 ? n17883 : n32;
  assign n17885 = pi19 ? n17884 : n32;
  assign n17886 = pi18 ? n204 : n17885;
  assign n17887 = pi17 ? n204 : n17886;
  assign n17888 = pi16 ? n11804 : n17887;
  assign n17889 = pi15 ? n17882 : n17888;
  assign n17890 = pi14 ? n17455 : n17889;
  assign n17891 = pi13 ? n17876 : n17890;
  assign n17892 = pi21 ? n3763 : n1009;
  assign n17893 = pi20 ? n17892 : n32;
  assign n17894 = pi19 ? n17893 : n32;
  assign n17895 = pi18 ? n17479 : n17894;
  assign n17896 = pi17 ? n17477 : n17895;
  assign n17897 = pi16 ? n17474 : n17896;
  assign n17898 = pi21 ? n12635 : n32;
  assign n17899 = pi20 ? n17898 : n32;
  assign n17900 = pi19 ? n17899 : n32;
  assign n17901 = pi18 ? n17487 : n17900;
  assign n17902 = pi17 ? n17485 : n17901;
  assign n17903 = pi16 ? n439 : n17902;
  assign n17904 = pi15 ? n17897 : n17903;
  assign n17905 = pi21 ? n12659 : n32;
  assign n17906 = pi20 ? n17905 : n32;
  assign n17907 = pi19 ? n17906 : n32;
  assign n17908 = pi18 ? n17496 : n17907;
  assign n17909 = pi17 ? n17494 : n17908;
  assign n17910 = pi16 ? n439 : n17909;
  assign n17911 = pi18 ? n335 : n17907;
  assign n17912 = pi17 ? n17508 : n17911;
  assign n17913 = pi16 ? n17504 : n17912;
  assign n17914 = pi15 ? n17910 : n17913;
  assign n17915 = pi14 ? n17904 : n17914;
  assign n17916 = pi16 ? n10118 : n17537;
  assign n17917 = pi15 ? n17527 : n17916;
  assign n17918 = pi18 ? n17544 : n8919;
  assign n17919 = pi17 ? n17541 : n17918;
  assign n17920 = pi16 ? n10118 : n17919;
  assign n17921 = pi16 ? n12658 : n17555;
  assign n17922 = pi15 ? n17920 : n17921;
  assign n17923 = pi14 ? n17917 : n17922;
  assign n17924 = pi13 ? n17915 : n17923;
  assign n17925 = pi12 ? n17891 : n17924;
  assign n17926 = pi11 ? n17863 : n17925;
  assign n17927 = pi10 ? n17792 : n17926;
  assign n17928 = pi09 ? n16985 : n17927;
  assign n17929 = pi08 ? n17563 : n17928;
  assign n17930 = pi20 ? n37 : n4520;
  assign n17931 = pi19 ? n17930 : n32;
  assign n17932 = pi18 ? n37 : n17931;
  assign n17933 = pi17 ? n37 : n17932;
  assign n17934 = pi16 ? n11885 : n17933;
  assign n17935 = pi15 ? n32 : n17934;
  assign n17936 = pi16 ? n12689 : n17933;
  assign n17937 = pi15 ? n17934 : n17936;
  assign n17938 = pi14 ? n17935 : n17937;
  assign n17939 = pi13 ? n32 : n17938;
  assign n17940 = pi12 ? n32 : n17939;
  assign n17941 = pi11 ? n32 : n17940;
  assign n17942 = pi10 ? n32 : n17941;
  assign n17943 = pi20 ? n99 : n4560;
  assign n17944 = pi19 ? n17943 : n32;
  assign n17945 = pi18 ? n37 : n17944;
  assign n17946 = pi17 ? n37 : n17945;
  assign n17947 = pi16 ? n13561 : n17946;
  assign n17948 = pi21 ? n10453 : n32;
  assign n17949 = pi20 ? n99 : n17948;
  assign n17950 = pi19 ? n17949 : n32;
  assign n17951 = pi18 ? n37 : n17950;
  assign n17952 = pi17 ? n37 : n17951;
  assign n17953 = pi16 ? n14445 : n17952;
  assign n17954 = pi15 ? n17947 : n17953;
  assign n17955 = pi22 ? n39 : n112;
  assign n17956 = pi21 ? n17955 : n2175;
  assign n17957 = pi20 ? n32 : n17956;
  assign n17958 = pi19 ? n32 : n17957;
  assign n17959 = pi20 ? n2958 : n2973;
  assign n17960 = pi21 ? n2175 : n181;
  assign n17961 = pi20 ? n15960 : n17960;
  assign n17962 = pi19 ? n17959 : n17961;
  assign n17963 = pi18 ? n17958 : n17962;
  assign n17964 = pi17 ? n32 : n17963;
  assign n17965 = pi20 ? n2982 : n11415;
  assign n17966 = pi21 ? n99 : n2175;
  assign n17967 = pi20 ? n17966 : n2747;
  assign n17968 = pi19 ? n17965 : n17967;
  assign n17969 = pi20 ? n5405 : n2185;
  assign n17970 = pi19 ? n17969 : n2178;
  assign n17971 = pi18 ? n17968 : n17970;
  assign n17972 = pi20 ? n220 : n99;
  assign n17973 = pi20 ? n3042 : n14844;
  assign n17974 = pi19 ? n17972 : n17973;
  assign n17975 = pi21 ? n11393 : n32;
  assign n17976 = pi20 ? n226 : n17975;
  assign n17977 = pi19 ? n17976 : n32;
  assign n17978 = pi18 ? n17974 : n17977;
  assign n17979 = pi17 ? n17971 : n17978;
  assign n17980 = pi16 ? n17964 : n17979;
  assign n17981 = pi20 ? n2974 : n3814;
  assign n17982 = pi19 ? n37 : n17981;
  assign n17983 = pi18 ? n17008 : n17982;
  assign n17984 = pi17 ? n32 : n17983;
  assign n17985 = pi20 ? n17960 : n2967;
  assign n17986 = pi19 ? n5502 : n17985;
  assign n17987 = pi20 ? n3824 : n37;
  assign n17988 = pi20 ? n5496 : n2967;
  assign n17989 = pi19 ? n17987 : n17988;
  assign n17990 = pi18 ? n17986 : n17989;
  assign n17991 = pi20 ? n3824 : n2961;
  assign n17992 = pi20 ? n2163 : n5509;
  assign n17993 = pi19 ? n17991 : n17992;
  assign n17994 = pi22 ? n13918 : n32;
  assign n17995 = pi21 ? n17994 : n32;
  assign n17996 = pi20 ? n2749 : n17995;
  assign n17997 = pi19 ? n17996 : n32;
  assign n17998 = pi18 ? n17993 : n17997;
  assign n17999 = pi17 ? n17990 : n17998;
  assign n18000 = pi16 ? n17984 : n17999;
  assign n18001 = pi15 ? n17980 : n18000;
  assign n18002 = pi14 ? n17954 : n18001;
  assign n18003 = pi20 ? n37 : n17995;
  assign n18004 = pi19 ? n18003 : n32;
  assign n18005 = pi18 ? n37 : n18004;
  assign n18006 = pi17 ? n37 : n18005;
  assign n18007 = pi16 ? n439 : n18006;
  assign n18008 = pi22 ? n6027 : n32;
  assign n18009 = pi21 ? n18008 : n32;
  assign n18010 = pi20 ? n37 : n18009;
  assign n18011 = pi19 ? n18010 : n32;
  assign n18012 = pi18 ? n37 : n18011;
  assign n18013 = pi17 ? n37 : n18012;
  assign n18014 = pi16 ? n439 : n18013;
  assign n18015 = pi15 ? n18007 : n18014;
  assign n18016 = pi22 ? n13969 : n32;
  assign n18017 = pi21 ? n18016 : n32;
  assign n18018 = pi20 ? n7745 : n18017;
  assign n18019 = pi19 ? n18018 : n32;
  assign n18020 = pi18 ? n37 : n18019;
  assign n18021 = pi17 ? n37 : n18020;
  assign n18022 = pi16 ? n439 : n18021;
  assign n18023 = pi22 ? n6774 : n32;
  assign n18024 = pi21 ? n18023 : n32;
  assign n18025 = pi20 ? n7745 : n18024;
  assign n18026 = pi19 ? n18025 : n32;
  assign n18027 = pi18 ? n37 : n18026;
  assign n18028 = pi17 ? n37 : n18027;
  assign n18029 = pi16 ? n439 : n18028;
  assign n18030 = pi15 ? n18022 : n18029;
  assign n18031 = pi14 ? n18015 : n18030;
  assign n18032 = pi13 ? n18002 : n18031;
  assign n18033 = pi18 ? n99 : n16987;
  assign n18034 = pi17 ? n99 : n18033;
  assign n18035 = pi16 ? n201 : n18034;
  assign n18036 = pi16 ? n744 : n18034;
  assign n18037 = pi15 ? n18035 : n18036;
  assign n18038 = pi23 ? n139 : n260;
  assign n18039 = pi22 ? n18038 : n32;
  assign n18040 = pi21 ? n18039 : n32;
  assign n18041 = pi20 ? n139 : n18040;
  assign n18042 = pi19 ? n18041 : n32;
  assign n18043 = pi18 ? n139 : n18042;
  assign n18044 = pi17 ? n139 : n18043;
  assign n18045 = pi16 ? n17063 : n18044;
  assign n18046 = pi15 ? n18036 : n18045;
  assign n18047 = pi14 ? n18037 : n18046;
  assign n18048 = pi20 ? n37 : n3077;
  assign n18049 = pi19 ? n18048 : n139;
  assign n18050 = pi18 ? n18049 : n139;
  assign n18051 = pi22 ? n2026 : n32;
  assign n18052 = pi21 ? n18051 : n32;
  assign n18053 = pi20 ? n139 : n18052;
  assign n18054 = pi19 ? n18053 : n32;
  assign n18055 = pi18 ? n139 : n18054;
  assign n18056 = pi17 ? n18050 : n18055;
  assign n18057 = pi16 ? n439 : n18056;
  assign n18058 = pi20 ? n37 : n16058;
  assign n18059 = pi19 ? n37 : n18058;
  assign n18060 = pi20 ? n8729 : n139;
  assign n18061 = pi19 ? n18060 : n139;
  assign n18062 = pi18 ? n18059 : n18061;
  assign n18063 = pi21 ? n11083 : n32;
  assign n18064 = pi20 ? n139 : n18063;
  assign n18065 = pi19 ? n18064 : n32;
  assign n18066 = pi18 ? n139 : n18065;
  assign n18067 = pi17 ? n18062 : n18066;
  assign n18068 = pi16 ? n439 : n18067;
  assign n18069 = pi15 ? n18057 : n18068;
  assign n18070 = pi20 ? n3104 : n37;
  assign n18071 = pi19 ? n18070 : n139;
  assign n18072 = pi18 ? n37 : n18071;
  assign n18073 = pi17 ? n18072 : n18066;
  assign n18074 = pi16 ? n439 : n18073;
  assign n18075 = pi18 ? n37 : n9766;
  assign n18076 = pi17 ? n18075 : n18066;
  assign n18077 = pi16 ? n439 : n18076;
  assign n18078 = pi15 ? n18074 : n18077;
  assign n18079 = pi14 ? n18069 : n18078;
  assign n18080 = pi13 ? n18047 : n18079;
  assign n18081 = pi12 ? n18032 : n18080;
  assign n18082 = pi20 ? n37 : n997;
  assign n18083 = pi19 ? n37 : n18082;
  assign n18084 = pi18 ? n37 : n18083;
  assign n18085 = pi18 ? n10030 : n18065;
  assign n18086 = pi17 ? n18084 : n18085;
  assign n18087 = pi16 ? n439 : n18086;
  assign n18088 = pi20 ? n139 : n3176;
  assign n18089 = pi19 ? n18088 : n32;
  assign n18090 = pi18 ? n139 : n18089;
  assign n18091 = pi17 ? n37 : n18090;
  assign n18092 = pi16 ? n439 : n18091;
  assign n18093 = pi15 ? n18087 : n18092;
  assign n18094 = pi20 ? n939 : n3176;
  assign n18095 = pi19 ? n18094 : n32;
  assign n18096 = pi18 ? n9770 : n18095;
  assign n18097 = pi17 ? n37 : n18096;
  assign n18098 = pi16 ? n439 : n18097;
  assign n18099 = pi20 ? n1056 : n204;
  assign n18100 = pi19 ? n18099 : n204;
  assign n18101 = pi20 ? n204 : n3176;
  assign n18102 = pi19 ? n18101 : n32;
  assign n18103 = pi18 ? n18100 : n18102;
  assign n18104 = pi17 ? n37 : n18103;
  assign n18105 = pi16 ? n439 : n18104;
  assign n18106 = pi15 ? n18098 : n18105;
  assign n18107 = pi14 ? n18093 : n18106;
  assign n18108 = pi20 ? n37 : n204;
  assign n18109 = pi19 ? n18108 : n204;
  assign n18110 = pi18 ? n18109 : n18102;
  assign n18111 = pi17 ? n37 : n18110;
  assign n18112 = pi16 ? n439 : n18111;
  assign n18113 = pi19 ? n8928 : n233;
  assign n18114 = pi20 ? n233 : n4110;
  assign n18115 = pi19 ? n18114 : n32;
  assign n18116 = pi18 ? n18113 : n18115;
  assign n18117 = pi17 ? n37 : n18116;
  assign n18118 = pi16 ? n439 : n18117;
  assign n18119 = pi15 ? n18112 : n18118;
  assign n18120 = pi19 ? n7685 : n15469;
  assign n18121 = pi21 ? n335 : n6361;
  assign n18122 = pi20 ? n18121 : n4110;
  assign n18123 = pi19 ? n18122 : n32;
  assign n18124 = pi18 ? n18120 : n18123;
  assign n18125 = pi17 ? n37 : n18124;
  assign n18126 = pi16 ? n439 : n18125;
  assign n18127 = pi19 ? n6373 : n15470;
  assign n18128 = pi20 ? n335 : n4110;
  assign n18129 = pi19 ? n18128 : n32;
  assign n18130 = pi18 ? n18127 : n18129;
  assign n18131 = pi17 ? n37 : n18130;
  assign n18132 = pi16 ? n439 : n18131;
  assign n18133 = pi15 ? n18126 : n18132;
  assign n18134 = pi14 ? n18119 : n18133;
  assign n18135 = pi13 ? n18107 : n18134;
  assign n18136 = pi20 ? n13527 : n4110;
  assign n18137 = pi19 ? n18136 : n32;
  assign n18138 = pi18 ? n9856 : n18137;
  assign n18139 = pi17 ? n37 : n18138;
  assign n18140 = pi16 ? n439 : n18139;
  assign n18141 = pi20 ? n37 : n2004;
  assign n18142 = pi19 ? n37 : n18141;
  assign n18143 = pi20 ? n569 : n6417;
  assign n18144 = pi19 ? n18143 : n32;
  assign n18145 = pi18 ? n18142 : n18144;
  assign n18146 = pi17 ? n37 : n18145;
  assign n18147 = pi16 ? n439 : n18146;
  assign n18148 = pi15 ? n18140 : n18147;
  assign n18149 = pi18 ? n17216 : n18144;
  assign n18150 = pi17 ? n37 : n18149;
  assign n18151 = pi16 ? n439 : n18150;
  assign n18152 = pi20 ? n649 : n5830;
  assign n18153 = pi19 ? n18152 : n32;
  assign n18154 = pi18 ? n7677 : n18153;
  assign n18155 = pi17 ? n37 : n18154;
  assign n18156 = pi16 ? n439 : n18155;
  assign n18157 = pi15 ? n18151 : n18156;
  assign n18158 = pi14 ? n18148 : n18157;
  assign n18159 = pi21 ? n2091 : n3392;
  assign n18160 = pi20 ? n37 : n18159;
  assign n18161 = pi19 ? n37 : n18160;
  assign n18162 = pi21 ? n1920 : n3409;
  assign n18163 = pi20 ? n18162 : n10011;
  assign n18164 = pi19 ? n18163 : n32;
  assign n18165 = pi18 ? n18161 : n18164;
  assign n18166 = pi17 ? n37 : n18165;
  assign n18167 = pi16 ? n439 : n18166;
  assign n18168 = pi20 ? n18162 : n1822;
  assign n18169 = pi19 ? n18168 : n32;
  assign n18170 = pi18 ? n37 : n18169;
  assign n18171 = pi17 ? n37 : n18170;
  assign n18172 = pi16 ? n439 : n18171;
  assign n18173 = pi15 ? n18167 : n18172;
  assign n18174 = pi21 ? n233 : n2091;
  assign n18175 = pi20 ? n37 : n18174;
  assign n18176 = pi19 ? n37 : n18175;
  assign n18177 = pi20 ? n2091 : n2701;
  assign n18178 = pi19 ? n18177 : n32;
  assign n18179 = pi18 ? n18176 : n18178;
  assign n18180 = pi17 ? n37 : n18179;
  assign n18181 = pi16 ? n439 : n18180;
  assign n18182 = pi20 ? n2107 : n1822;
  assign n18183 = pi19 ? n18182 : n32;
  assign n18184 = pi18 ? n2109 : n18183;
  assign n18185 = pi17 ? n37 : n18184;
  assign n18186 = pi16 ? n439 : n18185;
  assign n18187 = pi15 ? n18181 : n18186;
  assign n18188 = pi14 ? n18173 : n18187;
  assign n18189 = pi13 ? n18158 : n18188;
  assign n18190 = pi12 ? n18135 : n18189;
  assign n18191 = pi11 ? n18081 : n18190;
  assign n18192 = pi20 ? n37 : n2106;
  assign n18193 = pi19 ? n37 : n18192;
  assign n18194 = pi21 ? n685 : n2721;
  assign n18195 = pi20 ? n18194 : n1822;
  assign n18196 = pi19 ? n18195 : n32;
  assign n18197 = pi18 ? n18193 : n18196;
  assign n18198 = pi17 ? n37 : n18197;
  assign n18199 = pi16 ? n439 : n18198;
  assign n18200 = pi20 ? n2106 : n32;
  assign n18201 = pi19 ? n18200 : n32;
  assign n18202 = pi18 ? n2109 : n18201;
  assign n18203 = pi17 ? n37 : n18202;
  assign n18204 = pi16 ? n439 : n18203;
  assign n18205 = pi15 ? n18199 : n18204;
  assign n18206 = pi21 ? n2106 : n2721;
  assign n18207 = pi20 ? n18206 : n32;
  assign n18208 = pi19 ? n18207 : n32;
  assign n18209 = pi18 ? n37 : n18208;
  assign n18210 = pi17 ? n37 : n18209;
  assign n18211 = pi16 ? n439 : n18210;
  assign n18212 = pi21 ? n37 : n11208;
  assign n18213 = pi20 ? n18212 : n32;
  assign n18214 = pi19 ? n18213 : n32;
  assign n18215 = pi18 ? n37 : n18214;
  assign n18216 = pi17 ? n37 : n18215;
  assign n18217 = pi16 ? n439 : n18216;
  assign n18218 = pi15 ? n18211 : n18217;
  assign n18219 = pi14 ? n18205 : n18218;
  assign n18220 = pi22 ? n893 : n685;
  assign n18221 = pi21 ? n37 : n18220;
  assign n18222 = pi20 ? n18221 : n32;
  assign n18223 = pi19 ? n18222 : n32;
  assign n18224 = pi18 ? n37 : n18223;
  assign n18225 = pi17 ? n37 : n18224;
  assign n18226 = pi16 ? n439 : n18225;
  assign n18227 = pi15 ? n18217 : n18226;
  assign n18228 = pi20 ? n5085 : n32;
  assign n18229 = pi19 ? n18228 : n32;
  assign n18230 = pi18 ? n99 : n18229;
  assign n18231 = pi17 ? n99 : n18230;
  assign n18232 = pi16 ? n721 : n18231;
  assign n18233 = pi21 ? n685 : n3445;
  assign n18234 = pi20 ? n18233 : n32;
  assign n18235 = pi19 ? n18234 : n32;
  assign n18236 = pi18 ? n5087 : n18235;
  assign n18237 = pi17 ? n99 : n18236;
  assign n18238 = pi16 ? n721 : n18237;
  assign n18239 = pi15 ? n18232 : n18238;
  assign n18240 = pi14 ? n18227 : n18239;
  assign n18241 = pi13 ? n18219 : n18240;
  assign n18242 = pi19 ? n99 : n11445;
  assign n18243 = pi18 ? n99 : n18242;
  assign n18244 = pi20 ? n15263 : n6090;
  assign n18245 = pi19 ? n16307 : n18244;
  assign n18246 = pi21 ? n6089 : n2147;
  assign n18247 = pi20 ? n18246 : n32;
  assign n18248 = pi19 ? n18247 : n32;
  assign n18249 = pi18 ? n18245 : n18248;
  assign n18250 = pi17 ? n18243 : n18249;
  assign n18251 = pi16 ? n721 : n18250;
  assign n18252 = pi21 ? n7815 : n99;
  assign n18253 = pi20 ? n99 : n18252;
  assign n18254 = pi19 ? n18253 : n99;
  assign n18255 = pi18 ? n18254 : n17340;
  assign n18256 = pi23 ? n2766 : n395;
  assign n18257 = pi22 ? n3443 : n18256;
  assign n18258 = pi21 ? n767 : n18257;
  assign n18259 = pi20 ? n18258 : n32;
  assign n18260 = pi19 ? n18259 : n32;
  assign n18261 = pi18 ? n17355 : n18260;
  assign n18262 = pi17 ? n18255 : n18261;
  assign n18263 = pi16 ? n721 : n18262;
  assign n18264 = pi15 ? n18251 : n18263;
  assign n18265 = pi21 ? n5899 : n157;
  assign n18266 = pi20 ? n7818 : n18265;
  assign n18267 = pi19 ? n157 : n18266;
  assign n18268 = pi18 ? n18267 : n157;
  assign n18269 = pi19 ? n157 : n16276;
  assign n18270 = pi21 ? n99 : n6535;
  assign n18271 = pi20 ? n18270 : n32;
  assign n18272 = pi19 ? n18271 : n32;
  assign n18273 = pi18 ? n18269 : n18272;
  assign n18274 = pi17 ? n18268 : n18273;
  assign n18275 = pi16 ? n9291 : n18274;
  assign n18276 = pi22 ? n1484 : n99;
  assign n18277 = pi21 ? n775 : n18276;
  assign n18278 = pi20 ? n157 : n18277;
  assign n18279 = pi19 ? n157 : n18278;
  assign n18280 = pi18 ? n18279 : n16320;
  assign n18281 = pi17 ? n157 : n18280;
  assign n18282 = pi16 ? n5910 : n18281;
  assign n18283 = pi15 ? n18275 : n18282;
  assign n18284 = pi14 ? n18264 : n18283;
  assign n18285 = pi21 ? n157 : n3523;
  assign n18286 = pi20 ? n18285 : n32;
  assign n18287 = pi19 ? n18286 : n32;
  assign n18288 = pi18 ? n17368 : n18287;
  assign n18289 = pi17 ? n157 : n18288;
  assign n18290 = pi16 ? n5910 : n18289;
  assign n18291 = pi21 ? n777 : n17375;
  assign n18292 = pi20 ? n157 : n18291;
  assign n18293 = pi19 ? n157 : n18292;
  assign n18294 = pi18 ? n18293 : n11500;
  assign n18295 = pi17 ? n157 : n18294;
  assign n18296 = pi16 ? n9291 : n18295;
  assign n18297 = pi15 ? n18290 : n18296;
  assign n18298 = pi21 ? n5168 : n204;
  assign n18299 = pi20 ? n32 : n18298;
  assign n18300 = pi19 ? n32 : n18299;
  assign n18301 = pi18 ? n18300 : n204;
  assign n18302 = pi17 ? n32 : n18301;
  assign n18303 = pi20 ? n17394 : n17390;
  assign n18304 = pi19 ? n204 : n18303;
  assign n18305 = pi18 ? n17389 : n18304;
  assign n18306 = pi20 ? n204 : n17366;
  assign n18307 = pi19 ? n17396 : n18306;
  assign n18308 = pi18 ? n18307 : n11500;
  assign n18309 = pi17 ? n18305 : n18308;
  assign n18310 = pi16 ? n18302 : n18309;
  assign n18311 = pi21 ? n139 : n3668;
  assign n18312 = pi20 ? n18311 : n204;
  assign n18313 = pi19 ? n204 : n18312;
  assign n18314 = pi20 ? n2318 : n316;
  assign n18315 = pi19 ? n204 : n18314;
  assign n18316 = pi18 ? n18313 : n18315;
  assign n18317 = pi21 ? n356 : n204;
  assign n18318 = pi20 ? n7909 : n18317;
  assign n18319 = pi19 ? n18318 : n17409;
  assign n18320 = pi18 ? n18319 : n11500;
  assign n18321 = pi17 ? n18316 : n18320;
  assign n18322 = pi16 ? n13833 : n18321;
  assign n18323 = pi15 ? n18310 : n18322;
  assign n18324 = pi14 ? n18297 : n18323;
  assign n18325 = pi13 ? n18284 : n18324;
  assign n18326 = pi12 ? n18241 : n18325;
  assign n18327 = pi20 ? n347 : n316;
  assign n18328 = pi19 ? n139 : n18327;
  assign n18329 = pi18 ? n139 : n18328;
  assign n18330 = pi20 ? n316 : n9773;
  assign n18331 = pi20 ? n1022 : n975;
  assign n18332 = pi19 ? n18330 : n18331;
  assign n18333 = pi18 ? n18332 : n11500;
  assign n18334 = pi17 ? n18329 : n18333;
  assign n18335 = pi16 ? n915 : n18334;
  assign n18336 = pi21 ? n2319 : n139;
  assign n18337 = pi20 ? n139 : n18336;
  assign n18338 = pi19 ? n18337 : n139;
  assign n18339 = pi18 ? n18338 : n17418;
  assign n18340 = pi18 ? n17429 : n11500;
  assign n18341 = pi17 ? n18339 : n18340;
  assign n18342 = pi16 ? n915 : n18341;
  assign n18343 = pi15 ? n18335 : n18342;
  assign n18344 = pi20 ? n7900 : n3702;
  assign n18345 = pi19 ? n316 : n18344;
  assign n18346 = pi18 ? n18345 : n316;
  assign n18347 = pi17 ? n18346 : n17430;
  assign n18348 = pi16 ? n6235 : n18347;
  assign n18349 = pi21 ? n1549 : n316;
  assign n18350 = pi20 ? n32 : n18349;
  assign n18351 = pi19 ? n32 : n18350;
  assign n18352 = pi18 ? n18351 : n316;
  assign n18353 = pi17 ? n32 : n18352;
  assign n18354 = pi20 ? n5286 : n4778;
  assign n18355 = pi19 ? n316 : n18354;
  assign n18356 = pi18 ? n18355 : n316;
  assign n18357 = pi17 ? n18356 : n10597;
  assign n18358 = pi16 ? n18353 : n18357;
  assign n18359 = pi15 ? n18348 : n18358;
  assign n18360 = pi14 ? n18343 : n18359;
  assign n18361 = pi20 ? n139 : n927;
  assign n18362 = pi19 ? n139 : n18361;
  assign n18363 = pi21 ? n916 : n5829;
  assign n18364 = pi20 ? n18363 : n32;
  assign n18365 = pi19 ? n18364 : n32;
  assign n18366 = pi18 ? n18362 : n18365;
  assign n18367 = pi17 ? n139 : n18366;
  assign n18368 = pi16 ? n1773 : n18367;
  assign n18369 = pi15 ? n18358 : n18368;
  assign n18370 = pi20 ? n954 : n32;
  assign n18371 = pi19 ? n18370 : n32;
  assign n18372 = pi18 ? n139 : n18371;
  assign n18373 = pi17 ? n139 : n18372;
  assign n18374 = pi16 ? n915 : n18373;
  assign n18375 = pi20 ? n6003 : n32;
  assign n18376 = pi19 ? n18375 : n32;
  assign n18377 = pi18 ? n204 : n18376;
  assign n18378 = pi17 ? n204 : n18377;
  assign n18379 = pi16 ? n11804 : n18378;
  assign n18380 = pi15 ? n18374 : n18379;
  assign n18381 = pi14 ? n18369 : n18380;
  assign n18382 = pi13 ? n18360 : n18381;
  assign n18383 = pi20 ? n603 : n647;
  assign n18384 = pi19 ? n18383 : n37;
  assign n18385 = pi18 ? n18384 : n17476;
  assign n18386 = pi21 ? n204 : n1009;
  assign n18387 = pi20 ? n18386 : n32;
  assign n18388 = pi19 ? n18387 : n32;
  assign n18389 = pi18 ? n17479 : n18388;
  assign n18390 = pi17 ? n18385 : n18389;
  assign n18391 = pi16 ? n439 : n18390;
  assign n18392 = pi21 ? n233 : n32;
  assign n18393 = pi20 ? n18392 : n32;
  assign n18394 = pi19 ? n18393 : n32;
  assign n18395 = pi18 ? n17487 : n18394;
  assign n18396 = pi17 ? n17485 : n18395;
  assign n18397 = pi16 ? n439 : n18396;
  assign n18398 = pi15 ? n18391 : n18397;
  assign n18399 = pi20 ? n577 : n7980;
  assign n18400 = pi19 ? n37 : n18399;
  assign n18401 = pi18 ? n37 : n18400;
  assign n18402 = pi19 ? n14394 : n17495;
  assign n18403 = pi18 ? n18402 : n18394;
  assign n18404 = pi17 ? n18401 : n18403;
  assign n18405 = pi16 ? n439 : n18404;
  assign n18406 = pi18 ? n374 : n17502;
  assign n18407 = pi17 ? n32 : n18406;
  assign n18408 = pi20 ? n642 : n335;
  assign n18409 = pi19 ? n335 : n18408;
  assign n18410 = pi18 ? n18409 : n335;
  assign n18411 = pi22 ? n233 : n685;
  assign n18412 = pi21 ? n18411 : n32;
  assign n18413 = pi20 ? n18412 : n32;
  assign n18414 = pi19 ? n18413 : n32;
  assign n18415 = pi18 ? n335 : n18414;
  assign n18416 = pi17 ? n18410 : n18415;
  assign n18417 = pi16 ? n18407 : n18416;
  assign n18418 = pi15 ? n18405 : n18417;
  assign n18419 = pi14 ? n18398 : n18418;
  assign n18420 = pi18 ? n374 : n7677;
  assign n18421 = pi17 ? n32 : n18420;
  assign n18422 = pi19 ? n335 : n17204;
  assign n18423 = pi18 ? n18422 : n17487;
  assign n18424 = pi22 ? n673 : n1070;
  assign n18425 = pi21 ? n18424 : n32;
  assign n18426 = pi20 ? n18425 : n32;
  assign n18427 = pi19 ? n18426 : n32;
  assign n18428 = pi18 ? n17487 : n18427;
  assign n18429 = pi17 ? n18423 : n18428;
  assign n18430 = pi16 ? n18421 : n18429;
  assign n18431 = pi21 ? n233 : n6376;
  assign n18432 = pi20 ? n335 : n18431;
  assign n18433 = pi19 ? n335 : n18432;
  assign n18434 = pi18 ? n335 : n18433;
  assign n18435 = pi20 ? n335 : n15469;
  assign n18436 = pi19 ? n18435 : n17486;
  assign n18437 = pi22 ? n673 : n6415;
  assign n18438 = pi21 ? n18437 : n32;
  assign n18439 = pi20 ? n18438 : n32;
  assign n18440 = pi19 ? n18439 : n32;
  assign n18441 = pi18 ? n18436 : n18440;
  assign n18442 = pi17 ? n18434 : n18441;
  assign n18443 = pi16 ? n10118 : n18442;
  assign n18444 = pi15 ? n18430 : n18443;
  assign n18445 = pi18 ? n335 : n15438;
  assign n18446 = pi20 ? n233 : n15469;
  assign n18447 = pi19 ? n18446 : n17543;
  assign n18448 = pi23 ? n157 : n204;
  assign n18449 = pi22 ? n18448 : n3338;
  assign n18450 = pi21 ? n18449 : n32;
  assign n18451 = pi20 ? n18450 : n32;
  assign n18452 = pi19 ? n18451 : n32;
  assign n18453 = pi18 ? n18447 : n18452;
  assign n18454 = pi17 ? n18445 : n18453;
  assign n18455 = pi16 ? n17532 : n18454;
  assign n18456 = pi23 ? n1590 : n139;
  assign n18457 = pi22 ? n18456 : n9827;
  assign n18458 = pi21 ? n18457 : n363;
  assign n18459 = pi20 ? n32 : n18458;
  assign n18460 = pi19 ? n32 : n18459;
  assign n18461 = pi23 ? n363 : n335;
  assign n18462 = pi22 ? n335 : n18461;
  assign n18463 = pi21 ? n18462 : n17548;
  assign n18464 = pi21 ? n7986 : n17548;
  assign n18465 = pi20 ? n18463 : n18464;
  assign n18466 = pi21 ? n18462 : n9143;
  assign n18467 = pi22 ? n363 : n18461;
  assign n18468 = pi21 ? n18467 : n17548;
  assign n18469 = pi20 ? n18466 : n18468;
  assign n18470 = pi19 ? n18465 : n18469;
  assign n18471 = pi18 ? n18460 : n18470;
  assign n18472 = pi17 ? n32 : n18471;
  assign n18473 = pi22 ? n18461 : n9827;
  assign n18474 = pi21 ? n18473 : n233;
  assign n18475 = pi21 ? n233 : n7986;
  assign n18476 = pi20 ? n18474 : n18475;
  assign n18477 = pi21 ? n17548 : n9836;
  assign n18478 = pi21 ? n363 : n18473;
  assign n18479 = pi20 ? n18477 : n18478;
  assign n18480 = pi19 ? n18476 : n18479;
  assign n18481 = pi21 ? n4902 : n233;
  assign n18482 = pi20 ? n13527 : n18481;
  assign n18483 = pi19 ? n18482 : n233;
  assign n18484 = pi18 ? n18480 : n18483;
  assign n18485 = pi18 ? n233 : n16946;
  assign n18486 = pi17 ? n18484 : n18485;
  assign n18487 = pi16 ? n18472 : n18486;
  assign n18488 = pi15 ? n18455 : n18487;
  assign n18489 = pi14 ? n18444 : n18488;
  assign n18490 = pi13 ? n18419 : n18489;
  assign n18491 = pi12 ? n18382 : n18490;
  assign n18492 = pi11 ? n18326 : n18491;
  assign n18493 = pi10 ? n18191 : n18492;
  assign n18494 = pi09 ? n17942 : n18493;
  assign n18495 = pi21 ? n17955 : n2160;
  assign n18496 = pi20 ? n32 : n18495;
  assign n18497 = pi19 ? n32 : n18496;
  assign n18498 = pi20 ? n3814 : n3817;
  assign n18499 = pi21 ? n2168 : n218;
  assign n18500 = pi21 ? n2160 : n1143;
  assign n18501 = pi20 ? n18499 : n18500;
  assign n18502 = pi19 ? n18498 : n18501;
  assign n18503 = pi18 ? n18497 : n18502;
  assign n18504 = pi17 ? n32 : n18503;
  assign n18505 = pi20 ? n5496 : n11418;
  assign n18506 = pi21 ? n99 : n2160;
  assign n18507 = pi20 ? n18506 : n5420;
  assign n18508 = pi19 ? n18505 : n18507;
  assign n18509 = pi20 ? n99 : n2755;
  assign n18510 = pi19 ? n18509 : n220;
  assign n18511 = pi18 ? n18508 : n18510;
  assign n18512 = pi20 ? n2749 : n99;
  assign n18513 = pi20 ? n2189 : n3825;
  assign n18514 = pi19 ? n18512 : n18513;
  assign n18515 = pi18 ? n18514 : n17977;
  assign n18516 = pi17 ? n18511 : n18515;
  assign n18517 = pi16 ? n18504 : n18516;
  assign n18518 = pi20 ? n2974 : n2970;
  assign n18519 = pi19 ? n37 : n18518;
  assign n18520 = pi18 ? n17008 : n18519;
  assign n18521 = pi17 ? n32 : n18520;
  assign n18522 = pi20 ? n14518 : n14510;
  assign n18523 = pi20 ? n5077 : n2983;
  assign n18524 = pi19 ? n18522 : n18523;
  assign n18525 = pi20 ? n5496 : n37;
  assign n18526 = pi19 ? n18525 : n2984;
  assign n18527 = pi18 ? n18524 : n18526;
  assign n18528 = pi20 ? n2961 : n14518;
  assign n18529 = pi19 ? n17991 : n18528;
  assign n18530 = pi20 ? n17966 : n17995;
  assign n18531 = pi19 ? n18530 : n32;
  assign n18532 = pi18 ? n18529 : n18531;
  assign n18533 = pi17 ? n18527 : n18532;
  assign n18534 = pi16 ? n18521 : n18533;
  assign n18535 = pi15 ? n18517 : n18534;
  assign n18536 = pi14 ? n17954 : n18535;
  assign n18537 = pi16 ? n439 : n16975;
  assign n18538 = pi15 ? n18007 : n18537;
  assign n18539 = pi22 ? n112 : n32;
  assign n18540 = pi21 ? n18539 : n32;
  assign n18541 = pi20 ? n7745 : n18540;
  assign n18542 = pi19 ? n18541 : n32;
  assign n18543 = pi18 ? n37 : n18542;
  assign n18544 = pi17 ? n37 : n18543;
  assign n18545 = pi16 ? n439 : n18544;
  assign n18546 = pi14 ? n18538 : n18545;
  assign n18547 = pi13 ? n18536 : n18546;
  assign n18548 = pi22 ? n1504 : n37;
  assign n18549 = pi21 ? n18548 : n99;
  assign n18550 = pi20 ? n32 : n18549;
  assign n18551 = pi19 ? n32 : n18550;
  assign n18552 = pi18 ? n18551 : n99;
  assign n18553 = pi17 ? n32 : n18552;
  assign n18554 = pi18 ? n99 : n17944;
  assign n18555 = pi17 ? n99 : n18554;
  assign n18556 = pi16 ? n18553 : n18555;
  assign n18557 = pi16 ? n721 : n18555;
  assign n18558 = pi15 ? n18556 : n18557;
  assign n18559 = pi16 ? n744 : n18555;
  assign n18560 = pi18 ? n374 : n17102;
  assign n18561 = pi17 ? n32 : n18560;
  assign n18562 = pi20 ? n139 : n17948;
  assign n18563 = pi19 ? n18562 : n32;
  assign n18564 = pi18 ? n139 : n18563;
  assign n18565 = pi17 ? n139 : n18564;
  assign n18566 = pi16 ? n18561 : n18565;
  assign n18567 = pi15 ? n18559 : n18566;
  assign n18568 = pi14 ? n18558 : n18567;
  assign n18569 = pi20 ? n376 : n3915;
  assign n18570 = pi19 ? n18569 : n139;
  assign n18571 = pi18 ? n18570 : n139;
  assign n18572 = pi22 ? n9827 : n32;
  assign n18573 = pi21 ? n18572 : n32;
  assign n18574 = pi20 ? n139 : n18573;
  assign n18575 = pi19 ? n18574 : n32;
  assign n18576 = pi18 ? n139 : n18575;
  assign n18577 = pi17 ? n18571 : n18576;
  assign n18578 = pi16 ? n439 : n18577;
  assign n18579 = pi20 ? n8742 : n14988;
  assign n18580 = pi19 ? n37 : n18579;
  assign n18581 = pi21 ? n297 : n295;
  assign n18582 = pi20 ? n18581 : n139;
  assign n18583 = pi19 ? n18582 : n139;
  assign n18584 = pi18 ? n18580 : n18583;
  assign n18585 = pi21 ? n11534 : n32;
  assign n18586 = pi20 ? n139 : n18585;
  assign n18587 = pi19 ? n18586 : n32;
  assign n18588 = pi18 ? n139 : n18587;
  assign n18589 = pi17 ? n18584 : n18588;
  assign n18590 = pi16 ? n439 : n18589;
  assign n18591 = pi15 ? n18578 : n18590;
  assign n18592 = pi17 ? n18072 : n18588;
  assign n18593 = pi16 ? n439 : n18592;
  assign n18594 = pi15 ? n18593 : n18077;
  assign n18595 = pi14 ? n18591 : n18594;
  assign n18596 = pi13 ? n18568 : n18595;
  assign n18597 = pi12 ? n18547 : n18596;
  assign n18598 = pi20 ? n569 : n4110;
  assign n18599 = pi19 ? n18598 : n32;
  assign n18600 = pi18 ? n18142 : n18599;
  assign n18601 = pi17 ? n37 : n18600;
  assign n18602 = pi16 ? n439 : n18601;
  assign n18603 = pi15 ? n18140 : n18602;
  assign n18604 = pi20 ? n649 : n4116;
  assign n18605 = pi19 ? n18604 : n32;
  assign n18606 = pi18 ? n7677 : n18605;
  assign n18607 = pi17 ? n37 : n18606;
  assign n18608 = pi16 ? n439 : n18607;
  assign n18609 = pi15 ? n18151 : n18608;
  assign n18610 = pi14 ? n18603 : n18609;
  assign n18611 = pi22 ? n15697 : n32;
  assign n18612 = pi21 ? n18611 : n32;
  assign n18613 = pi20 ? n18162 : n18612;
  assign n18614 = pi19 ? n18613 : n32;
  assign n18615 = pi18 ? n18161 : n18614;
  assign n18616 = pi17 ? n37 : n18615;
  assign n18617 = pi16 ? n439 : n18616;
  assign n18618 = pi20 ? n18162 : n3398;
  assign n18619 = pi19 ? n18618 : n32;
  assign n18620 = pi18 ? n37 : n18619;
  assign n18621 = pi17 ? n37 : n18620;
  assign n18622 = pi16 ? n439 : n18621;
  assign n18623 = pi15 ? n18617 : n18622;
  assign n18624 = pi20 ? n2091 : n2679;
  assign n18625 = pi19 ? n18624 : n32;
  assign n18626 = pi18 ? n18176 : n18625;
  assign n18627 = pi17 ? n37 : n18626;
  assign n18628 = pi16 ? n439 : n18627;
  assign n18629 = pi20 ? n2107 : n2701;
  assign n18630 = pi19 ? n18629 : n32;
  assign n18631 = pi18 ? n2109 : n18630;
  assign n18632 = pi17 ? n37 : n18631;
  assign n18633 = pi16 ? n439 : n18632;
  assign n18634 = pi15 ? n18628 : n18633;
  assign n18635 = pi14 ? n18623 : n18634;
  assign n18636 = pi13 ? n18610 : n18635;
  assign n18637 = pi12 ? n18135 : n18636;
  assign n18638 = pi11 ? n18597 : n18637;
  assign n18639 = pi20 ? n18194 : n2701;
  assign n18640 = pi19 ? n18639 : n32;
  assign n18641 = pi18 ? n18193 : n18640;
  assign n18642 = pi17 ? n37 : n18641;
  assign n18643 = pi16 ? n439 : n18642;
  assign n18644 = pi20 ? n2106 : n2701;
  assign n18645 = pi19 ? n18644 : n32;
  assign n18646 = pi18 ? n2109 : n18645;
  assign n18647 = pi17 ? n37 : n18646;
  assign n18648 = pi16 ? n439 : n18647;
  assign n18649 = pi15 ? n18643 : n18648;
  assign n18650 = pi20 ? n18206 : n2701;
  assign n18651 = pi19 ? n18650 : n32;
  assign n18652 = pi18 ? n37 : n18651;
  assign n18653 = pi17 ? n37 : n18652;
  assign n18654 = pi16 ? n439 : n18653;
  assign n18655 = pi20 ? n18212 : n2701;
  assign n18656 = pi19 ? n18655 : n32;
  assign n18657 = pi18 ? n37 : n18656;
  assign n18658 = pi17 ? n37 : n18657;
  assign n18659 = pi16 ? n439 : n18658;
  assign n18660 = pi15 ? n18654 : n18659;
  assign n18661 = pi14 ? n18649 : n18660;
  assign n18662 = pi20 ? n18221 : n2701;
  assign n18663 = pi19 ? n18662 : n32;
  assign n18664 = pi18 ? n37 : n18663;
  assign n18665 = pi17 ? n37 : n18664;
  assign n18666 = pi16 ? n439 : n18665;
  assign n18667 = pi15 ? n18659 : n18666;
  assign n18668 = pi20 ? n5085 : n2701;
  assign n18669 = pi19 ? n18668 : n32;
  assign n18670 = pi18 ? n99 : n18669;
  assign n18671 = pi17 ? n99 : n18670;
  assign n18672 = pi16 ? n744 : n18671;
  assign n18673 = pi20 ? n18233 : n1822;
  assign n18674 = pi19 ? n18673 : n32;
  assign n18675 = pi18 ? n5087 : n18674;
  assign n18676 = pi17 ? n99 : n18675;
  assign n18677 = pi16 ? n744 : n18676;
  assign n18678 = pi15 ? n18672 : n18677;
  assign n18679 = pi14 ? n18667 : n18678;
  assign n18680 = pi13 ? n18661 : n18679;
  assign n18681 = pi21 ? n6089 : n5113;
  assign n18682 = pi20 ? n18681 : n32;
  assign n18683 = pi19 ? n18682 : n32;
  assign n18684 = pi18 ? n18245 : n18683;
  assign n18685 = pi17 ? n18243 : n18684;
  assign n18686 = pi16 ? n744 : n18685;
  assign n18687 = pi23 ? n170 : n685;
  assign n18688 = pi22 ? n18687 : n1475;
  assign n18689 = pi21 ? n767 : n18688;
  assign n18690 = pi20 ? n18689 : n32;
  assign n18691 = pi19 ? n18690 : n32;
  assign n18692 = pi18 ? n17355 : n18691;
  assign n18693 = pi17 ? n18255 : n18692;
  assign n18694 = pi16 ? n744 : n18693;
  assign n18695 = pi15 ? n18686 : n18694;
  assign n18696 = pi18 ? n18279 : n16844;
  assign n18697 = pi17 ? n157 : n18696;
  assign n18698 = pi16 ? n5910 : n18697;
  assign n18699 = pi15 ? n18275 : n18698;
  assign n18700 = pi14 ? n18695 : n18699;
  assign n18701 = pi20 ? n5179 : n32;
  assign n18702 = pi19 ? n18701 : n32;
  assign n18703 = pi18 ? n17368 : n18702;
  assign n18704 = pi17 ? n157 : n18703;
  assign n18705 = pi16 ? n7793 : n18704;
  assign n18706 = pi18 ? n18293 : n12349;
  assign n18707 = pi17 ? n157 : n18706;
  assign n18708 = pi16 ? n8620 : n18707;
  assign n18709 = pi15 ? n18705 : n18708;
  assign n18710 = pi21 ? n7788 : n204;
  assign n18711 = pi20 ? n32 : n18710;
  assign n18712 = pi19 ? n32 : n18711;
  assign n18713 = pi18 ? n18712 : n204;
  assign n18714 = pi17 ? n32 : n18713;
  assign n18715 = pi21 ? n316 : n4788;
  assign n18716 = pi20 ? n18715 : n32;
  assign n18717 = pi19 ? n18716 : n32;
  assign n18718 = pi18 ? n18307 : n18717;
  assign n18719 = pi17 ? n18305 : n18718;
  assign n18720 = pi16 ? n18714 : n18719;
  assign n18721 = pi21 ? n316 : n4208;
  assign n18722 = pi20 ? n18721 : n32;
  assign n18723 = pi19 ? n18722 : n32;
  assign n18724 = pi18 ? n18319 : n18723;
  assign n18725 = pi17 ? n18316 : n18724;
  assign n18726 = pi16 ? n13833 : n18725;
  assign n18727 = pi15 ? n18720 : n18726;
  assign n18728 = pi14 ? n18709 : n18727;
  assign n18729 = pi13 ? n18700 : n18728;
  assign n18730 = pi12 ? n18680 : n18729;
  assign n18731 = pi18 ? n18332 : n11981;
  assign n18732 = pi17 ? n18329 : n18731;
  assign n18733 = pi16 ? n915 : n18732;
  assign n18734 = pi15 ? n18733 : n18342;
  assign n18735 = pi18 ? n10903 : n316;
  assign n18736 = pi17 ? n32 : n18735;
  assign n18737 = pi16 ? n18736 : n18357;
  assign n18738 = pi15 ? n18348 : n18737;
  assign n18739 = pi14 ? n18734 : n18738;
  assign n18740 = pi21 ? n916 : n7048;
  assign n18741 = pi20 ? n18740 : n32;
  assign n18742 = pi19 ? n18741 : n32;
  assign n18743 = pi18 ? n18362 : n18742;
  assign n18744 = pi17 ? n139 : n18743;
  assign n18745 = pi16 ? n1773 : n18744;
  assign n18746 = pi15 ? n18737 : n18745;
  assign n18747 = pi21 ? n916 : n882;
  assign n18748 = pi20 ? n18747 : n32;
  assign n18749 = pi19 ? n18748 : n32;
  assign n18750 = pi18 ? n139 : n18749;
  assign n18751 = pi17 ? n139 : n18750;
  assign n18752 = pi16 ? n915 : n18751;
  assign n18753 = pi15 ? n18752 : n18379;
  assign n18754 = pi14 ? n18746 : n18753;
  assign n18755 = pi13 ? n18739 : n18754;
  assign n18756 = pi21 ? n233 : n1009;
  assign n18757 = pi20 ? n18756 : n32;
  assign n18758 = pi19 ? n18757 : n32;
  assign n18759 = pi18 ? n17487 : n18758;
  assign n18760 = pi17 ? n17485 : n18759;
  assign n18761 = pi16 ? n439 : n18760;
  assign n18762 = pi15 ? n18391 : n18761;
  assign n18763 = pi14 ? n18762 : n18418;
  assign n18764 = pi22 ? n2060 : n1070;
  assign n18765 = pi21 ? n18764 : n32;
  assign n18766 = pi20 ? n18765 : n32;
  assign n18767 = pi19 ? n18766 : n32;
  assign n18768 = pi18 ? n17487 : n18767;
  assign n18769 = pi17 ? n18423 : n18768;
  assign n18770 = pi16 ? n18421 : n18769;
  assign n18771 = pi22 ? n2060 : n6415;
  assign n18772 = pi21 ? n18771 : n32;
  assign n18773 = pi20 ? n18772 : n32;
  assign n18774 = pi19 ? n18773 : n32;
  assign n18775 = pi18 ? n18436 : n18774;
  assign n18776 = pi17 ? n18434 : n18775;
  assign n18777 = pi16 ? n10118 : n18776;
  assign n18778 = pi15 ? n18770 : n18777;
  assign n18779 = pi22 ? n448 : n3338;
  assign n18780 = pi21 ? n18779 : n32;
  assign n18781 = pi20 ? n18780 : n32;
  assign n18782 = pi19 ? n18781 : n32;
  assign n18783 = pi18 ? n18447 : n18782;
  assign n18784 = pi17 ? n18445 : n18783;
  assign n18785 = pi16 ? n10118 : n18784;
  assign n18786 = pi22 ? n962 : n9827;
  assign n18787 = pi21 ? n18786 : n363;
  assign n18788 = pi20 ? n32 : n18787;
  assign n18789 = pi19 ? n32 : n18788;
  assign n18790 = pi22 ? n9827 : n18461;
  assign n18791 = pi21 ? n18790 : n17548;
  assign n18792 = pi22 ? n9827 : n363;
  assign n18793 = pi21 ? n18792 : n17548;
  assign n18794 = pi20 ? n18791 : n18793;
  assign n18795 = pi23 ? n363 : n139;
  assign n18796 = pi22 ? n18461 : n18795;
  assign n18797 = pi21 ? n18796 : n9143;
  assign n18798 = pi22 ? n363 : n18795;
  assign n18799 = pi21 ? n18798 : n17548;
  assign n18800 = pi20 ? n18797 : n18799;
  assign n18801 = pi19 ? n18794 : n18800;
  assign n18802 = pi18 ? n18789 : n18801;
  assign n18803 = pi17 ? n32 : n18802;
  assign n18804 = pi22 ? n18461 : n364;
  assign n18805 = pi21 ? n18804 : n233;
  assign n18806 = pi21 ? n233 : n18792;
  assign n18807 = pi20 ? n18805 : n18806;
  assign n18808 = pi22 ? n18461 : n139;
  assign n18809 = pi21 ? n17548 : n18808;
  assign n18810 = pi21 ? n363 : n18804;
  assign n18811 = pi20 ? n18809 : n18810;
  assign n18812 = pi19 ? n18807 : n18811;
  assign n18813 = pi21 ? n9836 : n233;
  assign n18814 = pi20 ? n18813 : n18481;
  assign n18815 = pi19 ? n18814 : n233;
  assign n18816 = pi18 ? n18812 : n18815;
  assign n18817 = pi17 ? n18816 : n18485;
  assign n18818 = pi16 ? n18803 : n18817;
  assign n18819 = pi15 ? n18785 : n18818;
  assign n18820 = pi14 ? n18778 : n18819;
  assign n18821 = pi13 ? n18763 : n18820;
  assign n18822 = pi12 ? n18755 : n18821;
  assign n18823 = pi11 ? n18730 : n18822;
  assign n18824 = pi10 ? n18638 : n18823;
  assign n18825 = pi09 ? n17942 : n18824;
  assign n18826 = pi08 ? n18494 : n18825;
  assign n18827 = pi07 ? n17929 : n18826;
  assign n18828 = pi06 ? n16971 : n18827;
  assign n18829 = pi20 ? n37 : n4528;
  assign n18830 = pi19 ? n18829 : n32;
  assign n18831 = pi18 ? n37 : n18830;
  assign n18832 = pi17 ? n37 : n18831;
  assign n18833 = pi16 ? n11885 : n18832;
  assign n18834 = pi15 ? n32 : n18833;
  assign n18835 = pi16 ? n12689 : n18832;
  assign n18836 = pi14 ? n18834 : n18835;
  assign n18837 = pi13 ? n32 : n18836;
  assign n18838 = pi12 ? n32 : n18837;
  assign n18839 = pi11 ? n32 : n18838;
  assign n18840 = pi10 ? n32 : n18839;
  assign n18841 = pi20 ? n37 : n4566;
  assign n18842 = pi19 ? n18841 : n32;
  assign n18843 = pi18 ? n37 : n18842;
  assign n18844 = pi17 ? n37 : n18843;
  assign n18845 = pi16 ? n13561 : n18844;
  assign n18846 = pi21 ? n303 : n32;
  assign n18847 = pi20 ? n37 : n18846;
  assign n18848 = pi19 ? n18847 : n32;
  assign n18849 = pi18 ? n37 : n18848;
  assign n18850 = pi17 ? n37 : n18849;
  assign n18851 = pi16 ? n14445 : n18850;
  assign n18852 = pi15 ? n18845 : n18851;
  assign n18853 = pi20 ? n226 : n99;
  assign n18854 = pi19 ? n18853 : n99;
  assign n18855 = pi18 ? n15515 : n18854;
  assign n18856 = pi17 ? n32 : n18855;
  assign n18857 = pi20 ? n99 : n5420;
  assign n18858 = pi19 ? n18857 : n99;
  assign n18859 = pi20 ? n99 : n5624;
  assign n18860 = pi19 ? n18859 : n32;
  assign n18861 = pi18 ? n18858 : n18860;
  assign n18862 = pi17 ? n99 : n18861;
  assign n18863 = pi16 ? n18856 : n18862;
  assign n18864 = pi20 ? n181 : n17975;
  assign n18865 = pi19 ? n18864 : n32;
  assign n18866 = pi18 ? n37 : n18865;
  assign n18867 = pi17 ? n37 : n18866;
  assign n18868 = pi16 ? n17010 : n18867;
  assign n18869 = pi15 ? n18863 : n18868;
  assign n18870 = pi14 ? n18852 : n18869;
  assign n18871 = pi16 ? n439 : n17933;
  assign n18872 = pi20 ? n7745 : n4560;
  assign n18873 = pi19 ? n18872 : n32;
  assign n18874 = pi18 ? n37 : n18873;
  assign n18875 = pi17 ? n37 : n18874;
  assign n18876 = pi16 ? n439 : n18875;
  assign n18877 = pi15 ? n18871 : n18876;
  assign n18878 = pi21 ? n11938 : n32;
  assign n18879 = pi20 ? n99 : n18878;
  assign n18880 = pi19 ? n18879 : n32;
  assign n18881 = pi18 ? n99 : n18880;
  assign n18882 = pi17 ? n99 : n18881;
  assign n18883 = pi16 ? n201 : n18882;
  assign n18884 = pi21 ? n11945 : n32;
  assign n18885 = pi20 ? n99 : n18884;
  assign n18886 = pi19 ? n18885 : n32;
  assign n18887 = pi18 ? n99 : n18886;
  assign n18888 = pi17 ? n99 : n18887;
  assign n18889 = pi16 ? n801 : n18888;
  assign n18890 = pi15 ? n18883 : n18889;
  assign n18891 = pi14 ? n18877 : n18890;
  assign n18892 = pi13 ? n18870 : n18891;
  assign n18893 = pi16 ? n744 : n18888;
  assign n18894 = pi22 ? n99 : n625;
  assign n18895 = pi21 ? n18894 : n32;
  assign n18896 = pi20 ? n99 : n18895;
  assign n18897 = pi19 ? n18896 : n32;
  assign n18898 = pi18 ? n99 : n18897;
  assign n18899 = pi17 ? n99 : n18898;
  assign n18900 = pi16 ? n721 : n18899;
  assign n18901 = pi15 ? n18893 : n18900;
  assign n18902 = pi19 ? n37 : n15004;
  assign n18903 = pi18 ? n374 : n18902;
  assign n18904 = pi17 ? n32 : n18903;
  assign n18905 = pi22 ? n139 : n625;
  assign n18906 = pi21 ? n18905 : n32;
  assign n18907 = pi20 ? n139 : n18906;
  assign n18908 = pi19 ? n18907 : n32;
  assign n18909 = pi18 ? n139 : n18908;
  assign n18910 = pi17 ? n139 : n18909;
  assign n18911 = pi16 ? n18904 : n18910;
  assign n18912 = pi20 ? n37 : n1761;
  assign n18913 = pi19 ? n37 : n18912;
  assign n18914 = pi18 ? n374 : n18913;
  assign n18915 = pi17 ? n32 : n18914;
  assign n18916 = pi22 ? n139 : n688;
  assign n18917 = pi21 ? n18916 : n32;
  assign n18918 = pi20 ? n139 : n18917;
  assign n18919 = pi19 ? n18918 : n32;
  assign n18920 = pi18 ? n139 : n18919;
  assign n18921 = pi17 ? n139 : n18920;
  assign n18922 = pi16 ? n18915 : n18921;
  assign n18923 = pi15 ? n18911 : n18922;
  assign n18924 = pi14 ? n18901 : n18923;
  assign n18925 = pi19 ? n9765 : n9769;
  assign n18926 = pi18 ? n18925 : n139;
  assign n18927 = pi22 ? n335 : n688;
  assign n18928 = pi21 ? n18927 : n32;
  assign n18929 = pi20 ? n139 : n18928;
  assign n18930 = pi19 ? n18929 : n32;
  assign n18931 = pi18 ? n139 : n18930;
  assign n18932 = pi17 ? n18926 : n18931;
  assign n18933 = pi16 ? n439 : n18932;
  assign n18934 = pi20 ? n37 : n297;
  assign n18935 = pi19 ? n37 : n18934;
  assign n18936 = pi18 ? n18935 : n6598;
  assign n18937 = pi21 ? n365 : n32;
  assign n18938 = pi20 ? n139 : n18937;
  assign n18939 = pi19 ? n18938 : n32;
  assign n18940 = pi18 ? n139 : n18939;
  assign n18941 = pi17 ? n18936 : n18940;
  assign n18942 = pi16 ? n439 : n18941;
  assign n18943 = pi15 ? n18933 : n18942;
  assign n18944 = pi19 ? n9824 : n2374;
  assign n18945 = pi18 ? n37 : n18944;
  assign n18946 = pi21 ? n12389 : n32;
  assign n18947 = pi20 ? n139 : n18946;
  assign n18948 = pi19 ? n18947 : n32;
  assign n18949 = pi18 ? n139 : n18948;
  assign n18950 = pi17 ? n18945 : n18949;
  assign n18951 = pi16 ? n439 : n18950;
  assign n18952 = pi21 ? n3073 : n1211;
  assign n18953 = pi20 ? n18952 : n14043;
  assign n18954 = pi19 ? n18953 : n14045;
  assign n18955 = pi20 ? n14061 : n4749;
  assign n18956 = pi19 ? n18955 : n32;
  assign n18957 = pi18 ? n18954 : n18956;
  assign n18958 = pi17 ? n37 : n18957;
  assign n18959 = pi16 ? n439 : n18958;
  assign n18960 = pi15 ? n18951 : n18959;
  assign n18961 = pi14 ? n18943 : n18960;
  assign n18962 = pi13 ? n18924 : n18961;
  assign n18963 = pi12 ? n18892 : n18962;
  assign n18964 = pi20 ? n37 : n14352;
  assign n18965 = pi19 ? n18964 : n32;
  assign n18966 = pi18 ? n37 : n18965;
  assign n18967 = pi17 ? n37 : n18966;
  assign n18968 = pi16 ? n439 : n18967;
  assign n18969 = pi20 ? n1057 : n204;
  assign n18970 = pi19 ? n18969 : n204;
  assign n18971 = pi21 ? n12404 : n32;
  assign n18972 = pi20 ? n204 : n18971;
  assign n18973 = pi19 ? n18972 : n32;
  assign n18974 = pi18 ? n18970 : n18973;
  assign n18975 = pi17 ? n37 : n18974;
  assign n18976 = pi16 ? n439 : n18975;
  assign n18977 = pi15 ? n18968 : n18976;
  assign n18978 = pi21 ? n1056 : n139;
  assign n18979 = pi20 ? n18978 : n204;
  assign n18980 = pi19 ? n18979 : n204;
  assign n18981 = pi18 ? n18980 : n18973;
  assign n18982 = pi17 ? n37 : n18981;
  assign n18983 = pi16 ? n439 : n18982;
  assign n18984 = pi20 ? n37 : n1057;
  assign n18985 = pi19 ? n18984 : n204;
  assign n18986 = pi18 ? n18985 : n18973;
  assign n18987 = pi17 ? n37 : n18986;
  assign n18988 = pi16 ? n439 : n18987;
  assign n18989 = pi15 ? n18983 : n18988;
  assign n18990 = pi14 ? n18977 : n18989;
  assign n18991 = pi21 ? n37 : n9871;
  assign n18992 = pi20 ? n37 : n18991;
  assign n18993 = pi23 ? n233 : n204;
  assign n18994 = pi22 ? n4079 : n18993;
  assign n18995 = pi22 ? n18993 : n233;
  assign n18996 = pi21 ? n18994 : n18995;
  assign n18997 = pi22 ? n4079 : n204;
  assign n18998 = pi21 ? n18997 : n18995;
  assign n18999 = pi20 ? n18996 : n18998;
  assign n19000 = pi19 ? n18992 : n18999;
  assign n19001 = pi21 ? n18993 : n204;
  assign n19002 = pi20 ? n19001 : n18971;
  assign n19003 = pi19 ? n19002 : n32;
  assign n19004 = pi18 ? n19000 : n19003;
  assign n19005 = pi17 ? n37 : n19004;
  assign n19006 = pi16 ? n439 : n19005;
  assign n19007 = pi20 ? n335 : n7035;
  assign n19008 = pi19 ? n19007 : n32;
  assign n19009 = pi18 ? n15099 : n19008;
  assign n19010 = pi17 ? n37 : n19009;
  assign n19011 = pi16 ? n439 : n19010;
  assign n19012 = pi15 ? n19006 : n19011;
  assign n19013 = pi18 ? n16138 : n19008;
  assign n19014 = pi17 ? n37 : n19013;
  assign n19015 = pi16 ? n439 : n19014;
  assign n19016 = pi18 ? n9856 : n19008;
  assign n19017 = pi17 ? n37 : n19016;
  assign n19018 = pi16 ? n439 : n19017;
  assign n19019 = pi15 ? n19015 : n19018;
  assign n19020 = pi14 ? n19012 : n19019;
  assign n19021 = pi13 ? n18990 : n19020;
  assign n19022 = pi20 ? n605 : n7035;
  assign n19023 = pi19 ? n19022 : n32;
  assign n19024 = pi18 ? n10682 : n19023;
  assign n19025 = pi17 ? n37 : n19024;
  assign n19026 = pi16 ? n439 : n19025;
  assign n19027 = pi20 ? n569 : n7724;
  assign n19028 = pi19 ? n19027 : n32;
  assign n19029 = pi18 ? n7677 : n19028;
  assign n19030 = pi17 ? n37 : n19029;
  assign n19031 = pi16 ? n439 : n19030;
  assign n19032 = pi15 ? n19026 : n19031;
  assign n19033 = pi20 ? n2094 : n7724;
  assign n19034 = pi19 ? n19033 : n32;
  assign n19035 = pi18 ? n37 : n19034;
  assign n19036 = pi17 ? n37 : n19035;
  assign n19037 = pi16 ? n439 : n19036;
  assign n19038 = pi20 ? n37 : n2091;
  assign n19039 = pi19 ? n37 : n19038;
  assign n19040 = pi20 ? n18162 : n4102;
  assign n19041 = pi19 ? n19040 : n32;
  assign n19042 = pi18 ? n19039 : n19041;
  assign n19043 = pi17 ? n37 : n19042;
  assign n19044 = pi16 ? n439 : n19043;
  assign n19045 = pi15 ? n19037 : n19044;
  assign n19046 = pi14 ? n19032 : n19045;
  assign n19047 = pi20 ? n233 : n3340;
  assign n19048 = pi19 ? n19047 : n32;
  assign n19049 = pi18 ? n16209 : n19048;
  assign n19050 = pi17 ? n37 : n19049;
  assign n19051 = pi16 ? n439 : n19050;
  assign n19052 = pi21 ? n233 : n11635;
  assign n19053 = pi20 ? n6402 : n19052;
  assign n19054 = pi19 ? n37 : n19053;
  assign n19055 = pi20 ? n15177 : n2638;
  assign n19056 = pi19 ? n19055 : n32;
  assign n19057 = pi18 ? n19054 : n19056;
  assign n19058 = pi17 ? n37 : n19057;
  assign n19059 = pi16 ? n439 : n19058;
  assign n19060 = pi15 ? n19051 : n19059;
  assign n19061 = pi20 ? n2106 : n2638;
  assign n19062 = pi19 ? n19061 : n32;
  assign n19063 = pi18 ? n2109 : n19062;
  assign n19064 = pi17 ? n37 : n19063;
  assign n19065 = pi16 ? n439 : n19064;
  assign n19066 = pi20 ? n2107 : n2653;
  assign n19067 = pi19 ? n19066 : n32;
  assign n19068 = pi18 ? n2109 : n19067;
  assign n19069 = pi17 ? n37 : n19068;
  assign n19070 = pi16 ? n439 : n19069;
  assign n19071 = pi15 ? n19065 : n19070;
  assign n19072 = pi14 ? n19060 : n19071;
  assign n19073 = pi13 ? n19046 : n19072;
  assign n19074 = pi12 ? n19021 : n19073;
  assign n19075 = pi11 ? n18963 : n19074;
  assign n19076 = pi21 ? n685 : n2106;
  assign n19077 = pi20 ? n37 : n19076;
  assign n19078 = pi19 ? n37 : n19077;
  assign n19079 = pi20 ? n2106 : n2470;
  assign n19080 = pi19 ? n19079 : n32;
  assign n19081 = pi18 ? n19078 : n19080;
  assign n19082 = pi17 ? n37 : n19081;
  assign n19083 = pi16 ? n439 : n19082;
  assign n19084 = pi21 ? n363 : n2721;
  assign n19085 = pi20 ? n19084 : n2470;
  assign n19086 = pi19 ? n19085 : n32;
  assign n19087 = pi18 ? n2731 : n19086;
  assign n19088 = pi17 ? n37 : n19087;
  assign n19089 = pi16 ? n439 : n19088;
  assign n19090 = pi15 ? n19083 : n19089;
  assign n19091 = pi21 ? n37 : n5015;
  assign n19092 = pi20 ? n37 : n19091;
  assign n19093 = pi19 ? n37 : n19092;
  assign n19094 = pi20 ? n18212 : n2554;
  assign n19095 = pi19 ? n19094 : n32;
  assign n19096 = pi18 ? n19093 : n19095;
  assign n19097 = pi17 ? n37 : n19096;
  assign n19098 = pi16 ? n439 : n19097;
  assign n19099 = pi20 ? n2107 : n2554;
  assign n19100 = pi19 ? n19099 : n32;
  assign n19101 = pi18 ? n37 : n19100;
  assign n19102 = pi17 ? n37 : n19101;
  assign n19103 = pi16 ? n439 : n19102;
  assign n19104 = pi15 ? n19098 : n19103;
  assign n19105 = pi14 ? n19090 : n19104;
  assign n19106 = pi21 ? n37 : n14246;
  assign n19107 = pi20 ? n99 : n19106;
  assign n19108 = pi19 ? n99 : n19107;
  assign n19109 = pi21 ? n99 : n2106;
  assign n19110 = pi20 ? n19109 : n2679;
  assign n19111 = pi19 ? n19110 : n32;
  assign n19112 = pi18 ? n19108 : n19111;
  assign n19113 = pi17 ? n99 : n19112;
  assign n19114 = pi16 ? n201 : n19113;
  assign n19115 = pi20 ? n5085 : n2679;
  assign n19116 = pi19 ? n19115 : n32;
  assign n19117 = pi18 ? n13377 : n19116;
  assign n19118 = pi17 ? n99 : n19117;
  assign n19119 = pi16 ? n801 : n19118;
  assign n19120 = pi15 ? n19114 : n19119;
  assign n19121 = pi18 ? n13377 : n18669;
  assign n19122 = pi17 ? n99 : n19121;
  assign n19123 = pi16 ? n721 : n19122;
  assign n19124 = pi19 ? n99 : n2255;
  assign n19125 = pi18 ? n99 : n19124;
  assign n19126 = pi20 ? n685 : n1822;
  assign n19127 = pi19 ? n19126 : n32;
  assign n19128 = pi18 ? n5087 : n19127;
  assign n19129 = pi17 ? n19125 : n19128;
  assign n19130 = pi16 ? n721 : n19129;
  assign n19131 = pi15 ? n19123 : n19130;
  assign n19132 = pi14 ? n19120 : n19131;
  assign n19133 = pi13 ? n19105 : n19132;
  assign n19134 = pi20 ? n99 : n157;
  assign n19135 = pi19 ? n99 : n19134;
  assign n19136 = pi18 ? n99 : n19135;
  assign n19137 = pi20 ? n157 : n15263;
  assign n19138 = pi20 ? n157 : n685;
  assign n19139 = pi19 ? n19137 : n19138;
  assign n19140 = pi20 ? n685 : n32;
  assign n19141 = pi19 ? n19140 : n32;
  assign n19142 = pi18 ? n19139 : n19141;
  assign n19143 = pi17 ? n19136 : n19142;
  assign n19144 = pi16 ? n721 : n19143;
  assign n19145 = pi19 ? n7845 : n99;
  assign n19146 = pi18 ? n719 : n19145;
  assign n19147 = pi17 ? n32 : n19146;
  assign n19148 = pi19 ? n161 : n2265;
  assign n19149 = pi20 ? n802 : n15263;
  assign n19150 = pi19 ? n19149 : n157;
  assign n19151 = pi18 ? n19148 : n19150;
  assign n19152 = pi19 ? n157 : n6512;
  assign n19153 = pi22 ? n157 : n5452;
  assign n19154 = pi21 ? n19153 : n3562;
  assign n19155 = pi20 ? n19154 : n32;
  assign n19156 = pi19 ? n19155 : n32;
  assign n19157 = pi18 ? n19152 : n19156;
  assign n19158 = pi17 ? n19151 : n19157;
  assign n19159 = pi16 ? n19147 : n19158;
  assign n19160 = pi15 ? n19144 : n19159;
  assign n19161 = pi22 ? n1504 : n157;
  assign n19162 = pi21 ? n19161 : n157;
  assign n19163 = pi20 ? n32 : n19162;
  assign n19164 = pi19 ? n32 : n19163;
  assign n19165 = pi18 ? n19164 : n157;
  assign n19166 = pi17 ? n32 : n19165;
  assign n19167 = pi18 ? n16324 : n157;
  assign n19168 = pi21 ? n99 : n18276;
  assign n19169 = pi20 ? n157 : n19168;
  assign n19170 = pi19 ? n157 : n19169;
  assign n19171 = pi21 ? n99 : n3562;
  assign n19172 = pi20 ? n19171 : n32;
  assign n19173 = pi19 ? n19172 : n32;
  assign n19174 = pi18 ? n19170 : n19173;
  assign n19175 = pi17 ? n19167 : n19174;
  assign n19176 = pi16 ? n19166 : n19175;
  assign n19177 = pi23 ? n99 : n316;
  assign n19178 = pi22 ? n19177 : n157;
  assign n19179 = pi21 ? n157 : n19178;
  assign n19180 = pi20 ? n157 : n19179;
  assign n19181 = pi19 ? n157 : n19180;
  assign n19182 = pi20 ? n5161 : n32;
  assign n19183 = pi19 ? n19182 : n32;
  assign n19184 = pi18 ? n19181 : n19183;
  assign n19185 = pi17 ? n157 : n19184;
  assign n19186 = pi16 ? n12535 : n19185;
  assign n19187 = pi15 ? n19176 : n19186;
  assign n19188 = pi14 ? n19160 : n19187;
  assign n19189 = pi18 ? n157 : n16324;
  assign n19190 = pi18 ? n17368 : n12349;
  assign n19191 = pi17 ? n19189 : n19190;
  assign n19192 = pi16 ? n12535 : n19191;
  assign n19193 = pi21 ? n3759 : n99;
  assign n19194 = pi22 ? n204 : n99;
  assign n19195 = pi21 ? n19194 : n99;
  assign n19196 = pi19 ? n19193 : n19195;
  assign n19197 = pi18 ? n742 : n19196;
  assign n19198 = pi17 ? n32 : n19197;
  assign n19199 = pi21 ? n19194 : n3759;
  assign n19200 = pi20 ? n19195 : n19199;
  assign n19201 = pi21 ? n99 : n19194;
  assign n19202 = pi19 ? n19200 : n19201;
  assign n19203 = pi20 ? n19201 : n19193;
  assign n19204 = pi20 ? n19193 : n3760;
  assign n19205 = pi19 ? n19203 : n19204;
  assign n19206 = pi18 ? n19202 : n19205;
  assign n19207 = pi20 ? n19201 : n19194;
  assign n19208 = pi21 ? n99 : n316;
  assign n19209 = pi20 ? n3759 : n19208;
  assign n19210 = pi19 ? n19207 : n19209;
  assign n19211 = pi18 ? n19210 : n12349;
  assign n19212 = pi17 ? n19206 : n19211;
  assign n19213 = pi16 ? n19198 : n19212;
  assign n19214 = pi15 ? n19192 : n19213;
  assign n19215 = pi21 ? n5186 : n204;
  assign n19216 = pi20 ? n32 : n19215;
  assign n19217 = pi19 ? n32 : n19216;
  assign n19218 = pi18 ? n19217 : n204;
  assign n19219 = pi17 ? n32 : n19218;
  assign n19220 = pi20 ? n204 : n1001;
  assign n19221 = pi19 ? n204 : n19220;
  assign n19222 = pi18 ? n204 : n19221;
  assign n19223 = pi19 ? n7454 : n3727;
  assign n19224 = pi18 ? n19223 : n12349;
  assign n19225 = pi17 ? n19222 : n19224;
  assign n19226 = pi16 ? n19219 : n19225;
  assign n19227 = pi20 ? n204 : n3087;
  assign n19228 = pi19 ? n204 : n19227;
  assign n19229 = pi19 ? n204 : n17409;
  assign n19230 = pi18 ? n19228 : n19229;
  assign n19231 = pi20 ? n204 : n316;
  assign n19232 = pi19 ? n10892 : n19231;
  assign n19233 = pi18 ? n19232 : n12349;
  assign n19234 = pi17 ? n19230 : n19233;
  assign n19235 = pi16 ? n11804 : n19234;
  assign n19236 = pi15 ? n19226 : n19235;
  assign n19237 = pi14 ? n19214 : n19236;
  assign n19238 = pi13 ? n19188 : n19237;
  assign n19239 = pi12 ? n19133 : n19238;
  assign n19240 = pi18 ? n139 : n11798;
  assign n19241 = pi20 ? n316 : n1022;
  assign n19242 = pi19 ? n19241 : n999;
  assign n19243 = pi18 ? n19242 : n12349;
  assign n19244 = pi17 ? n19240 : n19243;
  assign n19245 = pi16 ? n915 : n19244;
  assign n19246 = pi20 ? n139 : n6923;
  assign n19247 = pi19 ? n19246 : n139;
  assign n19248 = pi18 ? n19247 : n9111;
  assign n19249 = pi21 ? n356 : n5178;
  assign n19250 = pi20 ? n19249 : n32;
  assign n19251 = pi19 ? n19250 : n32;
  assign n19252 = pi18 ? n316 : n19251;
  assign n19253 = pi17 ? n19248 : n19252;
  assign n19254 = pi16 ? n915 : n19253;
  assign n19255 = pi15 ? n19245 : n19254;
  assign n19256 = pi18 ? n990 : n316;
  assign n19257 = pi17 ? n32 : n19256;
  assign n19258 = pi21 ? n356 : n4015;
  assign n19259 = pi20 ? n316 : n19258;
  assign n19260 = pi19 ? n316 : n19259;
  assign n19261 = pi18 ? n19260 : n316;
  assign n19262 = pi17 ? n19261 : n11501;
  assign n19263 = pi16 ? n19257 : n19262;
  assign n19264 = pi19 ? n2353 : n347;
  assign n19265 = pi18 ? n913 : n19264;
  assign n19266 = pi17 ? n32 : n19265;
  assign n19267 = pi20 ? n347 : n1001;
  assign n19268 = pi19 ? n19267 : n7557;
  assign n19269 = pi20 ? n4766 : n5317;
  assign n19270 = pi19 ? n19269 : n316;
  assign n19271 = pi18 ? n19268 : n19270;
  assign n19272 = pi21 ? n316 : n921;
  assign n19273 = pi20 ? n316 : n19272;
  assign n19274 = pi19 ? n316 : n19273;
  assign n19275 = pi21 ? n204 : n3523;
  assign n19276 = pi20 ? n19275 : n32;
  assign n19277 = pi19 ? n19276 : n32;
  assign n19278 = pi18 ? n19274 : n19277;
  assign n19279 = pi17 ? n19271 : n19278;
  assign n19280 = pi16 ? n19266 : n19279;
  assign n19281 = pi15 ? n19263 : n19280;
  assign n19282 = pi14 ? n19255 : n19281;
  assign n19283 = pi21 ? n1777 : n921;
  assign n19284 = pi21 ? n1777 : n2402;
  assign n19285 = pi20 ? n19283 : n19284;
  assign n19286 = pi22 ? n37 : n2401;
  assign n19287 = pi21 ? n139 : n19286;
  assign n19288 = pi19 ? n19285 : n19287;
  assign n19289 = pi18 ? n913 : n19288;
  assign n19290 = pi17 ? n32 : n19289;
  assign n19291 = pi20 ? n19287 : n19283;
  assign n19292 = pi22 ? n383 : n204;
  assign n19293 = pi22 ? n348 : n2299;
  assign n19294 = pi21 ? n19292 : n19293;
  assign n19295 = pi21 ? n921 : n19293;
  assign n19296 = pi20 ? n19294 : n19295;
  assign n19297 = pi19 ? n19291 : n19296;
  assign n19298 = pi21 ? n921 : n1777;
  assign n19299 = pi21 ? n8431 : n2876;
  assign n19300 = pi20 ? n19298 : n19299;
  assign n19301 = pi21 ? n5705 : n2402;
  assign n19302 = pi22 ? n1784 : n204;
  assign n19303 = pi21 ? n19292 : n19302;
  assign n19304 = pi20 ? n19301 : n19303;
  assign n19305 = pi19 ? n19300 : n19304;
  assign n19306 = pi18 ? n19297 : n19305;
  assign n19307 = pi21 ? n19302 : n19292;
  assign n19308 = pi22 ? n348 : n204;
  assign n19309 = pi21 ? n19308 : n19293;
  assign n19310 = pi20 ? n19307 : n19309;
  assign n19311 = pi22 ? n204 : n383;
  assign n19312 = pi21 ? n19311 : n8431;
  assign n19313 = pi20 ? n19312 : n204;
  assign n19314 = pi19 ? n19310 : n19313;
  assign n19315 = pi18 ? n19314 : n19277;
  assign n19316 = pi17 ? n19306 : n19315;
  assign n19317 = pi16 ? n19290 : n19316;
  assign n19318 = pi19 ? n204 : n1919;
  assign n19319 = pi18 ? n19318 : n204;
  assign n19320 = pi21 ? n204 : n7048;
  assign n19321 = pi20 ? n19320 : n32;
  assign n19322 = pi19 ? n19321 : n32;
  assign n19323 = pi18 ? n204 : n19322;
  assign n19324 = pi17 ? n19319 : n19323;
  assign n19325 = pi16 ? n13846 : n19324;
  assign n19326 = pi15 ? n19317 : n19325;
  assign n19327 = pi23 ? n8133 : n395;
  assign n19328 = pi22 ? n19327 : n32;
  assign n19329 = pi21 ? n204 : n19328;
  assign n19330 = pi20 ? n19329 : n32;
  assign n19331 = pi19 ? n19330 : n32;
  assign n19332 = pi18 ? n204 : n19331;
  assign n19333 = pi17 ? n204 : n19332;
  assign n19334 = pi16 ? n13477 : n19333;
  assign n19335 = pi18 ? n374 : n233;
  assign n19336 = pi17 ? n32 : n19335;
  assign n19337 = pi22 ? n233 : n204;
  assign n19338 = pi21 ? n233 : n19337;
  assign n19339 = pi20 ? n233 : n19338;
  assign n19340 = pi19 ? n19339 : n233;
  assign n19341 = pi21 ? n19337 : n882;
  assign n19342 = pi20 ? n19341 : n32;
  assign n19343 = pi19 ? n19342 : n32;
  assign n19344 = pi18 ? n19340 : n19343;
  assign n19345 = pi17 ? n233 : n19344;
  assign n19346 = pi16 ? n19336 : n19345;
  assign n19347 = pi15 ? n19334 : n19346;
  assign n19348 = pi14 ? n19326 : n19347;
  assign n19349 = pi13 ? n19282 : n19348;
  assign n19350 = pi19 ? n13337 : n37;
  assign n19351 = pi18 ? n19350 : n18113;
  assign n19352 = pi21 ? n233 : n928;
  assign n19353 = pi20 ? n19352 : n32;
  assign n19354 = pi19 ? n19353 : n32;
  assign n19355 = pi18 ? n233 : n19354;
  assign n19356 = pi17 ? n19351 : n19355;
  assign n19357 = pi16 ? n439 : n19356;
  assign n19358 = pi20 ? n8927 : n233;
  assign n19359 = pi19 ? n37 : n19358;
  assign n19360 = pi18 ? n37 : n19359;
  assign n19361 = pi21 ? n233 : n2678;
  assign n19362 = pi20 ? n19361 : n32;
  assign n19363 = pi19 ? n19362 : n32;
  assign n19364 = pi18 ? n233 : n19363;
  assign n19365 = pi17 ? n19360 : n19364;
  assign n19366 = pi16 ? n439 : n19365;
  assign n19367 = pi15 ? n19357 : n19366;
  assign n19368 = pi21 ? n569 : n574;
  assign n19369 = pi20 ? n37 : n19368;
  assign n19370 = pi19 ? n19369 : n37;
  assign n19371 = pi18 ? n19370 : n10682;
  assign n19372 = pi22 ? n10400 : n233;
  assign n19373 = pi21 ? n19372 : n2678;
  assign n19374 = pi20 ? n19373 : n32;
  assign n19375 = pi19 ? n19374 : n32;
  assign n19376 = pi18 ? n335 : n19375;
  assign n19377 = pi17 ? n19371 : n19376;
  assign n19378 = pi16 ? n439 : n19377;
  assign n19379 = pi20 ? n577 : n639;
  assign n19380 = pi19 ? n19379 : n37;
  assign n19381 = pi18 ? n374 : n19380;
  assign n19382 = pi17 ? n32 : n19381;
  assign n19383 = pi20 ? n335 : n8857;
  assign n19384 = pi19 ? n335 : n19383;
  assign n19385 = pi18 ? n19384 : n335;
  assign n19386 = pi22 ? n2060 : n233;
  assign n19387 = pi21 ? n19386 : n2700;
  assign n19388 = pi20 ? n19387 : n32;
  assign n19389 = pi19 ? n19388 : n32;
  assign n19390 = pi18 ? n335 : n19389;
  assign n19391 = pi17 ? n19385 : n19390;
  assign n19392 = pi16 ? n19382 : n19391;
  assign n19393 = pi15 ? n19378 : n19392;
  assign n19394 = pi14 ? n19367 : n19393;
  assign n19395 = pi21 ? n796 : n37;
  assign n19396 = pi20 ? n32 : n19395;
  assign n19397 = pi19 ? n32 : n19396;
  assign n19398 = pi20 ? n569 : n647;
  assign n19399 = pi19 ? n19398 : n37;
  assign n19400 = pi18 ? n19397 : n19399;
  assign n19401 = pi17 ? n32 : n19400;
  assign n19402 = pi21 ? n218 : n569;
  assign n19403 = pi20 ? n335 : n19402;
  assign n19404 = pi19 ? n10681 : n19403;
  assign n19405 = pi20 ? n335 : n16544;
  assign n19406 = pi19 ? n335 : n19405;
  assign n19407 = pi18 ? n19404 : n19406;
  assign n19408 = pi22 ? n2060 : n6365;
  assign n19409 = pi21 ? n19408 : n1009;
  assign n19410 = pi20 ? n19409 : n32;
  assign n19411 = pi19 ? n19410 : n32;
  assign n19412 = pi18 ? n335 : n19411;
  assign n19413 = pi17 ? n19407 : n19412;
  assign n19414 = pi16 ? n19401 : n19413;
  assign n19415 = pi18 ? n335 : n19406;
  assign n19416 = pi20 ? n233 : n15465;
  assign n19417 = pi19 ? n19416 : n335;
  assign n19418 = pi18 ? n19417 : n17900;
  assign n19419 = pi17 ? n19415 : n19418;
  assign n19420 = pi16 ? n10980 : n19419;
  assign n19421 = pi15 ? n19414 : n19420;
  assign n19422 = pi21 ? n363 : n233;
  assign n19423 = pi20 ? n19422 : n233;
  assign n19424 = pi19 ? n335 : n19423;
  assign n19425 = pi18 ? n335 : n19424;
  assign n19426 = pi18 ? n233 : n17907;
  assign n19427 = pi17 ? n19425 : n19426;
  assign n19428 = pi16 ? n10980 : n19427;
  assign n19429 = pi23 ? n961 : n363;
  assign n19430 = pi22 ? n19429 : n363;
  assign n19431 = pi21 ? n19430 : n363;
  assign n19432 = pi20 ? n32 : n19431;
  assign n19433 = pi19 ? n32 : n19432;
  assign n19434 = pi20 ? n15177 : n233;
  assign n19435 = pi19 ? n233 : n19434;
  assign n19436 = pi18 ? n19433 : n19435;
  assign n19437 = pi17 ? n32 : n19436;
  assign n19438 = pi22 ? n233 : n1475;
  assign n19439 = pi21 ? n19438 : n32;
  assign n19440 = pi20 ? n19439 : n32;
  assign n19441 = pi19 ? n19440 : n32;
  assign n19442 = pi18 ? n233 : n19441;
  assign n19443 = pi17 ? n233 : n19442;
  assign n19444 = pi16 ? n19437 : n19443;
  assign n19445 = pi15 ? n19428 : n19444;
  assign n19446 = pi14 ? n19421 : n19445;
  assign n19447 = pi13 ? n19394 : n19446;
  assign n19448 = pi12 ? n19349 : n19447;
  assign n19449 = pi11 ? n19239 : n19448;
  assign n19450 = pi10 ? n19075 : n19449;
  assign n19451 = pi09 ? n18840 : n19450;
  assign n19452 = pi21 ? n12224 : n32;
  assign n19453 = pi20 ? n37 : n19452;
  assign n19454 = pi19 ? n19453 : n32;
  assign n19455 = pi18 ? n37 : n19454;
  assign n19456 = pi17 ? n37 : n19455;
  assign n19457 = pi16 ? n12689 : n19456;
  assign n19458 = pi15 ? n19457 : n18835;
  assign n19459 = pi14 ? n18834 : n19458;
  assign n19460 = pi13 ? n32 : n19459;
  assign n19461 = pi12 ? n32 : n19460;
  assign n19462 = pi11 ? n32 : n19461;
  assign n19463 = pi10 ? n32 : n19462;
  assign n19464 = pi20 ? n37 : n5438;
  assign n19465 = pi19 ? n19464 : n32;
  assign n19466 = pi18 ? n37 : n19465;
  assign n19467 = pi17 ? n37 : n19466;
  assign n19468 = pi16 ? n13561 : n19467;
  assign n19469 = pi15 ? n19468 : n18851;
  assign n19470 = pi20 ? n99 : n221;
  assign n19471 = pi19 ? n19470 : n99;
  assign n19472 = pi18 ? n19471 : n18860;
  assign n19473 = pi17 ? n99 : n19472;
  assign n19474 = pi16 ? n18856 : n19473;
  assign n19475 = pi15 ? n19474 : n18868;
  assign n19476 = pi14 ? n19469 : n19475;
  assign n19477 = pi22 ? n37 : n5631;
  assign n19478 = pi21 ? n19477 : n32;
  assign n19479 = pi20 ? n37 : n19478;
  assign n19480 = pi19 ? n19479 : n32;
  assign n19481 = pi18 ? n37 : n19480;
  assign n19482 = pi17 ? n37 : n19481;
  assign n19483 = pi16 ? n439 : n19482;
  assign n19484 = pi20 ? n7745 : n5483;
  assign n19485 = pi19 ? n19484 : n32;
  assign n19486 = pi18 ? n37 : n19485;
  assign n19487 = pi17 ? n37 : n19486;
  assign n19488 = pi16 ? n439 : n19487;
  assign n19489 = pi15 ? n19483 : n19488;
  assign n19490 = pi20 ? n99 : n5483;
  assign n19491 = pi19 ? n19490 : n32;
  assign n19492 = pi18 ? n99 : n19491;
  assign n19493 = pi17 ? n99 : n19492;
  assign n19494 = pi16 ? n201 : n19493;
  assign n19495 = pi21 ? n12747 : n32;
  assign n19496 = pi20 ? n99 : n19495;
  assign n19497 = pi19 ? n19496 : n32;
  assign n19498 = pi18 ? n99 : n19497;
  assign n19499 = pi17 ? n99 : n19498;
  assign n19500 = pi16 ? n801 : n19499;
  assign n19501 = pi15 ? n19494 : n19500;
  assign n19502 = pi14 ? n19489 : n19501;
  assign n19503 = pi13 ? n19476 : n19502;
  assign n19504 = pi16 ? n744 : n19499;
  assign n19505 = pi21 ? n13086 : n32;
  assign n19506 = pi20 ? n99 : n19505;
  assign n19507 = pi19 ? n19506 : n32;
  assign n19508 = pi18 ? n99 : n19507;
  assign n19509 = pi17 ? n99 : n19508;
  assign n19510 = pi16 ? n744 : n19509;
  assign n19511 = pi15 ? n19504 : n19510;
  assign n19512 = pi20 ? n8707 : n1708;
  assign n19513 = pi19 ? n37 : n19512;
  assign n19514 = pi18 ? n374 : n19513;
  assign n19515 = pi17 ? n32 : n19514;
  assign n19516 = pi21 ? n13102 : n32;
  assign n19517 = pi20 ? n139 : n19516;
  assign n19518 = pi19 ? n19517 : n32;
  assign n19519 = pi18 ? n139 : n19518;
  assign n19520 = pi17 ? n139 : n19519;
  assign n19521 = pi16 ? n19515 : n19520;
  assign n19522 = pi22 ? n139 : n1407;
  assign n19523 = pi21 ? n19522 : n32;
  assign n19524 = pi20 ? n139 : n19523;
  assign n19525 = pi19 ? n19524 : n32;
  assign n19526 = pi18 ? n139 : n19525;
  assign n19527 = pi17 ? n139 : n19526;
  assign n19528 = pi16 ? n18915 : n19527;
  assign n19529 = pi15 ? n19521 : n19528;
  assign n19530 = pi14 ? n19511 : n19529;
  assign n19531 = pi20 ? n139 : n8261;
  assign n19532 = pi19 ? n19531 : n32;
  assign n19533 = pi18 ? n139 : n19532;
  assign n19534 = pi17 ? n18926 : n19533;
  assign n19535 = pi16 ? n439 : n19534;
  assign n19536 = pi20 ? n139 : n5585;
  assign n19537 = pi19 ? n19536 : n32;
  assign n19538 = pi18 ? n139 : n19537;
  assign n19539 = pi17 ? n18936 : n19538;
  assign n19540 = pi16 ? n439 : n19539;
  assign n19541 = pi15 ? n19535 : n19540;
  assign n19542 = pi17 ? n18945 : n19538;
  assign n19543 = pi16 ? n439 : n19542;
  assign n19544 = pi15 ? n19543 : n18959;
  assign n19545 = pi14 ? n19541 : n19544;
  assign n19546 = pi13 ? n19530 : n19545;
  assign n19547 = pi12 ? n19503 : n19546;
  assign n19548 = pi22 ? n204 : n625;
  assign n19549 = pi21 ? n19548 : n32;
  assign n19550 = pi20 ? n37 : n19549;
  assign n19551 = pi19 ? n19550 : n32;
  assign n19552 = pi18 ? n37 : n19551;
  assign n19553 = pi17 ? n37 : n19552;
  assign n19554 = pi16 ? n439 : n19553;
  assign n19555 = pi20 ? n204 : n5747;
  assign n19556 = pi19 ? n19555 : n32;
  assign n19557 = pi18 ? n18970 : n19556;
  assign n19558 = pi17 ? n37 : n19557;
  assign n19559 = pi16 ? n439 : n19558;
  assign n19560 = pi15 ? n19554 : n19559;
  assign n19561 = pi20 ? n204 : n14352;
  assign n19562 = pi19 ? n19561 : n32;
  assign n19563 = pi18 ? n18980 : n19562;
  assign n19564 = pi17 ? n37 : n19563;
  assign n19565 = pi16 ? n439 : n19564;
  assign n19566 = pi15 ? n19565 : n18988;
  assign n19567 = pi14 ? n19560 : n19566;
  assign n19568 = pi21 ? n18994 : n3409;
  assign n19569 = pi22 ? n4079 : n456;
  assign n19570 = pi21 ? n19569 : n3409;
  assign n19571 = pi20 ? n19568 : n19570;
  assign n19572 = pi19 ? n18992 : n19571;
  assign n19573 = pi22 ? n18993 : n2116;
  assign n19574 = pi21 ? n19573 : n522;
  assign n19575 = pi20 ? n19574 : n18971;
  assign n19576 = pi19 ? n19575 : n32;
  assign n19577 = pi18 ? n19572 : n19576;
  assign n19578 = pi17 ? n37 : n19577;
  assign n19579 = pi16 ? n439 : n19578;
  assign n19580 = pi15 ? n19579 : n19011;
  assign n19581 = pi14 ? n19580 : n19019;
  assign n19582 = pi13 ? n19567 : n19581;
  assign n19583 = pi20 ? n233 : n4102;
  assign n19584 = pi19 ? n19583 : n32;
  assign n19585 = pi18 ? n16209 : n19584;
  assign n19586 = pi17 ? n37 : n19585;
  assign n19587 = pi16 ? n439 : n19586;
  assign n19588 = pi15 ? n19587 : n19059;
  assign n19589 = pi14 ? n19588 : n19071;
  assign n19590 = pi13 ? n19046 : n19589;
  assign n19591 = pi12 ? n19582 : n19590;
  assign n19592 = pi11 ? n19547 : n19591;
  assign n19593 = pi18 ? n19078 : n19062;
  assign n19594 = pi17 ? n37 : n19593;
  assign n19595 = pi16 ? n439 : n19594;
  assign n19596 = pi20 ? n19084 : n2638;
  assign n19597 = pi19 ? n19596 : n32;
  assign n19598 = pi18 ? n2731 : n19597;
  assign n19599 = pi17 ? n37 : n19598;
  assign n19600 = pi16 ? n439 : n19599;
  assign n19601 = pi15 ? n19595 : n19600;
  assign n19602 = pi20 ? n18212 : n2638;
  assign n19603 = pi19 ? n19602 : n32;
  assign n19604 = pi18 ? n19093 : n19603;
  assign n19605 = pi17 ? n37 : n19604;
  assign n19606 = pi16 ? n439 : n19605;
  assign n19607 = pi20 ? n2107 : n2638;
  assign n19608 = pi19 ? n19607 : n32;
  assign n19609 = pi18 ? n37 : n19608;
  assign n19610 = pi17 ? n37 : n19609;
  assign n19611 = pi16 ? n439 : n19610;
  assign n19612 = pi15 ? n19606 : n19611;
  assign n19613 = pi14 ? n19601 : n19612;
  assign n19614 = pi20 ? n19109 : n2638;
  assign n19615 = pi19 ? n19614 : n32;
  assign n19616 = pi18 ? n19108 : n19615;
  assign n19617 = pi17 ? n99 : n19616;
  assign n19618 = pi16 ? n201 : n19617;
  assign n19619 = pi20 ? n5085 : n2638;
  assign n19620 = pi19 ? n19619 : n32;
  assign n19621 = pi18 ? n13377 : n19620;
  assign n19622 = pi17 ? n99 : n19621;
  assign n19623 = pi16 ? n801 : n19622;
  assign n19624 = pi15 ? n19618 : n19623;
  assign n19625 = pi16 ? n744 : n19622;
  assign n19626 = pi20 ? n685 : n2653;
  assign n19627 = pi19 ? n19626 : n32;
  assign n19628 = pi18 ? n5087 : n19627;
  assign n19629 = pi17 ? n19125 : n19628;
  assign n19630 = pi16 ? n744 : n19629;
  assign n19631 = pi15 ? n19625 : n19630;
  assign n19632 = pi14 ? n19624 : n19631;
  assign n19633 = pi13 ? n19613 : n19632;
  assign n19634 = pi18 ? n19139 : n19127;
  assign n19635 = pi17 ? n19136 : n19634;
  assign n19636 = pi16 ? n744 : n19635;
  assign n19637 = pi18 ? n742 : n19145;
  assign n19638 = pi17 ? n32 : n19637;
  assign n19639 = pi21 ? n775 : n3562;
  assign n19640 = pi20 ? n19639 : n32;
  assign n19641 = pi19 ? n19640 : n32;
  assign n19642 = pi18 ? n19152 : n19641;
  assign n19643 = pi17 ? n19151 : n19642;
  assign n19644 = pi16 ? n19638 : n19643;
  assign n19645 = pi15 ? n19636 : n19644;
  assign n19646 = pi22 ? n55 : n157;
  assign n19647 = pi21 ? n19646 : n157;
  assign n19648 = pi20 ? n32 : n19647;
  assign n19649 = pi19 ? n32 : n19648;
  assign n19650 = pi18 ? n19649 : n157;
  assign n19651 = pi17 ? n32 : n19650;
  assign n19652 = pi18 ? n19170 : n18272;
  assign n19653 = pi17 ? n19167 : n19652;
  assign n19654 = pi16 ? n19651 : n19653;
  assign n19655 = pi20 ? n6543 : n32;
  assign n19656 = pi19 ? n19655 : n32;
  assign n19657 = pi18 ? n19181 : n19656;
  assign n19658 = pi17 ? n157 : n19657;
  assign n19659 = pi16 ? n12535 : n19658;
  assign n19660 = pi15 ? n19654 : n19659;
  assign n19661 = pi14 ? n19645 : n19660;
  assign n19662 = pi13 ? n19661 : n19237;
  assign n19663 = pi12 ? n19633 : n19662;
  assign n19664 = pi16 ? n2291 : n19244;
  assign n19665 = pi16 ? n2291 : n19253;
  assign n19666 = pi15 ? n19664 : n19665;
  assign n19667 = pi14 ? n19666 : n19281;
  assign n19668 = pi21 ? n820 : n921;
  assign n19669 = pi20 ? n19287 : n19668;
  assign n19670 = pi21 ? n1056 : n7217;
  assign n19671 = pi21 ? n921 : n7217;
  assign n19672 = pi20 ? n19670 : n19671;
  assign n19673 = pi19 ? n19669 : n19672;
  assign n19674 = pi21 ? n921 : n820;
  assign n19675 = pi21 ? n5559 : n2876;
  assign n19676 = pi20 ? n19674 : n19675;
  assign n19677 = pi21 ? n19292 : n1049;
  assign n19678 = pi20 ? n19301 : n19677;
  assign n19679 = pi19 ? n19676 : n19678;
  assign n19680 = pi18 ? n19673 : n19679;
  assign n19681 = pi21 ? n1049 : n19292;
  assign n19682 = pi21 ? n6676 : n7217;
  assign n19683 = pi20 ? n19681 : n19682;
  assign n19684 = pi21 ? n19311 : n5559;
  assign n19685 = pi20 ? n19684 : n204;
  assign n19686 = pi19 ? n19683 : n19685;
  assign n19687 = pi18 ? n19686 : n19277;
  assign n19688 = pi17 ? n19680 : n19687;
  assign n19689 = pi16 ? n19290 : n19688;
  assign n19690 = pi15 ? n19689 : n19325;
  assign n19691 = pi20 ? n5990 : n32;
  assign n19692 = pi19 ? n19691 : n32;
  assign n19693 = pi18 ? n204 : n19692;
  assign n19694 = pi17 ? n204 : n19693;
  assign n19695 = pi16 ? n13846 : n19694;
  assign n19696 = pi23 ? n316 : n14362;
  assign n19697 = pi22 ? n19696 : n32;
  assign n19698 = pi21 ? n19337 : n19697;
  assign n19699 = pi20 ? n19698 : n32;
  assign n19700 = pi19 ? n19699 : n32;
  assign n19701 = pi18 ? n19340 : n19700;
  assign n19702 = pi17 ? n233 : n19701;
  assign n19703 = pi16 ? n19336 : n19702;
  assign n19704 = pi15 ? n19695 : n19703;
  assign n19705 = pi14 ? n19690 : n19704;
  assign n19706 = pi13 ? n19667 : n19705;
  assign n19707 = pi21 ? n233 : n2553;
  assign n19708 = pi20 ? n19707 : n32;
  assign n19709 = pi19 ? n19708 : n32;
  assign n19710 = pi18 ? n233 : n19709;
  assign n19711 = pi17 ? n19360 : n19710;
  assign n19712 = pi16 ? n439 : n19711;
  assign n19713 = pi15 ? n19357 : n19712;
  assign n19714 = pi24 ? n335 : n363;
  assign n19715 = pi23 ? n335 : n19714;
  assign n19716 = pi22 ? n19715 : n233;
  assign n19717 = pi21 ? n19716 : n2678;
  assign n19718 = pi20 ? n19717 : n32;
  assign n19719 = pi19 ? n19718 : n32;
  assign n19720 = pi18 ? n335 : n19719;
  assign n19721 = pi17 ? n19371 : n19720;
  assign n19722 = pi16 ? n439 : n19721;
  assign n19723 = pi15 ? n19722 : n19392;
  assign n19724 = pi14 ? n19713 : n19723;
  assign n19725 = pi16 ? n12658 : n19427;
  assign n19726 = pi22 ? n233 : n759;
  assign n19727 = pi21 ? n19726 : n32;
  assign n19728 = pi20 ? n19727 : n32;
  assign n19729 = pi19 ? n19728 : n32;
  assign n19730 = pi18 ? n233 : n19729;
  assign n19731 = pi17 ? n233 : n19730;
  assign n19732 = pi16 ? n19437 : n19731;
  assign n19733 = pi15 ? n19725 : n19732;
  assign n19734 = pi14 ? n19421 : n19733;
  assign n19735 = pi13 ? n19724 : n19734;
  assign n19736 = pi12 ? n19706 : n19735;
  assign n19737 = pi11 ? n19663 : n19736;
  assign n19738 = pi10 ? n19592 : n19737;
  assign n19739 = pi09 ? n19463 : n19738;
  assign n19740 = pi08 ? n19451 : n19739;
  assign n19741 = pi20 ? n37 : n5396;
  assign n19742 = pi19 ? n19741 : n32;
  assign n19743 = pi18 ? n37 : n19742;
  assign n19744 = pi17 ? n37 : n19743;
  assign n19745 = pi16 ? n11885 : n19744;
  assign n19746 = pi15 ? n32 : n19745;
  assign n19747 = pi20 ? n37 : n6776;
  assign n19748 = pi19 ? n19747 : n32;
  assign n19749 = pi18 ? n37 : n19748;
  assign n19750 = pi17 ? n37 : n19749;
  assign n19751 = pi16 ? n12689 : n19750;
  assign n19752 = pi16 ? n13561 : n19744;
  assign n19753 = pi15 ? n19751 : n19752;
  assign n19754 = pi14 ? n19746 : n19753;
  assign n19755 = pi13 ? n32 : n19754;
  assign n19756 = pi12 ? n32 : n19755;
  assign n19757 = pi11 ? n32 : n19756;
  assign n19758 = pi10 ? n32 : n19757;
  assign n19759 = pi22 ? n99 : n9628;
  assign n19760 = pi21 ? n19759 : n32;
  assign n19761 = pi20 ? n37 : n19760;
  assign n19762 = pi19 ? n19761 : n32;
  assign n19763 = pi18 ? n37 : n19762;
  assign n19764 = pi17 ? n37 : n19763;
  assign n19765 = pi16 ? n13561 : n19764;
  assign n19766 = pi21 ? n13039 : n32;
  assign n19767 = pi20 ? n37 : n19766;
  assign n19768 = pi19 ? n19767 : n32;
  assign n19769 = pi18 ? n37 : n19768;
  assign n19770 = pi17 ? n37 : n19769;
  assign n19771 = pi16 ? n14445 : n19770;
  assign n19772 = pi15 ? n19765 : n19771;
  assign n19773 = pi20 ? n5077 : n99;
  assign n19774 = pi19 ? n19773 : n99;
  assign n19775 = pi18 ? n16593 : n19774;
  assign n19776 = pi17 ? n32 : n19775;
  assign n19777 = pi22 ? n139 : n1344;
  assign n19778 = pi21 ? n19777 : n32;
  assign n19779 = pi20 ? n99 : n19778;
  assign n19780 = pi19 ? n19779 : n32;
  assign n19781 = pi18 ? n99 : n19780;
  assign n19782 = pi17 ? n99 : n19781;
  assign n19783 = pi16 ? n19776 : n19782;
  assign n19784 = pi22 ? n37 : n103;
  assign n19785 = pi21 ? n19784 : n32;
  assign n19786 = pi20 ? n37 : n19785;
  assign n19787 = pi19 ? n19786 : n32;
  assign n19788 = pi18 ? n37 : n19787;
  assign n19789 = pi17 ? n37 : n19788;
  assign n19790 = pi16 ? n17010 : n19789;
  assign n19791 = pi15 ? n19783 : n19790;
  assign n19792 = pi14 ? n19772 : n19791;
  assign n19793 = pi22 ? n37 : n1370;
  assign n19794 = pi21 ? n19793 : n32;
  assign n19795 = pi20 ? n37 : n19794;
  assign n19796 = pi19 ? n19795 : n32;
  assign n19797 = pi18 ? n37 : n19796;
  assign n19798 = pi17 ? n37 : n19797;
  assign n19799 = pi16 ? n439 : n19798;
  assign n19800 = pi15 ? n19799 : n19488;
  assign n19801 = pi16 ? n801 : n19493;
  assign n19802 = pi15 ? n19494 : n19801;
  assign n19803 = pi14 ? n19800 : n19802;
  assign n19804 = pi13 ? n19792 : n19803;
  assign n19805 = pi16 ? n721 : n19499;
  assign n19806 = pi18 ? n374 : n16093;
  assign n19807 = pi17 ? n32 : n19806;
  assign n19808 = pi16 ? n19807 : n19520;
  assign n19809 = pi20 ? n13121 : n139;
  assign n19810 = pi19 ? n19809 : n139;
  assign n19811 = pi18 ? n19810 : n139;
  assign n19812 = pi17 ? n19811 : n19519;
  assign n19813 = pi16 ? n17063 : n19812;
  assign n19814 = pi15 ? n19808 : n19813;
  assign n19815 = pi14 ? n19805 : n19814;
  assign n19816 = pi20 ? n3083 : n139;
  assign n19817 = pi19 ? n37 : n19816;
  assign n19818 = pi18 ? n19817 : n6598;
  assign n19819 = pi17 ? n19818 : n19533;
  assign n19820 = pi16 ? n439 : n19819;
  assign n19821 = pi20 ? n3579 : n942;
  assign n19822 = pi19 ? n19821 : n139;
  assign n19823 = pi18 ? n37 : n19822;
  assign n19824 = pi20 ? n139 : n5552;
  assign n19825 = pi19 ? n19824 : n32;
  assign n19826 = pi18 ? n139 : n19825;
  assign n19827 = pi17 ? n19823 : n19826;
  assign n19828 = pi16 ? n439 : n19827;
  assign n19829 = pi15 ? n19820 : n19828;
  assign n19830 = pi18 ? n37 : n16056;
  assign n19831 = pi19 ? n16062 : n14045;
  assign n19832 = pi20 ? n14062 : n5552;
  assign n19833 = pi19 ? n19832 : n32;
  assign n19834 = pi18 ? n19831 : n19833;
  assign n19835 = pi17 ? n19830 : n19834;
  assign n19836 = pi16 ? n439 : n19835;
  assign n19837 = pi20 ? n37 : n13429;
  assign n19838 = pi19 ? n19837 : n32;
  assign n19839 = pi18 ? n37 : n19838;
  assign n19840 = pi17 ? n37 : n19839;
  assign n19841 = pi16 ? n439 : n19840;
  assign n19842 = pi15 ? n19836 : n19841;
  assign n19843 = pi14 ? n19829 : n19842;
  assign n19844 = pi13 ? n19815 : n19843;
  assign n19845 = pi12 ? n19804 : n19844;
  assign n19846 = pi20 ? n1912 : n1057;
  assign n19847 = pi19 ? n37 : n19846;
  assign n19848 = pi18 ? n37 : n19847;
  assign n19849 = pi20 ? n204 : n4749;
  assign n19850 = pi19 ? n19849 : n32;
  assign n19851 = pi18 ? n18100 : n19850;
  assign n19852 = pi17 ? n19848 : n19851;
  assign n19853 = pi16 ? n439 : n19852;
  assign n19854 = pi20 ? n13613 : n37;
  assign n19855 = pi19 ? n19854 : n37;
  assign n19856 = pi18 ? n37 : n19855;
  assign n19857 = pi21 ? n37 : n921;
  assign n19858 = pi20 ? n19857 : n204;
  assign n19859 = pi19 ? n19858 : n204;
  assign n19860 = pi18 ? n19859 : n19850;
  assign n19861 = pi17 ? n19856 : n19860;
  assign n19862 = pi16 ? n439 : n19861;
  assign n19863 = pi15 ? n19853 : n19862;
  assign n19864 = pi18 ? n18985 : n19850;
  assign n19865 = pi17 ? n37 : n19864;
  assign n19866 = pi16 ? n439 : n19865;
  assign n19867 = pi20 ? n37 : n14358;
  assign n19868 = pi19 ? n19867 : n204;
  assign n19869 = pi18 ? n19868 : n19850;
  assign n19870 = pi17 ? n37 : n19869;
  assign n19871 = pi16 ? n439 : n19870;
  assign n19872 = pi15 ? n19866 : n19871;
  assign n19873 = pi14 ? n19863 : n19872;
  assign n19874 = pi20 ? n335 : n6984;
  assign n19875 = pi19 ? n19874 : n32;
  assign n19876 = pi18 ? n15099 : n19875;
  assign n19877 = pi17 ? n37 : n19876;
  assign n19878 = pi16 ? n439 : n19877;
  assign n19879 = pi20 ? n335 : n4852;
  assign n19880 = pi19 ? n19879 : n32;
  assign n19881 = pi18 ? n16147 : n19880;
  assign n19882 = pi17 ? n37 : n19881;
  assign n19883 = pi16 ? n439 : n19882;
  assign n19884 = pi15 ? n19878 : n19883;
  assign n19885 = pi18 ? n16138 : n19880;
  assign n19886 = pi17 ? n37 : n19885;
  assign n19887 = pi16 ? n439 : n19886;
  assign n19888 = pi18 ? n9856 : n19880;
  assign n19889 = pi17 ? n37 : n19888;
  assign n19890 = pi16 ? n439 : n19889;
  assign n19891 = pi15 ? n19887 : n19890;
  assign n19892 = pi14 ? n19884 : n19891;
  assign n19893 = pi13 ? n19873 : n19892;
  assign n19894 = pi20 ? n605 : n4852;
  assign n19895 = pi19 ? n19894 : n32;
  assign n19896 = pi18 ? n10682 : n19895;
  assign n19897 = pi17 ? n37 : n19896;
  assign n19898 = pi16 ? n439 : n19897;
  assign n19899 = pi20 ? n3299 : n15446;
  assign n19900 = pi19 ? n19899 : n32;
  assign n19901 = pi18 ? n7677 : n19900;
  assign n19902 = pi17 ? n37 : n19901;
  assign n19903 = pi16 ? n439 : n19902;
  assign n19904 = pi15 ? n19898 : n19903;
  assign n19905 = pi20 ? n18162 : n5759;
  assign n19906 = pi19 ? n19905 : n32;
  assign n19907 = pi18 ? n17255 : n19906;
  assign n19908 = pi17 ? n37 : n19907;
  assign n19909 = pi16 ? n439 : n19908;
  assign n19910 = pi19 ? n37 : n6391;
  assign n19911 = pi20 ? n2091 : n6367;
  assign n19912 = pi19 ? n19911 : n32;
  assign n19913 = pi18 ? n19910 : n19912;
  assign n19914 = pi17 ? n37 : n19913;
  assign n19915 = pi16 ? n439 : n19914;
  assign n19916 = pi15 ? n19909 : n19915;
  assign n19917 = pi14 ? n19904 : n19916;
  assign n19918 = pi20 ? n37 : n19052;
  assign n19919 = pi19 ? n37 : n19918;
  assign n19920 = pi22 ? n673 : n233;
  assign n19921 = pi21 ? n19920 : n233;
  assign n19922 = pi20 ? n19921 : n6417;
  assign n19923 = pi19 ? n19922 : n32;
  assign n19924 = pi18 ? n19919 : n19923;
  assign n19925 = pi17 ? n37 : n19924;
  assign n19926 = pi16 ? n439 : n19925;
  assign n19927 = pi15 ? n19587 : n19926;
  assign n19928 = pi20 ? n2106 : n5830;
  assign n19929 = pi19 ? n19928 : n32;
  assign n19930 = pi18 ? n2724 : n19929;
  assign n19931 = pi17 ? n37 : n19930;
  assign n19932 = pi16 ? n439 : n19931;
  assign n19933 = pi22 ? n37 : n14245;
  assign n19934 = pi21 ? n37 : n19933;
  assign n19935 = pi20 ? n19934 : n5830;
  assign n19936 = pi19 ? n19935 : n32;
  assign n19937 = pi18 ? n2109 : n19936;
  assign n19938 = pi17 ? n37 : n19937;
  assign n19939 = pi16 ? n439 : n19938;
  assign n19940 = pi15 ? n19932 : n19939;
  assign n19941 = pi14 ? n19927 : n19940;
  assign n19942 = pi13 ? n19917 : n19941;
  assign n19943 = pi12 ? n19893 : n19942;
  assign n19944 = pi11 ? n19845 : n19943;
  assign n19945 = pi20 ? n685 : n2638;
  assign n19946 = pi19 ? n19945 : n32;
  assign n19947 = pi18 ? n16239 : n19946;
  assign n19948 = pi17 ? n37 : n19947;
  assign n19949 = pi16 ? n439 : n19948;
  assign n19950 = pi15 ? n19949 : n19600;
  assign n19951 = pi20 ? n37 : n5013;
  assign n19952 = pi19 ? n37 : n19951;
  assign n19953 = pi18 ? n19952 : n19603;
  assign n19954 = pi17 ? n37 : n19953;
  assign n19955 = pi16 ? n439 : n19954;
  assign n19956 = pi15 ? n19955 : n19611;
  assign n19957 = pi14 ? n19950 : n19956;
  assign n19958 = pi22 ? n685 : n37;
  assign n19959 = pi21 ? n37 : n19958;
  assign n19960 = pi20 ? n99 : n19959;
  assign n19961 = pi19 ? n99 : n19960;
  assign n19962 = pi18 ? n19961 : n19615;
  assign n19963 = pi17 ? n99 : n19962;
  assign n19964 = pi16 ? n201 : n19963;
  assign n19965 = pi15 ? n19964 : n19625;
  assign n19966 = pi18 ? n99 : n9985;
  assign n19967 = pi17 ? n19966 : n19628;
  assign n19968 = pi16 ? n744 : n19967;
  assign n19969 = pi15 ? n19625 : n19968;
  assign n19970 = pi14 ? n19965 : n19969;
  assign n19971 = pi13 ? n19957 : n19970;
  assign n19972 = pi20 ? n2999 : n99;
  assign n19973 = pi19 ? n2242 : n19972;
  assign n19974 = pi18 ? n19973 : n19135;
  assign n19975 = pi22 ? n2244 : n7780;
  assign n19976 = pi21 ? n685 : n19975;
  assign n19977 = pi20 ? n157 : n19976;
  assign n19978 = pi19 ? n12525 : n19977;
  assign n19979 = pi21 ? n685 : n6132;
  assign n19980 = pi20 ? n19979 : n1822;
  assign n19981 = pi19 ? n19980 : n32;
  assign n19982 = pi18 ? n19978 : n19981;
  assign n19983 = pi17 ? n19974 : n19982;
  assign n19984 = pi16 ? n744 : n19983;
  assign n19985 = pi19 ? n2243 : n15263;
  assign n19986 = pi18 ? n742 : n19985;
  assign n19987 = pi17 ? n32 : n19986;
  assign n19988 = pi20 ? n2243 : n9997;
  assign n19989 = pi19 ? n15264 : n19988;
  assign n19990 = pi19 ? n16311 : n157;
  assign n19991 = pi18 ? n19989 : n19990;
  assign n19992 = pi20 ? n19639 : n1822;
  assign n19993 = pi19 ? n19992 : n32;
  assign n19994 = pi18 ? n19152 : n19993;
  assign n19995 = pi17 ? n19991 : n19994;
  assign n19996 = pi16 ? n19987 : n19995;
  assign n19997 = pi15 ? n19984 : n19996;
  assign n19998 = pi22 ? n6890 : n157;
  assign n19999 = pi21 ? n19998 : n157;
  assign n20000 = pi20 ? n32 : n19999;
  assign n20001 = pi19 ? n32 : n20000;
  assign n20002 = pi18 ? n20001 : n157;
  assign n20003 = pi17 ? n32 : n20002;
  assign n20004 = pi24 ? n316 : n13481;
  assign n20005 = pi23 ? n157 : n20004;
  assign n20006 = pi22 ? n157 : n20005;
  assign n20007 = pi21 ? n99 : n20006;
  assign n20008 = pi20 ? n20007 : n32;
  assign n20009 = pi19 ? n20008 : n32;
  assign n20010 = pi18 ? n12526 : n20009;
  assign n20011 = pi17 ? n157 : n20010;
  assign n20012 = pi16 ? n20003 : n20011;
  assign n20013 = pi21 ? n157 : n6147;
  assign n20014 = pi20 ? n20013 : n32;
  assign n20015 = pi19 ? n20014 : n32;
  assign n20016 = pi18 ? n157 : n20015;
  assign n20017 = pi17 ? n157 : n20016;
  assign n20018 = pi16 ? n7419 : n20017;
  assign n20019 = pi15 ? n20012 : n20018;
  assign n20020 = pi14 ? n19997 : n20019;
  assign n20021 = pi20 ? n6582 : n32;
  assign n20022 = pi19 ? n20021 : n32;
  assign n20023 = pi18 ? n17368 : n20022;
  assign n20024 = pi17 ? n19189 : n20023;
  assign n20025 = pi16 ? n16349 : n20024;
  assign n20026 = pi23 ? n961 : n204;
  assign n20027 = pi22 ? n20026 : n204;
  assign n20028 = pi21 ? n20027 : n204;
  assign n20029 = pi20 ? n32 : n20028;
  assign n20030 = pi19 ? n32 : n20029;
  assign n20031 = pi18 ? n20030 : n204;
  assign n20032 = pi17 ? n32 : n20031;
  assign n20033 = pi20 ? n204 : n7909;
  assign n20034 = pi19 ? n204 : n20033;
  assign n20035 = pi18 ? n20034 : n20022;
  assign n20036 = pi17 ? n204 : n20035;
  assign n20037 = pi16 ? n20032 : n20036;
  assign n20038 = pi15 ? n20025 : n20037;
  assign n20039 = pi20 ? n204 : n3172;
  assign n20040 = pi19 ? n204 : n20039;
  assign n20041 = pi18 ? n204 : n20040;
  assign n20042 = pi21 ? n204 : n346;
  assign n20043 = pi20 ? n204 : n20042;
  assign n20044 = pi19 ? n20043 : n3727;
  assign n20045 = pi18 ? n20044 : n20022;
  assign n20046 = pi17 ? n20041 : n20045;
  assign n20047 = pi16 ? n19219 : n20046;
  assign n20048 = pi20 ? n204 : n9348;
  assign n20049 = pi19 ? n204 : n20048;
  assign n20050 = pi20 ? n204 : n347;
  assign n20051 = pi19 ? n204 : n20050;
  assign n20052 = pi18 ? n20049 : n20051;
  assign n20053 = pi19 ? n316 : n19231;
  assign n20054 = pi18 ? n20053 : n20022;
  assign n20055 = pi17 ? n20052 : n20054;
  assign n20056 = pi16 ? n11804 : n20055;
  assign n20057 = pi15 ? n20047 : n20056;
  assign n20058 = pi14 ? n20038 : n20057;
  assign n20059 = pi13 ? n20020 : n20058;
  assign n20060 = pi12 ? n19971 : n20059;
  assign n20061 = pi18 ? n139 : n10078;
  assign n20062 = pi19 ? n10892 : n999;
  assign n20063 = pi18 ? n20062 : n20022;
  assign n20064 = pi17 ? n20061 : n20063;
  assign n20065 = pi16 ? n915 : n20064;
  assign n20066 = pi19 ? n1787 : n15339;
  assign n20067 = pi18 ? n20066 : n9111;
  assign n20068 = pi21 ? n356 : n397;
  assign n20069 = pi20 ? n20068 : n32;
  assign n20070 = pi19 ? n20069 : n32;
  assign n20071 = pi18 ? n316 : n20070;
  assign n20072 = pi17 ? n20067 : n20071;
  assign n20073 = pi16 ? n915 : n20072;
  assign n20074 = pi15 ? n20065 : n20073;
  assign n20075 = pi21 ? n356 : n297;
  assign n20076 = pi20 ? n316 : n20075;
  assign n20077 = pi19 ? n316 : n20076;
  assign n20078 = pi18 ? n20077 : n316;
  assign n20079 = pi18 ? n316 : n12349;
  assign n20080 = pi17 ? n20078 : n20079;
  assign n20081 = pi16 ? n19257 : n20080;
  assign n20082 = pi19 ? n347 : n6208;
  assign n20083 = pi18 ? n913 : n20082;
  assign n20084 = pi17 ? n32 : n20083;
  assign n20085 = pi22 ? n139 : n2401;
  assign n20086 = pi21 ? n3617 : n20085;
  assign n20087 = pi20 ? n6208 : n20086;
  assign n20088 = pi21 ? n921 : n4429;
  assign n20089 = pi21 ? n1774 : n1785;
  assign n20090 = pi20 ? n20088 : n20089;
  assign n20091 = pi19 ? n20087 : n20090;
  assign n20092 = pi20 ? n350 : n5961;
  assign n20093 = pi21 ? n1785 : n346;
  assign n20094 = pi21 ? n3617 : n1018;
  assign n20095 = pi20 ? n20093 : n20094;
  assign n20096 = pi19 ? n20092 : n20095;
  assign n20097 = pi18 ? n20091 : n20096;
  assign n20098 = pi22 ? n204 : n1784;
  assign n20099 = pi21 ? n3990 : n20098;
  assign n20100 = pi20 ? n2427 : n20099;
  assign n20101 = pi21 ? n20085 : n1027;
  assign n20102 = pi22 ? n2299 : n204;
  assign n20103 = pi21 ? n20102 : n3617;
  assign n20104 = pi20 ? n20101 : n20103;
  assign n20105 = pi19 ? n20100 : n20104;
  assign n20106 = pi21 ? n204 : n5178;
  assign n20107 = pi20 ? n20106 : n32;
  assign n20108 = pi19 ? n20107 : n32;
  assign n20109 = pi18 ? n20105 : n20108;
  assign n20110 = pi17 ? n20097 : n20109;
  assign n20111 = pi16 ? n20084 : n20110;
  assign n20112 = pi15 ? n20081 : n20111;
  assign n20113 = pi14 ? n20074 : n20112;
  assign n20114 = pi21 ? n820 : n204;
  assign n20115 = pi19 ? n20114 : n15421;
  assign n20116 = pi18 ? n329 : n20115;
  assign n20117 = pi17 ? n32 : n20116;
  assign n20118 = pi20 ? n15421 : n204;
  assign n20119 = pi21 ? n204 : n457;
  assign n20120 = pi20 ? n204 : n20119;
  assign n20121 = pi19 ? n20118 : n20120;
  assign n20122 = pi19 ? n7633 : n18969;
  assign n20123 = pi18 ? n20121 : n20122;
  assign n20124 = pi20 ? n9187 : n32;
  assign n20125 = pi19 ? n20124 : n32;
  assign n20126 = pi18 ? n204 : n20125;
  assign n20127 = pi17 ? n20123 : n20126;
  assign n20128 = pi16 ? n20117 : n20127;
  assign n20129 = pi22 ? n2299 : n14363;
  assign n20130 = pi21 ? n204 : n20129;
  assign n20131 = pi20 ? n20130 : n32;
  assign n20132 = pi19 ? n20131 : n32;
  assign n20133 = pi18 ? n204 : n20132;
  assign n20134 = pi17 ? n204 : n20133;
  assign n20135 = pi16 ? n13493 : n20134;
  assign n20136 = pi15 ? n20128 : n20135;
  assign n20137 = pi20 ? n7969 : n32;
  assign n20138 = pi19 ? n20137 : n32;
  assign n20139 = pi18 ? n204 : n20138;
  assign n20140 = pi17 ? n204 : n20139;
  assign n20141 = pi16 ? n13846 : n20140;
  assign n20142 = pi21 ? n233 : n16358;
  assign n20143 = pi20 ? n20142 : n32;
  assign n20144 = pi19 ? n20143 : n32;
  assign n20145 = pi18 ? n19340 : n20144;
  assign n20146 = pi17 ? n233 : n20145;
  assign n20147 = pi16 ? n19336 : n20146;
  assign n20148 = pi15 ? n20141 : n20147;
  assign n20149 = pi14 ? n20136 : n20148;
  assign n20150 = pi13 ? n20113 : n20149;
  assign n20151 = pi18 ? n233 : n13341;
  assign n20152 = pi17 ? n19351 : n20151;
  assign n20153 = pi16 ? n439 : n20152;
  assign n20154 = pi17 ? n19360 : n20151;
  assign n20155 = pi16 ? n439 : n20154;
  assign n20156 = pi15 ? n20153 : n20155;
  assign n20157 = pi21 ? n37 : n4938;
  assign n20158 = pi20 ? n37 : n20157;
  assign n20159 = pi19 ? n20158 : n37;
  assign n20160 = pi18 ? n20159 : n10682;
  assign n20161 = pi21 ? n6376 : n2578;
  assign n20162 = pi20 ? n20161 : n32;
  assign n20163 = pi19 ? n20162 : n32;
  assign n20164 = pi18 ? n14411 : n20163;
  assign n20165 = pi17 ? n20160 : n20164;
  assign n20166 = pi16 ? n439 : n20165;
  assign n20167 = pi19 ? n577 : n642;
  assign n20168 = pi18 ? n374 : n20167;
  assign n20169 = pi17 ? n32 : n20168;
  assign n20170 = pi19 ? n335 : n17500;
  assign n20171 = pi18 ? n20170 : n335;
  assign n20172 = pi21 ? n19386 : n2637;
  assign n20173 = pi20 ? n20172 : n32;
  assign n20174 = pi19 ? n20173 : n32;
  assign n20175 = pi18 ? n335 : n20174;
  assign n20176 = pi17 ? n20171 : n20175;
  assign n20177 = pi16 ? n20169 : n20176;
  assign n20178 = pi15 ? n20166 : n20177;
  assign n20179 = pi14 ? n20156 : n20178;
  assign n20180 = pi21 ? n796 : n2746;
  assign n20181 = pi20 ? n32 : n20180;
  assign n20182 = pi19 ? n32 : n20181;
  assign n20183 = pi22 ? n2160 : n335;
  assign n20184 = pi21 ? n20183 : n335;
  assign n20185 = pi20 ? n20184 : n335;
  assign n20186 = pi22 ? n335 : n112;
  assign n20187 = pi21 ? n20186 : n1143;
  assign n20188 = pi22 ? n112 : n335;
  assign n20189 = pi21 ? n20186 : n20188;
  assign n20190 = pi20 ? n20187 : n20189;
  assign n20191 = pi19 ? n20185 : n20190;
  assign n20192 = pi18 ? n20182 : n20191;
  assign n20193 = pi17 ? n32 : n20192;
  assign n20194 = pi21 ? n20186 : n335;
  assign n20195 = pi20 ? n20194 : n335;
  assign n20196 = pi20 ? n335 : n14866;
  assign n20197 = pi19 ? n20195 : n20196;
  assign n20198 = pi18 ? n20197 : n12631;
  assign n20199 = pi21 ? n2707 : n928;
  assign n20200 = pi20 ? n20199 : n32;
  assign n20201 = pi19 ? n20200 : n32;
  assign n20202 = pi18 ? n14411 : n20201;
  assign n20203 = pi17 ? n20198 : n20202;
  assign n20204 = pi16 ? n20193 : n20203;
  assign n20205 = pi18 ? n335 : n12631;
  assign n20206 = pi19 ? n233 : n335;
  assign n20207 = pi21 ? n12635 : n2700;
  assign n20208 = pi20 ? n20207 : n32;
  assign n20209 = pi19 ? n20208 : n32;
  assign n20210 = pi18 ? n20206 : n20209;
  assign n20211 = pi17 ? n20205 : n20210;
  assign n20212 = pi16 ? n10980 : n20211;
  assign n20213 = pi15 ? n20204 : n20212;
  assign n20214 = pi22 ? n9827 : n139;
  assign n20215 = pi21 ? n20214 : n335;
  assign n20216 = pi21 ? n20214 : n18467;
  assign n20217 = pi20 ? n20215 : n20216;
  assign n20218 = pi22 ? n9827 : n335;
  assign n20219 = pi22 ? n9123 : n9827;
  assign n20220 = pi21 ? n20218 : n20219;
  assign n20221 = pi19 ? n20217 : n20220;
  assign n20222 = pi18 ? n12656 : n20221;
  assign n20223 = pi17 ? n32 : n20222;
  assign n20224 = pi21 ? n17548 : n363;
  assign n20225 = pi20 ? n20220 : n20224;
  assign n20226 = pi22 ? n18461 : n363;
  assign n20227 = pi21 ? n7986 : n20226;
  assign n20228 = pi22 ? n139 : n363;
  assign n20229 = pi21 ? n9836 : n20228;
  assign n20230 = pi20 ? n20227 : n20229;
  assign n20231 = pi19 ? n20225 : n20230;
  assign n20232 = pi22 ? n363 : n9123;
  assign n20233 = pi21 ? n18467 : n20232;
  assign n20234 = pi20 ? n18466 : n20233;
  assign n20235 = pi19 ? n20234 : n19423;
  assign n20236 = pi18 ? n20231 : n20235;
  assign n20237 = pi21 ? n18411 : n1009;
  assign n20238 = pi20 ? n20237 : n32;
  assign n20239 = pi19 ? n20238 : n32;
  assign n20240 = pi18 ? n233 : n20239;
  assign n20241 = pi17 ? n20236 : n20240;
  assign n20242 = pi16 ? n20223 : n20241;
  assign n20243 = pi18 ? n19433 : n233;
  assign n20244 = pi17 ? n32 : n20243;
  assign n20245 = pi17 ? n233 : n19426;
  assign n20246 = pi16 ? n20244 : n20245;
  assign n20247 = pi15 ? n20242 : n20246;
  assign n20248 = pi14 ? n20213 : n20247;
  assign n20249 = pi13 ? n20179 : n20248;
  assign n20250 = pi12 ? n20150 : n20249;
  assign n20251 = pi11 ? n20060 : n20250;
  assign n20252 = pi10 ? n19944 : n20251;
  assign n20253 = pi09 ? n19758 : n20252;
  assign n20254 = pi20 ? n37 : n7294;
  assign n20255 = pi19 ? n20254 : n32;
  assign n20256 = pi18 ? n37 : n20255;
  assign n20257 = pi17 ? n37 : n20256;
  assign n20258 = pi16 ? n11885 : n20257;
  assign n20259 = pi15 ? n32 : n20258;
  assign n20260 = pi16 ? n13561 : n19750;
  assign n20261 = pi15 ? n19751 : n20260;
  assign n20262 = pi14 ? n20259 : n20261;
  assign n20263 = pi13 ? n32 : n20262;
  assign n20264 = pi12 ? n32 : n20263;
  assign n20265 = pi11 ? n32 : n20264;
  assign n20266 = pi10 ? n32 : n20265;
  assign n20267 = pi21 ? n13049 : n32;
  assign n20268 = pi20 ? n37 : n20267;
  assign n20269 = pi19 ? n20268 : n32;
  assign n20270 = pi18 ? n37 : n20269;
  assign n20271 = pi17 ? n37 : n20270;
  assign n20272 = pi16 ? n17010 : n20271;
  assign n20273 = pi15 ? n19783 : n20272;
  assign n20274 = pi14 ? n19772 : n20273;
  assign n20275 = pi21 ? n13576 : n32;
  assign n20276 = pi20 ? n7745 : n20275;
  assign n20277 = pi19 ? n20276 : n32;
  assign n20278 = pi18 ? n37 : n20277;
  assign n20279 = pi17 ? n37 : n20278;
  assign n20280 = pi16 ? n439 : n20279;
  assign n20281 = pi15 ? n19799 : n20280;
  assign n20282 = pi20 ? n99 : n20275;
  assign n20283 = pi19 ? n20282 : n32;
  assign n20284 = pi18 ? n99 : n20283;
  assign n20285 = pi17 ? n99 : n20284;
  assign n20286 = pi16 ? n201 : n20285;
  assign n20287 = pi20 ? n99 : n6050;
  assign n20288 = pi19 ? n20287 : n32;
  assign n20289 = pi18 ? n99 : n20288;
  assign n20290 = pi17 ? n99 : n20289;
  assign n20291 = pi16 ? n801 : n20290;
  assign n20292 = pi15 ? n20286 : n20291;
  assign n20293 = pi14 ? n20281 : n20292;
  assign n20294 = pi13 ? n20274 : n20293;
  assign n20295 = pi20 ? n99 : n6060;
  assign n20296 = pi19 ? n20295 : n32;
  assign n20297 = pi18 ? n99 : n20296;
  assign n20298 = pi17 ? n99 : n20297;
  assign n20299 = pi16 ? n744 : n20298;
  assign n20300 = pi22 ? n139 : n6069;
  assign n20301 = pi21 ? n20300 : n32;
  assign n20302 = pi20 ? n139 : n20301;
  assign n20303 = pi19 ? n20302 : n32;
  assign n20304 = pi18 ? n139 : n20303;
  assign n20305 = pi17 ? n139 : n20304;
  assign n20306 = pi16 ? n19807 : n20305;
  assign n20307 = pi23 ? n139 : n687;
  assign n20308 = pi22 ? n139 : n20307;
  assign n20309 = pi21 ? n20308 : n32;
  assign n20310 = pi20 ? n139 : n20309;
  assign n20311 = pi19 ? n20310 : n32;
  assign n20312 = pi18 ? n139 : n20311;
  assign n20313 = pi17 ? n19811 : n20312;
  assign n20314 = pi16 ? n17063 : n20313;
  assign n20315 = pi15 ? n20306 : n20314;
  assign n20316 = pi14 ? n20299 : n20315;
  assign n20317 = pi23 ? n335 : n687;
  assign n20318 = pi22 ? n335 : n20317;
  assign n20319 = pi21 ? n20318 : n32;
  assign n20320 = pi20 ? n139 : n20319;
  assign n20321 = pi19 ? n20320 : n32;
  assign n20322 = pi18 ? n139 : n20321;
  assign n20323 = pi17 ? n19818 : n20322;
  assign n20324 = pi16 ? n439 : n20323;
  assign n20325 = pi15 ? n20324 : n19828;
  assign n20326 = pi14 ? n20325 : n19842;
  assign n20327 = pi13 ? n20316 : n20326;
  assign n20328 = pi12 ? n20294 : n20327;
  assign n20329 = pi20 ? n204 : n6271;
  assign n20330 = pi19 ? n20329 : n32;
  assign n20331 = pi18 ? n18100 : n20330;
  assign n20332 = pi17 ? n19848 : n20331;
  assign n20333 = pi16 ? n439 : n20332;
  assign n20334 = pi20 ? n204 : n10335;
  assign n20335 = pi19 ? n20334 : n32;
  assign n20336 = pi18 ? n19859 : n20335;
  assign n20337 = pi17 ? n19856 : n20336;
  assign n20338 = pi16 ? n439 : n20337;
  assign n20339 = pi15 ? n20333 : n20338;
  assign n20340 = pi23 ? n10750 : n32;
  assign n20341 = pi22 ? n204 : n20340;
  assign n20342 = pi21 ? n20341 : n32;
  assign n20343 = pi20 ? n204 : n20342;
  assign n20344 = pi19 ? n20343 : n32;
  assign n20345 = pi18 ? n18985 : n20344;
  assign n20346 = pi17 ? n37 : n20345;
  assign n20347 = pi16 ? n439 : n20346;
  assign n20348 = pi22 ? n204 : n2468;
  assign n20349 = pi21 ? n20348 : n32;
  assign n20350 = pi20 ? n204 : n20349;
  assign n20351 = pi19 ? n20350 : n32;
  assign n20352 = pi18 ? n19868 : n20351;
  assign n20353 = pi17 ? n37 : n20352;
  assign n20354 = pi16 ? n439 : n20353;
  assign n20355 = pi15 ? n20347 : n20354;
  assign n20356 = pi14 ? n20339 : n20355;
  assign n20357 = pi22 ? n2060 : n2468;
  assign n20358 = pi21 ? n20357 : n32;
  assign n20359 = pi20 ? n335 : n20358;
  assign n20360 = pi19 ? n20359 : n32;
  assign n20361 = pi18 ? n15099 : n20360;
  assign n20362 = pi17 ? n37 : n20361;
  assign n20363 = pi16 ? n439 : n20362;
  assign n20364 = pi20 ? n335 : n8947;
  assign n20365 = pi19 ? n20364 : n32;
  assign n20366 = pi18 ? n16147 : n20365;
  assign n20367 = pi17 ? n37 : n20366;
  assign n20368 = pi16 ? n439 : n20367;
  assign n20369 = pi15 ? n20363 : n20368;
  assign n20370 = pi18 ? n16138 : n20365;
  assign n20371 = pi17 ? n37 : n20370;
  assign n20372 = pi16 ? n439 : n20371;
  assign n20373 = pi15 ? n20372 : n19890;
  assign n20374 = pi14 ? n20369 : n20373;
  assign n20375 = pi13 ? n20356 : n20374;
  assign n20376 = pi22 ? n37 : n11889;
  assign n20377 = pi21 ? n37 : n20376;
  assign n20378 = pi20 ? n20377 : n4852;
  assign n20379 = pi19 ? n20378 : n32;
  assign n20380 = pi18 ? n7677 : n20379;
  assign n20381 = pi17 ? n37 : n20380;
  assign n20382 = pi16 ? n439 : n20381;
  assign n20383 = pi15 ? n19898 : n20382;
  assign n20384 = pi20 ? n18162 : n15446;
  assign n20385 = pi19 ? n20384 : n32;
  assign n20386 = pi18 ? n17255 : n20385;
  assign n20387 = pi17 ? n37 : n20386;
  assign n20388 = pi16 ? n439 : n20387;
  assign n20389 = pi15 ? n20388 : n19915;
  assign n20390 = pi14 ? n20383 : n20389;
  assign n20391 = pi21 ? n9202 : n32;
  assign n20392 = pi20 ? n233 : n20391;
  assign n20393 = pi19 ? n20392 : n32;
  assign n20394 = pi18 ? n16209 : n20393;
  assign n20395 = pi17 ? n37 : n20394;
  assign n20396 = pi16 ? n439 : n20395;
  assign n20397 = pi20 ? n19921 : n4110;
  assign n20398 = pi19 ? n20397 : n32;
  assign n20399 = pi18 ? n19919 : n20398;
  assign n20400 = pi17 ? n37 : n20399;
  assign n20401 = pi16 ? n439 : n20400;
  assign n20402 = pi15 ? n20396 : n20401;
  assign n20403 = pi20 ? n2106 : n4116;
  assign n20404 = pi19 ? n20403 : n32;
  assign n20405 = pi18 ? n2724 : n20404;
  assign n20406 = pi17 ? n37 : n20405;
  assign n20407 = pi16 ? n439 : n20406;
  assign n20408 = pi20 ? n19934 : n4116;
  assign n20409 = pi19 ? n20408 : n32;
  assign n20410 = pi18 ? n2109 : n20409;
  assign n20411 = pi17 ? n37 : n20410;
  assign n20412 = pi16 ? n439 : n20411;
  assign n20413 = pi15 ? n20407 : n20412;
  assign n20414 = pi14 ? n20402 : n20413;
  assign n20415 = pi13 ? n20390 : n20414;
  assign n20416 = pi12 ? n20375 : n20415;
  assign n20417 = pi11 ? n20328 : n20416;
  assign n20418 = pi20 ? n685 : n4116;
  assign n20419 = pi19 ? n20418 : n32;
  assign n20420 = pi18 ? n16239 : n20419;
  assign n20421 = pi17 ? n37 : n20420;
  assign n20422 = pi16 ? n439 : n20421;
  assign n20423 = pi20 ? n19084 : n4116;
  assign n20424 = pi19 ? n20423 : n32;
  assign n20425 = pi18 ? n2731 : n20424;
  assign n20426 = pi17 ? n37 : n20425;
  assign n20427 = pi16 ? n439 : n20426;
  assign n20428 = pi15 ? n20422 : n20427;
  assign n20429 = pi20 ? n18212 : n4116;
  assign n20430 = pi19 ? n20429 : n32;
  assign n20431 = pi18 ? n19952 : n20430;
  assign n20432 = pi17 ? n37 : n20431;
  assign n20433 = pi16 ? n439 : n20432;
  assign n20434 = pi20 ? n2107 : n4116;
  assign n20435 = pi19 ? n20434 : n32;
  assign n20436 = pi18 ? n37 : n20435;
  assign n20437 = pi17 ? n37 : n20436;
  assign n20438 = pi16 ? n439 : n20437;
  assign n20439 = pi15 ? n20433 : n20438;
  assign n20440 = pi14 ? n20428 : n20439;
  assign n20441 = pi20 ? n19109 : n4116;
  assign n20442 = pi19 ? n20441 : n32;
  assign n20443 = pi18 ? n19961 : n20442;
  assign n20444 = pi17 ? n99 : n20443;
  assign n20445 = pi16 ? n201 : n20444;
  assign n20446 = pi20 ? n5085 : n4116;
  assign n20447 = pi19 ? n20446 : n32;
  assign n20448 = pi18 ? n13377 : n20447;
  assign n20449 = pi17 ? n99 : n20448;
  assign n20450 = pi16 ? n721 : n20449;
  assign n20451 = pi15 ? n20445 : n20450;
  assign n20452 = pi20 ? n685 : n10011;
  assign n20453 = pi19 ? n20452 : n32;
  assign n20454 = pi18 ? n5087 : n20453;
  assign n20455 = pi17 ? n19966 : n20454;
  assign n20456 = pi16 ? n721 : n20455;
  assign n20457 = pi15 ? n20450 : n20456;
  assign n20458 = pi14 ? n20451 : n20457;
  assign n20459 = pi13 ? n20440 : n20458;
  assign n20460 = pi22 ? n157 : n2244;
  assign n20461 = pi21 ? n685 : n20460;
  assign n20462 = pi20 ? n20461 : n2653;
  assign n20463 = pi19 ? n20462 : n32;
  assign n20464 = pi18 ? n19978 : n20463;
  assign n20465 = pi17 ? n19974 : n20464;
  assign n20466 = pi16 ? n721 : n20465;
  assign n20467 = pi15 ? n20466 : n19996;
  assign n20468 = pi21 ? n99 : n6132;
  assign n20469 = pi20 ? n20468 : n32;
  assign n20470 = pi19 ? n20469 : n32;
  assign n20471 = pi18 ? n12526 : n20470;
  assign n20472 = pi17 ? n157 : n20471;
  assign n20473 = pi16 ? n19651 : n20472;
  assign n20474 = pi20 ? n7838 : n32;
  assign n20475 = pi19 ? n20474 : n32;
  assign n20476 = pi18 ? n157 : n20475;
  assign n20477 = pi17 ? n157 : n20476;
  assign n20478 = pi16 ? n5910 : n20477;
  assign n20479 = pi15 ? n20473 : n20478;
  assign n20480 = pi14 ? n20467 : n20479;
  assign n20481 = pi21 ? n316 : n8229;
  assign n20482 = pi20 ? n20481 : n32;
  assign n20483 = pi19 ? n20482 : n32;
  assign n20484 = pi18 ? n17368 : n20483;
  assign n20485 = pi17 ? n19189 : n20484;
  assign n20486 = pi16 ? n12535 : n20485;
  assign n20487 = pi16 ? n13493 : n20036;
  assign n20488 = pi15 ? n20486 : n20487;
  assign n20489 = pi20 ? n204 : n2365;
  assign n20490 = pi19 ? n204 : n20489;
  assign n20491 = pi18 ? n204 : n20490;
  assign n20492 = pi21 ? n316 : n1246;
  assign n20493 = pi20 ? n20492 : n32;
  assign n20494 = pi19 ? n20493 : n32;
  assign n20495 = pi18 ? n20044 : n20494;
  assign n20496 = pi17 ? n20491 : n20495;
  assign n20497 = pi16 ? n19219 : n20496;
  assign n20498 = pi15 ? n20497 : n20056;
  assign n20499 = pi14 ? n20488 : n20498;
  assign n20500 = pi13 ? n20480 : n20499;
  assign n20501 = pi12 ? n20459 : n20500;
  assign n20502 = pi18 ? n966 : n20082;
  assign n20503 = pi17 ? n32 : n20502;
  assign n20504 = pi21 ? n3617 : n1810;
  assign n20505 = pi20 ? n6208 : n20504;
  assign n20506 = pi21 ? n921 : n1529;
  assign n20507 = pi21 ? n820 : n1711;
  assign n20508 = pi20 ? n20506 : n20507;
  assign n20509 = pi19 ? n20505 : n20508;
  assign n20510 = pi19 ? n2540 : n20095;
  assign n20511 = pi18 ? n20509 : n20510;
  assign n20512 = pi22 ? n316 : n455;
  assign n20513 = pi21 ? n20512 : n1044;
  assign n20514 = pi20 ? n1578 : n20513;
  assign n20515 = pi21 ? n1810 : n1027;
  assign n20516 = pi21 ? n516 : n3617;
  assign n20517 = pi20 ? n20515 : n20516;
  assign n20518 = pi19 ? n20514 : n20517;
  assign n20519 = pi18 ? n20518 : n20108;
  assign n20520 = pi17 ? n20511 : n20519;
  assign n20521 = pi16 ? n20503 : n20520;
  assign n20522 = pi15 ? n20081 : n20521;
  assign n20523 = pi14 ? n20074 : n20522;
  assign n20524 = pi22 ? n3762 : n317;
  assign n20525 = pi21 ? n204 : n20524;
  assign n20526 = pi20 ? n20525 : n32;
  assign n20527 = pi19 ? n20526 : n32;
  assign n20528 = pi18 ? n204 : n20527;
  assign n20529 = pi17 ? n20123 : n20528;
  assign n20530 = pi16 ? n20117 : n20529;
  assign n20531 = pi21 ? n204 : n13465;
  assign n20532 = pi20 ? n20531 : n32;
  assign n20533 = pi19 ? n20532 : n32;
  assign n20534 = pi18 ? n204 : n20533;
  assign n20535 = pi17 ? n204 : n20534;
  assign n20536 = pi16 ? n13493 : n20535;
  assign n20537 = pi15 ? n20530 : n20536;
  assign n20538 = pi22 ? n233 : n448;
  assign n20539 = pi21 ? n233 : n20538;
  assign n20540 = pi20 ? n233 : n20539;
  assign n20541 = pi19 ? n20540 : n233;
  assign n20542 = pi18 ? n20541 : n20144;
  assign n20543 = pi17 ? n233 : n20542;
  assign n20544 = pi16 ? n19336 : n20543;
  assign n20545 = pi15 ? n20141 : n20544;
  assign n20546 = pi14 ? n20537 : n20545;
  assign n20547 = pi13 ? n20523 : n20546;
  assign n20548 = pi21 ? n233 : n3339;
  assign n20549 = pi20 ? n20548 : n32;
  assign n20550 = pi19 ? n20549 : n32;
  assign n20551 = pi18 ? n233 : n20550;
  assign n20552 = pi17 ? n19351 : n20551;
  assign n20553 = pi16 ? n439 : n20552;
  assign n20554 = pi15 ? n20553 : n20155;
  assign n20555 = pi21 ? n19386 : n4147;
  assign n20556 = pi20 ? n20555 : n32;
  assign n20557 = pi19 ? n20556 : n32;
  assign n20558 = pi18 ? n335 : n20557;
  assign n20559 = pi17 ? n20171 : n20558;
  assign n20560 = pi16 ? n20169 : n20559;
  assign n20561 = pi15 ? n20166 : n20560;
  assign n20562 = pi14 ? n20554 : n20561;
  assign n20563 = pi25 ? n36 : n32;
  assign n20564 = pi24 ? n32 : n20563;
  assign n20565 = pi23 ? n20564 : n99;
  assign n20566 = pi22 ? n20565 : n99;
  assign n20567 = pi21 ? n20566 : n99;
  assign n20568 = pi20 ? n32 : n20567;
  assign n20569 = pi19 ? n32 : n20568;
  assign n20570 = pi21 ? n14865 : n335;
  assign n20571 = pi20 ? n20570 : n335;
  assign n20572 = pi21 ? n3746 : n99;
  assign n20573 = pi21 ? n3746 : n14865;
  assign n20574 = pi20 ? n20572 : n20573;
  assign n20575 = pi19 ? n20571 : n20574;
  assign n20576 = pi18 ? n20569 : n20575;
  assign n20577 = pi17 ? n32 : n20576;
  assign n20578 = pi21 ? n3746 : n335;
  assign n20579 = pi20 ? n20578 : n335;
  assign n20580 = pi19 ? n20579 : n20196;
  assign n20581 = pi18 ? n20580 : n12631;
  assign n20582 = pi17 ? n20581 : n20202;
  assign n20583 = pi16 ? n20577 : n20582;
  assign n20584 = pi21 ? n12635 : n1009;
  assign n20585 = pi20 ? n20584 : n32;
  assign n20586 = pi19 ? n20585 : n32;
  assign n20587 = pi18 ? n20206 : n20586;
  assign n20588 = pi17 ? n20205 : n20587;
  assign n20589 = pi16 ? n10980 : n20588;
  assign n20590 = pi15 ? n20583 : n20589;
  assign n20591 = pi21 ? n139 : n18462;
  assign n20592 = pi21 ? n139 : n18467;
  assign n20593 = pi20 ? n20591 : n20592;
  assign n20594 = pi22 ? n364 : n335;
  assign n20595 = pi21 ? n20594 : n9828;
  assign n20596 = pi19 ? n20593 : n20595;
  assign n20597 = pi18 ? n12656 : n20596;
  assign n20598 = pi17 ? n32 : n20597;
  assign n20599 = pi20 ? n20595 : n20224;
  assign n20600 = pi22 ? n18795 : n363;
  assign n20601 = pi21 ? n7986 : n20600;
  assign n20602 = pi20 ? n20601 : n20229;
  assign n20603 = pi19 ? n20599 : n20602;
  assign n20604 = pi21 ? n18790 : n9143;
  assign n20605 = pi22 ? n363 : n139;
  assign n20606 = pi21 ? n18798 : n20605;
  assign n20607 = pi20 ? n20604 : n20606;
  assign n20608 = pi19 ? n20607 : n19423;
  assign n20609 = pi18 ? n20603 : n20608;
  assign n20610 = pi17 ? n20609 : n20240;
  assign n20611 = pi16 ? n20598 : n20610;
  assign n20612 = pi15 ? n20611 : n20246;
  assign n20613 = pi14 ? n20590 : n20612;
  assign n20614 = pi13 ? n20562 : n20613;
  assign n20615 = pi12 ? n20547 : n20614;
  assign n20616 = pi11 ? n20501 : n20615;
  assign n20617 = pi10 ? n20417 : n20616;
  assign n20618 = pi09 ? n20266 : n20617;
  assign n20619 = pi08 ? n20253 : n20618;
  assign n20620 = pi07 ? n19740 : n20619;
  assign n20621 = pi20 ? n37 : n6761;
  assign n20622 = pi19 ? n20621 : n32;
  assign n20623 = pi18 ? n37 : n20622;
  assign n20624 = pi17 ? n37 : n20623;
  assign n20625 = pi16 ? n12689 : n20624;
  assign n20626 = pi15 ? n32 : n20625;
  assign n20627 = pi24 ? n37 : n99;
  assign n20628 = pi23 ? n37 : n20627;
  assign n20629 = pi22 ? n37 : n20628;
  assign n20630 = pi21 ? n20629 : n32;
  assign n20631 = pi20 ? n37 : n20630;
  assign n20632 = pi19 ? n20631 : n32;
  assign n20633 = pi18 ? n37 : n20632;
  assign n20634 = pi17 ? n37 : n20633;
  assign n20635 = pi16 ? n12689 : n20634;
  assign n20636 = pi16 ? n13561 : n20634;
  assign n20637 = pi15 ? n20635 : n20636;
  assign n20638 = pi14 ? n20626 : n20637;
  assign n20639 = pi13 ? n32 : n20638;
  assign n20640 = pi12 ? n32 : n20639;
  assign n20641 = pi11 ? n32 : n20640;
  assign n20642 = pi10 ? n32 : n20641;
  assign n20643 = pi23 ? n37 : n3491;
  assign n20644 = pi22 ? n37 : n20643;
  assign n20645 = pi21 ? n20644 : n32;
  assign n20646 = pi20 ? n37 : n20645;
  assign n20647 = pi19 ? n20646 : n32;
  assign n20648 = pi18 ? n37 : n20647;
  assign n20649 = pi17 ? n37 : n20648;
  assign n20650 = pi16 ? n14445 : n20649;
  assign n20651 = pi20 ? n99 : n19760;
  assign n20652 = pi19 ? n20651 : n32;
  assign n20653 = pi18 ? n99 : n20652;
  assign n20654 = pi17 ? n99 : n20653;
  assign n20655 = pi16 ? n14857 : n20654;
  assign n20656 = pi15 ? n20650 : n20655;
  assign n20657 = pi20 ? n2973 : n37;
  assign n20658 = pi19 ? n20657 : n37;
  assign n20659 = pi18 ? n37 : n20658;
  assign n20660 = pi21 ? n218 : n2981;
  assign n20661 = pi20 ? n2974 : n20660;
  assign n20662 = pi20 ? n2982 : n37;
  assign n20663 = pi19 ? n20661 : n20662;
  assign n20664 = pi21 ? n2162 : n181;
  assign n20665 = pi22 ? n37 : n13918;
  assign n20666 = pi21 ? n20665 : n32;
  assign n20667 = pi20 ? n20664 : n20666;
  assign n20668 = pi19 ? n20667 : n32;
  assign n20669 = pi18 ? n20663 : n20668;
  assign n20670 = pi17 ? n20659 : n20669;
  assign n20671 = pi16 ? n16595 : n20670;
  assign n20672 = pi20 ? n14887 : n20666;
  assign n20673 = pi19 ? n20672 : n32;
  assign n20674 = pi18 ? n37 : n20673;
  assign n20675 = pi17 ? n37 : n20674;
  assign n20676 = pi16 ? n17010 : n20675;
  assign n20677 = pi15 ? n20671 : n20676;
  assign n20678 = pi14 ? n20656 : n20677;
  assign n20679 = pi22 ? n112 : n10510;
  assign n20680 = pi21 ? n20679 : n32;
  assign n20681 = pi20 ? n14887 : n20680;
  assign n20682 = pi19 ? n20681 : n32;
  assign n20683 = pi18 ? n37 : n20682;
  assign n20684 = pi17 ? n37 : n20683;
  assign n20685 = pi16 ? n439 : n20684;
  assign n20686 = pi22 ? n99 : n6027;
  assign n20687 = pi21 ? n20686 : n32;
  assign n20688 = pi20 ? n99 : n20687;
  assign n20689 = pi19 ? n20688 : n32;
  assign n20690 = pi18 ? n99 : n20689;
  assign n20691 = pi17 ? n99 : n20690;
  assign n20692 = pi16 ? n801 : n20691;
  assign n20693 = pi15 ? n20685 : n20692;
  assign n20694 = pi16 ? n721 : n20290;
  assign n20695 = pi15 ? n20291 : n20694;
  assign n20696 = pi14 ? n20693 : n20695;
  assign n20697 = pi13 ? n20678 : n20696;
  assign n20698 = pi16 ? n721 : n20298;
  assign n20699 = pi19 ? n1806 : n7867;
  assign n20700 = pi18 ? n1692 : n20699;
  assign n20701 = pi17 ? n32 : n20700;
  assign n20702 = pi20 ? n139 : n7502;
  assign n20703 = pi19 ? n20702 : n32;
  assign n20704 = pi18 ? n139 : n20703;
  assign n20705 = pi17 ? n139 : n20704;
  assign n20706 = pi16 ? n20701 : n20705;
  assign n20707 = pi15 ? n20698 : n20706;
  assign n20708 = pi20 ? n13612 : n3075;
  assign n20709 = pi20 ? n37 : n3656;
  assign n20710 = pi19 ? n20708 : n20709;
  assign n20711 = pi18 ? n8706 : n20710;
  assign n20712 = pi17 ? n32 : n20711;
  assign n20713 = pi16 ? n20712 : n20305;
  assign n20714 = pi20 ? n37 : n13612;
  assign n20715 = pi20 ? n5258 : n939;
  assign n20716 = pi19 ? n20714 : n20715;
  assign n20717 = pi18 ? n20716 : n139;
  assign n20718 = pi17 ? n20717 : n20312;
  assign n20719 = pi16 ? n439 : n20718;
  assign n20720 = pi15 ? n20713 : n20719;
  assign n20721 = pi14 ? n20707 : n20720;
  assign n20722 = pi20 ? n37 : n947;
  assign n20723 = pi19 ? n20722 : n139;
  assign n20724 = pi18 ? n37 : n20723;
  assign n20725 = pi17 ? n20724 : n20322;
  assign n20726 = pi16 ? n439 : n20725;
  assign n20727 = pi20 ? n3075 : n3645;
  assign n20728 = pi19 ? n20727 : n139;
  assign n20729 = pi21 ? n3436 : n32;
  assign n20730 = pi20 ? n139 : n20729;
  assign n20731 = pi19 ? n20730 : n32;
  assign n20732 = pi18 ? n20728 : n20731;
  assign n20733 = pi17 ? n19830 : n20732;
  assign n20734 = pi16 ? n439 : n20733;
  assign n20735 = pi15 ? n20726 : n20734;
  assign n20736 = pi22 ? n456 : n316;
  assign n20737 = pi21 ? n20736 : n32;
  assign n20738 = pi20 ? n37 : n20737;
  assign n20739 = pi19 ? n20738 : n32;
  assign n20740 = pi18 ? n37 : n20739;
  assign n20741 = pi17 ? n37 : n20740;
  assign n20742 = pi16 ? n439 : n20741;
  assign n20743 = pi20 ? n37 : n1912;
  assign n20744 = pi21 ? n1056 : n516;
  assign n20745 = pi20 ? n1912 : n20744;
  assign n20746 = pi19 ? n20743 : n20745;
  assign n20747 = pi18 ? n37 : n20746;
  assign n20748 = pi20 ? n1906 : n204;
  assign n20749 = pi19 ? n20748 : n204;
  assign n20750 = pi20 ? n204 : n7622;
  assign n20751 = pi19 ? n20750 : n32;
  assign n20752 = pi18 ? n20749 : n20751;
  assign n20753 = pi17 ? n20747 : n20752;
  assign n20754 = pi16 ? n439 : n20753;
  assign n20755 = pi15 ? n20742 : n20754;
  assign n20756 = pi14 ? n20735 : n20755;
  assign n20757 = pi13 ? n20721 : n20756;
  assign n20758 = pi12 ? n20697 : n20757;
  assign n20759 = pi20 ? n37 : n9354;
  assign n20760 = pi19 ? n37 : n20759;
  assign n20761 = pi18 ? n20760 : n37;
  assign n20762 = pi20 ? n37 : n20114;
  assign n20763 = pi19 ? n20762 : n204;
  assign n20764 = pi20 ? n204 : n6195;
  assign n20765 = pi19 ? n20764 : n32;
  assign n20766 = pi18 ? n20763 : n20765;
  assign n20767 = pi17 ? n20761 : n20766;
  assign n20768 = pi16 ? n439 : n20767;
  assign n20769 = pi21 ? n180 : n3073;
  assign n20770 = pi20 ? n32 : n20769;
  assign n20771 = pi19 ? n32 : n20770;
  assign n20772 = pi20 ? n13613 : n3932;
  assign n20773 = pi19 ? n37 : n20772;
  assign n20774 = pi18 ? n20771 : n20773;
  assign n20775 = pi17 ? n32 : n20774;
  assign n20776 = pi20 ? n9354 : n1003;
  assign n20777 = pi19 ? n9354 : n20776;
  assign n20778 = pi20 ? n939 : n297;
  assign n20779 = pi20 ? n8707 : n3090;
  assign n20780 = pi19 ? n20778 : n20779;
  assign n20781 = pi18 ? n20777 : n20780;
  assign n20782 = pi20 ? n820 : n139;
  assign n20783 = pi19 ? n20782 : n139;
  assign n20784 = pi20 ? n139 : n6185;
  assign n20785 = pi19 ? n20784 : n32;
  assign n20786 = pi18 ? n20783 : n20785;
  assign n20787 = pi17 ? n20781 : n20786;
  assign n20788 = pi16 ? n20775 : n20787;
  assign n20789 = pi15 ? n20768 : n20788;
  assign n20790 = pi21 ? n1936 : n1943;
  assign n20791 = pi20 ? n13300 : n20790;
  assign n20792 = pi19 ? n37 : n20791;
  assign n20793 = pi22 ? n335 : n2564;
  assign n20794 = pi21 ? n20793 : n32;
  assign n20795 = pi20 ? n4870 : n20794;
  assign n20796 = pi19 ? n20795 : n32;
  assign n20797 = pi18 ? n20792 : n20796;
  assign n20798 = pi17 ? n37 : n20797;
  assign n20799 = pi16 ? n439 : n20798;
  assign n20800 = pi22 ? n335 : n664;
  assign n20801 = pi21 ? n20800 : n32;
  assign n20802 = pi20 ? n335 : n20801;
  assign n20803 = pi19 ? n20802 : n32;
  assign n20804 = pi18 ? n9856 : n20803;
  assign n20805 = pi17 ? n37 : n20804;
  assign n20806 = pi16 ? n439 : n20805;
  assign n20807 = pi15 ? n20799 : n20806;
  assign n20808 = pi14 ? n20789 : n20807;
  assign n20809 = pi20 ? n3299 : n20157;
  assign n20810 = pi19 ? n20809 : n335;
  assign n20811 = pi18 ? n20810 : n20803;
  assign n20812 = pi17 ? n37 : n20811;
  assign n20813 = pi16 ? n439 : n20812;
  assign n20814 = pi18 ? n10682 : n20803;
  assign n20815 = pi17 ? n37 : n20814;
  assign n20816 = pi16 ? n439 : n20815;
  assign n20817 = pi15 ? n20813 : n20816;
  assign n20818 = pi19 ? n37 : n16516;
  assign n20819 = pi18 ? n20818 : n20803;
  assign n20820 = pi17 ? n37 : n20819;
  assign n20821 = pi16 ? n439 : n20820;
  assign n20822 = pi20 ? n335 : n9943;
  assign n20823 = pi19 ? n20822 : n32;
  assign n20824 = pi18 ? n10682 : n20823;
  assign n20825 = pi17 ? n37 : n20824;
  assign n20826 = pi16 ? n439 : n20825;
  assign n20827 = pi15 ? n20821 : n20826;
  assign n20828 = pi14 ? n20817 : n20827;
  assign n20829 = pi13 ? n20808 : n20828;
  assign n20830 = pi20 ? n638 : n335;
  assign n20831 = pi19 ? n37 : n20830;
  assign n20832 = pi20 ? n335 : n9957;
  assign n20833 = pi19 ? n20832 : n32;
  assign n20834 = pi18 ? n20831 : n20833;
  assign n20835 = pi17 ? n37 : n20834;
  assign n20836 = pi16 ? n439 : n20835;
  assign n20837 = pi20 ? n37 : n10335;
  assign n20838 = pi19 ? n20837 : n32;
  assign n20839 = pi18 ? n37 : n20838;
  assign n20840 = pi17 ? n37 : n20839;
  assign n20841 = pi16 ? n439 : n20840;
  assign n20842 = pi15 ? n20836 : n20841;
  assign n20843 = pi20 ? n233 : n8917;
  assign n20844 = pi19 ? n20843 : n32;
  assign n20845 = pi18 ? n16209 : n20844;
  assign n20846 = pi17 ? n37 : n20845;
  assign n20847 = pi16 ? n439 : n20846;
  assign n20848 = pi22 ? n4925 : n317;
  assign n20849 = pi21 ? n20848 : n32;
  assign n20850 = pi20 ? n233 : n20849;
  assign n20851 = pi19 ? n20850 : n32;
  assign n20852 = pi18 ? n16209 : n20851;
  assign n20853 = pi17 ? n37 : n20852;
  assign n20854 = pi16 ? n439 : n20853;
  assign n20855 = pi15 ? n20847 : n20854;
  assign n20856 = pi14 ? n20842 : n20855;
  assign n20857 = pi21 ? n5015 : n2707;
  assign n20858 = pi20 ? n37 : n20857;
  assign n20859 = pi19 ? n37 : n20858;
  assign n20860 = pi21 ? n2707 : n363;
  assign n20861 = pi20 ? n20860 : n9482;
  assign n20862 = pi19 ? n20861 : n32;
  assign n20863 = pi18 ? n20859 : n20862;
  assign n20864 = pi17 ? n37 : n20863;
  assign n20865 = pi16 ? n439 : n20864;
  assign n20866 = pi21 ? n2721 : n363;
  assign n20867 = pi20 ? n20866 : n14397;
  assign n20868 = pi19 ? n20867 : n32;
  assign n20869 = pi18 ? n2724 : n20868;
  assign n20870 = pi17 ? n37 : n20869;
  assign n20871 = pi16 ? n439 : n20870;
  assign n20872 = pi15 ? n20865 : n20871;
  assign n20873 = pi21 ? n2106 : n3392;
  assign n20874 = pi20 ? n20873 : n3210;
  assign n20875 = pi19 ? n20874 : n32;
  assign n20876 = pi18 ? n2724 : n20875;
  assign n20877 = pi17 ? n37 : n20876;
  assign n20878 = pi16 ? n439 : n20877;
  assign n20879 = pi20 ? n7730 : n4116;
  assign n20880 = pi19 ? n20879 : n32;
  assign n20881 = pi18 ? n2109 : n20880;
  assign n20882 = pi17 ? n37 : n20881;
  assign n20883 = pi16 ? n439 : n20882;
  assign n20884 = pi15 ? n20878 : n20883;
  assign n20885 = pi14 ? n20872 : n20884;
  assign n20886 = pi13 ? n20856 : n20885;
  assign n20887 = pi12 ? n20829 : n20886;
  assign n20888 = pi11 ? n20758 : n20887;
  assign n20889 = pi22 ? n16771 : n32;
  assign n20890 = pi21 ? n20889 : n32;
  assign n20891 = pi20 ? n363 : n20890;
  assign n20892 = pi19 ? n20891 : n32;
  assign n20893 = pi18 ? n7732 : n20892;
  assign n20894 = pi17 ? n37 : n20893;
  assign n20895 = pi16 ? n439 : n20894;
  assign n20896 = pi20 ? n363 : n4116;
  assign n20897 = pi19 ? n20896 : n32;
  assign n20898 = pi18 ? n19952 : n20897;
  assign n20899 = pi17 ? n37 : n20898;
  assign n20900 = pi16 ? n439 : n20899;
  assign n20901 = pi15 ? n20895 : n20900;
  assign n20902 = pi21 ? n1512 : n32;
  assign n20903 = pi20 ? n7730 : n20902;
  assign n20904 = pi19 ? n20903 : n32;
  assign n20905 = pi18 ? n37 : n20904;
  assign n20906 = pi17 ? n37 : n20905;
  assign n20907 = pi16 ? n439 : n20906;
  assign n20908 = pi15 ? n20907 : n20438;
  assign n20909 = pi14 ? n20901 : n20908;
  assign n20910 = pi18 ? n99 : n20447;
  assign n20911 = pi17 ? n99 : n20910;
  assign n20912 = pi16 ? n801 : n20911;
  assign n20913 = pi16 ? n744 : n20911;
  assign n20914 = pi15 ? n20912 : n20913;
  assign n20915 = pi20 ? n802 : n7754;
  assign n20916 = pi19 ? n20915 : n6091;
  assign n20917 = pi21 ? n6089 : n685;
  assign n20918 = pi20 ? n20917 : n5830;
  assign n20919 = pi19 ? n20918 : n32;
  assign n20920 = pi18 ? n20916 : n20919;
  assign n20921 = pi17 ? n99 : n20920;
  assign n20922 = pi16 ? n744 : n20921;
  assign n20923 = pi15 ? n20913 : n20922;
  assign n20924 = pi14 ? n20914 : n20923;
  assign n20925 = pi13 ? n20909 : n20924;
  assign n20926 = pi21 ? n5899 : n99;
  assign n20927 = pi20 ? n20926 : n99;
  assign n20928 = pi19 ? n99 : n20927;
  assign n20929 = pi18 ? n20928 : n10010;
  assign n20930 = pi21 ? n157 : n20460;
  assign n20931 = pi20 ? n20930 : n2653;
  assign n20932 = pi19 ? n20931 : n32;
  assign n20933 = pi18 ? n157 : n20932;
  assign n20934 = pi17 ? n20929 : n20933;
  assign n20935 = pi16 ? n744 : n20934;
  assign n20936 = pi20 ? n99 : n15263;
  assign n20937 = pi20 ? n7818 : n6500;
  assign n20938 = pi19 ? n20936 : n20937;
  assign n20939 = pi18 ? n742 : n20938;
  assign n20940 = pi17 ? n32 : n20939;
  assign n20941 = pi20 ? n157 : n10529;
  assign n20942 = pi19 ? n6500 : n20941;
  assign n20943 = pi19 ? n6524 : n6532;
  assign n20944 = pi18 ? n20942 : n20943;
  assign n20945 = pi21 ? n775 : n20460;
  assign n20946 = pi20 ? n20945 : n2653;
  assign n20947 = pi19 ? n20946 : n32;
  assign n20948 = pi18 ? n157 : n20947;
  assign n20949 = pi17 ? n20944 : n20948;
  assign n20950 = pi16 ? n20940 : n20949;
  assign n20951 = pi15 ? n20935 : n20950;
  assign n20952 = pi22 ? n14363 : n32;
  assign n20953 = pi21 ? n20952 : n32;
  assign n20954 = pi20 ? n7435 : n20953;
  assign n20955 = pi19 ? n20954 : n32;
  assign n20956 = pi18 ? n157 : n20955;
  assign n20957 = pi17 ? n157 : n20956;
  assign n20958 = pi16 ? n5910 : n20957;
  assign n20959 = pi20 ? n7435 : n32;
  assign n20960 = pi19 ? n20959 : n32;
  assign n20961 = pi18 ? n157 : n20960;
  assign n20962 = pi17 ? n157 : n20961;
  assign n20963 = pi16 ? n16338 : n20962;
  assign n20964 = pi15 ? n20958 : n20963;
  assign n20965 = pi14 ? n20951 : n20964;
  assign n20966 = pi21 ? n716 : n777;
  assign n20967 = pi20 ? n32 : n20966;
  assign n20968 = pi19 ? n32 : n20967;
  assign n20969 = pi19 ? n9715 : n14285;
  assign n20970 = pi18 ? n20968 : n20969;
  assign n20971 = pi17 ? n32 : n20970;
  assign n20972 = pi20 ? n6500 : n13948;
  assign n20973 = pi20 ? n13948 : n99;
  assign n20974 = pi19 ? n20972 : n20973;
  assign n20975 = pi18 ? n19124 : n20974;
  assign n20976 = pi19 ? n99 : n13944;
  assign n20977 = pi22 ? n99 : n316;
  assign n20978 = pi21 ? n20977 : n316;
  assign n20979 = pi20 ? n20978 : n32;
  assign n20980 = pi19 ? n20979 : n32;
  assign n20981 = pi18 ? n20976 : n20980;
  assign n20982 = pi17 ? n20975 : n20981;
  assign n20983 = pi16 ? n20971 : n20982;
  assign n20984 = pi21 ? n13441 : n204;
  assign n20985 = pi20 ? n32 : n20984;
  assign n20986 = pi19 ? n32 : n20985;
  assign n20987 = pi18 ? n20986 : n204;
  assign n20988 = pi17 ? n32 : n20987;
  assign n20989 = pi20 ? n1060 : n204;
  assign n20990 = pi19 ? n204 : n20989;
  assign n20991 = pi20 ? n7909 : n32;
  assign n20992 = pi19 ? n20991 : n32;
  assign n20993 = pi18 ? n20990 : n20992;
  assign n20994 = pi17 ? n204 : n20993;
  assign n20995 = pi16 ? n20988 : n20994;
  assign n20996 = pi15 ? n20983 : n20995;
  assign n20997 = pi22 ? n1519 : n204;
  assign n20998 = pi21 ? n20997 : n204;
  assign n20999 = pi20 ? n32 : n20998;
  assign n21000 = pi19 ? n32 : n20999;
  assign n21001 = pi18 ? n21000 : n204;
  assign n21002 = pi17 ? n32 : n21001;
  assign n21003 = pi20 ? n3731 : n7909;
  assign n21004 = pi19 ? n19231 : n21003;
  assign n21005 = pi20 ? n316 : n32;
  assign n21006 = pi19 ? n21005 : n32;
  assign n21007 = pi18 ? n21004 : n21006;
  assign n21008 = pi17 ? n204 : n21007;
  assign n21009 = pi16 ? n21002 : n21008;
  assign n21010 = pi19 ? n204 : n1064;
  assign n21011 = pi21 ? n1721 : n204;
  assign n21012 = pi20 ? n21011 : n204;
  assign n21013 = pi19 ? n21012 : n204;
  assign n21014 = pi18 ? n21010 : n21013;
  assign n21015 = pi20 ? n3731 : n316;
  assign n21016 = pi19 ? n19231 : n21015;
  assign n21017 = pi18 ? n21016 : n21006;
  assign n21018 = pi17 ? n21014 : n21017;
  assign n21019 = pi16 ? n13846 : n21018;
  assign n21020 = pi15 ? n21009 : n21019;
  assign n21021 = pi14 ? n20996 : n21020;
  assign n21022 = pi13 ? n20965 : n21021;
  assign n21023 = pi12 ? n20925 : n21022;
  assign n21024 = pi20 ? n356 : n316;
  assign n21025 = pi20 ? n356 : n975;
  assign n21026 = pi19 ? n21024 : n21025;
  assign n21027 = pi18 ? n21026 : n21006;
  assign n21028 = pi17 ? n139 : n21027;
  assign n21029 = pi16 ? n915 : n21028;
  assign n21030 = pi20 ? n6930 : n139;
  assign n21031 = pi19 ? n139 : n21030;
  assign n21032 = pi18 ? n21031 : n139;
  assign n21033 = pi18 ? n316 : n21006;
  assign n21034 = pi17 ? n21032 : n21033;
  assign n21035 = pi16 ? n915 : n21034;
  assign n21036 = pi15 ? n21029 : n21035;
  assign n21037 = pi21 ? n6609 : n139;
  assign n21038 = pi20 ? n32 : n21037;
  assign n21039 = pi19 ? n32 : n21038;
  assign n21040 = pi20 ? n139 : n1022;
  assign n21041 = pi19 ? n21040 : n16401;
  assign n21042 = pi18 ? n21039 : n21041;
  assign n21043 = pi17 ? n32 : n21042;
  assign n21044 = pi20 ? n1001 : n5317;
  assign n21045 = pi19 ? n975 : n21044;
  assign n21046 = pi20 ? n9082 : n347;
  assign n21047 = pi19 ? n21046 : n9066;
  assign n21048 = pi18 ? n21045 : n21047;
  assign n21049 = pi20 ? n316 : n356;
  assign n21050 = pi19 ? n10039 : n21049;
  assign n21051 = pi18 ? n21050 : n20070;
  assign n21052 = pi17 ? n21048 : n21051;
  assign n21053 = pi16 ? n21043 : n21052;
  assign n21054 = pi19 ? n139 : n6576;
  assign n21055 = pi18 ? n21054 : n1796;
  assign n21056 = pi17 ? n21055 : n20528;
  assign n21057 = pi16 ? n915 : n21056;
  assign n21058 = pi15 ? n21053 : n21057;
  assign n21059 = pi14 ? n21036 : n21058;
  assign n21060 = pi20 ? n139 : n2318;
  assign n21061 = pi20 ? n5204 : n6568;
  assign n21062 = pi19 ? n21060 : n21061;
  assign n21063 = pi18 ? n913 : n21062;
  assign n21064 = pi17 ? n32 : n21063;
  assign n21065 = pi20 ? n6158 : n204;
  assign n21066 = pi19 ? n6568 : n21065;
  assign n21067 = pi20 ? n2316 : n1016;
  assign n21068 = pi19 ? n21067 : n21065;
  assign n21069 = pi18 ? n21066 : n21068;
  assign n21070 = pi17 ? n21069 : n20528;
  assign n21071 = pi16 ? n21064 : n21070;
  assign n21072 = pi19 ? n7964 : n204;
  assign n21073 = pi18 ? n16488 : n21072;
  assign n21074 = pi17 ? n32 : n21073;
  assign n21075 = pi20 ? n3749 : n204;
  assign n21076 = pi19 ? n21075 : n204;
  assign n21077 = pi18 ? n204 : n21076;
  assign n21078 = pi23 ? n20004 : n32;
  assign n21079 = pi22 ? n705 : n21078;
  assign n21080 = pi21 ? n204 : n21079;
  assign n21081 = pi20 ? n21080 : n32;
  assign n21082 = pi19 ? n21081 : n32;
  assign n21083 = pi18 ? n204 : n21082;
  assign n21084 = pi17 ? n21077 : n21083;
  assign n21085 = pi16 ? n21074 : n21084;
  assign n21086 = pi15 ? n21071 : n21085;
  assign n21087 = pi18 ? n12968 : n21072;
  assign n21088 = pi17 ? n32 : n21087;
  assign n21089 = pi21 ? n204 : n19337;
  assign n21090 = pi20 ? n21089 : n3749;
  assign n21091 = pi21 ? n19337 : n204;
  assign n21092 = pi21 ? n11808 : n204;
  assign n21093 = pi20 ? n21091 : n21092;
  assign n21094 = pi19 ? n21090 : n21093;
  assign n21095 = pi21 ? n19337 : n13465;
  assign n21096 = pi20 ? n21095 : n32;
  assign n21097 = pi19 ? n21096 : n32;
  assign n21098 = pi18 ? n21094 : n21097;
  assign n21099 = pi17 ? n21077 : n21098;
  assign n21100 = pi16 ? n21088 : n21099;
  assign n21101 = pi21 ? n559 : n2091;
  assign n21102 = pi20 ? n21101 : n18431;
  assign n21103 = pi19 ? n21102 : n233;
  assign n21104 = pi18 ? n374 : n21103;
  assign n21105 = pi17 ? n32 : n21104;
  assign n21106 = pi19 ? n233 : n19416;
  assign n21107 = pi20 ? n16544 : n233;
  assign n21108 = pi19 ? n21107 : n233;
  assign n21109 = pi18 ? n21106 : n21108;
  assign n21110 = pi20 ? n233 : n16544;
  assign n21111 = pi19 ? n21110 : n233;
  assign n21112 = pi24 ? n233 : n13481;
  assign n21113 = pi23 ? n157 : n21112;
  assign n21114 = pi22 ? n21113 : n32;
  assign n21115 = pi21 ? n6376 : n21114;
  assign n21116 = pi20 ? n21115 : n32;
  assign n21117 = pi19 ? n21116 : n32;
  assign n21118 = pi18 ? n21111 : n21117;
  assign n21119 = pi17 ? n21109 : n21118;
  assign n21120 = pi16 ? n21105 : n21119;
  assign n21121 = pi15 ? n21100 : n21120;
  assign n21122 = pi14 ? n21086 : n21121;
  assign n21123 = pi13 ? n21059 : n21122;
  assign n21124 = pi21 ? n2048 : n37;
  assign n21125 = pi20 ? n21124 : n37;
  assign n21126 = pi19 ? n37 : n21125;
  assign n21127 = pi18 ? n374 : n21126;
  assign n21128 = pi17 ? n32 : n21127;
  assign n21129 = pi21 ? n4920 : n1920;
  assign n21130 = pi20 ? n21129 : n37;
  assign n21131 = pi19 ? n12476 : n21130;
  assign n21132 = pi20 ? n2092 : n561;
  assign n21133 = pi21 ? n2048 : n4893;
  assign n21134 = pi20 ? n21133 : n18431;
  assign n21135 = pi19 ? n21132 : n21134;
  assign n21136 = pi18 ? n21131 : n21135;
  assign n21137 = pi20 ? n7980 : n16544;
  assign n21138 = pi20 ? n13527 : n6362;
  assign n21139 = pi19 ? n21137 : n21138;
  assign n21140 = pi18 ? n21139 : n13745;
  assign n21141 = pi17 ? n21136 : n21140;
  assign n21142 = pi16 ? n21128 : n21141;
  assign n21143 = pi19 ? n37 : n7695;
  assign n21144 = pi18 ? n374 : n21143;
  assign n21145 = pi17 ? n32 : n21144;
  assign n21146 = pi20 ? n16530 : n21124;
  assign n21147 = pi19 ? n6355 : n21146;
  assign n21148 = pi21 ? n37 : n6376;
  assign n21149 = pi20 ? n2092 : n21148;
  assign n21150 = pi21 ? n2048 : n6376;
  assign n21151 = pi20 ? n21150 : n16544;
  assign n21152 = pi19 ? n21149 : n21151;
  assign n21153 = pi18 ? n21147 : n21152;
  assign n21154 = pi20 ? n233 : n13527;
  assign n21155 = pi19 ? n21154 : n233;
  assign n21156 = pi18 ? n21155 : n13745;
  assign n21157 = pi17 ? n21153 : n21156;
  assign n21158 = pi16 ? n21145 : n21157;
  assign n21159 = pi15 ? n21142 : n21158;
  assign n21160 = pi21 ? n6376 : n37;
  assign n21161 = pi20 ? n21160 : n21124;
  assign n21162 = pi19 ? n37 : n21161;
  assign n21163 = pi18 ? n21162 : n19910;
  assign n21164 = pi19 ? n233 : n21154;
  assign n21165 = pi18 ? n21164 : n13745;
  assign n21166 = pi17 ? n21163 : n21165;
  assign n21167 = pi16 ? n439 : n21166;
  assign n21168 = pi20 ? n37 : n575;
  assign n21169 = pi20 ? n568 : n638;
  assign n21170 = pi19 ? n21168 : n21169;
  assign n21171 = pi18 ? n374 : n21170;
  assign n21172 = pi17 ? n32 : n21171;
  assign n21173 = pi20 ? n638 : n647;
  assign n21174 = pi20 ? n604 : n647;
  assign n21175 = pi19 ? n21173 : n21174;
  assign n21176 = pi20 ? n610 : n577;
  assign n21177 = pi19 ? n21176 : n10681;
  assign n21178 = pi18 ? n21175 : n21177;
  assign n21179 = pi20 ? n15469 : n16544;
  assign n21180 = pi20 ? n7980 : n6376;
  assign n21181 = pi19 ? n21179 : n21180;
  assign n21182 = pi21 ? n233 : n6416;
  assign n21183 = pi20 ? n21182 : n32;
  assign n21184 = pi19 ? n21183 : n32;
  assign n21185 = pi18 ? n21181 : n21184;
  assign n21186 = pi17 ? n21178 : n21185;
  assign n21187 = pi16 ? n21172 : n21186;
  assign n21188 = pi15 ? n21167 : n21187;
  assign n21189 = pi14 ? n21159 : n21188;
  assign n21190 = pi18 ? n15459 : n15438;
  assign n21191 = pi20 ? n6362 : n6376;
  assign n21192 = pi19 ? n21110 : n21191;
  assign n21193 = pi21 ? n8860 : n5829;
  assign n21194 = pi20 ? n21193 : n32;
  assign n21195 = pi19 ? n21194 : n32;
  assign n21196 = pi18 ? n21192 : n21195;
  assign n21197 = pi17 ? n21190 : n21196;
  assign n21198 = pi16 ? n12648 : n21197;
  assign n21199 = pi21 ? n335 : n7986;
  assign n21200 = pi20 ? n335 : n21199;
  assign n21201 = pi22 ? n363 : n4899;
  assign n21202 = pi21 ? n21201 : n335;
  assign n21203 = pi20 ? n21202 : n335;
  assign n21204 = pi19 ? n21200 : n21203;
  assign n21205 = pi20 ? n335 : n18464;
  assign n21206 = pi20 ? n20224 : n233;
  assign n21207 = pi19 ? n21205 : n21206;
  assign n21208 = pi18 ? n21204 : n21207;
  assign n21209 = pi20 ? n18431 : n6376;
  assign n21210 = pi19 ? n233 : n21209;
  assign n21211 = pi21 ? n18411 : n928;
  assign n21212 = pi20 ? n21211 : n32;
  assign n21213 = pi19 ? n21212 : n32;
  assign n21214 = pi18 ? n21210 : n21213;
  assign n21215 = pi17 ? n21208 : n21214;
  assign n21216 = pi16 ? n10980 : n21215;
  assign n21217 = pi15 ? n21198 : n21216;
  assign n21218 = pi18 ? n19433 : n363;
  assign n21219 = pi17 ? n32 : n21218;
  assign n21220 = pi21 ? n363 : n5014;
  assign n21221 = pi20 ? n363 : n21220;
  assign n21222 = pi21 ? n233 : n363;
  assign n21223 = pi20 ? n21222 : n363;
  assign n21224 = pi19 ? n21221 : n21223;
  assign n21225 = pi20 ? n363 : n19422;
  assign n21226 = pi20 ? n5020 : n233;
  assign n21227 = pi19 ? n21225 : n21226;
  assign n21228 = pi18 ? n21224 : n21227;
  assign n21229 = pi21 ? n12659 : n928;
  assign n21230 = pi20 ? n21229 : n32;
  assign n21231 = pi19 ? n21230 : n32;
  assign n21232 = pi18 ? n233 : n21231;
  assign n21233 = pi17 ? n21228 : n21232;
  assign n21234 = pi16 ? n21219 : n21233;
  assign n21235 = pi22 ? n363 : n673;
  assign n21236 = pi21 ? n233 : n21235;
  assign n21237 = pi21 ? n2707 : n21235;
  assign n21238 = pi20 ? n21236 : n21237;
  assign n21239 = pi19 ? n19423 : n21238;
  assign n21240 = pi18 ? n19433 : n21239;
  assign n21241 = pi17 ? n32 : n21240;
  assign n21242 = pi20 ? n233 : n21222;
  assign n21243 = pi19 ? n233 : n21242;
  assign n21244 = pi18 ? n21243 : n233;
  assign n21245 = pi21 ? n12659 : n20952;
  assign n21246 = pi20 ? n21245 : n32;
  assign n21247 = pi19 ? n21246 : n32;
  assign n21248 = pi18 ? n233 : n21247;
  assign n21249 = pi17 ? n21244 : n21248;
  assign n21250 = pi16 ? n21241 : n21249;
  assign n21251 = pi15 ? n21234 : n21250;
  assign n21252 = pi14 ? n21217 : n21251;
  assign n21253 = pi13 ? n21189 : n21252;
  assign n21254 = pi12 ? n21123 : n21253;
  assign n21255 = pi11 ? n21023 : n21254;
  assign n21256 = pi10 ? n20888 : n21255;
  assign n21257 = pi09 ? n20642 : n21256;
  assign n21258 = pi21 ? n2957 : n32;
  assign n21259 = pi20 ? n37 : n21258;
  assign n21260 = pi19 ? n21259 : n32;
  assign n21261 = pi18 ? n37 : n21260;
  assign n21262 = pi17 ? n37 : n21261;
  assign n21263 = pi16 ? n12689 : n21262;
  assign n21264 = pi16 ? n13561 : n21262;
  assign n21265 = pi15 ? n21263 : n21264;
  assign n21266 = pi14 ? n20626 : n21265;
  assign n21267 = pi13 ? n32 : n21266;
  assign n21268 = pi12 ? n32 : n21267;
  assign n21269 = pi11 ? n32 : n21268;
  assign n21270 = pi10 ? n32 : n21269;
  assign n21271 = pi20 ? n37 : n8028;
  assign n21272 = pi19 ? n21271 : n32;
  assign n21273 = pi18 ? n37 : n21272;
  assign n21274 = pi17 ? n37 : n21273;
  assign n21275 = pi16 ? n14445 : n21274;
  assign n21276 = pi21 ? n1657 : n32;
  assign n21277 = pi20 ? n99 : n21276;
  assign n21278 = pi19 ? n21277 : n32;
  assign n21279 = pi18 ? n99 : n21278;
  assign n21280 = pi17 ? n99 : n21279;
  assign n21281 = pi16 ? n14857 : n21280;
  assign n21282 = pi15 ? n21275 : n21281;
  assign n21283 = pi14 ? n21282 : n20677;
  assign n21284 = pi21 ? n14477 : n32;
  assign n21285 = pi20 ? n99 : n21284;
  assign n21286 = pi19 ? n21285 : n32;
  assign n21287 = pi18 ? n99 : n21286;
  assign n21288 = pi17 ? n99 : n21287;
  assign n21289 = pi16 ? n801 : n21288;
  assign n21290 = pi15 ? n20685 : n21289;
  assign n21291 = pi20 ? n99 : n6815;
  assign n21292 = pi19 ? n21291 : n32;
  assign n21293 = pi18 ? n99 : n21292;
  assign n21294 = pi17 ? n99 : n21293;
  assign n21295 = pi16 ? n801 : n21294;
  assign n21296 = pi16 ? n744 : n21294;
  assign n21297 = pi15 ? n21295 : n21296;
  assign n21298 = pi14 ? n21290 : n21297;
  assign n21299 = pi13 ? n21283 : n21298;
  assign n21300 = pi20 ? n99 : n6824;
  assign n21301 = pi19 ? n21300 : n32;
  assign n21302 = pi18 ? n99 : n21301;
  assign n21303 = pi17 ? n99 : n21302;
  assign n21304 = pi16 ? n721 : n21303;
  assign n21305 = pi21 ? n14952 : n32;
  assign n21306 = pi20 ? n139 : n21305;
  assign n21307 = pi19 ? n21306 : n32;
  assign n21308 = pi18 ? n139 : n21307;
  assign n21309 = pi17 ? n139 : n21308;
  assign n21310 = pi16 ? n20701 : n21309;
  assign n21311 = pi15 ? n21304 : n21310;
  assign n21312 = pi21 ? n1564 : n1696;
  assign n21313 = pi20 ? n32 : n21312;
  assign n21314 = pi19 ? n32 : n21313;
  assign n21315 = pi20 ? n3606 : n1699;
  assign n21316 = pi19 ? n21315 : n20709;
  assign n21317 = pi18 ? n21314 : n21316;
  assign n21318 = pi17 ? n32 : n21317;
  assign n21319 = pi16 ? n21318 : n21309;
  assign n21320 = pi21 ? n14541 : n32;
  assign n21321 = pi20 ? n139 : n21320;
  assign n21322 = pi19 ? n21321 : n32;
  assign n21323 = pi18 ? n139 : n21322;
  assign n21324 = pi17 ? n20717 : n21323;
  assign n21325 = pi16 ? n439 : n21324;
  assign n21326 = pi15 ? n21319 : n21325;
  assign n21327 = pi14 ? n21311 : n21326;
  assign n21328 = pi20 ? n139 : n10262;
  assign n21329 = pi19 ? n21328 : n32;
  assign n21330 = pi18 ? n139 : n21329;
  assign n21331 = pi17 ? n20724 : n21330;
  assign n21332 = pi16 ? n439 : n21331;
  assign n21333 = pi15 ? n21332 : n20734;
  assign n21334 = pi14 ? n21333 : n20755;
  assign n21335 = pi13 ? n21327 : n21334;
  assign n21336 = pi12 ? n21299 : n21335;
  assign n21337 = pi22 ? n204 : n3301;
  assign n21338 = pi21 ? n21337 : n32;
  assign n21339 = pi20 ? n204 : n21338;
  assign n21340 = pi19 ? n21339 : n32;
  assign n21341 = pi18 ? n20763 : n21340;
  assign n21342 = pi17 ? n20761 : n21341;
  assign n21343 = pi16 ? n439 : n21342;
  assign n21344 = pi22 ? n139 : n3318;
  assign n21345 = pi21 ? n21344 : n32;
  assign n21346 = pi20 ? n139 : n21345;
  assign n21347 = pi19 ? n21346 : n32;
  assign n21348 = pi18 ? n20783 : n21347;
  assign n21349 = pi17 ? n20781 : n21348;
  assign n21350 = pi16 ? n20775 : n21349;
  assign n21351 = pi15 ? n21343 : n21350;
  assign n21352 = pi21 ? n1936 : n335;
  assign n21353 = pi20 ? n7591 : n21352;
  assign n21354 = pi19 ? n37 : n21353;
  assign n21355 = pi22 ? n335 : n430;
  assign n21356 = pi21 ? n21355 : n32;
  assign n21357 = pi20 ? n6724 : n21356;
  assign n21358 = pi19 ? n21357 : n32;
  assign n21359 = pi18 ? n21354 : n21358;
  assign n21360 = pi17 ? n37 : n21359;
  assign n21361 = pi16 ? n439 : n21360;
  assign n21362 = pi15 ? n21361 : n20806;
  assign n21363 = pi14 ? n21351 : n21362;
  assign n21364 = pi13 ? n21363 : n20828;
  assign n21365 = pi14 ? n20842 : n20847;
  assign n21366 = pi20 ? n20860 : n9963;
  assign n21367 = pi19 ? n21366 : n32;
  assign n21368 = pi18 ? n20859 : n21367;
  assign n21369 = pi17 ? n37 : n21368;
  assign n21370 = pi16 ? n439 : n21369;
  assign n21371 = pi20 ? n20866 : n7042;
  assign n21372 = pi19 ? n21371 : n32;
  assign n21373 = pi18 ? n2724 : n21372;
  assign n21374 = pi17 ? n37 : n21373;
  assign n21375 = pi16 ? n439 : n21374;
  assign n21376 = pi15 ? n21370 : n21375;
  assign n21377 = pi20 ? n7730 : n7724;
  assign n21378 = pi19 ? n21377 : n32;
  assign n21379 = pi18 ? n2109 : n21378;
  assign n21380 = pi17 ? n37 : n21379;
  assign n21381 = pi16 ? n439 : n21380;
  assign n21382 = pi15 ? n20878 : n21381;
  assign n21383 = pi14 ? n21376 : n21382;
  assign n21384 = pi13 ? n21365 : n21383;
  assign n21385 = pi12 ? n21364 : n21384;
  assign n21386 = pi11 ? n21336 : n21385;
  assign n21387 = pi22 ? n686 : n32;
  assign n21388 = pi21 ? n21387 : n32;
  assign n21389 = pi20 ? n363 : n21388;
  assign n21390 = pi19 ? n21389 : n32;
  assign n21391 = pi18 ? n7732 : n21390;
  assign n21392 = pi17 ? n37 : n21391;
  assign n21393 = pi16 ? n439 : n21392;
  assign n21394 = pi20 ? n363 : n7724;
  assign n21395 = pi19 ? n21394 : n32;
  assign n21396 = pi18 ? n19952 : n21395;
  assign n21397 = pi17 ? n37 : n21396;
  assign n21398 = pi16 ? n439 : n21397;
  assign n21399 = pi15 ? n21393 : n21398;
  assign n21400 = pi20 ? n7730 : n8967;
  assign n21401 = pi19 ? n21400 : n32;
  assign n21402 = pi18 ? n37 : n21401;
  assign n21403 = pi17 ? n37 : n21402;
  assign n21404 = pi16 ? n439 : n21403;
  assign n21405 = pi20 ? n2107 : n7724;
  assign n21406 = pi19 ? n21405 : n32;
  assign n21407 = pi18 ? n37 : n21406;
  assign n21408 = pi17 ? n37 : n21407;
  assign n21409 = pi16 ? n439 : n21408;
  assign n21410 = pi15 ? n21404 : n21409;
  assign n21411 = pi14 ? n21399 : n21410;
  assign n21412 = pi20 ? n5085 : n7724;
  assign n21413 = pi19 ? n21412 : n32;
  assign n21414 = pi18 ? n99 : n21413;
  assign n21415 = pi17 ? n99 : n21414;
  assign n21416 = pi16 ? n801 : n21415;
  assign n21417 = pi16 ? n721 : n21415;
  assign n21418 = pi15 ? n21416 : n21417;
  assign n21419 = pi20 ? n20917 : n7049;
  assign n21420 = pi19 ? n21419 : n32;
  assign n21421 = pi18 ? n20916 : n21420;
  assign n21422 = pi17 ? n99 : n21421;
  assign n21423 = pi16 ? n721 : n21422;
  assign n21424 = pi15 ? n21417 : n21423;
  assign n21425 = pi14 ? n21418 : n21424;
  assign n21426 = pi13 ? n21411 : n21425;
  assign n21427 = pi20 ? n157 : n10011;
  assign n21428 = pi19 ? n21427 : n32;
  assign n21429 = pi18 ? n157 : n21428;
  assign n21430 = pi17 ? n20929 : n21429;
  assign n21431 = pi16 ? n721 : n21430;
  assign n21432 = pi18 ? n719 : n20938;
  assign n21433 = pi17 ? n32 : n21432;
  assign n21434 = pi20 ? n6523 : n2653;
  assign n21435 = pi19 ? n21434 : n32;
  assign n21436 = pi18 ? n157 : n21435;
  assign n21437 = pi17 ? n20944 : n21436;
  assign n21438 = pi16 ? n21433 : n21437;
  assign n21439 = pi15 ? n21431 : n21438;
  assign n21440 = pi20 ? n7435 : n1822;
  assign n21441 = pi19 ? n21440 : n32;
  assign n21442 = pi18 ? n157 : n21441;
  assign n21443 = pi17 ? n157 : n21442;
  assign n21444 = pi16 ? n5910 : n21443;
  assign n21445 = pi16 ? n12535 : n21443;
  assign n21446 = pi15 ? n21444 : n21445;
  assign n21447 = pi14 ? n21439 : n21446;
  assign n21448 = pi21 ? n739 : n777;
  assign n21449 = pi20 ? n32 : n21448;
  assign n21450 = pi19 ? n32 : n21449;
  assign n21451 = pi18 ? n21450 : n20969;
  assign n21452 = pi17 ? n32 : n21451;
  assign n21453 = pi16 ? n21452 : n20982;
  assign n21454 = pi16 ? n19219 : n20994;
  assign n21455 = pi15 ? n21453 : n21454;
  assign n21456 = pi16 ? n13846 : n21008;
  assign n21457 = pi15 ? n21456 : n21019;
  assign n21458 = pi14 ? n21455 : n21457;
  assign n21459 = pi13 ? n21447 : n21458;
  assign n21460 = pi12 ? n21426 : n21459;
  assign n21461 = pi21 ? n4017 : n356;
  assign n21462 = pi20 ? n21461 : n316;
  assign n21463 = pi19 ? n21462 : n21025;
  assign n21464 = pi18 ? n21463 : n21006;
  assign n21465 = pi17 ? n139 : n21464;
  assign n21466 = pi16 ? n915 : n21465;
  assign n21467 = pi15 ? n21466 : n21035;
  assign n21468 = pi21 ? n356 : n7137;
  assign n21469 = pi20 ? n21468 : n32;
  assign n21470 = pi19 ? n21469 : n32;
  assign n21471 = pi18 ? n21050 : n21470;
  assign n21472 = pi17 ? n21048 : n21471;
  assign n21473 = pi16 ? n21043 : n21472;
  assign n21474 = pi21 ? n204 : n491;
  assign n21475 = pi20 ? n21474 : n32;
  assign n21476 = pi19 ? n21475 : n32;
  assign n21477 = pi18 ? n204 : n21476;
  assign n21478 = pi17 ? n21055 : n21477;
  assign n21479 = pi16 ? n915 : n21478;
  assign n21480 = pi15 ? n21473 : n21479;
  assign n21481 = pi14 ? n21467 : n21480;
  assign n21482 = pi21 ? n4339 : n139;
  assign n21483 = pi20 ? n32 : n21482;
  assign n21484 = pi19 ? n32 : n21483;
  assign n21485 = pi18 ? n21484 : n21062;
  assign n21486 = pi17 ? n32 : n21485;
  assign n21487 = pi22 ? n4883 : n396;
  assign n21488 = pi21 ? n204 : n21487;
  assign n21489 = pi20 ? n21488 : n32;
  assign n21490 = pi19 ? n21489 : n32;
  assign n21491 = pi18 ? n204 : n21490;
  assign n21492 = pi17 ? n21069 : n21491;
  assign n21493 = pi16 ? n21486 : n21492;
  assign n21494 = pi23 ? n3719 : n204;
  assign n21495 = pi22 ? n21494 : n335;
  assign n21496 = pi21 ? n21495 : n204;
  assign n21497 = pi20 ? n32 : n21496;
  assign n21498 = pi19 ? n32 : n21497;
  assign n21499 = pi18 ? n21498 : n21072;
  assign n21500 = pi17 ? n32 : n21499;
  assign n21501 = pi23 ? n363 : n1598;
  assign n21502 = pi23 ? n13481 : n32;
  assign n21503 = pi22 ? n21501 : n21502;
  assign n21504 = pi21 ? n204 : n21503;
  assign n21505 = pi20 ? n21504 : n32;
  assign n21506 = pi19 ? n21505 : n32;
  assign n21507 = pi18 ? n204 : n21506;
  assign n21508 = pi17 ? n21077 : n21507;
  assign n21509 = pi16 ? n21500 : n21508;
  assign n21510 = pi15 ? n21493 : n21509;
  assign n21511 = pi23 ? n204 : n1598;
  assign n21512 = pi22 ? n21511 : n706;
  assign n21513 = pi21 ? n19337 : n21512;
  assign n21514 = pi20 ? n21513 : n32;
  assign n21515 = pi19 ? n21514 : n32;
  assign n21516 = pi18 ? n21094 : n21515;
  assign n21517 = pi17 ? n21077 : n21516;
  assign n21518 = pi16 ? n21088 : n21517;
  assign n21519 = pi23 ? n157 : n2120;
  assign n21520 = pi22 ? n21519 : n32;
  assign n21521 = pi21 ? n6376 : n21520;
  assign n21522 = pi20 ? n21521 : n32;
  assign n21523 = pi19 ? n21522 : n32;
  assign n21524 = pi18 ? n21111 : n21523;
  assign n21525 = pi17 ? n21109 : n21524;
  assign n21526 = pi16 ? n21105 : n21525;
  assign n21527 = pi15 ? n21518 : n21526;
  assign n21528 = pi14 ? n21510 : n21527;
  assign n21529 = pi13 ? n21481 : n21528;
  assign n21530 = pi21 ? n233 : n12825;
  assign n21531 = pi20 ? n21530 : n32;
  assign n21532 = pi19 ? n21531 : n32;
  assign n21533 = pi18 ? n21139 : n21532;
  assign n21534 = pi17 ? n21136 : n21533;
  assign n21535 = pi16 ? n21128 : n21534;
  assign n21536 = pi15 ? n21535 : n21158;
  assign n21537 = pi23 ? n4145 : n687;
  assign n21538 = pi22 ? n21537 : n32;
  assign n21539 = pi21 ? n233 : n21538;
  assign n21540 = pi20 ? n21539 : n32;
  assign n21541 = pi19 ? n21540 : n32;
  assign n21542 = pi18 ? n21181 : n21541;
  assign n21543 = pi17 ? n21178 : n21542;
  assign n21544 = pi16 ? n21172 : n21543;
  assign n21545 = pi15 ? n21167 : n21544;
  assign n21546 = pi14 ? n21536 : n21545;
  assign n21547 = pi21 ? n18411 : n5370;
  assign n21548 = pi20 ? n21547 : n32;
  assign n21549 = pi19 ? n21548 : n32;
  assign n21550 = pi18 ? n21210 : n21549;
  assign n21551 = pi17 ? n21208 : n21550;
  assign n21552 = pi16 ? n2425 : n21551;
  assign n21553 = pi15 ? n21198 : n21552;
  assign n21554 = pi24 ? n32 : n363;
  assign n21555 = pi23 ? n21554 : n363;
  assign n21556 = pi22 ? n21555 : n363;
  assign n21557 = pi21 ? n21556 : n363;
  assign n21558 = pi20 ? n32 : n21557;
  assign n21559 = pi19 ? n32 : n21558;
  assign n21560 = pi18 ? n21559 : n363;
  assign n21561 = pi17 ? n32 : n21560;
  assign n21562 = pi16 ? n21561 : n21233;
  assign n21563 = pi18 ? n21559 : n21239;
  assign n21564 = pi17 ? n32 : n21563;
  assign n21565 = pi21 ? n12659 : n1009;
  assign n21566 = pi20 ? n21565 : n32;
  assign n21567 = pi19 ? n21566 : n32;
  assign n21568 = pi18 ? n233 : n21567;
  assign n21569 = pi17 ? n21244 : n21568;
  assign n21570 = pi16 ? n21564 : n21569;
  assign n21571 = pi15 ? n21562 : n21570;
  assign n21572 = pi14 ? n21553 : n21571;
  assign n21573 = pi13 ? n21546 : n21572;
  assign n21574 = pi12 ? n21529 : n21573;
  assign n21575 = pi11 ? n21460 : n21574;
  assign n21576 = pi10 ? n21386 : n21575;
  assign n21577 = pi09 ? n21270 : n21576;
  assign n21578 = pi08 ? n21257 : n21577;
  assign n21579 = pi20 ? n37 : n7282;
  assign n21580 = pi19 ? n21579 : n32;
  assign n21581 = pi18 ? n37 : n21580;
  assign n21582 = pi17 ? n37 : n21581;
  assign n21583 = pi16 ? n12689 : n21582;
  assign n21584 = pi15 ? n32 : n21583;
  assign n21585 = pi21 ? n37 : n8008;
  assign n21586 = pi20 ? n37 : n21585;
  assign n21587 = pi19 ? n21586 : n32;
  assign n21588 = pi18 ? n37 : n21587;
  assign n21589 = pi17 ? n37 : n21588;
  assign n21590 = pi16 ? n13561 : n21589;
  assign n21591 = pi20 ? n37 : n8009;
  assign n21592 = pi19 ? n21591 : n32;
  assign n21593 = pi18 ? n37 : n21592;
  assign n21594 = pi17 ? n37 : n21593;
  assign n21595 = pi16 ? n13561 : n21594;
  assign n21596 = pi15 ? n21590 : n21595;
  assign n21597 = pi14 ? n21584 : n21596;
  assign n21598 = pi13 ? n32 : n21597;
  assign n21599 = pi12 ? n32 : n21598;
  assign n21600 = pi11 ? n32 : n21599;
  assign n21601 = pi10 ? n32 : n21600;
  assign n21602 = pi21 ? n3073 : n8015;
  assign n21603 = pi20 ? n37 : n21602;
  assign n21604 = pi19 ? n21603 : n32;
  assign n21605 = pi18 ? n37 : n21604;
  assign n21606 = pi17 ? n37 : n21605;
  assign n21607 = pi16 ? n14445 : n21606;
  assign n21608 = pi21 ? n3779 : n218;
  assign n21609 = pi20 ? n32 : n21608;
  assign n21610 = pi19 ? n32 : n21609;
  assign n21611 = pi20 ? n14844 : n99;
  assign n21612 = pi19 ? n21611 : n99;
  assign n21613 = pi18 ? n21610 : n21612;
  assign n21614 = pi17 ? n32 : n21613;
  assign n21615 = pi21 ? n746 : n8557;
  assign n21616 = pi20 ? n99 : n21615;
  assign n21617 = pi19 ? n21616 : n32;
  assign n21618 = pi18 ? n99 : n21617;
  assign n21619 = pi17 ? n99 : n21618;
  assign n21620 = pi16 ? n21614 : n21619;
  assign n21621 = pi15 ? n21607 : n21620;
  assign n21622 = pi22 ? n37 : n1656;
  assign n21623 = pi21 ? n21622 : n32;
  assign n21624 = pi20 ? n37 : n21623;
  assign n21625 = pi19 ? n21624 : n32;
  assign n21626 = pi18 ? n37 : n21625;
  assign n21627 = pi17 ? n37 : n21626;
  assign n21628 = pi16 ? n16595 : n21627;
  assign n21629 = pi20 ? n5077 : n3814;
  assign n21630 = pi19 ? n37 : n21629;
  assign n21631 = pi18 ? n17008 : n21630;
  assign n21632 = pi17 ? n32 : n21631;
  assign n21633 = pi21 ? n2164 : n2156;
  assign n21634 = pi20 ? n21633 : n6044;
  assign n21635 = pi21 ? n37 : n2957;
  assign n21636 = pi20 ? n21635 : n3038;
  assign n21637 = pi19 ? n21634 : n21636;
  assign n21638 = pi21 ? n181 : n2156;
  assign n21639 = pi20 ? n21638 : n37;
  assign n21640 = pi20 ? n2176 : n3824;
  assign n21641 = pi19 ? n21639 : n21640;
  assign n21642 = pi18 ? n21637 : n21641;
  assign n21643 = pi21 ? n2164 : n37;
  assign n21644 = pi20 ? n21638 : n21643;
  assign n21645 = pi19 ? n21644 : n2185;
  assign n21646 = pi20 ? n218 : n21623;
  assign n21647 = pi19 ? n21646 : n32;
  assign n21648 = pi18 ? n21645 : n21647;
  assign n21649 = pi17 ? n21642 : n21648;
  assign n21650 = pi16 ? n21632 : n21649;
  assign n21651 = pi15 ? n21628 : n21650;
  assign n21652 = pi14 ? n21621 : n21651;
  assign n21653 = pi22 ? n37 : n4537;
  assign n21654 = pi21 ? n21653 : n32;
  assign n21655 = pi20 ? n14887 : n21654;
  assign n21656 = pi19 ? n21655 : n32;
  assign n21657 = pi18 ? n37 : n21656;
  assign n21658 = pi17 ? n37 : n21657;
  assign n21659 = pi16 ? n439 : n21658;
  assign n21660 = pi15 ? n21659 : n21289;
  assign n21661 = pi14 ? n21660 : n21296;
  assign n21662 = pi13 ? n21652 : n21661;
  assign n21663 = pi16 ? n744 : n21303;
  assign n21664 = pi21 ? n935 : n1211;
  assign n21665 = pi20 ? n32 : n21664;
  assign n21666 = pi19 ? n32 : n21665;
  assign n21667 = pi19 ? n6596 : n139;
  assign n21668 = pi18 ? n21666 : n21667;
  assign n21669 = pi17 ? n32 : n21668;
  assign n21670 = pi16 ? n21669 : n21309;
  assign n21671 = pi15 ? n21663 : n21670;
  assign n21672 = pi16 ? n439 : n21309;
  assign n21673 = pi19 ? n37 : n1003;
  assign n21674 = pi18 ? n21673 : n2350;
  assign n21675 = pi17 ? n21674 : n21323;
  assign n21676 = pi16 ? n439 : n21675;
  assign n21677 = pi15 ? n21672 : n21676;
  assign n21678 = pi14 ? n21671 : n21677;
  assign n21679 = pi20 ? n139 : n3645;
  assign n21680 = pi19 ? n21679 : n139;
  assign n21681 = pi18 ? n21680 : n21329;
  assign n21682 = pi17 ? n9826 : n21681;
  assign n21683 = pi16 ? n439 : n21682;
  assign n21684 = pi22 ? n363 : n1784;
  assign n21685 = pi21 ? n21684 : n1009;
  assign n21686 = pi20 ? n139 : n21685;
  assign n21687 = pi19 ? n21686 : n32;
  assign n21688 = pi18 ? n9825 : n21687;
  assign n21689 = pi17 ? n37 : n21688;
  assign n21690 = pi16 ? n439 : n21689;
  assign n21691 = pi15 ? n21683 : n21690;
  assign n21692 = pi19 ? n12415 : n204;
  assign n21693 = pi21 ? n16438 : n1009;
  assign n21694 = pi20 ? n204 : n21693;
  assign n21695 = pi19 ? n21694 : n32;
  assign n21696 = pi18 ? n21692 : n21695;
  assign n21697 = pi17 ? n37 : n21696;
  assign n21698 = pi16 ? n439 : n21697;
  assign n21699 = pi19 ? n37 : n204;
  assign n21700 = pi20 ? n204 : n9390;
  assign n21701 = pi19 ? n21700 : n32;
  assign n21702 = pi18 ? n21699 : n21701;
  assign n21703 = pi17 ? n37 : n21702;
  assign n21704 = pi16 ? n439 : n21703;
  assign n21705 = pi15 ? n21698 : n21704;
  assign n21706 = pi14 ? n21691 : n21705;
  assign n21707 = pi13 ? n21678 : n21706;
  assign n21708 = pi12 ? n21662 : n21707;
  assign n21709 = pi21 ? n296 : n37;
  assign n21710 = pi20 ? n32 : n21709;
  assign n21711 = pi19 ? n32 : n21710;
  assign n21712 = pi20 ? n3075 : n37;
  assign n21713 = pi19 ? n21712 : n376;
  assign n21714 = pi18 ? n21711 : n21713;
  assign n21715 = pi17 ? n32 : n21714;
  assign n21716 = pi20 ? n13179 : n14034;
  assign n21717 = pi19 ? n13179 : n21716;
  assign n21718 = pi20 ? n3075 : n13613;
  assign n21719 = pi20 ? n9354 : n8742;
  assign n21720 = pi19 ? n21718 : n21719;
  assign n21721 = pi18 ? n21717 : n21720;
  assign n21722 = pi20 ? n16058 : n139;
  assign n21723 = pi21 ? n2876 : n919;
  assign n21724 = pi19 ? n21722 : n21723;
  assign n21725 = pi22 ? n139 : n3174;
  assign n21726 = pi21 ? n21725 : n32;
  assign n21727 = pi20 ? n5199 : n21726;
  assign n21728 = pi19 ? n21727 : n32;
  assign n21729 = pi18 ? n21724 : n21728;
  assign n21730 = pi17 ? n21721 : n21729;
  assign n21731 = pi16 ? n21715 : n21730;
  assign n21732 = pi21 ? n37 : n204;
  assign n21733 = pi20 ? n21732 : n204;
  assign n21734 = pi19 ? n37 : n21733;
  assign n21735 = pi18 ? n21734 : n20751;
  assign n21736 = pi17 ? n37 : n21735;
  assign n21737 = pi16 ? n439 : n21736;
  assign n21738 = pi15 ? n21731 : n21737;
  assign n21739 = pi20 ? n335 : n7598;
  assign n21740 = pi19 ? n21739 : n32;
  assign n21741 = pi18 ? n20818 : n21740;
  assign n21742 = pi17 ? n37 : n21741;
  assign n21743 = pi16 ? n439 : n21742;
  assign n21744 = pi23 ? n6960 : n624;
  assign n21745 = pi22 ? n335 : n21744;
  assign n21746 = pi21 ? n21745 : n32;
  assign n21747 = pi20 ? n335 : n21746;
  assign n21748 = pi19 ? n21747 : n32;
  assign n21749 = pi18 ? n9856 : n21748;
  assign n21750 = pi17 ? n37 : n21749;
  assign n21751 = pi16 ? n439 : n21750;
  assign n21752 = pi15 ? n21743 : n21751;
  assign n21753 = pi14 ? n21738 : n21752;
  assign n21754 = pi18 ? n37 : n3286;
  assign n21755 = pi20 ? n37 : n3335;
  assign n21756 = pi19 ? n21755 : n335;
  assign n21757 = pi18 ? n21756 : n21748;
  assign n21758 = pi17 ? n21754 : n21757;
  assign n21759 = pi16 ? n439 : n21758;
  assign n21760 = pi21 ? n15100 : n32;
  assign n21761 = pi20 ? n335 : n21760;
  assign n21762 = pi19 ? n21761 : n32;
  assign n21763 = pi18 ? n10682 : n21762;
  assign n21764 = pi17 ? n37 : n21763;
  assign n21765 = pi16 ? n439 : n21764;
  assign n21766 = pi15 ? n21759 : n21765;
  assign n21767 = pi18 ? n20818 : n21762;
  assign n21768 = pi17 ? n37 : n21767;
  assign n21769 = pi16 ? n439 : n21768;
  assign n21770 = pi19 ? n37 : n12628;
  assign n21771 = pi18 ? n21770 : n21762;
  assign n21772 = pi17 ? n37 : n21771;
  assign n21773 = pi16 ? n439 : n21772;
  assign n21774 = pi15 ? n21769 : n21773;
  assign n21775 = pi14 ? n21766 : n21774;
  assign n21776 = pi13 ? n21753 : n21775;
  assign n21777 = pi20 ? n335 : n7659;
  assign n21778 = pi19 ? n21777 : n32;
  assign n21779 = pi18 ? n20831 : n21778;
  assign n21780 = pi17 ? n37 : n21779;
  assign n21781 = pi16 ? n439 : n21780;
  assign n21782 = pi20 ? n37 : n7659;
  assign n21783 = pi19 ? n21782 : n32;
  assign n21784 = pi18 ? n37 : n21783;
  assign n21785 = pi17 ? n37 : n21784;
  assign n21786 = pi16 ? n439 : n21785;
  assign n21787 = pi15 ? n21781 : n21786;
  assign n21788 = pi20 ? n233 : n9431;
  assign n21789 = pi19 ? n21788 : n32;
  assign n21790 = pi18 ? n16209 : n21789;
  assign n21791 = pi17 ? n37 : n21790;
  assign n21792 = pi16 ? n439 : n21791;
  assign n21793 = pi20 ? n233 : n16944;
  assign n21794 = pi19 ? n21793 : n32;
  assign n21795 = pi18 ? n16209 : n21794;
  assign n21796 = pi17 ? n37 : n21795;
  assign n21797 = pi16 ? n439 : n21796;
  assign n21798 = pi15 ? n21792 : n21797;
  assign n21799 = pi14 ? n21787 : n21798;
  assign n21800 = pi18 ? n2717 : n21367;
  assign n21801 = pi17 ? n37 : n21800;
  assign n21802 = pi16 ? n439 : n21801;
  assign n21803 = pi21 ? n2106 : n363;
  assign n21804 = pi20 ? n21803 : n9482;
  assign n21805 = pi19 ? n21804 : n32;
  assign n21806 = pi18 ? n2109 : n21805;
  assign n21807 = pi17 ? n37 : n21806;
  assign n21808 = pi16 ? n439 : n21807;
  assign n21809 = pi15 ? n21802 : n21808;
  assign n21810 = pi20 ? n17274 : n4008;
  assign n21811 = pi19 ? n21810 : n32;
  assign n21812 = pi18 ? n2109 : n21811;
  assign n21813 = pi17 ? n37 : n21812;
  assign n21814 = pi16 ? n439 : n21813;
  assign n21815 = pi21 ? n11015 : n32;
  assign n21816 = pi20 ? n7730 : n21815;
  assign n21817 = pi19 ? n21816 : n32;
  assign n21818 = pi18 ? n37 : n21817;
  assign n21819 = pi17 ? n37 : n21818;
  assign n21820 = pi16 ? n439 : n21819;
  assign n21821 = pi15 ? n21814 : n21820;
  assign n21822 = pi14 ? n21809 : n21821;
  assign n21823 = pi13 ? n21799 : n21822;
  assign n21824 = pi12 ? n21776 : n21823;
  assign n21825 = pi11 ? n21708 : n21824;
  assign n21826 = pi21 ? n37 : n10488;
  assign n21827 = pi20 ? n37 : n21826;
  assign n21828 = pi19 ? n37 : n21827;
  assign n21829 = pi18 ? n21828 : n21395;
  assign n21830 = pi17 ? n37 : n21829;
  assign n21831 = pi16 ? n439 : n21830;
  assign n21832 = pi18 ? n37 : n21395;
  assign n21833 = pi17 ? n37 : n21832;
  assign n21834 = pi16 ? n439 : n21833;
  assign n21835 = pi15 ? n21831 : n21834;
  assign n21836 = pi18 ? n37 : n21378;
  assign n21837 = pi17 ? n37 : n21836;
  assign n21838 = pi16 ? n439 : n21837;
  assign n21839 = pi15 ? n21838 : n21409;
  assign n21840 = pi14 ? n21835 : n21839;
  assign n21841 = pi16 ? n744 : n21415;
  assign n21842 = pi22 ? n99 : n2244;
  assign n21843 = pi21 ? n21842 : n99;
  assign n21844 = pi20 ? n21843 : n99;
  assign n21845 = pi19 ? n99 : n21844;
  assign n21846 = pi18 ? n21845 : n21413;
  assign n21847 = pi17 ? n99 : n21846;
  assign n21848 = pi16 ? n744 : n21847;
  assign n21849 = pi20 ? n99 : n5453;
  assign n21850 = pi22 ? n3443 : n157;
  assign n21851 = pi21 ? n21850 : n99;
  assign n21852 = pi21 ? n99 : n8341;
  assign n21853 = pi20 ? n21851 : n21852;
  assign n21854 = pi19 ? n21849 : n21853;
  assign n21855 = pi21 ? n8341 : n767;
  assign n21856 = pi20 ? n21855 : n7049;
  assign n21857 = pi19 ? n21856 : n32;
  assign n21858 = pi18 ? n21854 : n21857;
  assign n21859 = pi17 ? n99 : n21858;
  assign n21860 = pi16 ? n744 : n21859;
  assign n21861 = pi15 ? n21848 : n21860;
  assign n21862 = pi14 ? n21841 : n21861;
  assign n21863 = pi13 ? n21840 : n21862;
  assign n21864 = pi20 ? n7818 : n157;
  assign n21865 = pi19 ? n15271 : n21864;
  assign n21866 = pi18 ? n21865 : n21428;
  assign n21867 = pi17 ? n99 : n21866;
  assign n21868 = pi16 ? n744 : n21867;
  assign n21869 = pi22 ? n5167 : n99;
  assign n21870 = pi21 ? n21869 : n99;
  assign n21871 = pi20 ? n32 : n21870;
  assign n21872 = pi19 ? n32 : n21871;
  assign n21873 = pi19 ? n161 : n9708;
  assign n21874 = pi18 ? n21872 : n21873;
  assign n21875 = pi17 ? n32 : n21874;
  assign n21876 = pi20 ? n776 : n3006;
  assign n21877 = pi19 ? n166 : n21876;
  assign n21878 = pi21 ? n775 : n168;
  assign n21879 = pi20 ? n21878 : n802;
  assign n21880 = pi20 ? n3014 : n7104;
  assign n21881 = pi19 ? n21879 : n21880;
  assign n21882 = pi18 ? n21877 : n21881;
  assign n21883 = pi20 ? n7111 : n157;
  assign n21884 = pi19 ? n21883 : n157;
  assign n21885 = pi20 ? n7435 : n10011;
  assign n21886 = pi19 ? n21885 : n32;
  assign n21887 = pi18 ? n21884 : n21886;
  assign n21888 = pi17 ? n21882 : n21887;
  assign n21889 = pi16 ? n21875 : n21888;
  assign n21890 = pi15 ? n21868 : n21889;
  assign n21891 = pi16 ? n16338 : n21443;
  assign n21892 = pi15 ? n21444 : n21891;
  assign n21893 = pi14 ? n21890 : n21892;
  assign n21894 = pi23 ? n204 : n157;
  assign n21895 = pi22 ? n16332 : n21894;
  assign n21896 = pi21 ? n21895 : n5176;
  assign n21897 = pi20 ? n32 : n21896;
  assign n21898 = pi19 ? n32 : n21897;
  assign n21899 = pi22 ? n164 : n21894;
  assign n21900 = pi22 ? n893 : n204;
  assign n21901 = pi21 ? n21899 : n21900;
  assign n21902 = pi22 ? n21894 : n204;
  assign n21903 = pi21 ? n7815 : n21902;
  assign n21904 = pi20 ? n21901 : n21903;
  assign n21905 = pi20 ? n21903 : n21901;
  assign n21906 = pi19 ? n21904 : n21905;
  assign n21907 = pi18 ? n21898 : n21906;
  assign n21908 = pi17 ? n32 : n21907;
  assign n21909 = pi22 ? n204 : n164;
  assign n21910 = pi21 ? n21899 : n21909;
  assign n21911 = pi22 ? n157 : n21894;
  assign n21912 = pi21 ? n21902 : n21911;
  assign n21913 = pi20 ? n21910 : n21912;
  assign n21914 = pi19 ? n21901 : n21913;
  assign n21915 = pi21 ? n5176 : n21911;
  assign n21916 = pi21 ? n5176 : n21899;
  assign n21917 = pi20 ? n21915 : n21916;
  assign n21918 = pi22 ? n21894 : n893;
  assign n21919 = pi21 ? n5176 : n21918;
  assign n21920 = pi21 ? n21909 : n21902;
  assign n21921 = pi20 ? n21919 : n21920;
  assign n21922 = pi19 ? n21917 : n21921;
  assign n21923 = pi18 ? n21914 : n21922;
  assign n21924 = pi22 ? n164 : n204;
  assign n21925 = pi22 ? n861 : n204;
  assign n21926 = pi21 ? n21924 : n21925;
  assign n21927 = pi21 ? n4268 : n20977;
  assign n21928 = pi20 ? n21926 : n21927;
  assign n21929 = pi22 ? n19177 : n204;
  assign n21930 = pi21 ? n21929 : n4281;
  assign n21931 = pi21 ? n21909 : n5176;
  assign n21932 = pi20 ? n21930 : n21931;
  assign n21933 = pi19 ? n21928 : n21932;
  assign n21934 = pi22 ? n21894 : n316;
  assign n21935 = pi21 ? n21934 : n316;
  assign n21936 = pi20 ? n21935 : n1822;
  assign n21937 = pi19 ? n21936 : n32;
  assign n21938 = pi18 ? n21933 : n21937;
  assign n21939 = pi17 ? n21923 : n21938;
  assign n21940 = pi16 ? n21908 : n21939;
  assign n21941 = pi20 ? n7909 : n1822;
  assign n21942 = pi19 ? n21941 : n32;
  assign n21943 = pi18 ? n20990 : n21942;
  assign n21944 = pi17 ? n204 : n21943;
  assign n21945 = pi16 ? n20988 : n21944;
  assign n21946 = pi15 ? n21940 : n21945;
  assign n21947 = pi20 ? n316 : n1822;
  assign n21948 = pi19 ? n21947 : n32;
  assign n21949 = pi18 ? n21004 : n21948;
  assign n21950 = pi17 ? n204 : n21949;
  assign n21951 = pi16 ? n20988 : n21950;
  assign n21952 = pi21 ? n1309 : n204;
  assign n21953 = pi20 ? n21952 : n204;
  assign n21954 = pi19 ? n21953 : n204;
  assign n21955 = pi18 ? n204 : n21954;
  assign n21956 = pi18 ? n21016 : n21948;
  assign n21957 = pi17 ? n21955 : n21956;
  assign n21958 = pi16 ? n13477 : n21957;
  assign n21959 = pi15 ? n21951 : n21958;
  assign n21960 = pi14 ? n21946 : n21959;
  assign n21961 = pi13 ? n21893 : n21960;
  assign n21962 = pi12 ? n21863 : n21961;
  assign n21963 = pi20 ? n1008 : n316;
  assign n21964 = pi19 ? n21963 : n15347;
  assign n21965 = pi18 ? n21964 : n21948;
  assign n21966 = pi17 ? n139 : n21965;
  assign n21967 = pi16 ? n2291 : n21966;
  assign n21968 = pi20 ? n6568 : n316;
  assign n21969 = pi19 ? n21968 : n316;
  assign n21970 = pi18 ? n21969 : n21948;
  assign n21971 = pi17 ? n139 : n21970;
  assign n21972 = pi16 ? n2291 : n21971;
  assign n21973 = pi15 ? n21967 : n21972;
  assign n21974 = pi19 ? n1809 : n9769;
  assign n21975 = pi18 ? n2364 : n21974;
  assign n21976 = pi17 ? n32 : n21975;
  assign n21977 = pi20 ? n6568 : n922;
  assign n21978 = pi20 ? n1016 : n139;
  assign n21979 = pi19 ? n21977 : n21978;
  assign n21980 = pi22 ? n204 : n6415;
  assign n21981 = pi21 ? n139 : n21980;
  assign n21982 = pi20 ? n21981 : n32;
  assign n21983 = pi19 ? n21982 : n32;
  assign n21984 = pi18 ? n21979 : n21983;
  assign n21985 = pi17 ? n139 : n21984;
  assign n21986 = pi16 ? n21976 : n21985;
  assign n21987 = pi20 ? n2316 : n204;
  assign n21988 = pi19 ? n21987 : n204;
  assign n21989 = pi21 ? n204 : n10417;
  assign n21990 = pi20 ? n21989 : n32;
  assign n21991 = pi19 ? n21990 : n32;
  assign n21992 = pi18 ? n21988 : n21991;
  assign n21993 = pi17 ? n139 : n21992;
  assign n21994 = pi16 ? n915 : n21993;
  assign n21995 = pi15 ? n21986 : n21994;
  assign n21996 = pi14 ? n21973 : n21995;
  assign n21997 = pi19 ? n16516 : n612;
  assign n21998 = pi18 ? n7941 : n21997;
  assign n21999 = pi17 ? n32 : n21998;
  assign n22000 = pi21 ? n569 : n1046;
  assign n22001 = pi20 ? n22000 : n335;
  assign n22002 = pi19 ? n603 : n22001;
  assign n22003 = pi19 ? n3384 : n335;
  assign n22004 = pi18 ? n22002 : n22003;
  assign n22005 = pi21 ? n204 : n12381;
  assign n22006 = pi20 ? n22005 : n32;
  assign n22007 = pi19 ? n22006 : n32;
  assign n22008 = pi18 ? n21076 : n22007;
  assign n22009 = pi17 ? n22004 : n22008;
  assign n22010 = pi16 ? n21999 : n22009;
  assign n22011 = pi15 ? n21994 : n22010;
  assign n22012 = pi19 ? n610 : n335;
  assign n22013 = pi18 ? n374 : n22012;
  assign n22014 = pi17 ? n32 : n22013;
  assign n22015 = pi19 ? n612 : n335;
  assign n22016 = pi18 ? n335 : n22015;
  assign n22017 = pi20 ? n18121 : n335;
  assign n22018 = pi20 ? n15469 : n15457;
  assign n22019 = pi19 ? n22017 : n22018;
  assign n22020 = pi21 ? n233 : n8916;
  assign n22021 = pi20 ? n22020 : n32;
  assign n22022 = pi19 ? n22021 : n32;
  assign n22023 = pi18 ? n22019 : n22022;
  assign n22024 = pi17 ? n22016 : n22023;
  assign n22025 = pi16 ? n22014 : n22024;
  assign n22026 = pi20 ? n37 : n610;
  assign n22027 = pi20 ? n610 : n639;
  assign n22028 = pi19 ? n22026 : n22027;
  assign n22029 = pi18 ? n374 : n22028;
  assign n22030 = pi17 ? n32 : n22029;
  assign n22031 = pi20 ? n639 : n335;
  assign n22032 = pi19 ? n22031 : n335;
  assign n22033 = pi18 ? n22032 : n335;
  assign n22034 = pi20 ? n15457 : n18121;
  assign n22035 = pi20 ? n15465 : n6376;
  assign n22036 = pi19 ? n22034 : n22035;
  assign n22037 = pi21 ? n6376 : n7034;
  assign n22038 = pi20 ? n22037 : n32;
  assign n22039 = pi19 ? n22038 : n32;
  assign n22040 = pi18 ? n22036 : n22039;
  assign n22041 = pi17 ? n22033 : n22040;
  assign n22042 = pi16 ? n22030 : n22041;
  assign n22043 = pi15 ? n22025 : n22042;
  assign n22044 = pi14 ? n22011 : n22043;
  assign n22045 = pi13 ? n21996 : n22044;
  assign n22046 = pi20 ? n638 : n37;
  assign n22047 = pi19 ? n37 : n22046;
  assign n22048 = pi20 ? n649 : n571;
  assign n22049 = pi19 ? n37 : n22048;
  assign n22050 = pi18 ? n22047 : n22049;
  assign n22051 = pi20 ? n15457 : n16544;
  assign n22052 = pi20 ? n16544 : n13527;
  assign n22053 = pi19 ? n22051 : n22052;
  assign n22054 = pi18 ? n22053 : n14676;
  assign n22055 = pi17 ? n22050 : n22054;
  assign n22056 = pi16 ? n439 : n22055;
  assign n22057 = pi19 ? n37 : n2050;
  assign n22058 = pi21 ? n2117 : n2091;
  assign n22059 = pi20 ? n37 : n22058;
  assign n22060 = pi19 ? n37 : n22059;
  assign n22061 = pi18 ? n22057 : n22060;
  assign n22062 = pi20 ? n4921 : n13527;
  assign n22063 = pi19 ? n22062 : n233;
  assign n22064 = pi18 ? n22063 : n14676;
  assign n22065 = pi17 ? n22061 : n22064;
  assign n22066 = pi16 ? n439 : n22065;
  assign n22067 = pi15 ? n22056 : n22066;
  assign n22068 = pi19 ? n37 : n6340;
  assign n22069 = pi18 ? n22068 : n16209;
  assign n22070 = pi18 ? n21164 : n14676;
  assign n22071 = pi17 ? n22069 : n22070;
  assign n22072 = pi16 ? n439 : n22071;
  assign n22073 = pi21 ? n180 : n569;
  assign n22074 = pi20 ? n32 : n22073;
  assign n22075 = pi19 ? n32 : n22074;
  assign n22076 = pi21 ? n335 : n574;
  assign n22077 = pi20 ? n22076 : n19368;
  assign n22078 = pi19 ? n644 : n22077;
  assign n22079 = pi18 ? n22075 : n22078;
  assign n22080 = pi17 ? n32 : n22079;
  assign n22081 = pi20 ? n19368 : n610;
  assign n22082 = pi19 ? n22081 : n10957;
  assign n22083 = pi20 ? n603 : n577;
  assign n22084 = pi19 ? n22083 : n14166;
  assign n22085 = pi18 ? n22082 : n22084;
  assign n22086 = pi20 ? n7980 : n13527;
  assign n22087 = pi20 ? n7980 : n6377;
  assign n22088 = pi19 ? n22086 : n22087;
  assign n22089 = pi21 ? n233 : n7723;
  assign n22090 = pi20 ? n22089 : n32;
  assign n22091 = pi19 ? n22090 : n32;
  assign n22092 = pi18 ? n22088 : n22091;
  assign n22093 = pi17 ? n22085 : n22092;
  assign n22094 = pi16 ? n22080 : n22093;
  assign n22095 = pi15 ? n22072 : n22094;
  assign n22096 = pi14 ? n22067 : n22095;
  assign n22097 = pi21 ? n2061 : n6361;
  assign n22098 = pi20 ? n22097 : n335;
  assign n22099 = pi19 ? n335 : n22098;
  assign n22100 = pi18 ? n22099 : n15438;
  assign n22101 = pi20 ? n6362 : n6377;
  assign n22102 = pi19 ? n21110 : n22101;
  assign n22103 = pi21 ? n6376 : n2320;
  assign n22104 = pi20 ? n22103 : n32;
  assign n22105 = pi19 ? n22104 : n32;
  assign n22106 = pi18 ? n22102 : n22105;
  assign n22107 = pi17 ? n22100 : n22106;
  assign n22108 = pi16 ? n12648 : n22107;
  assign n22109 = pi21 ? n716 : n1657;
  assign n22110 = pi20 ? n32 : n22109;
  assign n22111 = pi19 ? n32 : n22110;
  assign n22112 = pi21 ? n335 : n1657;
  assign n22113 = pi22 ? n1656 : n99;
  assign n22114 = pi21 ? n17548 : n22113;
  assign n22115 = pi20 ? n22112 : n22114;
  assign n22116 = pi23 ? n335 : n99;
  assign n22117 = pi22 ? n363 : n22116;
  assign n22118 = pi22 ? n18461 : n99;
  assign n22119 = pi21 ? n22117 : n22118;
  assign n22120 = pi22 ? n335 : n22116;
  assign n22121 = pi21 ? n22120 : n22118;
  assign n22122 = pi20 ? n22119 : n22121;
  assign n22123 = pi19 ? n22115 : n22122;
  assign n22124 = pi18 ? n22111 : n22123;
  assign n22125 = pi17 ? n32 : n22124;
  assign n22126 = pi21 ? n335 : n20226;
  assign n22127 = pi20 ? n22121 : n22126;
  assign n22128 = pi22 ? n233 : n99;
  assign n22129 = pi21 ? n21235 : n22128;
  assign n22130 = pi22 ? n18461 : n1656;
  assign n22131 = pi21 ? n22130 : n22120;
  assign n22132 = pi20 ? n22129 : n22131;
  assign n22133 = pi19 ? n22127 : n22132;
  assign n22134 = pi21 ? n722 : n335;
  assign n22135 = pi22 ? n1656 : n363;
  assign n22136 = pi21 ? n22135 : n18467;
  assign n22137 = pi20 ? n22134 : n22136;
  assign n22138 = pi19 ? n22137 : n21206;
  assign n22139 = pi18 ? n22133 : n22138;
  assign n22140 = pi22 ? n233 : n18461;
  assign n22141 = pi21 ? n22140 : n233;
  assign n22142 = pi22 ? n18461 : n233;
  assign n22143 = pi21 ? n2707 : n22142;
  assign n22144 = pi20 ? n22141 : n22143;
  assign n22145 = pi19 ? n21110 : n22144;
  assign n22146 = pi21 ? n22142 : n882;
  assign n22147 = pi20 ? n22146 : n32;
  assign n22148 = pi19 ? n22147 : n32;
  assign n22149 = pi18 ? n22145 : n22148;
  assign n22150 = pi17 ? n22139 : n22149;
  assign n22151 = pi16 ? n22125 : n22150;
  assign n22152 = pi15 ? n22108 : n22151;
  assign n22153 = pi21 ? n233 : n5014;
  assign n22154 = pi20 ? n22153 : n363;
  assign n22155 = pi19 ? n21225 : n22154;
  assign n22156 = pi19 ? n21225 : n233;
  assign n22157 = pi18 ? n22155 : n22156;
  assign n22158 = pi21 ? n12635 : n882;
  assign n22159 = pi20 ? n22158 : n32;
  assign n22160 = pi19 ? n22159 : n32;
  assign n22161 = pi18 ? n233 : n22160;
  assign n22162 = pi17 ? n22157 : n22161;
  assign n22163 = pi16 ? n21219 : n22162;
  assign n22164 = pi20 ? n21222 : n20860;
  assign n22165 = pi19 ? n19423 : n22164;
  assign n22166 = pi18 ? n19433 : n22165;
  assign n22167 = pi17 ? n32 : n22166;
  assign n22168 = pi18 ? n233 : n20209;
  assign n22169 = pi17 ? n21244 : n22168;
  assign n22170 = pi16 ? n22167 : n22169;
  assign n22171 = pi15 ? n22163 : n22170;
  assign n22172 = pi14 ? n22152 : n22171;
  assign n22173 = pi13 ? n22096 : n22172;
  assign n22174 = pi12 ? n22045 : n22173;
  assign n22175 = pi11 ? n21962 : n22174;
  assign n22176 = pi10 ? n21825 : n22175;
  assign n22177 = pi09 ? n21601 : n22176;
  assign n22178 = pi16 ? n13561 : n21582;
  assign n22179 = pi15 ? n32 : n22178;
  assign n22180 = pi14 ? n22179 : n21596;
  assign n22181 = pi13 ? n32 : n22180;
  assign n22182 = pi12 ? n32 : n22181;
  assign n22183 = pi11 ? n32 : n22182;
  assign n22184 = pi10 ? n32 : n22183;
  assign n22185 = pi16 ? n17010 : n21627;
  assign n22186 = pi15 ? n22185 : n21650;
  assign n22187 = pi14 ? n21621 : n22186;
  assign n22188 = pi21 ? n14477 : n2469;
  assign n22189 = pi20 ? n99 : n22188;
  assign n22190 = pi19 ? n22189 : n32;
  assign n22191 = pi18 ? n99 : n22190;
  assign n22192 = pi17 ? n99 : n22191;
  assign n22193 = pi16 ? n801 : n22192;
  assign n22194 = pi15 ? n21659 : n22193;
  assign n22195 = pi20 ? n99 : n8088;
  assign n22196 = pi19 ? n22195 : n32;
  assign n22197 = pi18 ? n99 : n22196;
  assign n22198 = pi17 ? n99 : n22197;
  assign n22199 = pi16 ? n744 : n22198;
  assign n22200 = pi20 ? n99 : n8095;
  assign n22201 = pi19 ? n22200 : n32;
  assign n22202 = pi18 ? n99 : n22201;
  assign n22203 = pi17 ? n99 : n22202;
  assign n22204 = pi16 ? n721 : n22203;
  assign n22205 = pi15 ? n22199 : n22204;
  assign n22206 = pi14 ? n22194 : n22205;
  assign n22207 = pi13 ? n22187 : n22206;
  assign n22208 = pi22 ? n962 : n295;
  assign n22209 = pi21 ? n22208 : n1211;
  assign n22210 = pi20 ? n32 : n22209;
  assign n22211 = pi19 ? n32 : n22210;
  assign n22212 = pi18 ? n22211 : n21667;
  assign n22213 = pi17 ? n32 : n22212;
  assign n22214 = pi21 ? n139 : n2678;
  assign n22215 = pi20 ? n139 : n22214;
  assign n22216 = pi19 ? n22215 : n32;
  assign n22217 = pi18 ? n139 : n22216;
  assign n22218 = pi17 ? n139 : n22217;
  assign n22219 = pi16 ? n22213 : n22218;
  assign n22220 = pi15 ? n22204 : n22219;
  assign n22221 = pi16 ? n439 : n22218;
  assign n22222 = pi21 ? n139 : n2700;
  assign n22223 = pi20 ? n139 : n22222;
  assign n22224 = pi19 ? n22223 : n32;
  assign n22225 = pi18 ? n139 : n22224;
  assign n22226 = pi17 ? n21674 : n22225;
  assign n22227 = pi16 ? n439 : n22226;
  assign n22228 = pi15 ? n22221 : n22227;
  assign n22229 = pi14 ? n22220 : n22228;
  assign n22230 = pi21 ? n335 : n2700;
  assign n22231 = pi20 ? n139 : n22230;
  assign n22232 = pi19 ? n22231 : n32;
  assign n22233 = pi18 ? n21680 : n22232;
  assign n22234 = pi17 ? n9826 : n22233;
  assign n22235 = pi16 ? n439 : n22234;
  assign n22236 = pi22 ? n363 : n364;
  assign n22237 = pi21 ? n22236 : n1009;
  assign n22238 = pi20 ? n139 : n22237;
  assign n22239 = pi19 ? n22238 : n32;
  assign n22240 = pi18 ? n9825 : n22239;
  assign n22241 = pi17 ? n37 : n22240;
  assign n22242 = pi16 ? n439 : n22241;
  assign n22243 = pi15 ? n22235 : n22242;
  assign n22244 = pi22 ? n204 : n21894;
  assign n22245 = pi21 ? n22244 : n1009;
  assign n22246 = pi20 ? n204 : n22245;
  assign n22247 = pi19 ? n22246 : n32;
  assign n22248 = pi18 ? n21692 : n22247;
  assign n22249 = pi17 ? n37 : n22248;
  assign n22250 = pi16 ? n439 : n22249;
  assign n22251 = pi15 ? n22250 : n21704;
  assign n22252 = pi14 ? n22243 : n22251;
  assign n22253 = pi13 ? n22229 : n22252;
  assign n22254 = pi12 ? n22207 : n22253;
  assign n22255 = pi20 ? n14061 : n13179;
  assign n22256 = pi21 ? n3668 : n1529;
  assign n22257 = pi20 ? n13179 : n22256;
  assign n22258 = pi19 ? n22255 : n22257;
  assign n22259 = pi20 ? n3606 : n17681;
  assign n22260 = pi20 ? n13138 : n14076;
  assign n22261 = pi19 ? n22259 : n22260;
  assign n22262 = pi18 ? n22258 : n22261;
  assign n22263 = pi19 ? n18582 : n5215;
  assign n22264 = pi22 ? n139 : n4079;
  assign n22265 = pi21 ? n22264 : n32;
  assign n22266 = pi20 ? n5229 : n22265;
  assign n22267 = pi19 ? n22266 : n32;
  assign n22268 = pi18 ? n22263 : n22267;
  assign n22269 = pi17 ? n22262 : n22268;
  assign n22270 = pi16 ? n21715 : n22269;
  assign n22271 = pi21 ? n3763 : n32;
  assign n22272 = pi20 ? n204 : n22271;
  assign n22273 = pi19 ? n22272 : n32;
  assign n22274 = pi18 ? n21734 : n22273;
  assign n22275 = pi17 ? n37 : n22274;
  assign n22276 = pi16 ? n439 : n22275;
  assign n22277 = pi15 ? n22270 : n22276;
  assign n22278 = pi22 ? n335 : n6077;
  assign n22279 = pi21 ? n22278 : n32;
  assign n22280 = pi20 ? n335 : n22279;
  assign n22281 = pi19 ? n22280 : n32;
  assign n22282 = pi18 ? n9856 : n22281;
  assign n22283 = pi17 ? n37 : n22282;
  assign n22284 = pi16 ? n439 : n22283;
  assign n22285 = pi15 ? n21743 : n22284;
  assign n22286 = pi14 ? n22277 : n22285;
  assign n22287 = pi21 ? n15647 : n32;
  assign n22288 = pi20 ? n335 : n22287;
  assign n22289 = pi19 ? n22288 : n32;
  assign n22290 = pi18 ? n21756 : n22289;
  assign n22291 = pi17 ? n21754 : n22290;
  assign n22292 = pi16 ? n439 : n22291;
  assign n22293 = pi15 ? n22292 : n21765;
  assign n22294 = pi14 ? n22293 : n21774;
  assign n22295 = pi13 ? n22286 : n22294;
  assign n22296 = pi18 ? n20831 : n21762;
  assign n22297 = pi17 ? n37 : n22296;
  assign n22298 = pi16 ? n439 : n22297;
  assign n22299 = pi15 ? n22298 : n21786;
  assign n22300 = pi20 ? n233 : n17510;
  assign n22301 = pi19 ? n22300 : n32;
  assign n22302 = pi18 ? n16209 : n22301;
  assign n22303 = pi17 ? n37 : n22302;
  assign n22304 = pi16 ? n439 : n22303;
  assign n22305 = pi22 ? n233 : n10098;
  assign n22306 = pi21 ? n22305 : n32;
  assign n22307 = pi20 ? n233 : n22306;
  assign n22308 = pi19 ? n22307 : n32;
  assign n22309 = pi18 ? n16209 : n22308;
  assign n22310 = pi17 ? n37 : n22309;
  assign n22311 = pi16 ? n439 : n22310;
  assign n22312 = pi15 ? n22304 : n22311;
  assign n22313 = pi14 ? n22299 : n22312;
  assign n22314 = pi22 ? n685 : n15697;
  assign n22315 = pi21 ? n22314 : n32;
  assign n22316 = pi20 ? n20860 : n22315;
  assign n22317 = pi19 ? n22316 : n32;
  assign n22318 = pi18 ? n2717 : n22317;
  assign n22319 = pi17 ? n37 : n22318;
  assign n22320 = pi16 ? n439 : n22319;
  assign n22321 = pi20 ? n21803 : n8295;
  assign n22322 = pi19 ? n22321 : n32;
  assign n22323 = pi18 ? n2109 : n22322;
  assign n22324 = pi17 ? n37 : n22323;
  assign n22325 = pi16 ? n439 : n22324;
  assign n22326 = pi15 ? n22320 : n22325;
  assign n22327 = pi20 ? n17274 : n12149;
  assign n22328 = pi19 ? n22327 : n32;
  assign n22329 = pi18 ? n2109 : n22328;
  assign n22330 = pi17 ? n37 : n22329;
  assign n22331 = pi16 ? n439 : n22330;
  assign n22332 = pi22 ? n363 : n688;
  assign n22333 = pi21 ? n22332 : n32;
  assign n22334 = pi20 ? n7730 : n22333;
  assign n22335 = pi19 ? n22334 : n32;
  assign n22336 = pi18 ? n37 : n22335;
  assign n22337 = pi17 ? n37 : n22336;
  assign n22338 = pi16 ? n439 : n22337;
  assign n22339 = pi15 ? n22331 : n22338;
  assign n22340 = pi14 ? n22326 : n22339;
  assign n22341 = pi13 ? n22313 : n22340;
  assign n22342 = pi12 ? n22295 : n22341;
  assign n22343 = pi11 ? n22254 : n22342;
  assign n22344 = pi20 ? n363 : n8295;
  assign n22345 = pi19 ? n22344 : n32;
  assign n22346 = pi18 ? n21828 : n22345;
  assign n22347 = pi17 ? n37 : n22346;
  assign n22348 = pi16 ? n439 : n22347;
  assign n22349 = pi18 ? n37 : n22345;
  assign n22350 = pi17 ? n37 : n22349;
  assign n22351 = pi16 ? n439 : n22350;
  assign n22352 = pi15 ? n22348 : n22351;
  assign n22353 = pi20 ? n7730 : n8295;
  assign n22354 = pi19 ? n22353 : n32;
  assign n22355 = pi18 ? n37 : n22354;
  assign n22356 = pi17 ? n37 : n22355;
  assign n22357 = pi16 ? n439 : n22356;
  assign n22358 = pi20 ? n2107 : n8295;
  assign n22359 = pi19 ? n22358 : n32;
  assign n22360 = pi18 ? n37 : n22359;
  assign n22361 = pi17 ? n37 : n22360;
  assign n22362 = pi16 ? n439 : n22361;
  assign n22363 = pi15 ? n22357 : n22362;
  assign n22364 = pi14 ? n22352 : n22363;
  assign n22365 = pi20 ? n5085 : n8295;
  assign n22366 = pi19 ? n22365 : n32;
  assign n22367 = pi18 ? n99 : n22366;
  assign n22368 = pi17 ? n99 : n22367;
  assign n22369 = pi16 ? n721 : n22368;
  assign n22370 = pi20 ? n5085 : n9482;
  assign n22371 = pi19 ? n22370 : n32;
  assign n22372 = pi18 ? n21845 : n22371;
  assign n22373 = pi17 ? n99 : n22372;
  assign n22374 = pi16 ? n721 : n22373;
  assign n22375 = pi21 ? n2164 : n5453;
  assign n22376 = pi20 ? n99 : n22375;
  assign n22377 = pi22 ? n2160 : n157;
  assign n22378 = pi21 ? n22377 : n99;
  assign n22379 = pi22 ? n157 : n2160;
  assign n22380 = pi21 ? n99 : n22379;
  assign n22381 = pi20 ? n22378 : n22380;
  assign n22382 = pi19 ? n22376 : n22381;
  assign n22383 = pi23 ? n842 : n316;
  assign n22384 = pi22 ? n22383 : n706;
  assign n22385 = pi21 ? n22384 : n32;
  assign n22386 = pi20 ? n21855 : n22385;
  assign n22387 = pi19 ? n22386 : n32;
  assign n22388 = pi18 ? n22382 : n22387;
  assign n22389 = pi17 ? n99 : n22388;
  assign n22390 = pi16 ? n721 : n22389;
  assign n22391 = pi15 ? n22374 : n22390;
  assign n22392 = pi14 ? n22369 : n22391;
  assign n22393 = pi13 ? n22364 : n22392;
  assign n22394 = pi21 ? n844 : n32;
  assign n22395 = pi20 ? n157 : n22394;
  assign n22396 = pi19 ? n22395 : n32;
  assign n22397 = pi18 ? n21865 : n22396;
  assign n22398 = pi17 ? n99 : n22397;
  assign n22399 = pi16 ? n721 : n22398;
  assign n22400 = pi20 ? n99 : n4617;
  assign n22401 = pi20 ? n4616 : n4625;
  assign n22402 = pi19 ? n22400 : n22401;
  assign n22403 = pi18 ? n1508 : n22402;
  assign n22404 = pi17 ? n32 : n22403;
  assign n22405 = pi19 ? n4625 : n21876;
  assign n22406 = pi20 ? n3014 : n2174;
  assign n22407 = pi19 ? n21879 : n22406;
  assign n22408 = pi18 ? n22405 : n22407;
  assign n22409 = pi21 ? n22377 : n777;
  assign n22410 = pi20 ? n22409 : n157;
  assign n22411 = pi19 ? n22410 : n157;
  assign n22412 = pi18 ? n22411 : n21886;
  assign n22413 = pi17 ? n22408 : n22412;
  assign n22414 = pi16 ? n22404 : n22413;
  assign n22415 = pi15 ? n22399 : n22414;
  assign n22416 = pi20 ? n7435 : n2653;
  assign n22417 = pi19 ? n22416 : n32;
  assign n22418 = pi18 ? n157 : n22417;
  assign n22419 = pi17 ? n157 : n22418;
  assign n22420 = pi16 ? n7419 : n22419;
  assign n22421 = pi16 ? n16349 : n22419;
  assign n22422 = pi15 ? n22420 : n22421;
  assign n22423 = pi14 ? n22415 : n22422;
  assign n22424 = pi22 ? n738 : n204;
  assign n22425 = pi21 ? n22424 : n5176;
  assign n22426 = pi20 ? n32 : n22425;
  assign n22427 = pi19 ? n32 : n22426;
  assign n22428 = pi23 ? n204 : n99;
  assign n22429 = pi22 ? n22428 : n21894;
  assign n22430 = pi21 ? n22429 : n1578;
  assign n22431 = pi22 ? n157 : n22428;
  assign n22432 = pi21 ? n22431 : n204;
  assign n22433 = pi20 ? n22430 : n22432;
  assign n22434 = pi20 ? n22432 : n22430;
  assign n22435 = pi19 ? n22433 : n22434;
  assign n22436 = pi18 ? n22427 : n22435;
  assign n22437 = pi17 ? n32 : n22436;
  assign n22438 = pi22 ? n204 : n22428;
  assign n22439 = pi21 ? n22429 : n22438;
  assign n22440 = pi20 ? n22439 : n21912;
  assign n22441 = pi19 ? n22430 : n22440;
  assign n22442 = pi21 ? n5176 : n22429;
  assign n22443 = pi20 ? n21915 : n22442;
  assign n22444 = pi22 ? n21894 : n456;
  assign n22445 = pi21 ? n5176 : n22444;
  assign n22446 = pi21 ? n22438 : n204;
  assign n22447 = pi20 ? n22445 : n22446;
  assign n22448 = pi19 ? n22443 : n22447;
  assign n22449 = pi18 ? n22441 : n22448;
  assign n22450 = pi22 ? n22428 : n204;
  assign n22451 = pi21 ? n22450 : n21925;
  assign n22452 = pi22 ? n812 : n316;
  assign n22453 = pi21 ? n4268 : n22452;
  assign n22454 = pi20 ? n22451 : n22453;
  assign n22455 = pi22 ? n204 : n812;
  assign n22456 = pi21 ? n22455 : n5176;
  assign n22457 = pi20 ? n21930 : n22456;
  assign n22458 = pi19 ? n22454 : n22457;
  assign n22459 = pi20 ? n7187 : n2554;
  assign n22460 = pi19 ? n22459 : n32;
  assign n22461 = pi18 ? n22458 : n22460;
  assign n22462 = pi17 ? n22449 : n22461;
  assign n22463 = pi16 ? n22437 : n22462;
  assign n22464 = pi20 ? n7909 : n2554;
  assign n22465 = pi19 ? n22464 : n32;
  assign n22466 = pi18 ? n20990 : n22465;
  assign n22467 = pi17 ? n204 : n22466;
  assign n22468 = pi16 ? n19219 : n22467;
  assign n22469 = pi15 ? n22463 : n22468;
  assign n22470 = pi20 ? n316 : n2554;
  assign n22471 = pi19 ? n22470 : n32;
  assign n22472 = pi18 ? n21004 : n22471;
  assign n22473 = pi17 ? n204 : n22472;
  assign n22474 = pi16 ? n19219 : n22473;
  assign n22475 = pi20 ? n316 : n2679;
  assign n22476 = pi19 ? n22475 : n32;
  assign n22477 = pi18 ? n21016 : n22476;
  assign n22478 = pi17 ? n21955 : n22477;
  assign n22479 = pi16 ? n13846 : n22478;
  assign n22480 = pi15 ? n22474 : n22479;
  assign n22481 = pi14 ? n22469 : n22480;
  assign n22482 = pi13 ? n22423 : n22481;
  assign n22483 = pi12 ? n22393 : n22482;
  assign n22484 = pi20 ? n316 : n2701;
  assign n22485 = pi19 ? n22484 : n32;
  assign n22486 = pi18 ? n21964 : n22485;
  assign n22487 = pi17 ? n139 : n22486;
  assign n22488 = pi16 ? n915 : n22487;
  assign n22489 = pi16 ? n915 : n21971;
  assign n22490 = pi15 ? n22488 : n22489;
  assign n22491 = pi22 ? n204 : n6365;
  assign n22492 = pi21 ? n139 : n22491;
  assign n22493 = pi20 ? n22492 : n32;
  assign n22494 = pi19 ? n22493 : n32;
  assign n22495 = pi18 ? n21979 : n22494;
  assign n22496 = pi17 ? n139 : n22495;
  assign n22497 = pi16 ? n21976 : n22496;
  assign n22498 = pi23 ? n4145 : n316;
  assign n22499 = pi22 ? n204 : n22498;
  assign n22500 = pi21 ? n204 : n22499;
  assign n22501 = pi20 ? n22500 : n32;
  assign n22502 = pi19 ? n22501 : n32;
  assign n22503 = pi18 ? n21988 : n22502;
  assign n22504 = pi17 ? n139 : n22503;
  assign n22505 = pi16 ? n915 : n22504;
  assign n22506 = pi15 ? n22497 : n22505;
  assign n22507 = pi14 ? n22490 : n22506;
  assign n22508 = pi21 ? n204 : n10410;
  assign n22509 = pi20 ? n22508 : n32;
  assign n22510 = pi19 ? n22509 : n32;
  assign n22511 = pi18 ? n21988 : n22510;
  assign n22512 = pi17 ? n139 : n22511;
  assign n22513 = pi16 ? n915 : n22512;
  assign n22514 = pi22 ? n204 : n5369;
  assign n22515 = pi21 ? n204 : n22514;
  assign n22516 = pi20 ? n22515 : n32;
  assign n22517 = pi19 ? n22516 : n32;
  assign n22518 = pi18 ? n21076 : n22517;
  assign n22519 = pi17 ? n22004 : n22518;
  assign n22520 = pi16 ? n21999 : n22519;
  assign n22521 = pi15 ? n22513 : n22520;
  assign n22522 = pi18 ? n8884 : n22012;
  assign n22523 = pi17 ? n32 : n22522;
  assign n22524 = pi16 ? n22523 : n22024;
  assign n22525 = pi21 ? n6376 : n5758;
  assign n22526 = pi20 ? n22525 : n32;
  assign n22527 = pi19 ? n22526 : n32;
  assign n22528 = pi18 ? n22036 : n22527;
  assign n22529 = pi17 ? n22033 : n22528;
  assign n22530 = pi16 ? n22030 : n22529;
  assign n22531 = pi15 ? n22524 : n22530;
  assign n22532 = pi14 ? n22521 : n22531;
  assign n22533 = pi13 ? n22507 : n22532;
  assign n22534 = pi18 ? n22053 : n15164;
  assign n22535 = pi17 ? n22050 : n22534;
  assign n22536 = pi16 ? n439 : n22535;
  assign n22537 = pi20 ? n37 : n17777;
  assign n22538 = pi19 ? n37 : n22537;
  assign n22539 = pi18 ? n22057 : n22538;
  assign n22540 = pi17 ? n22539 : n22064;
  assign n22541 = pi16 ? n439 : n22540;
  assign n22542 = pi15 ? n22536 : n22541;
  assign n22543 = pi14 ? n22542 : n22095;
  assign n22544 = pi21 ? n716 : n4548;
  assign n22545 = pi20 ? n32 : n22544;
  assign n22546 = pi19 ? n32 : n22545;
  assign n22547 = pi21 ? n335 : n99;
  assign n22548 = pi20 ? n22547 : n22114;
  assign n22549 = pi22 ? n363 : n99;
  assign n22550 = pi21 ? n22549 : n22118;
  assign n22551 = pi21 ? n3746 : n22118;
  assign n22552 = pi20 ? n22550 : n22551;
  assign n22553 = pi19 ? n22548 : n22552;
  assign n22554 = pi18 ? n22546 : n22553;
  assign n22555 = pi17 ? n32 : n22554;
  assign n22556 = pi22 ? n335 : n1656;
  assign n22557 = pi22 ? n4543 : n363;
  assign n22558 = pi21 ? n22556 : n22557;
  assign n22559 = pi20 ? n22551 : n22558;
  assign n22560 = pi22 ? n18461 : n4537;
  assign n22561 = pi21 ? n22560 : n3746;
  assign n22562 = pi20 ? n22129 : n22561;
  assign n22563 = pi19 ? n22559 : n22562;
  assign n22564 = pi21 ? n722 : n18462;
  assign n22565 = pi21 ? n722 : n18467;
  assign n22566 = pi20 ? n22564 : n22565;
  assign n22567 = pi19 ? n22566 : n21206;
  assign n22568 = pi18 ? n22563 : n22567;
  assign n22569 = pi22 ? n1656 : n233;
  assign n22570 = pi21 ? n22569 : n233;
  assign n22571 = pi20 ? n233 : n22570;
  assign n22572 = pi22 ? n233 : n4543;
  assign n22573 = pi21 ? n22572 : n233;
  assign n22574 = pi22 ? n4543 : n233;
  assign n22575 = pi21 ? n2707 : n22574;
  assign n22576 = pi20 ? n22573 : n22575;
  assign n22577 = pi19 ? n22571 : n22576;
  assign n22578 = pi18 ? n22577 : n22148;
  assign n22579 = pi17 ? n22568 : n22578;
  assign n22580 = pi16 ? n22555 : n22579;
  assign n22581 = pi15 ? n22108 : n22580;
  assign n22582 = pi21 ? n12635 : n2637;
  assign n22583 = pi20 ? n22582 : n32;
  assign n22584 = pi19 ? n22583 : n32;
  assign n22585 = pi18 ? n233 : n22584;
  assign n22586 = pi17 ? n21244 : n22585;
  assign n22587 = pi16 ? n22167 : n22586;
  assign n22588 = pi15 ? n22163 : n22587;
  assign n22589 = pi14 ? n22581 : n22588;
  assign n22590 = pi13 ? n22543 : n22589;
  assign n22591 = pi12 ? n22533 : n22590;
  assign n22592 = pi11 ? n22483 : n22591;
  assign n22593 = pi10 ? n22343 : n22592;
  assign n22594 = pi09 ? n22184 : n22593;
  assign n22595 = pi08 ? n22177 : n22594;
  assign n22596 = pi07 ? n21578 : n22595;
  assign n22597 = pi06 ? n20620 : n22596;
  assign n22598 = pi05 ? n18828 : n22597;
  assign n22599 = pi04 ? n14814 : n22598;
  assign n22600 = pi03 ? n7281 : n22599;
  assign n22601 = pi20 ? n37 : n8517;
  assign n22602 = pi19 ? n22601 : n32;
  assign n22603 = pi18 ? n37 : n22602;
  assign n22604 = pi17 ? n37 : n22603;
  assign n22605 = pi16 ? n13561 : n22604;
  assign n22606 = pi15 ? n32 : n22605;
  assign n22607 = pi20 ? n37 : n8530;
  assign n22608 = pi19 ? n22607 : n32;
  assign n22609 = pi18 ? n37 : n22608;
  assign n22610 = pi17 ? n37 : n22609;
  assign n22611 = pi16 ? n13561 : n22610;
  assign n22612 = pi16 ? n14445 : n22610;
  assign n22613 = pi15 ? n22611 : n22612;
  assign n22614 = pi14 ? n22606 : n22613;
  assign n22615 = pi13 ? n32 : n22614;
  assign n22616 = pi12 ? n32 : n22615;
  assign n22617 = pi11 ? n32 : n22616;
  assign n22618 = pi10 ? n32 : n22617;
  assign n22619 = pi21 ? n92 : n2168;
  assign n22620 = pi20 ? n32 : n22619;
  assign n22621 = pi19 ? n32 : n22620;
  assign n22622 = pi20 ? n2968 : n2185;
  assign n22623 = pi19 ? n22622 : n2963;
  assign n22624 = pi18 ? n22621 : n22623;
  assign n22625 = pi17 ? n32 : n22624;
  assign n22626 = pi19 ? n2969 : n2755;
  assign n22627 = pi20 ? n11424 : n3805;
  assign n22628 = pi19 ? n22627 : n2185;
  assign n22629 = pi18 ? n22626 : n22628;
  assign n22630 = pi20 ? n11424 : n3824;
  assign n22631 = pi19 ? n22630 : n3824;
  assign n22632 = pi21 ? n181 : n2162;
  assign n22633 = pi21 ? n218 : n3022;
  assign n22634 = pi20 ? n22632 : n22633;
  assign n22635 = pi19 ? n22634 : n32;
  assign n22636 = pi18 ? n22631 : n22635;
  assign n22637 = pi17 ? n22629 : n22636;
  assign n22638 = pi16 ? n22625 : n22637;
  assign n22639 = pi20 ? n14513 : n21633;
  assign n22640 = pi20 ? n6044 : n3824;
  assign n22641 = pi19 ? n22639 : n22640;
  assign n22642 = pi18 ? n21610 : n22641;
  assign n22643 = pi17 ? n32 : n22642;
  assign n22644 = pi21 ? n2156 : n2161;
  assign n22645 = pi20 ? n22644 : n3814;
  assign n22646 = pi19 ? n22645 : n21643;
  assign n22647 = pi20 ? n3884 : n2970;
  assign n22648 = pi19 ? n22647 : n21633;
  assign n22649 = pi18 ? n22646 : n22648;
  assign n22650 = pi20 ? n3884 : n3041;
  assign n22651 = pi21 ? n2156 : n2164;
  assign n22652 = pi19 ? n22650 : n22651;
  assign n22653 = pi21 ? n2164 : n3066;
  assign n22654 = pi20 ? n21638 : n22653;
  assign n22655 = pi19 ? n22654 : n32;
  assign n22656 = pi18 ? n22652 : n22655;
  assign n22657 = pi17 ? n22649 : n22656;
  assign n22658 = pi16 ? n22643 : n22657;
  assign n22659 = pi15 ? n22638 : n22658;
  assign n22660 = pi20 ? n14524 : n14510;
  assign n22661 = pi20 ? n2982 : n14513;
  assign n22662 = pi19 ? n22660 : n22661;
  assign n22663 = pi18 ? n17008 : n22662;
  assign n22664 = pi17 ? n32 : n22663;
  assign n22665 = pi19 ? n14519 : n16999;
  assign n22666 = pi21 ? n2175 : n37;
  assign n22667 = pi19 ? n21639 : n22666;
  assign n22668 = pi18 ? n22665 : n22667;
  assign n22669 = pi20 ? n14524 : n21643;
  assign n22670 = pi19 ? n22669 : n2958;
  assign n22671 = pi21 ? n181 : n8557;
  assign n22672 = pi20 ? n3041 : n22671;
  assign n22673 = pi19 ? n22672 : n32;
  assign n22674 = pi18 ? n22670 : n22673;
  assign n22675 = pi17 ? n22668 : n22674;
  assign n22676 = pi16 ? n22664 : n22675;
  assign n22677 = pi20 ? n37 : n22671;
  assign n22678 = pi19 ? n22677 : n32;
  assign n22679 = pi18 ? n37 : n22678;
  assign n22680 = pi17 ? n37 : n22679;
  assign n22681 = pi16 ? n439 : n22680;
  assign n22682 = pi15 ? n22676 : n22681;
  assign n22683 = pi14 ? n22659 : n22682;
  assign n22684 = pi20 ? n2961 : n6044;
  assign n22685 = pi20 ? n3825 : n99;
  assign n22686 = pi19 ? n22684 : n22685;
  assign n22687 = pi18 ? n2159 : n22686;
  assign n22688 = pi17 ? n32 : n22687;
  assign n22689 = pi21 ? n99 : n8044;
  assign n22690 = pi20 ? n99 : n22689;
  assign n22691 = pi19 ? n22690 : n32;
  assign n22692 = pi18 ? n99 : n22691;
  assign n22693 = pi17 ? n99 : n22692;
  assign n22694 = pi16 ? n22688 : n22693;
  assign n22695 = pi21 ? n180 : n2957;
  assign n22696 = pi20 ? n32 : n22695;
  assign n22697 = pi19 ? n32 : n22696;
  assign n22698 = pi18 ? n22697 : n21612;
  assign n22699 = pi17 ? n32 : n22698;
  assign n22700 = pi16 ? n22699 : n22693;
  assign n22701 = pi15 ? n22694 : n22700;
  assign n22702 = pi20 ? n99 : n14846;
  assign n22703 = pi19 ? n22702 : n139;
  assign n22704 = pi20 ? n14846 : n139;
  assign n22705 = pi19 ? n22704 : n139;
  assign n22706 = pi18 ? n22703 : n22705;
  assign n22707 = pi20 ? n139 : n8088;
  assign n22708 = pi19 ? n22707 : n32;
  assign n22709 = pi18 ? n139 : n22708;
  assign n22710 = pi17 ? n22706 : n22709;
  assign n22711 = pi16 ? n744 : n22710;
  assign n22712 = pi20 ? n139 : n8095;
  assign n22713 = pi19 ? n22712 : n32;
  assign n22714 = pi18 ? n139 : n22713;
  assign n22715 = pi17 ? n22706 : n22714;
  assign n22716 = pi16 ? n744 : n22715;
  assign n22717 = pi15 ? n22711 : n22716;
  assign n22718 = pi14 ? n22701 : n22717;
  assign n22719 = pi13 ? n22683 : n22718;
  assign n22720 = pi21 ? n326 : n4221;
  assign n22721 = pi20 ? n32 : n22720;
  assign n22722 = pi19 ? n32 : n22721;
  assign n22723 = pi21 ? n4234 : n4236;
  assign n22724 = pi20 ? n11734 : n22723;
  assign n22725 = pi21 ? n4234 : n837;
  assign n22726 = pi21 ? n812 : n825;
  assign n22727 = pi20 ? n22725 : n22726;
  assign n22728 = pi19 ? n22724 : n22727;
  assign n22729 = pi18 ? n22722 : n22728;
  assign n22730 = pi17 ? n32 : n22729;
  assign n22731 = pi21 ? n4252 : n825;
  assign n22732 = pi20 ? n22731 : n139;
  assign n22733 = pi19 ? n22732 : n139;
  assign n22734 = pi18 ? n22733 : n139;
  assign n22735 = pi20 ? n139 : n9798;
  assign n22736 = pi19 ? n22735 : n32;
  assign n22737 = pi18 ? n139 : n22736;
  assign n22738 = pi17 ? n22734 : n22737;
  assign n22739 = pi16 ? n22730 : n22738;
  assign n22740 = pi16 ? n331 : n22218;
  assign n22741 = pi15 ? n22739 : n22740;
  assign n22742 = pi20 ? n297 : n997;
  assign n22743 = pi19 ? n22742 : n20722;
  assign n22744 = pi18 ? n1692 : n22743;
  assign n22745 = pi17 ? n32 : n22744;
  assign n22746 = pi19 ? n14962 : n139;
  assign n22747 = pi18 ? n22746 : n139;
  assign n22748 = pi17 ? n22747 : n22217;
  assign n22749 = pi16 ? n22745 : n22748;
  assign n22750 = pi18 ? n374 : n19855;
  assign n22751 = pi17 ? n32 : n22750;
  assign n22752 = pi18 ? n37 : n10642;
  assign n22753 = pi18 ? n13183 : n22224;
  assign n22754 = pi17 ? n22752 : n22753;
  assign n22755 = pi16 ? n22751 : n22754;
  assign n22756 = pi15 ? n22749 : n22755;
  assign n22757 = pi14 ? n22741 : n22756;
  assign n22758 = pi19 ? n37 : n4733;
  assign n22759 = pi21 ? n363 : n928;
  assign n22760 = pi20 ? n139 : n22759;
  assign n22761 = pi19 ? n22760 : n32;
  assign n22762 = pi18 ? n22758 : n22761;
  assign n22763 = pi17 ? n37 : n22762;
  assign n22764 = pi16 ? n439 : n22763;
  assign n22765 = pi18 ? n14115 : n22761;
  assign n22766 = pi17 ? n37 : n22765;
  assign n22767 = pi16 ? n439 : n22766;
  assign n22768 = pi15 ? n22764 : n22767;
  assign n22769 = pi19 ? n37 : n18969;
  assign n22770 = pi20 ? n204 : n18386;
  assign n22771 = pi19 ? n22770 : n32;
  assign n22772 = pi18 ? n22769 : n22771;
  assign n22773 = pi17 ? n37 : n22772;
  assign n22774 = pi16 ? n439 : n22773;
  assign n22775 = pi20 ? n1912 : n204;
  assign n22776 = pi19 ? n37 : n22775;
  assign n22777 = pi21 ? n204 : n2553;
  assign n22778 = pi20 ? n204 : n22777;
  assign n22779 = pi19 ? n22778 : n32;
  assign n22780 = pi18 ? n22776 : n22779;
  assign n22781 = pi17 ? n37 : n22780;
  assign n22782 = pi16 ? n439 : n22781;
  assign n22783 = pi15 ? n22774 : n22782;
  assign n22784 = pi14 ? n22768 : n22783;
  assign n22785 = pi13 ? n22757 : n22784;
  assign n22786 = pi12 ? n22719 : n22785;
  assign n22787 = pi20 ? n997 : n37;
  assign n22788 = pi19 ? n22787 : n3096;
  assign n22789 = pi18 ? n3597 : n22788;
  assign n22790 = pi17 ? n32 : n22789;
  assign n22791 = pi20 ? n992 : n941;
  assign n22792 = pi20 ? n941 : n939;
  assign n22793 = pi19 ? n22791 : n22792;
  assign n22794 = pi20 ? n939 : n942;
  assign n22795 = pi19 ? n940 : n22794;
  assign n22796 = pi18 ? n22793 : n22795;
  assign n22797 = pi20 ? n139 : n8748;
  assign n22798 = pi19 ? n22797 : n32;
  assign n22799 = pi18 ? n139 : n22798;
  assign n22800 = pi17 ? n22796 : n22799;
  assign n22801 = pi16 ? n22790 : n22800;
  assign n22802 = pi20 ? n1912 : n21092;
  assign n22803 = pi19 ? n37 : n22802;
  assign n22804 = pi21 ? n19337 : n11808;
  assign n22805 = pi21 ? n11808 : n32;
  assign n22806 = pi20 ? n22804 : n22805;
  assign n22807 = pi19 ? n22806 : n32;
  assign n22808 = pi18 ? n22803 : n22807;
  assign n22809 = pi17 ? n37 : n22808;
  assign n22810 = pi16 ? n439 : n22809;
  assign n22811 = pi15 ? n22801 : n22810;
  assign n22812 = pi20 ? n569 : n335;
  assign n22813 = pi19 ? n7685 : n22812;
  assign n22814 = pi21 ? n2061 : n32;
  assign n22815 = pi20 ? n335 : n22814;
  assign n22816 = pi19 ? n22815 : n32;
  assign n22817 = pi18 ? n22813 : n22816;
  assign n22818 = pi17 ? n37 : n22817;
  assign n22819 = pi16 ? n439 : n22818;
  assign n22820 = pi18 ? n21770 : n22816;
  assign n22821 = pi17 ? n37 : n22820;
  assign n22822 = pi16 ? n439 : n22821;
  assign n22823 = pi15 ? n22819 : n22822;
  assign n22824 = pi14 ? n22811 : n22823;
  assign n22825 = pi18 ? n17205 : n22816;
  assign n22826 = pi17 ? n37 : n22825;
  assign n22827 = pi16 ? n439 : n22826;
  assign n22828 = pi20 ? n335 : n8849;
  assign n22829 = pi19 ? n22828 : n32;
  assign n22830 = pi18 ? n10682 : n22829;
  assign n22831 = pi17 ? n37 : n22830;
  assign n22832 = pi16 ? n439 : n22831;
  assign n22833 = pi15 ? n22827 : n22832;
  assign n22834 = pi14 ? n22833 : n22832;
  assign n22835 = pi13 ? n22824 : n22834;
  assign n22836 = pi21 ? n11336 : n32;
  assign n22837 = pi20 ? n569 : n22836;
  assign n22838 = pi19 ? n22837 : n32;
  assign n22839 = pi18 ? n37 : n22838;
  assign n22840 = pi17 ? n37 : n22839;
  assign n22841 = pi16 ? n439 : n22840;
  assign n22842 = pi22 ? n583 : n685;
  assign n22843 = pi21 ? n22842 : n32;
  assign n22844 = pi20 ? n37 : n22843;
  assign n22845 = pi19 ? n22844 : n32;
  assign n22846 = pi18 ? n37 : n22845;
  assign n22847 = pi17 ? n37 : n22846;
  assign n22848 = pi16 ? n439 : n22847;
  assign n22849 = pi15 ? n22841 : n22848;
  assign n22850 = pi20 ? n2091 : n17905;
  assign n22851 = pi19 ? n22850 : n32;
  assign n22852 = pi18 ? n2102 : n22851;
  assign n22853 = pi17 ? n37 : n22852;
  assign n22854 = pi16 ? n439 : n22853;
  assign n22855 = pi20 ? n2091 : n19439;
  assign n22856 = pi19 ? n22855 : n32;
  assign n22857 = pi18 ? n2102 : n22856;
  assign n22858 = pi17 ? n37 : n22857;
  assign n22859 = pi16 ? n439 : n22858;
  assign n22860 = pi15 ? n22854 : n22859;
  assign n22861 = pi14 ? n22849 : n22860;
  assign n22862 = pi20 ? n3393 : n11243;
  assign n22863 = pi19 ? n22862 : n32;
  assign n22864 = pi18 ? n37 : n22863;
  assign n22865 = pi17 ? n37 : n22864;
  assign n22866 = pi16 ? n439 : n22865;
  assign n22867 = pi20 ? n9660 : n9963;
  assign n22868 = pi19 ? n22867 : n32;
  assign n22869 = pi18 ? n37 : n22868;
  assign n22870 = pi17 ? n37 : n22869;
  assign n22871 = pi16 ? n439 : n22870;
  assign n22872 = pi15 ? n22866 : n22871;
  assign n22873 = pi20 ? n37 : n9963;
  assign n22874 = pi19 ? n22873 : n32;
  assign n22875 = pi18 ? n37 : n22874;
  assign n22876 = pi17 ? n37 : n22875;
  assign n22877 = pi16 ? n439 : n22876;
  assign n22878 = pi20 ? n37 : n9660;
  assign n22879 = pi19 ? n37 : n22878;
  assign n22880 = pi18 ? n22879 : n37;
  assign n22881 = pi21 ? n363 : n37;
  assign n22882 = pi20 ? n3393 : n22881;
  assign n22883 = pi20 ? n7730 : n363;
  assign n22884 = pi19 ? n22882 : n22883;
  assign n22885 = pi22 ? n363 : n2468;
  assign n22886 = pi21 ? n22885 : n32;
  assign n22887 = pi20 ? n363 : n22886;
  assign n22888 = pi19 ? n22887 : n32;
  assign n22889 = pi18 ? n22884 : n22888;
  assign n22890 = pi17 ? n22880 : n22889;
  assign n22891 = pi16 ? n439 : n22890;
  assign n22892 = pi15 ? n22877 : n22891;
  assign n22893 = pi14 ? n22872 : n22892;
  assign n22894 = pi13 ? n22861 : n22893;
  assign n22895 = pi12 ? n22835 : n22894;
  assign n22896 = pi11 ? n22786 : n22895;
  assign n22897 = pi20 ? n3393 : n363;
  assign n22898 = pi19 ? n22897 : n363;
  assign n22899 = pi21 ? n13687 : n32;
  assign n22900 = pi20 ? n363 : n22899;
  assign n22901 = pi19 ? n22900 : n32;
  assign n22902 = pi18 ? n22898 : n22901;
  assign n22903 = pi17 ? n22880 : n22902;
  assign n22904 = pi16 ? n439 : n22903;
  assign n22905 = pi18 ? n8040 : n37;
  assign n22906 = pi21 ? n10488 : n363;
  assign n22907 = pi20 ? n7332 : n22906;
  assign n22908 = pi21 ? n9666 : n3392;
  assign n22909 = pi20 ? n363 : n22908;
  assign n22910 = pi19 ? n22907 : n22909;
  assign n22911 = pi22 ? n157 : n532;
  assign n22912 = pi21 ? n22911 : n32;
  assign n22913 = pi20 ? n363 : n22912;
  assign n22914 = pi19 ? n22913 : n32;
  assign n22915 = pi18 ? n22910 : n22914;
  assign n22916 = pi17 ? n22905 : n22915;
  assign n22917 = pi16 ? n439 : n22916;
  assign n22918 = pi15 ? n22904 : n22917;
  assign n22919 = pi22 ? n685 : n625;
  assign n22920 = pi21 ? n22919 : n32;
  assign n22921 = pi20 ? n2107 : n22920;
  assign n22922 = pi19 ? n22921 : n32;
  assign n22923 = pi18 ? n37 : n22922;
  assign n22924 = pi17 ? n37 : n22923;
  assign n22925 = pi16 ? n439 : n22924;
  assign n22926 = pi14 ? n22918 : n22925;
  assign n22927 = pi20 ? n7754 : n9482;
  assign n22928 = pi19 ? n22927 : n32;
  assign n22929 = pi18 ? n99 : n22928;
  assign n22930 = pi17 ? n99 : n22929;
  assign n22931 = pi16 ? n744 : n22930;
  assign n22932 = pi16 ? n744 : n22368;
  assign n22933 = pi15 ? n22931 : n22932;
  assign n22934 = pi21 ? n99 : n21842;
  assign n22935 = pi20 ? n22934 : n8295;
  assign n22936 = pi19 ? n22935 : n32;
  assign n22937 = pi18 ? n99 : n22936;
  assign n22938 = pi17 ? n99 : n22937;
  assign n22939 = pi16 ? n744 : n22938;
  assign n22940 = pi22 ? n99 : n19177;
  assign n22941 = pi21 ? n99 : n22940;
  assign n22942 = pi20 ? n22941 : n4008;
  assign n22943 = pi19 ? n22942 : n32;
  assign n22944 = pi18 ? n99 : n22943;
  assign n22945 = pi17 ? n99 : n22944;
  assign n22946 = pi16 ? n744 : n22945;
  assign n22947 = pi15 ? n22939 : n22946;
  assign n22948 = pi14 ? n22933 : n22947;
  assign n22949 = pi13 ? n22926 : n22948;
  assign n22950 = pi20 ? n802 : n2238;
  assign n22951 = pi19 ? n2255 : n22950;
  assign n22952 = pi21 ? n777 : n22940;
  assign n22953 = pi20 ? n22952 : n3210;
  assign n22954 = pi19 ? n22953 : n32;
  assign n22955 = pi18 ? n22951 : n22954;
  assign n22956 = pi17 ? n99 : n22955;
  assign n22957 = pi16 ? n744 : n22956;
  assign n22958 = pi19 ? n99 : n14285;
  assign n22959 = pi20 ? n2243 : n3210;
  assign n22960 = pi19 ? n22959 : n32;
  assign n22961 = pi18 ? n22958 : n22960;
  assign n22962 = pi17 ? n99 : n22961;
  assign n22963 = pi16 ? n744 : n22962;
  assign n22964 = pi15 ? n22957 : n22963;
  assign n22965 = pi21 ? n99 : n17375;
  assign n22966 = pi20 ? n22965 : n99;
  assign n22967 = pi19 ? n99 : n22966;
  assign n22968 = pi20 ? n19171 : n2653;
  assign n22969 = pi19 ? n22968 : n32;
  assign n22970 = pi18 ? n22967 : n22969;
  assign n22971 = pi17 ? n99 : n22970;
  assign n22972 = pi16 ? n744 : n22971;
  assign n22973 = pi20 ? n259 : n282;
  assign n22974 = pi21 ? n248 : n168;
  assign n22975 = pi20 ? n7429 : n22974;
  assign n22976 = pi19 ? n22973 : n22975;
  assign n22977 = pi21 ? n258 : n3562;
  assign n22978 = pi20 ? n22977 : n2653;
  assign n22979 = pi19 ? n22978 : n32;
  assign n22980 = pi18 ? n22976 : n22979;
  assign n22981 = pi17 ? n157 : n22980;
  assign n22982 = pi16 ? n5910 : n22981;
  assign n22983 = pi15 ? n22972 : n22982;
  assign n22984 = pi14 ? n22964 : n22983;
  assign n22985 = pi20 ? n1786 : n9773;
  assign n22986 = pi19 ? n139 : n22985;
  assign n22987 = pi18 ? n22986 : n139;
  assign n22988 = pi20 ? n316 : n2653;
  assign n22989 = pi19 ? n22988 : n32;
  assign n22990 = pi18 ? n10073 : n22989;
  assign n22991 = pi17 ? n22987 : n22990;
  assign n22992 = pi16 ? n915 : n22991;
  assign n22993 = pi20 ? n204 : n2884;
  assign n22994 = pi19 ? n204 : n22993;
  assign n22995 = pi18 ? n2394 : n22994;
  assign n22996 = pi17 ? n32 : n22995;
  assign n22997 = pi21 ? n2427 : n2402;
  assign n22998 = pi20 ? n2884 : n22997;
  assign n22999 = pi19 ? n2884 : n22998;
  assign n23000 = pi21 ? n20102 : n2427;
  assign n23001 = pi22 ? n2401 : n2299;
  assign n23002 = pi21 ? n204 : n23001;
  assign n23003 = pi21 ? n204 : n1578;
  assign n23004 = pi20 ? n23002 : n23003;
  assign n23005 = pi19 ? n23000 : n23004;
  assign n23006 = pi18 ? n22999 : n23005;
  assign n23007 = pi21 ? n522 : n1027;
  assign n23008 = pi20 ? n23007 : n2383;
  assign n23009 = pi19 ? n23008 : n316;
  assign n23010 = pi18 ? n23009 : n22989;
  assign n23011 = pi17 ? n23006 : n23010;
  assign n23012 = pi16 ? n22996 : n23011;
  assign n23013 = pi15 ? n22992 : n23012;
  assign n23014 = pi21 ? n921 : n316;
  assign n23015 = pi20 ? n204 : n23014;
  assign n23016 = pi19 ? n23015 : n6645;
  assign n23017 = pi20 ? n2353 : n2653;
  assign n23018 = pi19 ? n23017 : n32;
  assign n23019 = pi18 ? n23016 : n23018;
  assign n23020 = pi17 ? n204 : n23019;
  assign n23021 = pi16 ? n13493 : n23020;
  assign n23022 = pi21 ? n204 : n1313;
  assign n23023 = pi20 ? n23022 : n204;
  assign n23024 = pi19 ? n23023 : n204;
  assign n23025 = pi18 ? n204 : n23024;
  assign n23026 = pi19 ? n20033 : n316;
  assign n23027 = pi18 ? n23026 : n22989;
  assign n23028 = pi17 ? n23025 : n23027;
  assign n23029 = pi16 ? n13846 : n23028;
  assign n23030 = pi15 ? n23021 : n23029;
  assign n23031 = pi14 ? n23013 : n23030;
  assign n23032 = pi13 ? n22984 : n23031;
  assign n23033 = pi12 ? n22949 : n23032;
  assign n23034 = pi20 ? n975 : n2653;
  assign n23035 = pi19 ? n23034 : n32;
  assign n23036 = pi18 ? n139 : n23035;
  assign n23037 = pi17 ? n139 : n23036;
  assign n23038 = pi16 ? n1575 : n23037;
  assign n23039 = pi20 ? n1026 : n2318;
  assign n23040 = pi19 ? n23039 : n139;
  assign n23041 = pi21 ? n139 : n8869;
  assign n23042 = pi20 ? n23041 : n2653;
  assign n23043 = pi19 ? n23042 : n32;
  assign n23044 = pi18 ? n23040 : n23043;
  assign n23045 = pi17 ? n139 : n23044;
  assign n23046 = pi16 ? n331 : n23045;
  assign n23047 = pi15 ? n23038 : n23046;
  assign n23048 = pi21 ? n139 : n11336;
  assign n23049 = pi20 ? n23048 : n32;
  assign n23050 = pi19 ? n23049 : n32;
  assign n23051 = pi18 ? n139 : n23050;
  assign n23052 = pi17 ? n139 : n23051;
  assign n23053 = pi16 ? n915 : n23052;
  assign n23054 = pi19 ? n139 : n15402;
  assign n23055 = pi20 ? n7858 : n32;
  assign n23056 = pi19 ? n23055 : n32;
  assign n23057 = pi18 ? n23054 : n23056;
  assign n23058 = pi17 ? n139 : n23057;
  assign n23059 = pi16 ? n915 : n23058;
  assign n23060 = pi15 ? n23053 : n23059;
  assign n23061 = pi14 ? n23047 : n23060;
  assign n23062 = pi20 ? n3311 : n7980;
  assign n23063 = pi19 ? n23062 : n6749;
  assign n23064 = pi18 ? n23063 : n23056;
  assign n23065 = pi17 ? n335 : n23064;
  assign n23066 = pi16 ? n7943 : n23065;
  assign n23067 = pi21 ? n233 : n204;
  assign n23068 = pi20 ? n335 : n23067;
  assign n23069 = pi21 ? n204 : n233;
  assign n23070 = pi20 ? n23069 : n7980;
  assign n23071 = pi19 ? n23068 : n23070;
  assign n23072 = pi21 ? n233 : n12381;
  assign n23073 = pi20 ? n23072 : n32;
  assign n23074 = pi19 ? n23073 : n32;
  assign n23075 = pi18 ? n23071 : n23074;
  assign n23076 = pi17 ? n335 : n23075;
  assign n23077 = pi16 ? n2035 : n23076;
  assign n23078 = pi15 ? n23066 : n23077;
  assign n23079 = pi19 ? n335 : n15488;
  assign n23080 = pi18 ? n23079 : n22022;
  assign n23081 = pi17 ? n335 : n23080;
  assign n23082 = pi16 ? n7943 : n23081;
  assign n23083 = pi18 ? n374 : n17476;
  assign n23084 = pi17 ? n32 : n23083;
  assign n23085 = pi18 ? n335 : n13259;
  assign n23086 = pi17 ? n335 : n23085;
  assign n23087 = pi16 ? n23084 : n23086;
  assign n23088 = pi15 ? n23082 : n23087;
  assign n23089 = pi14 ? n23078 : n23088;
  assign n23090 = pi13 ? n23061 : n23089;
  assign n23091 = pi19 ? n37 : n10957;
  assign n23092 = pi18 ? n23091 : n10682;
  assign n23093 = pi21 ? n233 : n650;
  assign n23094 = pi20 ? n23093 : n32;
  assign n23095 = pi19 ? n23094 : n32;
  assign n23096 = pi18 ? n17552 : n23095;
  assign n23097 = pi17 ? n23092 : n23096;
  assign n23098 = pi16 ? n439 : n23097;
  assign n23099 = pi21 ? n335 : n4893;
  assign n23100 = pi20 ? n23099 : n13527;
  assign n23101 = pi19 ? n23100 : n233;
  assign n23102 = pi18 ? n23101 : n23095;
  assign n23103 = pi17 ? n14165 : n23102;
  assign n23104 = pi16 ? n439 : n23103;
  assign n23105 = pi15 ? n23098 : n23104;
  assign n23106 = pi18 ? n15128 : n7686;
  assign n23107 = pi21 ? n233 : n13280;
  assign n23108 = pi20 ? n23107 : n32;
  assign n23109 = pi19 ? n23108 : n32;
  assign n23110 = pi18 ? n233 : n23109;
  assign n23111 = pi17 ? n23106 : n23110;
  assign n23112 = pi16 ? n439 : n23111;
  assign n23113 = pi18 ? n335 : n15082;
  assign n23114 = pi19 ? n13527 : n17542;
  assign n23115 = pi21 ? n233 : n696;
  assign n23116 = pi20 ? n23115 : n32;
  assign n23117 = pi19 ? n23116 : n32;
  assign n23118 = pi18 ? n23114 : n23117;
  assign n23119 = pi17 ? n23113 : n23118;
  assign n23120 = pi16 ? n3351 : n23119;
  assign n23121 = pi15 ? n23112 : n23120;
  assign n23122 = pi14 ? n23105 : n23121;
  assign n23123 = pi21 ? n363 : n335;
  assign n23124 = pi20 ? n23123 : n335;
  assign n23125 = pi19 ? n335 : n23124;
  assign n23126 = pi18 ? n17530 : n23125;
  assign n23127 = pi17 ? n32 : n23126;
  assign n23128 = pi21 ? n363 : n6376;
  assign n23129 = pi21 ? n16562 : n335;
  assign n23130 = pi20 ? n23128 : n23129;
  assign n23131 = pi19 ? n21200 : n23130;
  assign n23132 = pi21 ? n3746 : n17548;
  assign n23133 = pi21 ? n335 : n722;
  assign n23134 = pi20 ? n23132 : n23133;
  assign n23135 = pi21 ? n17548 : n233;
  assign n23136 = pi20 ? n19422 : n23135;
  assign n23137 = pi19 ? n23134 : n23136;
  assign n23138 = pi18 ? n23131 : n23137;
  assign n23139 = pi20 ? n233 : n16530;
  assign n23140 = pi19 ? n233 : n23139;
  assign n23141 = pi21 ? n4900 : n3523;
  assign n23142 = pi20 ? n23141 : n32;
  assign n23143 = pi19 ? n23142 : n32;
  assign n23144 = pi18 ? n23140 : n23143;
  assign n23145 = pi17 ? n23138 : n23144;
  assign n23146 = pi16 ? n23127 : n23145;
  assign n23147 = pi21 ? n716 : n363;
  assign n23148 = pi20 ? n32 : n23147;
  assign n23149 = pi19 ? n32 : n23148;
  assign n23150 = pi21 ? n22549 : n363;
  assign n23151 = pi20 ? n363 : n23150;
  assign n23152 = pi19 ? n363 : n23151;
  assign n23153 = pi18 ? n23149 : n23152;
  assign n23154 = pi17 ? n32 : n23153;
  assign n23155 = pi21 ? n363 : n2707;
  assign n23156 = pi23 ? n233 : n363;
  assign n23157 = pi22 ? n23156 : n363;
  assign n23158 = pi21 ? n23157 : n363;
  assign n23159 = pi20 ? n23155 : n23158;
  assign n23160 = pi19 ? n363 : n23159;
  assign n23161 = pi21 ? n22128 : n363;
  assign n23162 = pi21 ? n363 : n722;
  assign n23163 = pi20 ? n23161 : n23162;
  assign n23164 = pi19 ? n23163 : n19422;
  assign n23165 = pi18 ? n23160 : n23164;
  assign n23166 = pi18 ? n233 : n14228;
  assign n23167 = pi17 ? n23165 : n23166;
  assign n23168 = pi16 ? n23154 : n23167;
  assign n23169 = pi15 ? n23146 : n23168;
  assign n23170 = pi23 ? n21554 : n139;
  assign n23171 = pi22 ? n23170 : n363;
  assign n23172 = pi21 ? n23171 : n363;
  assign n23173 = pi20 ? n32 : n23172;
  assign n23174 = pi19 ? n32 : n23173;
  assign n23175 = pi21 ? n5014 : n363;
  assign n23176 = pi19 ? n363 : n23175;
  assign n23177 = pi18 ? n23174 : n23176;
  assign n23178 = pi17 ? n32 : n23177;
  assign n23179 = pi21 ? n233 : n2707;
  assign n23180 = pi20 ? n23179 : n23175;
  assign n23181 = pi19 ? n363 : n23180;
  assign n23182 = pi21 ? n20605 : n363;
  assign n23183 = pi20 ? n23182 : n5021;
  assign n23184 = pi19 ? n23183 : n15177;
  assign n23185 = pi18 ? n23181 : n23184;
  assign n23186 = pi22 ? n233 : n673;
  assign n23187 = pi21 ? n23186 : n5829;
  assign n23188 = pi20 ? n23187 : n32;
  assign n23189 = pi19 ? n23188 : n32;
  assign n23190 = pi18 ? n233 : n23189;
  assign n23191 = pi17 ? n23185 : n23190;
  assign n23192 = pi16 ? n23178 : n23191;
  assign n23193 = pi20 ? n15177 : n363;
  assign n23194 = pi19 ? n363 : n23193;
  assign n23195 = pi18 ? n23174 : n23194;
  assign n23196 = pi17 ? n32 : n23195;
  assign n23197 = pi20 ? n233 : n22153;
  assign n23198 = pi19 ? n363 : n23197;
  assign n23199 = pi21 ? n5014 : n2707;
  assign n23200 = pi20 ? n19422 : n23199;
  assign n23201 = pi19 ? n23200 : n233;
  assign n23202 = pi18 ? n23198 : n23201;
  assign n23203 = pi21 ? n233 : n2637;
  assign n23204 = pi20 ? n23203 : n32;
  assign n23205 = pi19 ? n23204 : n32;
  assign n23206 = pi18 ? n233 : n23205;
  assign n23207 = pi17 ? n23202 : n23206;
  assign n23208 = pi16 ? n23196 : n23207;
  assign n23209 = pi15 ? n23192 : n23208;
  assign n23210 = pi14 ? n23169 : n23209;
  assign n23211 = pi13 ? n23122 : n23210;
  assign n23212 = pi12 ? n23090 : n23211;
  assign n23213 = pi11 ? n23033 : n23212;
  assign n23214 = pi10 ? n22896 : n23213;
  assign n23215 = pi09 ? n22618 : n23214;
  assign n23216 = pi23 ? n20627 : n32;
  assign n23217 = pi22 ? n23216 : n32;
  assign n23218 = pi21 ? n37 : n23217;
  assign n23219 = pi20 ? n37 : n23218;
  assign n23220 = pi19 ? n23219 : n32;
  assign n23221 = pi18 ? n37 : n23220;
  assign n23222 = pi17 ? n37 : n23221;
  assign n23223 = pi16 ? n14445 : n23222;
  assign n23224 = pi15 ? n23223 : n22612;
  assign n23225 = pi14 ? n22606 : n23224;
  assign n23226 = pi13 ? n32 : n23225;
  assign n23227 = pi12 ? n32 : n23226;
  assign n23228 = pi11 ? n32 : n23227;
  assign n23229 = pi10 ? n32 : n23228;
  assign n23230 = pi22 ? n32 : n2160;
  assign n23231 = pi21 ? n23230 : n2168;
  assign n23232 = pi20 ? n32 : n23231;
  assign n23233 = pi19 ? n32 : n23232;
  assign n23234 = pi20 ? n2167 : n2755;
  assign n23235 = pi19 ? n23234 : n3808;
  assign n23236 = pi18 ? n23233 : n23235;
  assign n23237 = pi17 ? n32 : n23236;
  assign n23238 = pi20 ? n2749 : n2165;
  assign n23239 = pi19 ? n3813 : n23238;
  assign n23240 = pi20 ? n11424 : n3506;
  assign n23241 = pi19 ? n23240 : n2165;
  assign n23242 = pi18 ? n23239 : n23241;
  assign n23243 = pi21 ? n2746 : n2161;
  assign n23244 = pi20 ? n23243 : n3824;
  assign n23245 = pi19 ? n23244 : n2962;
  assign n23246 = pi20 ? n2752 : n22633;
  assign n23247 = pi19 ? n23246 : n32;
  assign n23248 = pi18 ? n23245 : n23247;
  assign n23249 = pi17 ? n23242 : n23248;
  assign n23250 = pi16 ? n23237 : n23249;
  assign n23251 = pi23 ? n32 : n714;
  assign n23252 = pi22 ? n23251 : n112;
  assign n23253 = pi21 ? n23252 : n2746;
  assign n23254 = pi20 ? n32 : n23253;
  assign n23255 = pi19 ? n32 : n23254;
  assign n23256 = pi21 ? n99 : n112;
  assign n23257 = pi20 ? n6043 : n23256;
  assign n23258 = pi20 ? n3807 : n3824;
  assign n23259 = pi19 ? n23257 : n23258;
  assign n23260 = pi18 ? n23255 : n23259;
  assign n23261 = pi17 ? n32 : n23260;
  assign n23262 = pi19 ? n22645 : n21633;
  assign n23263 = pi20 ? n3884 : n3870;
  assign n23264 = pi19 ? n23263 : n21633;
  assign n23265 = pi18 ? n23262 : n23264;
  assign n23266 = pi20 ? n3884 : n3877;
  assign n23267 = pi19 ? n23266 : n22651;
  assign n23268 = pi23 ? n8184 : n32;
  assign n23269 = pi22 ? n23268 : n32;
  assign n23270 = pi21 ? n2164 : n23269;
  assign n23271 = pi20 ? n21638 : n23270;
  assign n23272 = pi19 ? n23271 : n32;
  assign n23273 = pi18 ? n23267 : n23272;
  assign n23274 = pi17 ? n23265 : n23273;
  assign n23275 = pi16 ? n23261 : n23274;
  assign n23276 = pi15 ? n23250 : n23275;
  assign n23277 = pi20 ? n7346 : n2167;
  assign n23278 = pi20 ? n3805 : n6043;
  assign n23279 = pi19 ? n23277 : n23278;
  assign n23280 = pi18 ? n17008 : n23279;
  assign n23281 = pi17 ? n32 : n23280;
  assign n23282 = pi20 ? n6044 : n2962;
  assign n23283 = pi21 ? n1143 : n2168;
  assign n23284 = pi20 ? n5496 : n23283;
  assign n23285 = pi19 ? n23282 : n23284;
  assign n23286 = pi21 ? n1143 : n2164;
  assign n23287 = pi20 ? n23286 : n5496;
  assign n23288 = pi19 ? n23287 : n2169;
  assign n23289 = pi18 ? n23285 : n23288;
  assign n23290 = pi21 ? n99 : n2156;
  assign n23291 = pi20 ? n3824 : n23290;
  assign n23292 = pi19 ? n23291 : n2163;
  assign n23293 = pi21 ? n1143 : n8557;
  assign n23294 = pi20 ? n2164 : n23293;
  assign n23295 = pi19 ? n23294 : n32;
  assign n23296 = pi18 ? n23292 : n23295;
  assign n23297 = pi17 ? n23289 : n23296;
  assign n23298 = pi16 ? n23281 : n23297;
  assign n23299 = pi21 ? n180 : n2160;
  assign n23300 = pi20 ? n32 : n23299;
  assign n23301 = pi19 ? n32 : n23300;
  assign n23302 = pi20 ? n16008 : n37;
  assign n23303 = pi19 ? n23302 : n37;
  assign n23304 = pi18 ? n23301 : n23303;
  assign n23305 = pi17 ? n32 : n23304;
  assign n23306 = pi16 ? n23305 : n22680;
  assign n23307 = pi15 ? n23298 : n23306;
  assign n23308 = pi14 ? n23276 : n23307;
  assign n23309 = pi20 ? n6044 : n3807;
  assign n23310 = pi20 ? n2189 : n99;
  assign n23311 = pi19 ? n23309 : n23310;
  assign n23312 = pi18 ? n15526 : n23311;
  assign n23313 = pi17 ? n32 : n23312;
  assign n23314 = pi16 ? n23313 : n22693;
  assign n23315 = pi21 ? n1671 : n2168;
  assign n23316 = pi20 ? n32 : n23315;
  assign n23317 = pi19 ? n32 : n23316;
  assign n23318 = pi20 ? n3042 : n99;
  assign n23319 = pi19 ? n23318 : n99;
  assign n23320 = pi18 ? n23317 : n23319;
  assign n23321 = pi17 ? n32 : n23320;
  assign n23322 = pi21 ? n99 : n17044;
  assign n23323 = pi20 ? n99 : n23322;
  assign n23324 = pi19 ? n23323 : n32;
  assign n23325 = pi18 ? n99 : n23324;
  assign n23326 = pi17 ? n99 : n23325;
  assign n23327 = pi16 ? n23321 : n23326;
  assign n23328 = pi15 ? n23314 : n23327;
  assign n23329 = pi20 ? n139 : n23322;
  assign n23330 = pi19 ? n23329 : n32;
  assign n23331 = pi18 ? n139 : n23330;
  assign n23332 = pi17 ? n22706 : n23331;
  assign n23333 = pi16 ? n721 : n23332;
  assign n23334 = pi22 ? n206 : n32;
  assign n23335 = pi21 ? n99 : n23334;
  assign n23336 = pi20 ? n139 : n23335;
  assign n23337 = pi19 ? n23336 : n32;
  assign n23338 = pi18 ? n139 : n23337;
  assign n23339 = pi17 ? n22706 : n23338;
  assign n23340 = pi16 ? n721 : n23339;
  assign n23341 = pi15 ? n23333 : n23340;
  assign n23342 = pi14 ? n23328 : n23341;
  assign n23343 = pi13 ? n23308 : n23342;
  assign n23344 = pi21 ? n1549 : n813;
  assign n23345 = pi20 ? n32 : n23344;
  assign n23346 = pi19 ? n32 : n23345;
  assign n23347 = pi21 ? n1211 : n813;
  assign n23348 = pi21 ? n1211 : n4236;
  assign n23349 = pi20 ? n23347 : n23348;
  assign n23350 = pi21 ? n1211 : n831;
  assign n23351 = pi22 ? n812 : n1043;
  assign n23352 = pi21 ? n23351 : n825;
  assign n23353 = pi20 ? n23350 : n23352;
  assign n23354 = pi19 ? n23349 : n23353;
  assign n23355 = pi18 ? n23346 : n23354;
  assign n23356 = pi17 ? n32 : n23355;
  assign n23357 = pi21 ? n1711 : n825;
  assign n23358 = pi20 ? n23357 : n139;
  assign n23359 = pi19 ? n23358 : n139;
  assign n23360 = pi18 ? n23359 : n139;
  assign n23361 = pi23 ? n16890 : n32;
  assign n23362 = pi22 ? n23361 : n32;
  assign n23363 = pi21 ? n139 : n23362;
  assign n23364 = pi20 ? n139 : n23363;
  assign n23365 = pi19 ? n23364 : n32;
  assign n23366 = pi18 ? n139 : n23365;
  assign n23367 = pi17 ? n23360 : n23366;
  assign n23368 = pi16 ? n23356 : n23367;
  assign n23369 = pi23 ? n7393 : n32;
  assign n23370 = pi22 ? n23369 : n32;
  assign n23371 = pi21 ? n139 : n23370;
  assign n23372 = pi20 ? n139 : n23371;
  assign n23373 = pi19 ? n23372 : n32;
  assign n23374 = pi18 ? n139 : n23373;
  assign n23375 = pi17 ? n139 : n23374;
  assign n23376 = pi16 ? n331 : n23375;
  assign n23377 = pi15 ? n23368 : n23376;
  assign n23378 = pi17 ? n22747 : n23374;
  assign n23379 = pi16 ? n22745 : n23378;
  assign n23380 = pi23 ? n1748 : n32;
  assign n23381 = pi22 ? n23380 : n32;
  assign n23382 = pi21 ? n139 : n23381;
  assign n23383 = pi20 ? n139 : n23382;
  assign n23384 = pi19 ? n23383 : n32;
  assign n23385 = pi18 ? n13183 : n23384;
  assign n23386 = pi17 ? n22752 : n23385;
  assign n23387 = pi16 ? n22751 : n23386;
  assign n23388 = pi15 ? n23379 : n23387;
  assign n23389 = pi14 ? n23377 : n23388;
  assign n23390 = pi21 ? n204 : n2531;
  assign n23391 = pi20 ? n204 : n23390;
  assign n23392 = pi19 ? n23391 : n32;
  assign n23393 = pi18 ? n22769 : n23392;
  assign n23394 = pi17 ? n37 : n23393;
  assign n23395 = pi16 ? n439 : n23394;
  assign n23396 = pi15 ? n23395 : n22782;
  assign n23397 = pi14 ? n22768 : n23396;
  assign n23398 = pi13 ? n23389 : n23397;
  assign n23399 = pi12 ? n23343 : n23398;
  assign n23400 = pi21 ? n1793 : n2678;
  assign n23401 = pi20 ? n139 : n23400;
  assign n23402 = pi19 ? n23401 : n32;
  assign n23403 = pi18 ? n139 : n23402;
  assign n23404 = pi17 ? n22796 : n23403;
  assign n23405 = pi16 ? n22790 : n23404;
  assign n23406 = pi21 ? n11808 : n1009;
  assign n23407 = pi20 ? n22804 : n23406;
  assign n23408 = pi19 ? n23407 : n32;
  assign n23409 = pi18 ? n22803 : n23408;
  assign n23410 = pi17 ? n37 : n23409;
  assign n23411 = pi16 ? n439 : n23410;
  assign n23412 = pi15 ? n23405 : n23411;
  assign n23413 = pi14 ? n23412 : n22823;
  assign n23414 = pi13 ? n23413 : n22834;
  assign n23415 = pi21 ? n12983 : n32;
  assign n23416 = pi20 ? n2091 : n23415;
  assign n23417 = pi19 ? n23416 : n32;
  assign n23418 = pi18 ? n2102 : n23417;
  assign n23419 = pi17 ? n37 : n23418;
  assign n23420 = pi16 ? n439 : n23419;
  assign n23421 = pi15 ? n23420 : n22854;
  assign n23422 = pi14 ? n22849 : n23421;
  assign n23423 = pi20 ? n3393 : n12128;
  assign n23424 = pi19 ? n23423 : n32;
  assign n23425 = pi18 ? n37 : n23424;
  assign n23426 = pi17 ? n37 : n23425;
  assign n23427 = pi16 ? n439 : n23426;
  assign n23428 = pi15 ? n23427 : n22871;
  assign n23429 = pi20 ? n363 : n9949;
  assign n23430 = pi19 ? n23429 : n32;
  assign n23431 = pi18 ? n22884 : n23430;
  assign n23432 = pi17 ? n22880 : n23431;
  assign n23433 = pi16 ? n439 : n23432;
  assign n23434 = pi15 ? n22877 : n23433;
  assign n23435 = pi14 ? n23428 : n23434;
  assign n23436 = pi13 ? n23422 : n23435;
  assign n23437 = pi12 ? n23414 : n23436;
  assign n23438 = pi11 ? n23399 : n23437;
  assign n23439 = pi20 ? n363 : n9456;
  assign n23440 = pi19 ? n23439 : n32;
  assign n23441 = pi18 ? n22898 : n23440;
  assign n23442 = pi17 ? n22880 : n23441;
  assign n23443 = pi16 ? n439 : n23442;
  assign n23444 = pi20 ? n363 : n9957;
  assign n23445 = pi19 ? n23444 : n32;
  assign n23446 = pi18 ? n22910 : n23445;
  assign n23447 = pi17 ? n22905 : n23446;
  assign n23448 = pi16 ? n439 : n23447;
  assign n23449 = pi15 ? n23443 : n23448;
  assign n23450 = pi20 ? n2107 : n9456;
  assign n23451 = pi19 ? n23450 : n32;
  assign n23452 = pi18 ? n37 : n23451;
  assign n23453 = pi17 ? n37 : n23452;
  assign n23454 = pi16 ? n439 : n23453;
  assign n23455 = pi14 ? n23449 : n23454;
  assign n23456 = pi20 ? n7754 : n9456;
  assign n23457 = pi19 ? n23456 : n32;
  assign n23458 = pi18 ? n99 : n23457;
  assign n23459 = pi17 ? n99 : n23458;
  assign n23460 = pi16 ? n744 : n23459;
  assign n23461 = pi20 ? n5085 : n9456;
  assign n23462 = pi19 ? n23461 : n32;
  assign n23463 = pi18 ? n99 : n23462;
  assign n23464 = pi17 ? n99 : n23463;
  assign n23465 = pi16 ? n744 : n23464;
  assign n23466 = pi15 ? n23460 : n23465;
  assign n23467 = pi20 ? n22934 : n9963;
  assign n23468 = pi19 ? n23467 : n32;
  assign n23469 = pi18 ? n99 : n23468;
  assign n23470 = pi17 ? n99 : n23469;
  assign n23471 = pi16 ? n744 : n23470;
  assign n23472 = pi20 ? n22941 : n5667;
  assign n23473 = pi19 ? n23472 : n32;
  assign n23474 = pi18 ? n99 : n23473;
  assign n23475 = pi17 ? n99 : n23474;
  assign n23476 = pi16 ? n744 : n23475;
  assign n23477 = pi15 ? n23471 : n23476;
  assign n23478 = pi14 ? n23466 : n23477;
  assign n23479 = pi13 ? n23455 : n23478;
  assign n23480 = pi20 ? n19171 : n10011;
  assign n23481 = pi19 ? n23480 : n32;
  assign n23482 = pi18 ? n22967 : n23481;
  assign n23483 = pi17 ? n99 : n23482;
  assign n23484 = pi16 ? n744 : n23483;
  assign n23485 = pi20 ? n22977 : n10011;
  assign n23486 = pi19 ? n23485 : n32;
  assign n23487 = pi18 ? n22976 : n23486;
  assign n23488 = pi17 ? n157 : n23487;
  assign n23489 = pi16 ? n5910 : n23488;
  assign n23490 = pi15 ? n23484 : n23489;
  assign n23491 = pi14 ? n22964 : n23490;
  assign n23492 = pi21 ? n2391 : n2402;
  assign n23493 = pi20 ? n32 : n23492;
  assign n23494 = pi19 ? n32 : n23493;
  assign n23495 = pi21 ? n2427 : n204;
  assign n23496 = pi21 ? n5705 : n204;
  assign n23497 = pi20 ? n23495 : n23496;
  assign n23498 = pi19 ? n204 : n23497;
  assign n23499 = pi18 ? n23494 : n23498;
  assign n23500 = pi17 ? n32 : n23499;
  assign n23501 = pi21 ? n19311 : n204;
  assign n23502 = pi21 ? n1018 : n2402;
  assign n23503 = pi20 ? n23501 : n23502;
  assign n23504 = pi19 ? n23501 : n23503;
  assign n23505 = pi21 ? n204 : n19292;
  assign n23506 = pi20 ? n23002 : n23505;
  assign n23507 = pi19 ? n23000 : n23506;
  assign n23508 = pi18 ? n23504 : n23507;
  assign n23509 = pi21 ? n5705 : n1027;
  assign n23510 = pi20 ? n23509 : n2383;
  assign n23511 = pi19 ? n23510 : n316;
  assign n23512 = pi18 ? n23511 : n22989;
  assign n23513 = pi17 ? n23508 : n23512;
  assign n23514 = pi16 ? n23500 : n23513;
  assign n23515 = pi15 ? n22992 : n23514;
  assign n23516 = pi14 ? n23515 : n23030;
  assign n23517 = pi13 ? n23491 : n23516;
  assign n23518 = pi12 ? n23479 : n23517;
  assign n23519 = pi16 ? n331 : n23037;
  assign n23520 = pi15 ? n23519 : n23046;
  assign n23521 = pi20 ? n23048 : n2701;
  assign n23522 = pi19 ? n23521 : n32;
  assign n23523 = pi18 ? n139 : n23522;
  assign n23524 = pi17 ? n139 : n23523;
  assign n23525 = pi16 ? n915 : n23524;
  assign n23526 = pi20 ? n7858 : n1822;
  assign n23527 = pi19 ? n23526 : n32;
  assign n23528 = pi18 ? n23054 : n23527;
  assign n23529 = pi17 ? n139 : n23528;
  assign n23530 = pi16 ? n915 : n23529;
  assign n23531 = pi15 ? n23525 : n23530;
  assign n23532 = pi14 ? n23520 : n23531;
  assign n23533 = pi18 ? n23063 : n23527;
  assign n23534 = pi17 ? n335 : n23533;
  assign n23535 = pi16 ? n7943 : n23534;
  assign n23536 = pi21 ? n233 : n491;
  assign n23537 = pi20 ? n23536 : n32;
  assign n23538 = pi19 ? n23537 : n32;
  assign n23539 = pi18 ? n23071 : n23538;
  assign n23540 = pi17 ? n335 : n23539;
  assign n23541 = pi16 ? n2035 : n23540;
  assign n23542 = pi15 ? n23535 : n23541;
  assign n23543 = pi22 ? n233 : n396;
  assign n23544 = pi21 ? n233 : n23543;
  assign n23545 = pi20 ? n23544 : n32;
  assign n23546 = pi19 ? n23545 : n32;
  assign n23547 = pi18 ? n23079 : n23546;
  assign n23548 = pi17 ? n335 : n23547;
  assign n23549 = pi16 ? n7943 : n23548;
  assign n23550 = pi20 ? n10126 : n32;
  assign n23551 = pi19 ? n23550 : n32;
  assign n23552 = pi18 ? n335 : n23551;
  assign n23553 = pi17 ? n335 : n23552;
  assign n23554 = pi16 ? n23084 : n23553;
  assign n23555 = pi15 ? n23549 : n23554;
  assign n23556 = pi14 ? n23542 : n23555;
  assign n23557 = pi13 ? n23532 : n23556;
  assign n23558 = pi18 ? n233 : n23095;
  assign n23559 = pi17 ? n23106 : n23558;
  assign n23560 = pi16 ? n439 : n23559;
  assign n23561 = pi15 ? n23560 : n23120;
  assign n23562 = pi14 ? n23105 : n23561;
  assign n23563 = pi18 ? n10116 : n23125;
  assign n23564 = pi17 ? n32 : n23563;
  assign n23565 = pi16 ? n23564 : n23145;
  assign n23566 = pi15 ? n23565 : n23168;
  assign n23567 = pi22 ? n962 : n363;
  assign n23568 = pi21 ? n23567 : n363;
  assign n23569 = pi20 ? n32 : n23568;
  assign n23570 = pi19 ? n32 : n23569;
  assign n23571 = pi18 ? n23570 : n23176;
  assign n23572 = pi17 ? n32 : n23571;
  assign n23573 = pi21 ? n23186 : n7048;
  assign n23574 = pi20 ? n23573 : n32;
  assign n23575 = pi19 ? n23574 : n32;
  assign n23576 = pi18 ? n233 : n23575;
  assign n23577 = pi17 ? n23185 : n23576;
  assign n23578 = pi16 ? n23572 : n23577;
  assign n23579 = pi18 ? n23570 : n23194;
  assign n23580 = pi17 ? n32 : n23579;
  assign n23581 = pi21 ? n233 : n5829;
  assign n23582 = pi20 ? n23581 : n32;
  assign n23583 = pi19 ? n23582 : n32;
  assign n23584 = pi18 ? n233 : n23583;
  assign n23585 = pi17 ? n23202 : n23584;
  assign n23586 = pi16 ? n23580 : n23585;
  assign n23587 = pi15 ? n23578 : n23586;
  assign n23588 = pi14 ? n23566 : n23587;
  assign n23589 = pi13 ? n23562 : n23588;
  assign n23590 = pi12 ? n23557 : n23589;
  assign n23591 = pi11 ? n23518 : n23590;
  assign n23592 = pi10 ? n23438 : n23591;
  assign n23593 = pi09 ? n23229 : n23592;
  assign n23594 = pi08 ? n23215 : n23593;
  assign n23595 = pi20 ? n37 : n9607;
  assign n23596 = pi19 ? n23595 : n32;
  assign n23597 = pi18 ? n37 : n23596;
  assign n23598 = pi17 ? n37 : n23597;
  assign n23599 = pi16 ? n13561 : n23598;
  assign n23600 = pi15 ? n32 : n23599;
  assign n23601 = pi21 ? n37 : n18023;
  assign n23602 = pi20 ? n37 : n23601;
  assign n23603 = pi19 ? n23602 : n32;
  assign n23604 = pi18 ? n37 : n23603;
  assign n23605 = pi17 ? n37 : n23604;
  assign n23606 = pi16 ? n14445 : n23605;
  assign n23607 = pi20 ? n37 : n9622;
  assign n23608 = pi19 ? n23607 : n32;
  assign n23609 = pi18 ? n37 : n23608;
  assign n23610 = pi17 ? n37 : n23609;
  assign n23611 = pi16 ? n14445 : n23610;
  assign n23612 = pi15 ? n23606 : n23611;
  assign n23613 = pi14 ? n23600 : n23612;
  assign n23614 = pi13 ? n32 : n23613;
  assign n23615 = pi12 ? n32 : n23614;
  assign n23616 = pi11 ? n32 : n23615;
  assign n23617 = pi10 ? n32 : n23616;
  assign n23618 = pi20 ? n7346 : n2967;
  assign n23619 = pi20 ? n22644 : n2755;
  assign n23620 = pi19 ? n23618 : n23619;
  assign n23621 = pi18 ? n16593 : n23620;
  assign n23622 = pi17 ? n32 : n23621;
  assign n23623 = pi19 ? n3808 : n18500;
  assign n23624 = pi21 ? n2161 : n218;
  assign n23625 = pi20 ? n23624 : n18500;
  assign n23626 = pi19 ? n23625 : n3825;
  assign n23627 = pi18 ? n23623 : n23626;
  assign n23628 = pi20 ? n2747 : n18506;
  assign n23629 = pi20 ? n18506 : n17966;
  assign n23630 = pi19 ? n23628 : n23629;
  assign n23631 = pi21 ? n181 : n18039;
  assign n23632 = pi20 ? n23243 : n23631;
  assign n23633 = pi19 ? n23632 : n32;
  assign n23634 = pi18 ? n23630 : n23633;
  assign n23635 = pi17 ? n23627 : n23634;
  assign n23636 = pi16 ? n23622 : n23635;
  assign n23637 = pi22 ? n39 : n2160;
  assign n23638 = pi21 ? n23637 : n99;
  assign n23639 = pi20 ? n32 : n23638;
  assign n23640 = pi19 ? n32 : n23639;
  assign n23641 = pi20 ? n22666 : n14887;
  assign n23642 = pi19 ? n23641 : n20657;
  assign n23643 = pi18 ? n23640 : n23642;
  assign n23644 = pi17 ? n32 : n23643;
  assign n23645 = pi20 ? n5077 : n37;
  assign n23646 = pi19 ? n23645 : n14887;
  assign n23647 = pi18 ? n37 : n23646;
  assign n23648 = pi20 ? n37 : n3039;
  assign n23649 = pi19 ? n37 : n23648;
  assign n23650 = pi21 ? n218 : n11994;
  assign n23651 = pi20 ? n37 : n23650;
  assign n23652 = pi19 ? n23651 : n32;
  assign n23653 = pi18 ? n23649 : n23652;
  assign n23654 = pi17 ? n23647 : n23653;
  assign n23655 = pi16 ? n23644 : n23654;
  assign n23656 = pi15 ? n23636 : n23655;
  assign n23657 = pi20 ? n2974 : n18499;
  assign n23658 = pi20 ? n18500 : n5496;
  assign n23659 = pi19 ? n23657 : n23658;
  assign n23660 = pi18 ? n17008 : n23659;
  assign n23661 = pi17 ? n32 : n23660;
  assign n23662 = pi20 ? n11418 : n3817;
  assign n23663 = pi20 ? n2740 : n2163;
  assign n23664 = pi19 ? n23662 : n23663;
  assign n23665 = pi20 ? n2184 : n2740;
  assign n23666 = pi21 ? n2168 : n2746;
  assign n23667 = pi19 ? n23665 : n23666;
  assign n23668 = pi18 ? n23664 : n23667;
  assign n23669 = pi20 ? n17966 : n11424;
  assign n23670 = pi19 ? n23669 : n12287;
  assign n23671 = pi21 ? n2175 : n2746;
  assign n23672 = pi21 ? n2161 : n17575;
  assign n23673 = pi20 ? n23671 : n23672;
  assign n23674 = pi19 ? n23673 : n32;
  assign n23675 = pi18 ? n23670 : n23674;
  assign n23676 = pi17 ? n23668 : n23675;
  assign n23677 = pi16 ? n23661 : n23676;
  assign n23678 = pi21 ? n2957 : n17575;
  assign n23679 = pi20 ? n37 : n23678;
  assign n23680 = pi19 ? n23679 : n32;
  assign n23681 = pi18 ? n37 : n23680;
  assign n23682 = pi17 ? n37 : n23681;
  assign n23683 = pi16 ? n439 : n23682;
  assign n23684 = pi15 ? n23677 : n23683;
  assign n23685 = pi14 ? n23656 : n23684;
  assign n23686 = pi21 ? n2957 : n99;
  assign n23687 = pi20 ? n23686 : n99;
  assign n23688 = pi19 ? n23687 : n99;
  assign n23689 = pi18 ? n374 : n23688;
  assign n23690 = pi17 ? n32 : n23689;
  assign n23691 = pi21 ? n99 : n17583;
  assign n23692 = pi20 ? n99 : n23691;
  assign n23693 = pi19 ? n23692 : n32;
  assign n23694 = pi18 ? n99 : n23693;
  assign n23695 = pi17 ? n99 : n23694;
  assign n23696 = pi16 ? n23690 : n23695;
  assign n23697 = pi18 ? n374 : n21612;
  assign n23698 = pi17 ? n32 : n23697;
  assign n23699 = pi20 ? n99 : n9247;
  assign n23700 = pi19 ? n23699 : n32;
  assign n23701 = pi18 ? n99 : n23700;
  assign n23702 = pi17 ? n99 : n23701;
  assign n23703 = pi16 ? n23698 : n23702;
  assign n23704 = pi15 ? n23696 : n23703;
  assign n23705 = pi20 ? n3824 : n5496;
  assign n23706 = pi20 ? n5496 : n2968;
  assign n23707 = pi19 ? n23705 : n23706;
  assign n23708 = pi18 ? n14509 : n23707;
  assign n23709 = pi17 ? n32 : n23708;
  assign n23710 = pi20 ? n2968 : n14846;
  assign n23711 = pi19 ? n23710 : n139;
  assign n23712 = pi18 ? n23711 : n22705;
  assign n23713 = pi20 ? n139 : n9247;
  assign n23714 = pi19 ? n23713 : n32;
  assign n23715 = pi18 ? n139 : n23714;
  assign n23716 = pi17 ? n23712 : n23715;
  assign n23717 = pi16 ? n23709 : n23716;
  assign n23718 = pi21 ? n16004 : n2161;
  assign n23719 = pi20 ? n32 : n23718;
  assign n23720 = pi19 ? n32 : n23719;
  assign n23721 = pi20 ? n11418 : n2185;
  assign n23722 = pi19 ? n22644 : n23721;
  assign n23723 = pi18 ? n23720 : n23722;
  assign n23724 = pi17 ? n32 : n23723;
  assign n23725 = pi20 ? n17966 : n14846;
  assign n23726 = pi19 ? n23725 : n139;
  assign n23727 = pi21 ? n2164 : n139;
  assign n23728 = pi20 ? n23727 : n139;
  assign n23729 = pi19 ? n23728 : n139;
  assign n23730 = pi18 ? n23726 : n23729;
  assign n23731 = pi20 ? n139 : n9256;
  assign n23732 = pi19 ? n23731 : n32;
  assign n23733 = pi18 ? n139 : n23732;
  assign n23734 = pi17 ? n23730 : n23733;
  assign n23735 = pi16 ? n23724 : n23734;
  assign n23736 = pi15 ? n23717 : n23735;
  assign n23737 = pi14 ? n23704 : n23736;
  assign n23738 = pi13 ? n23685 : n23737;
  assign n23739 = pi21 ? n297 : n1711;
  assign n23740 = pi21 ? n1211 : n1711;
  assign n23741 = pi20 ? n23739 : n23740;
  assign n23742 = pi19 ? n20714 : n23741;
  assign n23743 = pi20 ? n5255 : n139;
  assign n23744 = pi19 ? n23743 : n139;
  assign n23745 = pi18 ? n23742 : n23744;
  assign n23746 = pi20 ? n139 : n10644;
  assign n23747 = pi19 ? n23746 : n32;
  assign n23748 = pi18 ? n139 : n23747;
  assign n23749 = pi17 ? n23745 : n23748;
  assign n23750 = pi16 ? n439 : n23749;
  assign n23751 = pi19 ? n13125 : n1003;
  assign n23752 = pi18 ? n23751 : n10652;
  assign n23753 = pi19 ? n3554 : n139;
  assign n23754 = pi21 ? n139 : n2578;
  assign n23755 = pi20 ? n139 : n23754;
  assign n23756 = pi19 ? n23755 : n32;
  assign n23757 = pi18 ? n23753 : n23756;
  assign n23758 = pi17 ? n23752 : n23757;
  assign n23759 = pi16 ? n439 : n23758;
  assign n23760 = pi15 ? n23750 : n23759;
  assign n23761 = pi20 ? n1003 : n376;
  assign n23762 = pi19 ? n23761 : n8743;
  assign n23763 = pi18 ? n374 : n23762;
  assign n23764 = pi17 ? n32 : n23763;
  assign n23765 = pi20 ? n8742 : n3671;
  assign n23766 = pi19 ? n23765 : n3671;
  assign n23767 = pi20 ? n3671 : n3610;
  assign n23768 = pi19 ? n23767 : n16023;
  assign n23769 = pi18 ? n23766 : n23768;
  assign n23770 = pi20 ? n1715 : n3645;
  assign n23771 = pi20 ? n2518 : n139;
  assign n23772 = pi19 ? n23770 : n23771;
  assign n23773 = pi18 ? n23772 : n23756;
  assign n23774 = pi17 ? n23769 : n23773;
  assign n23775 = pi16 ? n23764 : n23774;
  assign n23776 = pi20 ? n997 : n23739;
  assign n23777 = pi19 ? n37 : n23776;
  assign n23778 = pi18 ? n37 : n23777;
  assign n23779 = pi19 ? n15002 : n8765;
  assign n23780 = pi21 ? n139 : n2637;
  assign n23781 = pi20 ? n139 : n23780;
  assign n23782 = pi19 ? n23781 : n32;
  assign n23783 = pi18 ? n23779 : n23782;
  assign n23784 = pi17 ? n23778 : n23783;
  assign n23785 = pi16 ? n439 : n23784;
  assign n23786 = pi15 ? n23775 : n23785;
  assign n23787 = pi14 ? n23760 : n23786;
  assign n23788 = pi21 ? n363 : n882;
  assign n23789 = pi20 ? n139 : n23788;
  assign n23790 = pi19 ? n23789 : n32;
  assign n23791 = pi18 ? n13193 : n23790;
  assign n23792 = pi17 ? n37 : n23791;
  assign n23793 = pi16 ? n439 : n23792;
  assign n23794 = pi15 ? n23793 : n22767;
  assign n23795 = pi22 ? n15863 : n32;
  assign n23796 = pi21 ? n204 : n23795;
  assign n23797 = pi20 ? n204 : n23796;
  assign n23798 = pi19 ? n23797 : n32;
  assign n23799 = pi18 ? n22776 : n23798;
  assign n23800 = pi17 ? n37 : n23799;
  assign n23801 = pi16 ? n439 : n23800;
  assign n23802 = pi19 ? n37 : n18108;
  assign n23803 = pi21 ? n204 : n2565;
  assign n23804 = pi20 ? n204 : n23803;
  assign n23805 = pi19 ? n23804 : n32;
  assign n23806 = pi18 ? n23802 : n23805;
  assign n23807 = pi17 ? n37 : n23806;
  assign n23808 = pi16 ? n439 : n23807;
  assign n23809 = pi15 ? n23801 : n23808;
  assign n23810 = pi14 ? n23794 : n23809;
  assign n23811 = pi13 ? n23787 : n23810;
  assign n23812 = pi12 ? n23738 : n23811;
  assign n23813 = pi18 ? n23802 : n22779;
  assign n23814 = pi17 ? n37 : n23813;
  assign n23815 = pi16 ? n439 : n23814;
  assign n23816 = pi21 ? n11199 : n1943;
  assign n23817 = pi20 ? n37 : n23816;
  assign n23818 = pi19 ? n37 : n23817;
  assign n23819 = pi22 ? n455 : n233;
  assign n23820 = pi21 ? n6361 : n23819;
  assign n23821 = pi21 ? n6376 : n2553;
  assign n23822 = pi20 ? n23820 : n23821;
  assign n23823 = pi19 ? n23822 : n32;
  assign n23824 = pi18 ? n23818 : n23823;
  assign n23825 = pi17 ? n37 : n23824;
  assign n23826 = pi16 ? n439 : n23825;
  assign n23827 = pi15 ? n23815 : n23826;
  assign n23828 = pi21 ? n2061 : n2678;
  assign n23829 = pi20 ? n335 : n23828;
  assign n23830 = pi19 ? n23829 : n32;
  assign n23831 = pi18 ? n21770 : n23830;
  assign n23832 = pi17 ? n37 : n23831;
  assign n23833 = pi16 ? n439 : n23832;
  assign n23834 = pi14 ? n23827 : n23833;
  assign n23835 = pi18 ? n17205 : n23830;
  assign n23836 = pi17 ? n37 : n23835;
  assign n23837 = pi16 ? n439 : n23836;
  assign n23838 = pi20 ? n649 : n603;
  assign n23839 = pi19 ? n37 : n23838;
  assign n23840 = pi18 ? n23839 : n23830;
  assign n23841 = pi17 ? n37 : n23840;
  assign n23842 = pi16 ? n439 : n23841;
  assign n23843 = pi15 ? n23837 : n23842;
  assign n23844 = pi20 ? n639 : n577;
  assign n23845 = pi19 ? n37 : n23844;
  assign n23846 = pi18 ? n23845 : n23830;
  assign n23847 = pi17 ? n37 : n23846;
  assign n23848 = pi16 ? n439 : n23847;
  assign n23849 = pi20 ? n577 : n3335;
  assign n23850 = pi19 ? n37 : n23849;
  assign n23851 = pi20 ? n569 : n10249;
  assign n23852 = pi19 ? n23851 : n32;
  assign n23853 = pi18 ? n23850 : n23852;
  assign n23854 = pi17 ? n37 : n23853;
  assign n23855 = pi16 ? n439 : n23854;
  assign n23856 = pi15 ? n23848 : n23855;
  assign n23857 = pi14 ? n23843 : n23856;
  assign n23858 = pi13 ? n23834 : n23857;
  assign n23859 = pi21 ? n11336 : n2700;
  assign n23860 = pi20 ? n649 : n23859;
  assign n23861 = pi19 ? n23860 : n32;
  assign n23862 = pi18 ? n37 : n23861;
  assign n23863 = pi17 ? n37 : n23862;
  assign n23864 = pi16 ? n439 : n23863;
  assign n23865 = pi20 ? n2094 : n18756;
  assign n23866 = pi19 ? n23865 : n32;
  assign n23867 = pi18 ? n37 : n23866;
  assign n23868 = pi17 ? n37 : n23867;
  assign n23869 = pi16 ? n439 : n23868;
  assign n23870 = pi15 ? n23864 : n23869;
  assign n23871 = pi20 ? n2094 : n20237;
  assign n23872 = pi19 ? n23871 : n32;
  assign n23873 = pi18 ? n37 : n23872;
  assign n23874 = pi17 ? n37 : n23873;
  assign n23875 = pi16 ? n439 : n23874;
  assign n23876 = pi20 ? n37 : n18412;
  assign n23877 = pi19 ? n23876 : n32;
  assign n23878 = pi18 ? n37 : n23877;
  assign n23879 = pi17 ? n37 : n23878;
  assign n23880 = pi16 ? n439 : n23879;
  assign n23881 = pi15 ? n23875 : n23880;
  assign n23882 = pi14 ? n23870 : n23881;
  assign n23883 = pi20 ? n37 : n12514;
  assign n23884 = pi19 ? n23883 : n32;
  assign n23885 = pi18 ? n37 : n23884;
  assign n23886 = pi17 ? n37 : n23885;
  assign n23887 = pi16 ? n439 : n23886;
  assign n23888 = pi22 ? n685 : n3124;
  assign n23889 = pi21 ? n23888 : n32;
  assign n23890 = pi20 ? n9660 : n23889;
  assign n23891 = pi19 ? n23890 : n32;
  assign n23892 = pi18 ? n37 : n23891;
  assign n23893 = pi17 ? n37 : n23892;
  assign n23894 = pi16 ? n439 : n23893;
  assign n23895 = pi15 ? n23887 : n23894;
  assign n23896 = pi22 ? n363 : n6146;
  assign n23897 = pi21 ? n23896 : n32;
  assign n23898 = pi20 ? n21826 : n23897;
  assign n23899 = pi19 ? n23898 : n32;
  assign n23900 = pi18 ? n37 : n23899;
  assign n23901 = pi17 ? n37 : n23900;
  assign n23902 = pi16 ? n439 : n23901;
  assign n23903 = pi20 ? n37 : n22881;
  assign n23904 = pi19 ? n23903 : n22883;
  assign n23905 = pi22 ? n363 : n1378;
  assign n23906 = pi21 ? n23905 : n32;
  assign n23907 = pi20 ? n363 : n23906;
  assign n23908 = pi19 ? n23907 : n32;
  assign n23909 = pi18 ? n23904 : n23908;
  assign n23910 = pi17 ? n37 : n23909;
  assign n23911 = pi16 ? n439 : n23910;
  assign n23912 = pi15 ? n23902 : n23911;
  assign n23913 = pi14 ? n23895 : n23912;
  assign n23914 = pi13 ? n23882 : n23913;
  assign n23915 = pi12 ? n23858 : n23914;
  assign n23916 = pi11 ? n23812 : n23915;
  assign n23917 = pi20 ? n37 : n363;
  assign n23918 = pi19 ? n23917 : n363;
  assign n23919 = pi18 ? n23918 : n23440;
  assign n23920 = pi17 ? n37 : n23919;
  assign n23921 = pi16 ? n439 : n23920;
  assign n23922 = pi18 ? n22898 : n23430;
  assign n23923 = pi17 ? n37 : n23922;
  assign n23924 = pi16 ? n439 : n23923;
  assign n23925 = pi15 ? n23921 : n23924;
  assign n23926 = pi21 ? n6433 : n244;
  assign n23927 = pi20 ? n37 : n23926;
  assign n23928 = pi21 ? n272 : n19958;
  assign n23929 = pi21 ? n19958 : n37;
  assign n23930 = pi20 ? n23928 : n23929;
  assign n23931 = pi19 ? n23927 : n23930;
  assign n23932 = pi22 ? n889 : n157;
  assign n23933 = pi21 ? n23932 : n2106;
  assign n23934 = pi20 ? n23933 : n9456;
  assign n23935 = pi19 ? n23934 : n32;
  assign n23936 = pi18 ? n23931 : n23935;
  assign n23937 = pi17 ? n37 : n23936;
  assign n23938 = pi16 ? n439 : n23937;
  assign n23939 = pi21 ? n37 : n23932;
  assign n23940 = pi20 ? n37 : n23939;
  assign n23941 = pi21 ? n22377 : n2106;
  assign n23942 = pi21 ? n37 : n8654;
  assign n23943 = pi20 ? n23941 : n23942;
  assign n23944 = pi19 ? n23940 : n23943;
  assign n23945 = pi21 ? n272 : n218;
  assign n23946 = pi20 ? n23945 : n9456;
  assign n23947 = pi19 ? n23946 : n32;
  assign n23948 = pi18 ? n23944 : n23947;
  assign n23949 = pi17 ? n37 : n23948;
  assign n23950 = pi16 ? n439 : n23949;
  assign n23951 = pi15 ? n23938 : n23950;
  assign n23952 = pi14 ? n23925 : n23951;
  assign n23953 = pi20 ? n5467 : n9456;
  assign n23954 = pi19 ? n23953 : n32;
  assign n23955 = pi18 ? n99 : n23954;
  assign n23956 = pi17 ? n99 : n23955;
  assign n23957 = pi16 ? n721 : n23956;
  assign n23958 = pi20 ? n16263 : n99;
  assign n23959 = pi19 ? n99 : n23958;
  assign n23960 = pi18 ? n23959 : n23462;
  assign n23961 = pi17 ? n99 : n23960;
  assign n23962 = pi16 ? n721 : n23961;
  assign n23963 = pi15 ? n23957 : n23962;
  assign n23964 = pi20 ? n2238 : n5667;
  assign n23965 = pi19 ? n23964 : n32;
  assign n23966 = pi18 ? n99 : n23965;
  assign n23967 = pi17 ? n99 : n23966;
  assign n23968 = pi16 ? n721 : n23967;
  assign n23969 = pi14 ? n23963 : n23968;
  assign n23970 = pi13 ? n23952 : n23969;
  assign n23971 = pi20 ? n777 : n3210;
  assign n23972 = pi19 ? n23971 : n32;
  assign n23973 = pi18 ? n99 : n23972;
  assign n23974 = pi17 ? n99 : n23973;
  assign n23975 = pi16 ? n721 : n23974;
  assign n23976 = pi18 ? n99 : n22960;
  assign n23977 = pi17 ? n99 : n23976;
  assign n23978 = pi16 ? n721 : n23977;
  assign n23979 = pi15 ? n23975 : n23978;
  assign n23980 = pi21 ? n16350 : n32;
  assign n23981 = pi20 ? n19171 : n23980;
  assign n23982 = pi19 ? n23981 : n32;
  assign n23983 = pi18 ? n22967 : n23982;
  assign n23984 = pi17 ? n99 : n23983;
  assign n23985 = pi16 ? n721 : n23984;
  assign n23986 = pi23 ? n714 : n139;
  assign n23987 = pi22 ? n23986 : n139;
  assign n23988 = pi21 ? n23987 : n139;
  assign n23989 = pi20 ? n32 : n23988;
  assign n23990 = pi19 ? n32 : n23989;
  assign n23991 = pi18 ? n23990 : n139;
  assign n23992 = pi17 ? n32 : n23991;
  assign n23993 = pi19 ? n1820 : n17420;
  assign n23994 = pi20 ? n10033 : n10011;
  assign n23995 = pi19 ? n23994 : n32;
  assign n23996 = pi18 ? n23993 : n23995;
  assign n23997 = pi17 ? n139 : n23996;
  assign n23998 = pi16 ? n23992 : n23997;
  assign n23999 = pi15 ? n23985 : n23998;
  assign n24000 = pi14 ? n23979 : n23999;
  assign n24001 = pi20 ? n139 : n6930;
  assign n24002 = pi19 ? n139 : n24001;
  assign n24003 = pi18 ? n24002 : n139;
  assign n24004 = pi20 ? n316 : n10011;
  assign n24005 = pi19 ? n24004 : n32;
  assign n24006 = pi18 ? n10073 : n24005;
  assign n24007 = pi17 ? n24003 : n24006;
  assign n24008 = pi16 ? n2291 : n24007;
  assign n24009 = pi21 ? n1037 : n19311;
  assign n24010 = pi20 ? n32 : n24009;
  assign n24011 = pi19 ? n32 : n24010;
  assign n24012 = pi21 ? n19292 : n204;
  assign n24013 = pi21 ? n384 : n1018;
  assign n24014 = pi20 ? n24012 : n24013;
  assign n24015 = pi19 ? n204 : n24014;
  assign n24016 = pi18 ? n24011 : n24015;
  assign n24017 = pi17 ? n32 : n24016;
  assign n24018 = pi21 ? n1046 : n1018;
  assign n24019 = pi21 ? n381 : n3258;
  assign n24020 = pi20 ? n24018 : n24019;
  assign n24021 = pi19 ? n24018 : n24020;
  assign n24022 = pi20 ? n5299 : n440;
  assign n24023 = pi21 ? n204 : n381;
  assign n24024 = pi21 ? n1018 : n381;
  assign n24025 = pi20 ? n24023 : n24024;
  assign n24026 = pi19 ? n24022 : n24025;
  assign n24027 = pi18 ? n24021 : n24026;
  assign n24028 = pi19 ? n5337 : n316;
  assign n24029 = pi18 ? n24028 : n24005;
  assign n24030 = pi17 ? n24027 : n24029;
  assign n24031 = pi16 ? n24017 : n24030;
  assign n24032 = pi15 ? n24008 : n24031;
  assign n24033 = pi21 ? n16358 : n32;
  assign n24034 = pi20 ? n316 : n24033;
  assign n24035 = pi19 ? n24034 : n32;
  assign n24036 = pi18 ? n23026 : n24035;
  assign n24037 = pi17 ? n204 : n24036;
  assign n24038 = pi16 ? n13493 : n24037;
  assign n24039 = pi18 ? n204 : n13479;
  assign n24040 = pi18 ? n23026 : n24005;
  assign n24041 = pi17 ? n24039 : n24040;
  assign n24042 = pi16 ? n13846 : n24041;
  assign n24043 = pi15 ? n24038 : n24042;
  assign n24044 = pi14 ? n24032 : n24043;
  assign n24045 = pi13 ? n24000 : n24044;
  assign n24046 = pi12 ? n23970 : n24045;
  assign n24047 = pi20 ? n347 : n139;
  assign n24048 = pi19 ? n139 : n24047;
  assign n24049 = pi20 ? n975 : n10011;
  assign n24050 = pi19 ? n24049 : n32;
  assign n24051 = pi18 ? n24048 : n24050;
  assign n24052 = pi17 ? n139 : n24051;
  assign n24053 = pi16 ? n915 : n24052;
  assign n24054 = pi19 ? n21060 : n139;
  assign n24055 = pi20 ? n23048 : n2653;
  assign n24056 = pi19 ? n24055 : n32;
  assign n24057 = pi18 ? n24054 : n24056;
  assign n24058 = pi17 ? n139 : n24057;
  assign n24059 = pi16 ? n331 : n24058;
  assign n24060 = pi15 ? n24053 : n24059;
  assign n24061 = pi21 ? n139 : n11818;
  assign n24062 = pi20 ? n24061 : n2701;
  assign n24063 = pi19 ? n24062 : n32;
  assign n24064 = pi18 ? n139 : n24063;
  assign n24065 = pi17 ? n139 : n24064;
  assign n24066 = pi16 ? n1575 : n24065;
  assign n24067 = pi21 ? n204 : n16438;
  assign n24068 = pi20 ? n24067 : n1822;
  assign n24069 = pi19 ? n24068 : n32;
  assign n24070 = pi18 ? n23054 : n24069;
  assign n24071 = pi17 ? n139 : n24070;
  assign n24072 = pi16 ? n1575 : n24071;
  assign n24073 = pi15 ? n24066 : n24072;
  assign n24074 = pi14 ? n24060 : n24073;
  assign n24075 = pi20 ? n335 : n7980;
  assign n24076 = pi19 ? n24075 : n6749;
  assign n24077 = pi18 ? n24076 : n24069;
  assign n24078 = pi17 ? n335 : n24077;
  assign n24079 = pi16 ? n10399 : n24078;
  assign n24080 = pi19 ? n24075 : n17533;
  assign n24081 = pi21 ? n233 : n9430;
  assign n24082 = pi20 ? n24081 : n32;
  assign n24083 = pi19 ? n24082 : n32;
  assign n24084 = pi18 ? n24080 : n24083;
  assign n24085 = pi17 ? n335 : n24084;
  assign n24086 = pi16 ? n2035 : n24085;
  assign n24087 = pi15 ? n24079 : n24086;
  assign n24088 = pi18 ? n23079 : n24083;
  assign n24089 = pi17 ? n335 : n24088;
  assign n24090 = pi16 ? n7943 : n24089;
  assign n24091 = pi19 ? n335 : n22017;
  assign n24092 = pi21 ? n335 : n665;
  assign n24093 = pi20 ? n24092 : n32;
  assign n24094 = pi19 ? n24093 : n32;
  assign n24095 = pi18 ? n24091 : n24094;
  assign n24096 = pi17 ? n335 : n24095;
  assign n24097 = pi16 ? n23084 : n24096;
  assign n24098 = pi15 ? n24090 : n24097;
  assign n24099 = pi14 ? n24087 : n24098;
  assign n24100 = pi13 ? n24074 : n24099;
  assign n24101 = pi19 ? n37 : n21168;
  assign n24102 = pi18 ? n374 : n24101;
  assign n24103 = pi17 ? n32 : n24102;
  assign n24104 = pi19 ? n37 : n3384;
  assign n24105 = pi21 ? n580 : n37;
  assign n24106 = pi20 ? n37 : n24105;
  assign n24107 = pi19 ? n24106 : n10681;
  assign n24108 = pi18 ? n24104 : n24107;
  assign n24109 = pi21 ? n233 : n665;
  assign n24110 = pi20 ? n24109 : n32;
  assign n24111 = pi19 ? n24110 : n32;
  assign n24112 = pi18 ? n17552 : n24111;
  assign n24113 = pi17 ? n24108 : n24112;
  assign n24114 = pi16 ? n24103 : n24113;
  assign n24115 = pi20 ? n605 : n13527;
  assign n24116 = pi19 ? n24115 : n233;
  assign n24117 = pi21 ? n233 : n14168;
  assign n24118 = pi20 ? n24117 : n32;
  assign n24119 = pi19 ? n24118 : n32;
  assign n24120 = pi18 ? n24116 : n24119;
  assign n24121 = pi17 ? n14165 : n24120;
  assign n24122 = pi16 ? n439 : n24121;
  assign n24123 = pi15 ? n24114 : n24122;
  assign n24124 = pi20 ? n3299 : n2092;
  assign n24125 = pi19 ? n37 : n24124;
  assign n24126 = pi20 ? n2094 : n577;
  assign n24127 = pi19 ? n37 : n24126;
  assign n24128 = pi18 ? n24125 : n24127;
  assign n24129 = pi18 ? n233 : n24119;
  assign n24130 = pi17 ? n24128 : n24129;
  assign n24131 = pi16 ? n439 : n24130;
  assign n24132 = pi18 ? n17487 : n15082;
  assign n24133 = pi20 ? n6377 : n6362;
  assign n24134 = pi19 ? n24133 : n17542;
  assign n24135 = pi21 ? n233 : n2230;
  assign n24136 = pi20 ? n24135 : n32;
  assign n24137 = pi19 ? n24136 : n32;
  assign n24138 = pi18 ? n24134 : n24137;
  assign n24139 = pi17 ? n24132 : n24138;
  assign n24140 = pi16 ? n3351 : n24139;
  assign n24141 = pi15 ? n24131 : n24140;
  assign n24142 = pi14 ? n24123 : n24141;
  assign n24143 = pi22 ? n2419 : n1656;
  assign n24144 = pi21 ? n24143 : n14865;
  assign n24145 = pi20 ? n32 : n24144;
  assign n24146 = pi19 ? n32 : n24145;
  assign n24147 = pi21 ? n18462 : n14865;
  assign n24148 = pi22 ? n22116 : n363;
  assign n24149 = pi21 ? n24148 : n14865;
  assign n24150 = pi20 ? n24147 : n24149;
  assign n24151 = pi21 ? n363 : n14865;
  assign n24152 = pi21 ? n21201 : n22549;
  assign n24153 = pi20 ? n24151 : n24152;
  assign n24154 = pi19 ? n24150 : n24153;
  assign n24155 = pi18 ? n24146 : n24154;
  assign n24156 = pi17 ? n32 : n24155;
  assign n24157 = pi22 ? n363 : n1656;
  assign n24158 = pi21 ? n24157 : n22549;
  assign n24159 = pi20 ? n24158 : n23150;
  assign n24160 = pi20 ? n21220 : n21222;
  assign n24161 = pi19 ? n24159 : n24160;
  assign n24162 = pi21 ? n722 : n5014;
  assign n24163 = pi20 ? n23161 : n24162;
  assign n24164 = pi21 ? n21201 : n233;
  assign n24165 = pi20 ? n19422 : n24164;
  assign n24166 = pi19 ? n24163 : n24165;
  assign n24167 = pi18 ? n24161 : n24166;
  assign n24168 = pi21 ? n4903 : n233;
  assign n24169 = pi20 ? n233 : n24168;
  assign n24170 = pi19 ? n233 : n24169;
  assign n24171 = pi21 ? n233 : n5178;
  assign n24172 = pi20 ? n24171 : n32;
  assign n24173 = pi19 ? n24172 : n32;
  assign n24174 = pi18 ? n24170 : n24173;
  assign n24175 = pi17 ? n24167 : n24174;
  assign n24176 = pi16 ? n24156 : n24175;
  assign n24177 = pi20 ? n363 : n20860;
  assign n24178 = pi19 ? n363 : n24177;
  assign n24179 = pi18 ? n23149 : n24178;
  assign n24180 = pi17 ? n32 : n24179;
  assign n24181 = pi19 ? n363 : n24160;
  assign n24182 = pi20 ? n23161 : n21220;
  assign n24183 = pi22 ? n363 : n23156;
  assign n24184 = pi21 ? n24183 : n233;
  assign n24185 = pi20 ? n19422 : n24184;
  assign n24186 = pi19 ? n24182 : n24185;
  assign n24187 = pi18 ? n24181 : n24186;
  assign n24188 = pi17 ? n24187 : n23166;
  assign n24189 = pi16 ? n24180 : n24188;
  assign n24190 = pi15 ? n24176 : n24189;
  assign n24191 = pi18 ? n21559 : n23176;
  assign n24192 = pi17 ? n32 : n24191;
  assign n24193 = pi21 ? n21235 : n363;
  assign n24194 = pi20 ? n363 : n24193;
  assign n24195 = pi21 ? n21235 : n2707;
  assign n24196 = pi22 ? n673 : n363;
  assign n24197 = pi21 ? n24196 : n21235;
  assign n24198 = pi20 ? n24195 : n24197;
  assign n24199 = pi19 ? n24194 : n24198;
  assign n24200 = pi21 ? n24183 : n363;
  assign n24201 = pi20 ? n24200 : n5021;
  assign n24202 = pi21 ? n2707 : n19920;
  assign n24203 = pi22 ? n23156 : n233;
  assign n24204 = pi21 ? n24203 : n19920;
  assign n24205 = pi20 ? n24202 : n24204;
  assign n24206 = pi19 ? n24201 : n24205;
  assign n24207 = pi18 ? n24199 : n24206;
  assign n24208 = pi22 ? n22498 : n32;
  assign n24209 = pi21 ? n233 : n24208;
  assign n24210 = pi20 ? n24209 : n32;
  assign n24211 = pi19 ? n24210 : n32;
  assign n24212 = pi18 ? n233 : n24211;
  assign n24213 = pi17 ? n24207 : n24212;
  assign n24214 = pi16 ? n24192 : n24213;
  assign n24215 = pi22 ? n686 : n363;
  assign n24216 = pi21 ? n24215 : n363;
  assign n24217 = pi20 ? n363 : n24216;
  assign n24218 = pi19 ? n363 : n24217;
  assign n24219 = pi18 ? n24218 : n363;
  assign n24220 = pi21 ? n2721 : n685;
  assign n24221 = pi20 ? n19084 : n24220;
  assign n24222 = pi22 ? n685 : n363;
  assign n24223 = pi21 ? n24222 : n2721;
  assign n24224 = pi20 ? n24223 : n19084;
  assign n24225 = pi19 ? n24221 : n24224;
  assign n24226 = pi18 ? n24225 : n14264;
  assign n24227 = pi17 ? n24219 : n24226;
  assign n24228 = pi16 ? n21561 : n24227;
  assign n24229 = pi15 ? n24214 : n24228;
  assign n24230 = pi14 ? n24190 : n24229;
  assign n24231 = pi13 ? n24142 : n24230;
  assign n24232 = pi12 ? n24100 : n24231;
  assign n24233 = pi11 ? n24046 : n24232;
  assign n24234 = pi10 ? n23916 : n24233;
  assign n24235 = pi09 ? n23617 : n24234;
  assign n24236 = pi16 ? n14445 : n23598;
  assign n24237 = pi15 ? n32 : n24236;
  assign n24238 = pi16 ? n16595 : n23610;
  assign n24239 = pi15 ? n23606 : n24238;
  assign n24240 = pi14 ? n24237 : n24239;
  assign n24241 = pi13 ? n32 : n24240;
  assign n24242 = pi12 ? n32 : n24241;
  assign n24243 = pi11 ? n32 : n24242;
  assign n24244 = pi10 ? n32 : n24243;
  assign n24245 = pi19 ? n23618 : n22622;
  assign n24246 = pi18 ? n16593 : n24245;
  assign n24247 = pi17 ? n32 : n24246;
  assign n24248 = pi19 ? n2963 : n17960;
  assign n24249 = pi20 ? n2176 : n17960;
  assign n24250 = pi19 ? n24249 : n2967;
  assign n24251 = pi18 ? n24248 : n24250;
  assign n24252 = pi20 ? n2176 : n2976;
  assign n24253 = pi19 ? n24252 : n2184;
  assign n24254 = pi21 ? n2175 : n18039;
  assign n24255 = pi20 ? n11424 : n24254;
  assign n24256 = pi19 ? n24255 : n32;
  assign n24257 = pi18 ? n24253 : n24256;
  assign n24258 = pi17 ? n24251 : n24257;
  assign n24259 = pi16 ? n24247 : n24258;
  assign n24260 = pi21 ? n65 : n2161;
  assign n24261 = pi20 ? n32 : n24260;
  assign n24262 = pi19 ? n32 : n24261;
  assign n24263 = pi20 ? n37 : n14887;
  assign n24264 = pi19 ? n24263 : n20657;
  assign n24265 = pi18 ? n24262 : n24264;
  assign n24266 = pi17 ? n32 : n24265;
  assign n24267 = pi16 ? n24266 : n23654;
  assign n24268 = pi15 ? n24259 : n24267;
  assign n24269 = pi20 ? n37 : n15960;
  assign n24270 = pi20 ? n17960 : n2982;
  assign n24271 = pi19 ? n24269 : n24270;
  assign n24272 = pi18 ? n17008 : n24271;
  assign n24273 = pi17 ? n32 : n24272;
  assign n24274 = pi20 ? n11415 : n2973;
  assign n24275 = pi19 ? n24274 : n2961;
  assign n24276 = pi20 ? n2184 : n2961;
  assign n24277 = pi19 ? n24276 : n15960;
  assign n24278 = pi18 ? n24275 : n24277;
  assign n24279 = pi20 ? n2184 : n11418;
  assign n24280 = pi19 ? n24279 : n20660;
  assign n24281 = pi21 ? n2161 : n3066;
  assign n24282 = pi20 ? n2176 : n24281;
  assign n24283 = pi19 ? n24282 : n32;
  assign n24284 = pi18 ? n24280 : n24283;
  assign n24285 = pi17 ? n24278 : n24284;
  assign n24286 = pi16 ? n24273 : n24285;
  assign n24287 = pi21 ? n2957 : n9238;
  assign n24288 = pi20 ? n37 : n24287;
  assign n24289 = pi19 ? n24288 : n32;
  assign n24290 = pi18 ? n37 : n24289;
  assign n24291 = pi17 ? n37 : n24290;
  assign n24292 = pi16 ? n439 : n24291;
  assign n24293 = pi15 ? n24286 : n24292;
  assign n24294 = pi14 ? n24268 : n24293;
  assign n24295 = pi23 ? n11910 : n32;
  assign n24296 = pi22 ? n24295 : n32;
  assign n24297 = pi21 ? n99 : n24296;
  assign n24298 = pi20 ? n99 : n24297;
  assign n24299 = pi19 ? n24298 : n32;
  assign n24300 = pi18 ? n99 : n24299;
  assign n24301 = pi17 ? n99 : n24300;
  assign n24302 = pi16 ? n23690 : n24301;
  assign n24303 = pi21 ? n99 : n3848;
  assign n24304 = pi20 ? n99 : n24303;
  assign n24305 = pi19 ? n24304 : n32;
  assign n24306 = pi18 ? n99 : n24305;
  assign n24307 = pi17 ? n99 : n24306;
  assign n24308 = pi16 ? n23698 : n24307;
  assign n24309 = pi15 ? n24302 : n24308;
  assign n24310 = pi20 ? n139 : n24303;
  assign n24311 = pi19 ? n24310 : n32;
  assign n24312 = pi18 ? n139 : n24311;
  assign n24313 = pi17 ? n23712 : n24312;
  assign n24314 = pi16 ? n23709 : n24313;
  assign n24315 = pi20 ? n139 : n10189;
  assign n24316 = pi19 ? n24315 : n32;
  assign n24317 = pi18 ? n139 : n24316;
  assign n24318 = pi17 ? n23730 : n24317;
  assign n24319 = pi16 ? n23724 : n24318;
  assign n24320 = pi15 ? n24314 : n24319;
  assign n24321 = pi14 ? n24309 : n24320;
  assign n24322 = pi13 ? n24294 : n24321;
  assign n24323 = pi20 ? n139 : n11559;
  assign n24324 = pi19 ? n24323 : n32;
  assign n24325 = pi18 ? n139 : n24324;
  assign n24326 = pi17 ? n23745 : n24325;
  assign n24327 = pi16 ? n439 : n24326;
  assign n24328 = pi21 ? n139 : n17618;
  assign n24329 = pi20 ? n139 : n24328;
  assign n24330 = pi19 ? n24329 : n32;
  assign n24331 = pi18 ? n23753 : n24330;
  assign n24332 = pi17 ? n23752 : n24331;
  assign n24333 = pi16 ? n439 : n24332;
  assign n24334 = pi15 ? n24327 : n24333;
  assign n24335 = pi18 ? n23772 : n24330;
  assign n24336 = pi17 ? n23769 : n24335;
  assign n24337 = pi16 ? n23764 : n24336;
  assign n24338 = pi22 ? n20307 : n32;
  assign n24339 = pi21 ? n139 : n24338;
  assign n24340 = pi20 ? n139 : n24339;
  assign n24341 = pi19 ? n24340 : n32;
  assign n24342 = pi18 ? n23779 : n24341;
  assign n24343 = pi17 ? n23778 : n24342;
  assign n24344 = pi16 ? n439 : n24343;
  assign n24345 = pi15 ? n24337 : n24344;
  assign n24346 = pi14 ? n24334 : n24345;
  assign n24347 = pi21 ? n363 : n2835;
  assign n24348 = pi20 ? n139 : n24347;
  assign n24349 = pi19 ? n24348 : n32;
  assign n24350 = pi18 ? n13193 : n24349;
  assign n24351 = pi17 ? n37 : n24350;
  assign n24352 = pi16 ? n439 : n24351;
  assign n24353 = pi21 ? n363 : n3125;
  assign n24354 = pi20 ? n139 : n24353;
  assign n24355 = pi19 ? n24354 : n32;
  assign n24356 = pi18 ? n14115 : n24355;
  assign n24357 = pi17 ? n37 : n24356;
  assign n24358 = pi16 ? n439 : n24357;
  assign n24359 = pi15 ? n24352 : n24358;
  assign n24360 = pi21 ? n204 : n16358;
  assign n24361 = pi20 ? n204 : n24360;
  assign n24362 = pi19 ? n24361 : n32;
  assign n24363 = pi18 ? n22776 : n24362;
  assign n24364 = pi17 ? n37 : n24363;
  assign n24365 = pi16 ? n439 : n24364;
  assign n24366 = pi15 ? n24365 : n23808;
  assign n24367 = pi14 ? n24359 : n24366;
  assign n24368 = pi13 ? n24346 : n24367;
  assign n24369 = pi12 ? n24322 : n24368;
  assign n24370 = pi19 ? n5357 : n32;
  assign n24371 = pi18 ? n23802 : n24370;
  assign n24372 = pi17 ? n37 : n24371;
  assign n24373 = pi16 ? n439 : n24372;
  assign n24374 = pi21 ? n11199 : n335;
  assign n24375 = pi20 ? n37 : n24374;
  assign n24376 = pi19 ? n37 : n24375;
  assign n24377 = pi22 ? n450 : n233;
  assign n24378 = pi21 ? n6361 : n24377;
  assign n24379 = pi21 ? n6376 : n928;
  assign n24380 = pi20 ? n24378 : n24379;
  assign n24381 = pi19 ? n24380 : n32;
  assign n24382 = pi18 ? n24376 : n24381;
  assign n24383 = pi17 ? n37 : n24382;
  assign n24384 = pi16 ? n439 : n24383;
  assign n24385 = pi15 ? n24373 : n24384;
  assign n24386 = pi21 ? n2061 : n2469;
  assign n24387 = pi20 ? n335 : n24386;
  assign n24388 = pi19 ? n24387 : n32;
  assign n24389 = pi18 ? n21770 : n24388;
  assign n24390 = pi17 ? n37 : n24389;
  assign n24391 = pi16 ? n439 : n24390;
  assign n24392 = pi21 ? n2061 : n2553;
  assign n24393 = pi20 ? n335 : n24392;
  assign n24394 = pi19 ? n24393 : n32;
  assign n24395 = pi18 ? n21770 : n24394;
  assign n24396 = pi17 ? n37 : n24395;
  assign n24397 = pi16 ? n439 : n24396;
  assign n24398 = pi15 ? n24391 : n24397;
  assign n24399 = pi14 ? n24385 : n24398;
  assign n24400 = pi18 ? n17205 : n24394;
  assign n24401 = pi17 ? n37 : n24400;
  assign n24402 = pi16 ? n439 : n24401;
  assign n24403 = pi22 ? n335 : n6961;
  assign n24404 = pi21 ? n24403 : n2678;
  assign n24405 = pi20 ? n335 : n24404;
  assign n24406 = pi19 ? n24405 : n32;
  assign n24407 = pi18 ? n23839 : n24406;
  assign n24408 = pi17 ? n37 : n24407;
  assign n24409 = pi16 ? n439 : n24408;
  assign n24410 = pi15 ? n24402 : n24409;
  assign n24411 = pi18 ? n23845 : n24406;
  assign n24412 = pi17 ? n37 : n24411;
  assign n24413 = pi16 ? n439 : n24412;
  assign n24414 = pi24 ? n363 : n233;
  assign n24415 = pi23 ? n335 : n24414;
  assign n24416 = pi22 ? n335 : n24415;
  assign n24417 = pi21 ? n24416 : n2678;
  assign n24418 = pi20 ? n569 : n24417;
  assign n24419 = pi19 ? n24418 : n32;
  assign n24420 = pi18 ? n23850 : n24419;
  assign n24421 = pi17 ? n37 : n24420;
  assign n24422 = pi16 ? n439 : n24421;
  assign n24423 = pi15 ? n24413 : n24422;
  assign n24424 = pi14 ? n24410 : n24423;
  assign n24425 = pi13 ? n24399 : n24424;
  assign n24426 = pi21 ? n11336 : n2678;
  assign n24427 = pi20 ? n649 : n24426;
  assign n24428 = pi19 ? n24427 : n32;
  assign n24429 = pi18 ? n37 : n24428;
  assign n24430 = pi17 ? n37 : n24429;
  assign n24431 = pi16 ? n439 : n24430;
  assign n24432 = pi21 ? n233 : n2700;
  assign n24433 = pi20 ? n2094 : n24432;
  assign n24434 = pi19 ? n24433 : n32;
  assign n24435 = pi18 ? n37 : n24434;
  assign n24436 = pi17 ? n37 : n24435;
  assign n24437 = pi16 ? n439 : n24436;
  assign n24438 = pi15 ? n24431 : n24437;
  assign n24439 = pi21 ? n18411 : n2700;
  assign n24440 = pi20 ? n2094 : n24439;
  assign n24441 = pi19 ? n24440 : n32;
  assign n24442 = pi18 ? n37 : n24441;
  assign n24443 = pi17 ? n37 : n24442;
  assign n24444 = pi16 ? n439 : n24443;
  assign n24445 = pi20 ? n37 : n20237;
  assign n24446 = pi19 ? n24445 : n32;
  assign n24447 = pi18 ? n37 : n24446;
  assign n24448 = pi17 ? n37 : n24447;
  assign n24449 = pi16 ? n439 : n24448;
  assign n24450 = pi15 ? n24444 : n24449;
  assign n24451 = pi14 ? n24438 : n24450;
  assign n24452 = pi20 ? n37 : n12925;
  assign n24453 = pi19 ? n24452 : n32;
  assign n24454 = pi18 ? n37 : n24453;
  assign n24455 = pi17 ? n37 : n24454;
  assign n24456 = pi16 ? n439 : n24455;
  assign n24457 = pi22 ? n685 : n16771;
  assign n24458 = pi21 ? n24457 : n32;
  assign n24459 = pi20 ? n9660 : n24458;
  assign n24460 = pi19 ? n24459 : n32;
  assign n24461 = pi18 ? n37 : n24460;
  assign n24462 = pi17 ? n37 : n24461;
  assign n24463 = pi16 ? n439 : n24462;
  assign n24464 = pi15 ? n24456 : n24463;
  assign n24465 = pi22 ? n363 : n1511;
  assign n24466 = pi21 ? n24465 : n32;
  assign n24467 = pi20 ? n21826 : n24466;
  assign n24468 = pi19 ? n24467 : n32;
  assign n24469 = pi18 ? n37 : n24468;
  assign n24470 = pi17 ? n37 : n24469;
  assign n24471 = pi16 ? n439 : n24470;
  assign n24472 = pi20 ? n363 : n24466;
  assign n24473 = pi19 ? n24472 : n32;
  assign n24474 = pi18 ? n23904 : n24473;
  assign n24475 = pi17 ? n37 : n24474;
  assign n24476 = pi16 ? n439 : n24475;
  assign n24477 = pi15 ? n24471 : n24476;
  assign n24478 = pi14 ? n24464 : n24477;
  assign n24479 = pi13 ? n24451 : n24478;
  assign n24480 = pi12 ? n24425 : n24479;
  assign n24481 = pi11 ? n24369 : n24480;
  assign n24482 = pi20 ? n363 : n11695;
  assign n24483 = pi19 ? n24482 : n32;
  assign n24484 = pi18 ? n23918 : n24483;
  assign n24485 = pi17 ? n37 : n24484;
  assign n24486 = pi16 ? n439 : n24485;
  assign n24487 = pi20 ? n363 : n10311;
  assign n24488 = pi19 ? n24487 : n32;
  assign n24489 = pi18 ? n22898 : n24488;
  assign n24490 = pi17 ? n37 : n24489;
  assign n24491 = pi16 ? n439 : n24490;
  assign n24492 = pi15 ? n24486 : n24491;
  assign n24493 = pi21 ? n37 : n244;
  assign n24494 = pi20 ? n37 : n24493;
  assign n24495 = pi19 ? n24494 : n23930;
  assign n24496 = pi20 ? n23933 : n11695;
  assign n24497 = pi19 ? n24496 : n32;
  assign n24498 = pi18 ? n24495 : n24497;
  assign n24499 = pi17 ? n37 : n24498;
  assign n24500 = pi16 ? n439 : n24499;
  assign n24501 = pi22 ? n893 : n37;
  assign n24502 = pi21 ? n24501 : n23932;
  assign n24503 = pi20 ? n37 : n24502;
  assign n24504 = pi21 ? n6433 : n8654;
  assign n24505 = pi20 ? n23941 : n24504;
  assign n24506 = pi19 ? n24503 : n24505;
  assign n24507 = pi21 ? n22379 : n218;
  assign n24508 = pi20 ? n24507 : n11695;
  assign n24509 = pi19 ? n24508 : n32;
  assign n24510 = pi18 ? n24506 : n24509;
  assign n24511 = pi17 ? n37 : n24510;
  assign n24512 = pi16 ? n439 : n24511;
  assign n24513 = pi15 ? n24500 : n24512;
  assign n24514 = pi14 ? n24492 : n24513;
  assign n24515 = pi20 ? n5467 : n11695;
  assign n24516 = pi19 ? n24515 : n32;
  assign n24517 = pi18 ? n99 : n24516;
  assign n24518 = pi17 ? n99 : n24517;
  assign n24519 = pi16 ? n744 : n24518;
  assign n24520 = pi20 ? n5085 : n11695;
  assign n24521 = pi19 ? n24520 : n32;
  assign n24522 = pi18 ? n23959 : n24521;
  assign n24523 = pi17 ? n99 : n24522;
  assign n24524 = pi16 ? n744 : n24523;
  assign n24525 = pi15 ? n24519 : n24524;
  assign n24526 = pi20 ? n2238 : n6935;
  assign n24527 = pi19 ? n24526 : n32;
  assign n24528 = pi18 ? n99 : n24527;
  assign n24529 = pi17 ? n99 : n24528;
  assign n24530 = pi16 ? n744 : n24529;
  assign n24531 = pi14 ? n24525 : n24530;
  assign n24532 = pi13 ? n24514 : n24531;
  assign n24533 = pi20 ? n777 : n4008;
  assign n24534 = pi19 ? n24533 : n32;
  assign n24535 = pi18 ? n99 : n24534;
  assign n24536 = pi17 ? n99 : n24535;
  assign n24537 = pi16 ? n744 : n24536;
  assign n24538 = pi20 ? n2243 : n4008;
  assign n24539 = pi19 ? n24538 : n32;
  assign n24540 = pi18 ? n99 : n24539;
  assign n24541 = pi17 ? n99 : n24540;
  assign n24542 = pi16 ? n744 : n24541;
  assign n24543 = pi15 ? n24537 : n24542;
  assign n24544 = pi20 ? n19171 : n7733;
  assign n24545 = pi19 ? n24544 : n32;
  assign n24546 = pi18 ? n22967 : n24545;
  assign n24547 = pi17 ? n99 : n24546;
  assign n24548 = pi16 ? n744 : n24547;
  assign n24549 = pi22 ? n1228 : n32;
  assign n24550 = pi21 ? n24549 : n32;
  assign n24551 = pi20 ? n10033 : n24550;
  assign n24552 = pi19 ? n24551 : n32;
  assign n24553 = pi18 ? n23993 : n24552;
  assign n24554 = pi17 ? n139 : n24553;
  assign n24555 = pi16 ? n915 : n24554;
  assign n24556 = pi15 ? n24548 : n24555;
  assign n24557 = pi14 ? n24543 : n24556;
  assign n24558 = pi16 ? n915 : n24007;
  assign n24559 = pi15 ? n24558 : n24031;
  assign n24560 = pi22 ? n21494 : n204;
  assign n24561 = pi21 ? n24560 : n204;
  assign n24562 = pi20 ? n32 : n24561;
  assign n24563 = pi19 ? n32 : n24562;
  assign n24564 = pi18 ? n24563 : n204;
  assign n24565 = pi17 ? n32 : n24564;
  assign n24566 = pi16 ? n24565 : n24037;
  assign n24567 = pi15 ? n24566 : n24042;
  assign n24568 = pi14 ? n24559 : n24567;
  assign n24569 = pi13 ? n24557 : n24568;
  assign n24570 = pi12 ? n24532 : n24569;
  assign n24571 = pi20 ? n23048 : n10011;
  assign n24572 = pi19 ? n24571 : n32;
  assign n24573 = pi18 ? n24054 : n24572;
  assign n24574 = pi17 ? n139 : n24573;
  assign n24575 = pi16 ? n331 : n24574;
  assign n24576 = pi15 ? n24053 : n24575;
  assign n24577 = pi20 ? n24061 : n2653;
  assign n24578 = pi19 ? n24577 : n32;
  assign n24579 = pi18 ? n139 : n24578;
  assign n24580 = pi17 ? n139 : n24579;
  assign n24581 = pi16 ? n331 : n24580;
  assign n24582 = pi20 ? n24067 : n2653;
  assign n24583 = pi19 ? n24582 : n32;
  assign n24584 = pi18 ? n23054 : n24583;
  assign n24585 = pi17 ? n139 : n24584;
  assign n24586 = pi16 ? n331 : n24585;
  assign n24587 = pi15 ? n24581 : n24586;
  assign n24588 = pi14 ? n24576 : n24587;
  assign n24589 = pi16 ? n2035 : n24078;
  assign n24590 = pi21 ? n233 : n12659;
  assign n24591 = pi20 ? n24590 : n32;
  assign n24592 = pi19 ? n24591 : n32;
  assign n24593 = pi18 ? n24080 : n24592;
  assign n24594 = pi17 ? n335 : n24593;
  assign n24595 = pi16 ? n2035 : n24594;
  assign n24596 = pi15 ? n24589 : n24595;
  assign n24597 = pi14 ? n24596 : n24098;
  assign n24598 = pi13 ? n24588 : n24597;
  assign n24599 = pi21 ? n12643 : n14865;
  assign n24600 = pi20 ? n32 : n24599;
  assign n24601 = pi19 ? n32 : n24600;
  assign n24602 = pi22 ? n1656 : n4543;
  assign n24603 = pi21 ? n24602 : n14865;
  assign n24604 = pi21 ? n722 : n14865;
  assign n24605 = pi20 ? n24603 : n24604;
  assign n24606 = pi23 ? n233 : n99;
  assign n24607 = pi22 ? n363 : n24606;
  assign n24608 = pi21 ? n24607 : n22549;
  assign n24609 = pi20 ? n24151 : n24608;
  assign n24610 = pi19 ? n24605 : n24609;
  assign n24611 = pi18 ? n24601 : n24610;
  assign n24612 = pi17 ? n32 : n24611;
  assign n24613 = pi20 ? n22549 : n23150;
  assign n24614 = pi19 ? n24613 : n24160;
  assign n24615 = pi18 ? n24614 : n24166;
  assign n24616 = pi22 ? n24606 : n233;
  assign n24617 = pi21 ? n24616 : n233;
  assign n24618 = pi20 ? n233 : n24617;
  assign n24619 = pi19 ? n233 : n24618;
  assign n24620 = pi18 ? n24619 : n24173;
  assign n24621 = pi17 ? n24615 : n24620;
  assign n24622 = pi16 ? n24612 : n24621;
  assign n24623 = pi18 ? n233 : n14659;
  assign n24624 = pi17 ? n24187 : n24623;
  assign n24625 = pi16 ? n24180 : n24624;
  assign n24626 = pi15 ? n24622 : n24625;
  assign n24627 = pi18 ? n19433 : n23176;
  assign n24628 = pi17 ? n32 : n24627;
  assign n24629 = pi21 ? n233 : n1476;
  assign n24630 = pi20 ? n24629 : n32;
  assign n24631 = pi19 ? n24630 : n32;
  assign n24632 = pi18 ? n233 : n24631;
  assign n24633 = pi17 ? n24207 : n24632;
  assign n24634 = pi16 ? n24628 : n24633;
  assign n24635 = pi18 ? n24225 : n14700;
  assign n24636 = pi17 ? n24219 : n24635;
  assign n24637 = pi16 ? n21219 : n24636;
  assign n24638 = pi15 ? n24634 : n24637;
  assign n24639 = pi14 ? n24626 : n24638;
  assign n24640 = pi13 ? n24142 : n24639;
  assign n24641 = pi12 ? n24598 : n24640;
  assign n24642 = pi11 ? n24570 : n24641;
  assign n24643 = pi10 ? n24481 : n24642;
  assign n24644 = pi09 ? n24244 : n24643;
  assign n24645 = pi08 ? n24235 : n24644;
  assign n24646 = pi07 ? n23594 : n24645;
  assign n24647 = pi20 ? n37 : n10432;
  assign n24648 = pi19 ? n24647 : n32;
  assign n24649 = pi18 ? n37 : n24648;
  assign n24650 = pi17 ? n37 : n24649;
  assign n24651 = pi16 ? n14445 : n24650;
  assign n24652 = pi15 ? n32 : n24651;
  assign n24653 = pi20 ? n37 : n10447;
  assign n24654 = pi19 ? n24653 : n32;
  assign n24655 = pi18 ? n37 : n24654;
  assign n24656 = pi17 ? n37 : n24655;
  assign n24657 = pi16 ? n14445 : n24656;
  assign n24658 = pi21 ? n2161 : n4559;
  assign n24659 = pi20 ? n2974 : n24658;
  assign n24660 = pi19 ? n24659 : n32;
  assign n24661 = pi18 ? n37 : n24660;
  assign n24662 = pi17 ? n37 : n24661;
  assign n24663 = pi16 ? n16595 : n24662;
  assign n24664 = pi15 ? n24657 : n24663;
  assign n24665 = pi14 ? n24652 : n24664;
  assign n24666 = pi13 ? n32 : n24665;
  assign n24667 = pi12 ? n32 : n24666;
  assign n24668 = pi11 ? n32 : n24667;
  assign n24669 = pi10 ? n32 : n24668;
  assign n24670 = pi21 ? n181 : n10453;
  assign n24671 = pi20 ? n5077 : n24670;
  assign n24672 = pi19 ? n24671 : n32;
  assign n24673 = pi18 ? n37 : n24672;
  assign n24674 = pi17 ? n37 : n24673;
  assign n24675 = pi16 ? n16595 : n24674;
  assign n24676 = pi21 ? n181 : n11393;
  assign n24677 = pi20 ? n37 : n24676;
  assign n24678 = pi19 ? n24677 : n32;
  assign n24679 = pi18 ? n37 : n24678;
  assign n24680 = pi17 ? n37 : n24679;
  assign n24681 = pi16 ? n17010 : n24680;
  assign n24682 = pi15 ? n24675 : n24681;
  assign n24683 = pi21 ? n37 : n17994;
  assign n24684 = pi20 ? n37 : n24683;
  assign n24685 = pi19 ? n24684 : n32;
  assign n24686 = pi18 ? n37 : n24685;
  assign n24687 = pi17 ? n37 : n24686;
  assign n24688 = pi16 ? n17010 : n24687;
  assign n24689 = pi21 ? n37 : n18008;
  assign n24690 = pi20 ? n37 : n24689;
  assign n24691 = pi19 ? n24690 : n32;
  assign n24692 = pi18 ? n37 : n24691;
  assign n24693 = pi17 ? n37 : n24692;
  assign n24694 = pi16 ? n439 : n24693;
  assign n24695 = pi15 ? n24688 : n24694;
  assign n24696 = pi14 ? n24682 : n24695;
  assign n24697 = pi18 ? n374 : n99;
  assign n24698 = pi17 ? n32 : n24697;
  assign n24699 = pi20 ? n99 : n10512;
  assign n24700 = pi19 ? n24699 : n32;
  assign n24701 = pi18 ? n99 : n24700;
  assign n24702 = pi17 ? n99 : n24701;
  assign n24703 = pi16 ? n24698 : n24702;
  assign n24704 = pi18 ? n3031 : n21612;
  assign n24705 = pi17 ? n32 : n24704;
  assign n24706 = pi16 ? n24705 : n24307;
  assign n24707 = pi15 ? n24703 : n24706;
  assign n24708 = pi20 ? n3882 : n14887;
  assign n24709 = pi20 ? n7745 : n2973;
  assign n24710 = pi19 ? n24708 : n24709;
  assign n24711 = pi18 ? n374 : n24710;
  assign n24712 = pi17 ? n32 : n24711;
  assign n24713 = pi20 ? n14844 : n14846;
  assign n24714 = pi19 ? n24713 : n139;
  assign n24715 = pi18 ? n24714 : n139;
  assign n24716 = pi21 ? n139 : n3848;
  assign n24717 = pi20 ? n139 : n24716;
  assign n24718 = pi19 ? n24717 : n32;
  assign n24719 = pi18 ? n139 : n24718;
  assign n24720 = pi17 ? n24715 : n24719;
  assign n24721 = pi16 ? n24712 : n24720;
  assign n24722 = pi18 ? n9815 : n139;
  assign n24723 = pi17 ? n24722 : n24325;
  assign n24724 = pi16 ? n439 : n24723;
  assign n24725 = pi15 ? n24721 : n24724;
  assign n24726 = pi14 ? n24707 : n24725;
  assign n24727 = pi13 ? n24696 : n24726;
  assign n24728 = pi17 ? n10653 : n24325;
  assign n24729 = pi16 ? n439 : n24728;
  assign n24730 = pi19 ? n13094 : n139;
  assign n24731 = pi18 ? n24730 : n24330;
  assign n24732 = pi17 ? n11568 : n24731;
  assign n24733 = pi16 ? n439 : n24732;
  assign n24734 = pi15 ? n24729 : n24733;
  assign n24735 = pi19 ? n37 : n3103;
  assign n24736 = pi18 ? n37 : n24735;
  assign n24737 = pi18 ? n13193 : n24330;
  assign n24738 = pi17 ? n24736 : n24737;
  assign n24739 = pi16 ? n439 : n24738;
  assign n24740 = pi18 ? n14115 : n24341;
  assign n24741 = pi17 ? n37 : n24740;
  assign n24742 = pi16 ? n439 : n24741;
  assign n24743 = pi15 ? n24739 : n24742;
  assign n24744 = pi14 ? n24734 : n24743;
  assign n24745 = pi21 ? n37 : n2320;
  assign n24746 = pi20 ? n1583 : n24745;
  assign n24747 = pi19 ? n24746 : n32;
  assign n24748 = pi18 ? n37 : n24747;
  assign n24749 = pi17 ? n37 : n24748;
  assign n24750 = pi16 ? n439 : n24749;
  assign n24751 = pi20 ? n2644 : n204;
  assign n24752 = pi19 ? n37 : n24751;
  assign n24753 = pi18 ? n24752 : n24362;
  assign n24754 = pi17 ? n37 : n24753;
  assign n24755 = pi16 ? n439 : n24754;
  assign n24756 = pi15 ? n24750 : n24755;
  assign n24757 = pi21 ? n204 : n3175;
  assign n24758 = pi20 ? n204 : n24757;
  assign n24759 = pi19 ? n24758 : n32;
  assign n24760 = pi18 ? n23802 : n24759;
  assign n24761 = pi17 ? n37 : n24760;
  assign n24762 = pi16 ? n439 : n24761;
  assign n24763 = pi20 ? n37 : n2316;
  assign n24764 = pi19 ? n37 : n24763;
  assign n24765 = pi18 ? n24764 : n24759;
  assign n24766 = pi17 ? n37 : n24765;
  assign n24767 = pi16 ? n439 : n24766;
  assign n24768 = pi15 ? n24762 : n24767;
  assign n24769 = pi14 ? n24756 : n24768;
  assign n24770 = pi13 ? n24744 : n24769;
  assign n24771 = pi12 ? n24727 : n24770;
  assign n24772 = pi21 ? n11808 : n233;
  assign n24773 = pi20 ? n37 : n24772;
  assign n24774 = pi19 ? n37 : n24773;
  assign n24775 = pi21 ? n233 : n2565;
  assign n24776 = pi20 ? n233 : n24775;
  assign n24777 = pi19 ? n24776 : n32;
  assign n24778 = pi18 ? n24774 : n24777;
  assign n24779 = pi17 ? n37 : n24778;
  assign n24780 = pi16 ? n439 : n24779;
  assign n24781 = pi21 ? n335 : n2578;
  assign n24782 = pi20 ? n335 : n24781;
  assign n24783 = pi19 ? n24782 : n32;
  assign n24784 = pi18 ? n17205 : n24783;
  assign n24785 = pi17 ? n37 : n24784;
  assign n24786 = pi16 ? n439 : n24785;
  assign n24787 = pi15 ? n24780 : n24786;
  assign n24788 = pi20 ? n37 : n603;
  assign n24789 = pi19 ? n37 : n24788;
  assign n24790 = pi18 ? n24789 : n24783;
  assign n24791 = pi17 ? n37 : n24790;
  assign n24792 = pi16 ? n439 : n24791;
  assign n24793 = pi20 ? n569 : n24781;
  assign n24794 = pi19 ? n24793 : n32;
  assign n24795 = pi18 ? n7686 : n24794;
  assign n24796 = pi17 ? n37 : n24795;
  assign n24797 = pi16 ? n439 : n24796;
  assign n24798 = pi15 ? n24792 : n24797;
  assign n24799 = pi14 ? n24787 : n24798;
  assign n24800 = pi18 ? n37 : n24794;
  assign n24801 = pi17 ? n37 : n24800;
  assign n24802 = pi16 ? n439 : n24801;
  assign n24803 = pi20 ? n37 : n24781;
  assign n24804 = pi19 ? n24803 : n32;
  assign n24805 = pi18 ? n37 : n24804;
  assign n24806 = pi17 ? n37 : n24805;
  assign n24807 = pi16 ? n439 : n24806;
  assign n24808 = pi21 ? n3392 : n2578;
  assign n24809 = pi20 ? n37 : n24808;
  assign n24810 = pi19 ? n24809 : n32;
  assign n24811 = pi18 ? n37 : n24810;
  assign n24812 = pi17 ? n37 : n24811;
  assign n24813 = pi16 ? n439 : n24812;
  assign n24814 = pi15 ? n24807 : n24813;
  assign n24815 = pi14 ? n24802 : n24814;
  assign n24816 = pi13 ? n24799 : n24815;
  assign n24817 = pi21 ? n233 : n4147;
  assign n24818 = pi20 ? n2091 : n24817;
  assign n24819 = pi19 ? n24818 : n32;
  assign n24820 = pi18 ? n2102 : n24819;
  assign n24821 = pi17 ? n37 : n24820;
  assign n24822 = pi16 ? n439 : n24821;
  assign n24823 = pi20 ? n37 : n23203;
  assign n24824 = pi19 ? n24823 : n32;
  assign n24825 = pi18 ? n37 : n24824;
  assign n24826 = pi17 ? n37 : n24825;
  assign n24827 = pi16 ? n439 : n24826;
  assign n24828 = pi15 ? n24822 : n24827;
  assign n24829 = pi20 ? n37 : n21547;
  assign n24830 = pi19 ? n24829 : n32;
  assign n24831 = pi18 ? n37 : n24830;
  assign n24832 = pi17 ? n37 : n24831;
  assign n24833 = pi16 ? n439 : n24832;
  assign n24834 = pi23 ? n685 : n37;
  assign n24835 = pi22 ? n24834 : n685;
  assign n24836 = pi21 ? n24835 : n928;
  assign n24837 = pi20 ? n37 : n24836;
  assign n24838 = pi19 ? n24837 : n32;
  assign n24839 = pi18 ? n37 : n24838;
  assign n24840 = pi17 ? n37 : n24839;
  assign n24841 = pi16 ? n439 : n24840;
  assign n24842 = pi15 ? n24833 : n24841;
  assign n24843 = pi14 ? n24828 : n24842;
  assign n24844 = pi21 ? n381 : n1009;
  assign n24845 = pi20 ? n37 : n24844;
  assign n24846 = pi19 ? n24845 : n32;
  assign n24847 = pi18 ? n37 : n24846;
  assign n24848 = pi17 ? n37 : n24847;
  assign n24849 = pi16 ? n439 : n24848;
  assign n24850 = pi21 ? n381 : n32;
  assign n24851 = pi20 ? n37 : n24850;
  assign n24852 = pi19 ? n24851 : n32;
  assign n24853 = pi18 ? n37 : n24852;
  assign n24854 = pi17 ? n37 : n24853;
  assign n24855 = pi16 ? n439 : n24854;
  assign n24856 = pi15 ? n24849 : n24855;
  assign n24857 = pi23 ? n363 : n2766;
  assign n24858 = pi22 ? n37 : n24857;
  assign n24859 = pi21 ? n24858 : n32;
  assign n24860 = pi20 ? n37 : n24859;
  assign n24861 = pi19 ? n24860 : n32;
  assign n24862 = pi18 ? n37 : n24861;
  assign n24863 = pi17 ? n37 : n24862;
  assign n24864 = pi16 ? n439 : n24863;
  assign n24865 = pi21 ? n3392 : n363;
  assign n24866 = pi20 ? n37 : n24865;
  assign n24867 = pi19 ? n24866 : n363;
  assign n24868 = pi22 ? n363 : n16771;
  assign n24869 = pi21 ? n24868 : n32;
  assign n24870 = pi20 ? n363 : n24869;
  assign n24871 = pi19 ? n24870 : n32;
  assign n24872 = pi18 ? n24867 : n24871;
  assign n24873 = pi17 ? n37 : n24872;
  assign n24874 = pi16 ? n439 : n24873;
  assign n24875 = pi15 ? n24864 : n24874;
  assign n24876 = pi14 ? n24856 : n24875;
  assign n24877 = pi13 ? n24843 : n24876;
  assign n24878 = pi12 ? n24816 : n24877;
  assign n24879 = pi11 ? n24771 : n24878;
  assign n24880 = pi20 ? n363 : n7730;
  assign n24881 = pi19 ? n7731 : n24880;
  assign n24882 = pi20 ? n7730 : n24466;
  assign n24883 = pi19 ? n24882 : n32;
  assign n24884 = pi18 ? n24881 : n24883;
  assign n24885 = pi17 ? n37 : n24884;
  assign n24886 = pi16 ? n439 : n24885;
  assign n24887 = pi20 ? n37 : n7327;
  assign n24888 = pi21 ? n5012 : n7334;
  assign n24889 = pi20 ? n24888 : n9670;
  assign n24890 = pi19 ? n24887 : n24889;
  assign n24891 = pi20 ? n3392 : n6898;
  assign n24892 = pi19 ? n24891 : n32;
  assign n24893 = pi18 ? n24890 : n24892;
  assign n24894 = pi17 ? n37 : n24893;
  assign n24895 = pi16 ? n439 : n24894;
  assign n24896 = pi15 ? n24886 : n24895;
  assign n24897 = pi20 ? n37 : n10319;
  assign n24898 = pi19 ? n24897 : n32;
  assign n24899 = pi18 ? n37 : n24898;
  assign n24900 = pi17 ? n37 : n24899;
  assign n24901 = pi16 ? n439 : n24900;
  assign n24902 = pi20 ? n37 : n278;
  assign n24903 = pi19 ? n24902 : n157;
  assign n24904 = pi22 ? n157 : n10784;
  assign n24905 = pi21 ? n24904 : n32;
  assign n24906 = pi20 ? n157 : n24905;
  assign n24907 = pi19 ? n24906 : n32;
  assign n24908 = pi18 ? n24903 : n24907;
  assign n24909 = pi17 ? n37 : n24908;
  assign n24910 = pi16 ? n439 : n24909;
  assign n24911 = pi15 ? n24901 : n24910;
  assign n24912 = pi14 ? n24896 : n24911;
  assign n24913 = pi20 ? n5085 : n99;
  assign n24914 = pi19 ? n99 : n24913;
  assign n24915 = pi20 ? n99 : n11695;
  assign n24916 = pi19 ? n24915 : n32;
  assign n24917 = pi18 ? n24914 : n24916;
  assign n24918 = pi17 ? n99 : n24917;
  assign n24919 = pi16 ? n721 : n24918;
  assign n24920 = pi21 ? n3444 : n99;
  assign n24921 = pi20 ? n24920 : n99;
  assign n24922 = pi19 ? n99 : n24921;
  assign n24923 = pi21 ? n3453 : n32;
  assign n24924 = pi20 ? n99 : n24923;
  assign n24925 = pi19 ? n24924 : n32;
  assign n24926 = pi18 ? n24922 : n24925;
  assign n24927 = pi17 ? n99 : n24926;
  assign n24928 = pi16 ? n721 : n24927;
  assign n24929 = pi15 ? n24919 : n24928;
  assign n24930 = pi20 ? n99 : n6935;
  assign n24931 = pi19 ? n24930 : n32;
  assign n24932 = pi18 ? n99 : n24931;
  assign n24933 = pi17 ? n99 : n24932;
  assign n24934 = pi16 ? n721 : n24933;
  assign n24935 = pi14 ? n24929 : n24934;
  assign n24936 = pi13 ? n24912 : n24935;
  assign n24937 = pi21 ? n16317 : n32;
  assign n24938 = pi20 ? n2238 : n24937;
  assign n24939 = pi19 ? n24938 : n32;
  assign n24940 = pi18 ? n99 : n24939;
  assign n24941 = pi17 ? n99 : n24940;
  assign n24942 = pi16 ? n721 : n24941;
  assign n24943 = pi20 ? n19208 : n99;
  assign n24944 = pi19 ? n99 : n24943;
  assign n24945 = pi18 ? n24944 : n24939;
  assign n24946 = pi17 ? n99 : n24945;
  assign n24947 = pi16 ? n721 : n24946;
  assign n24948 = pi15 ? n24942 : n24947;
  assign n24949 = pi21 ? n716 : n139;
  assign n24950 = pi20 ? n32 : n24949;
  assign n24951 = pi19 ? n32 : n24950;
  assign n24952 = pi18 ? n24951 : n139;
  assign n24953 = pi17 ? n32 : n24952;
  assign n24954 = pi21 ? n17375 : n139;
  assign n24955 = pi20 ? n19208 : n24954;
  assign n24956 = pi19 ? n139 : n24955;
  assign n24957 = pi21 ? n99 : n20977;
  assign n24958 = pi20 ? n24957 : n3210;
  assign n24959 = pi19 ? n24958 : n32;
  assign n24960 = pi18 ? n24956 : n24959;
  assign n24961 = pi17 ? n139 : n24960;
  assign n24962 = pi16 ? n24953 : n24961;
  assign n24963 = pi19 ? n139 : n18330;
  assign n24964 = pi20 ? n1026 : n3210;
  assign n24965 = pi19 ? n24964 : n32;
  assign n24966 = pi18 ? n24963 : n24965;
  assign n24967 = pi17 ? n139 : n24966;
  assign n24968 = pi16 ? n2291 : n24967;
  assign n24969 = pi15 ? n24962 : n24968;
  assign n24970 = pi14 ? n24948 : n24969;
  assign n24971 = pi21 ? n204 : n4015;
  assign n24972 = pi20 ? n204 : n24971;
  assign n24973 = pi19 ? n204 : n24972;
  assign n24974 = pi20 ? n21732 : n37;
  assign n24975 = pi19 ? n24974 : n204;
  assign n24976 = pi18 ? n24973 : n24975;
  assign n24977 = pi19 ? n19231 : n316;
  assign n24978 = pi20 ? n316 : n3210;
  assign n24979 = pi19 ? n24978 : n32;
  assign n24980 = pi18 ? n24977 : n24979;
  assign n24981 = pi17 ? n24976 : n24980;
  assign n24982 = pi16 ? n11804 : n24981;
  assign n24983 = pi20 ? n204 : n21732;
  assign n24984 = pi19 ? n24983 : n204;
  assign n24985 = pi18 ? n24973 : n24984;
  assign n24986 = pi19 ? n3727 : n316;
  assign n24987 = pi18 ? n24986 : n24979;
  assign n24988 = pi17 ? n24985 : n24987;
  assign n24989 = pi16 ? n13846 : n24988;
  assign n24990 = pi15 ? n24982 : n24989;
  assign n24991 = pi21 ? n1046 : n1578;
  assign n24992 = pi20 ? n204 : n24991;
  assign n24993 = pi19 ? n24992 : n204;
  assign n24994 = pi18 ? n204 : n24993;
  assign n24995 = pi19 ? n204 : n316;
  assign n24996 = pi18 ? n24995 : n24979;
  assign n24997 = pi17 ? n24994 : n24996;
  assign n24998 = pi16 ? n13493 : n24997;
  assign n24999 = pi19 ? n20033 : n6645;
  assign n25000 = pi18 ? n24999 : n24979;
  assign n25001 = pi17 ? n24994 : n25000;
  assign n25002 = pi16 ? n13493 : n25001;
  assign n25003 = pi15 ? n24998 : n25002;
  assign n25004 = pi14 ? n24990 : n25003;
  assign n25005 = pi13 ? n24970 : n25004;
  assign n25006 = pi12 ? n24936 : n25005;
  assign n25007 = pi20 ? n14953 : n4116;
  assign n25008 = pi19 ? n25007 : n32;
  assign n25009 = pi18 ? n139 : n25008;
  assign n25010 = pi17 ? n139 : n25009;
  assign n25011 = pi16 ? n915 : n25010;
  assign n25012 = pi20 ? n1026 : n139;
  assign n25013 = pi19 ? n139 : n25012;
  assign n25014 = pi22 ? n139 : n2060;
  assign n25015 = pi21 ? n139 : n25014;
  assign n25016 = pi20 ? n25015 : n5830;
  assign n25017 = pi19 ? n25016 : n32;
  assign n25018 = pi18 ? n25013 : n25017;
  assign n25019 = pi17 ? n139 : n25018;
  assign n25020 = pi16 ? n915 : n25019;
  assign n25021 = pi15 ? n25011 : n25020;
  assign n25022 = pi19 ? n139 : n21978;
  assign n25023 = pi21 ? n139 : n17456;
  assign n25024 = pi20 ? n25023 : n2653;
  assign n25025 = pi19 ? n25024 : n32;
  assign n25026 = pi18 ? n25022 : n25025;
  assign n25027 = pi17 ? n139 : n25026;
  assign n25028 = pi16 ? n2291 : n25027;
  assign n25029 = pi22 ? n962 : n9123;
  assign n25030 = pi21 ? n25029 : n9122;
  assign n25031 = pi20 ? n32 : n25030;
  assign n25032 = pi19 ? n32 : n25031;
  assign n25033 = pi22 ? n1043 : n566;
  assign n25034 = pi21 ? n25033 : n9122;
  assign n25035 = pi20 ? n25034 : n1699;
  assign n25036 = pi21 ? n139 : n9126;
  assign n25037 = pi19 ? n25035 : n25036;
  assign n25038 = pi18 ? n25032 : n25037;
  assign n25039 = pi17 ? n32 : n25038;
  assign n25040 = pi21 ? n1698 : n9119;
  assign n25041 = pi21 ? n1698 : n9146;
  assign n25042 = pi20 ? n25040 : n25041;
  assign n25043 = pi19 ? n25040 : n25042;
  assign n25044 = pi21 ? n9119 : n9144;
  assign n25045 = pi21 ? n375 : n9144;
  assign n25046 = pi20 ? n25044 : n25045;
  assign n25047 = pi21 ? n9122 : n1698;
  assign n25048 = pi22 ? n9123 : n295;
  assign n25049 = pi21 ? n9122 : n25048;
  assign n25050 = pi20 ? n25047 : n25049;
  assign n25051 = pi19 ? n25046 : n25050;
  assign n25052 = pi18 ? n25043 : n25051;
  assign n25053 = pi21 ? n9143 : n204;
  assign n25054 = pi20 ? n9141 : n25053;
  assign n25055 = pi19 ? n25054 : n204;
  assign n25056 = pi21 ? n204 : n3763;
  assign n25057 = pi20 ? n25056 : n2653;
  assign n25058 = pi19 ? n25057 : n32;
  assign n25059 = pi18 ? n25055 : n25058;
  assign n25060 = pi17 ? n25052 : n25059;
  assign n25061 = pi16 ? n25039 : n25060;
  assign n25062 = pi15 ? n25028 : n25061;
  assign n25063 = pi14 ? n25021 : n25062;
  assign n25064 = pi21 ? n4990 : n335;
  assign n25065 = pi20 ? n25064 : n335;
  assign n25066 = pi19 ? n25065 : n335;
  assign n25067 = pi18 ? n10397 : n25066;
  assign n25068 = pi17 ? n32 : n25067;
  assign n25069 = pi20 ? n335 : n18121;
  assign n25070 = pi20 ? n20539 : n233;
  assign n25071 = pi19 ? n25069 : n25070;
  assign n25072 = pi20 ? n24590 : n1822;
  assign n25073 = pi19 ? n25072 : n32;
  assign n25074 = pi18 ? n25071 : n25073;
  assign n25075 = pi17 ? n335 : n25074;
  assign n25076 = pi16 ? n25068 : n25075;
  assign n25077 = pi21 ? n4990 : n37;
  assign n25078 = pi20 ? n25077 : n335;
  assign n25079 = pi19 ? n25078 : n335;
  assign n25080 = pi18 ? n10397 : n25079;
  assign n25081 = pi17 ? n32 : n25080;
  assign n25082 = pi19 ? n335 : n7981;
  assign n25083 = pi18 ? n25082 : n24592;
  assign n25084 = pi17 ? n335 : n25083;
  assign n25085 = pi16 ? n25081 : n25084;
  assign n25086 = pi15 ? n25076 : n25085;
  assign n25087 = pi20 ? n37 : n647;
  assign n25088 = pi19 ? n37 : n25087;
  assign n25089 = pi18 ? n374 : n25088;
  assign n25090 = pi17 ? n32 : n25089;
  assign n25091 = pi19 ? n2068 : n577;
  assign n25092 = pi18 ? n25088 : n25091;
  assign n25093 = pi19 ? n335 : n7985;
  assign n25094 = pi21 ? n6376 : n1389;
  assign n25095 = pi20 ? n25094 : n32;
  assign n25096 = pi19 ? n25095 : n32;
  assign n25097 = pi18 ? n25093 : n25096;
  assign n25098 = pi17 ? n25092 : n25097;
  assign n25099 = pi16 ? n25090 : n25098;
  assign n25100 = pi20 ? n233 : n6362;
  assign n25101 = pi19 ? n10681 : n25100;
  assign n25102 = pi18 ? n25101 : n25096;
  assign n25103 = pi17 ? n37 : n25102;
  assign n25104 = pi16 ? n439 : n25103;
  assign n25105 = pi15 ? n25099 : n25104;
  assign n25106 = pi14 ? n25086 : n25105;
  assign n25107 = pi13 ? n25063 : n25106;
  assign n25108 = pi22 ? n335 : n2116;
  assign n25109 = pi21 ? n37 : n25108;
  assign n25110 = pi20 ? n37 : n25109;
  assign n25111 = pi19 ? n37 : n25110;
  assign n25112 = pi18 ? n374 : n25111;
  assign n25113 = pi17 ? n32 : n25112;
  assign n25114 = pi19 ? n37 : n644;
  assign n25115 = pi18 ? n37 : n25114;
  assign n25116 = pi20 ? n3412 : n4921;
  assign n25117 = pi19 ? n25116 : n233;
  assign n25118 = pi21 ? n233 : n1389;
  assign n25119 = pi20 ? n25118 : n32;
  assign n25120 = pi19 ? n25119 : n32;
  assign n25121 = pi18 ? n25117 : n25120;
  assign n25122 = pi17 ? n25115 : n25121;
  assign n25123 = pi16 ? n25113 : n25122;
  assign n25124 = pi18 ? n8929 : n37;
  assign n25125 = pi21 ? n560 : n233;
  assign n25126 = pi20 ? n25125 : n233;
  assign n25127 = pi19 ? n25126 : n233;
  assign n25128 = pi21 ? n233 : n17509;
  assign n25129 = pi20 ? n25128 : n32;
  assign n25130 = pi19 ? n25129 : n32;
  assign n25131 = pi18 ? n25127 : n25130;
  assign n25132 = pi17 ? n25124 : n25131;
  assign n25133 = pi16 ? n439 : n25132;
  assign n25134 = pi15 ? n25123 : n25133;
  assign n25135 = pi19 ? n19358 : n233;
  assign n25136 = pi18 ? n25135 : n25130;
  assign n25137 = pi17 ? n25124 : n25136;
  assign n25138 = pi16 ? n439 : n25137;
  assign n25139 = pi21 ? n570 : n2048;
  assign n25140 = pi20 ? n3335 : n25139;
  assign n25141 = pi19 ? n7676 : n25140;
  assign n25142 = pi18 ? n3349 : n25141;
  assign n25143 = pi17 ? n32 : n25142;
  assign n25144 = pi20 ? n605 : n5023;
  assign n25145 = pi19 ? n647 : n25144;
  assign n25146 = pi21 ? n570 : n233;
  assign n25147 = pi20 ? n6360 : n25146;
  assign n25148 = pi22 ? n37 : n4899;
  assign n25149 = pi21 ? n25148 : n2048;
  assign n25150 = pi20 ? n603 : n25149;
  assign n25151 = pi19 ? n25147 : n25150;
  assign n25152 = pi18 ? n25145 : n25151;
  assign n25153 = pi20 ? n6377 : n7980;
  assign n25154 = pi19 ? n19416 : n25153;
  assign n25155 = pi20 ? n10982 : n32;
  assign n25156 = pi19 ? n25155 : n32;
  assign n25157 = pi18 ? n25154 : n25156;
  assign n25158 = pi17 ? n25152 : n25157;
  assign n25159 = pi16 ? n25143 : n25158;
  assign n25160 = pi15 ? n25138 : n25159;
  assign n25161 = pi14 ? n25134 : n25160;
  assign n25162 = pi22 ? n715 : n233;
  assign n25163 = pi21 ? n25162 : n233;
  assign n25164 = pi20 ? n32 : n25163;
  assign n25165 = pi19 ? n32 : n25164;
  assign n25166 = pi21 ? n233 : n99;
  assign n25167 = pi21 ? n99 : n363;
  assign n25168 = pi20 ? n25166 : n25167;
  assign n25169 = pi19 ? n25168 : n19423;
  assign n25170 = pi18 ? n25165 : n25169;
  assign n25171 = pi17 ? n32 : n25170;
  assign n25172 = pi19 ? n21222 : n233;
  assign n25173 = pi18 ? n25172 : n233;
  assign n25174 = pi22 ? n6365 : n396;
  assign n25175 = pi21 ? n233 : n25174;
  assign n25176 = pi20 ? n25175 : n32;
  assign n25177 = pi19 ? n25176 : n32;
  assign n25178 = pi18 ? n233 : n25177;
  assign n25179 = pi17 ? n25173 : n25178;
  assign n25180 = pi16 ? n25171 : n25179;
  assign n25181 = pi21 ? n363 : n99;
  assign n25182 = pi20 ? n25181 : n25167;
  assign n25183 = pi19 ? n25182 : n21225;
  assign n25184 = pi18 ? n23149 : n25183;
  assign n25185 = pi17 ? n32 : n25184;
  assign n25186 = pi20 ? n363 : n233;
  assign n25187 = pi19 ? n363 : n25186;
  assign n25188 = pi20 ? n233 : n19422;
  assign n25189 = pi20 ? n23175 : n233;
  assign n25190 = pi19 ? n25188 : n25189;
  assign n25191 = pi18 ? n25187 : n25190;
  assign n25192 = pi21 ? n5014 : n6366;
  assign n25193 = pi20 ? n25192 : n32;
  assign n25194 = pi19 ? n25193 : n32;
  assign n25195 = pi18 ? n21243 : n25194;
  assign n25196 = pi17 ? n25191 : n25195;
  assign n25197 = pi16 ? n25185 : n25196;
  assign n25198 = pi15 ? n25180 : n25197;
  assign n25199 = pi21 ? n363 : n685;
  assign n25200 = pi20 ? n25199 : n20866;
  assign n25201 = pi19 ? n363 : n25200;
  assign n25202 = pi21 ? n363 : n1476;
  assign n25203 = pi20 ? n25202 : n32;
  assign n25204 = pi19 ? n25203 : n32;
  assign n25205 = pi18 ? n25201 : n25204;
  assign n25206 = pi17 ? n363 : n25205;
  assign n25207 = pi16 ? n21219 : n25206;
  assign n25208 = pi20 ? n25199 : n363;
  assign n25209 = pi19 ? n363 : n25208;
  assign n25210 = pi21 ? n363 : n7048;
  assign n25211 = pi20 ? n25210 : n32;
  assign n25212 = pi19 ? n25211 : n32;
  assign n25213 = pi18 ? n25209 : n25212;
  assign n25214 = pi17 ? n363 : n25213;
  assign n25215 = pi16 ? n21219 : n25214;
  assign n25216 = pi15 ? n25207 : n25215;
  assign n25217 = pi14 ? n25198 : n25216;
  assign n25218 = pi13 ? n25161 : n25217;
  assign n25219 = pi12 ? n25107 : n25218;
  assign n25220 = pi11 ? n25006 : n25219;
  assign n25221 = pi10 ? n24879 : n25220;
  assign n25222 = pi09 ? n24669 : n25221;
  assign n25223 = pi21 ? n99 : n4559;
  assign n25224 = pi20 ? n2974 : n25223;
  assign n25225 = pi19 ? n25224 : n32;
  assign n25226 = pi18 ? n37 : n25225;
  assign n25227 = pi17 ? n37 : n25226;
  assign n25228 = pi16 ? n16595 : n25227;
  assign n25229 = pi15 ? n24657 : n25228;
  assign n25230 = pi14 ? n24652 : n25229;
  assign n25231 = pi13 ? n32 : n25230;
  assign n25232 = pi12 ? n32 : n25231;
  assign n25233 = pi11 ? n32 : n25232;
  assign n25234 = pi10 ? n32 : n25233;
  assign n25235 = pi21 ? n99 : n3832;
  assign n25236 = pi20 ? n99 : n25235;
  assign n25237 = pi19 ? n25236 : n32;
  assign n25238 = pi18 ? n99 : n25237;
  assign n25239 = pi17 ? n99 : n25238;
  assign n25240 = pi16 ? n24698 : n25239;
  assign n25241 = pi22 ? n158 : n32;
  assign n25242 = pi21 ? n99 : n25241;
  assign n25243 = pi20 ? n99 : n25242;
  assign n25244 = pi19 ? n25243 : n32;
  assign n25245 = pi18 ? n99 : n25244;
  assign n25246 = pi17 ? n99 : n25245;
  assign n25247 = pi16 ? n24705 : n25246;
  assign n25248 = pi15 ? n25240 : n25247;
  assign n25249 = pi21 ? n139 : n25241;
  assign n25250 = pi20 ? n139 : n25249;
  assign n25251 = pi19 ? n25250 : n32;
  assign n25252 = pi18 ? n139 : n25251;
  assign n25253 = pi17 ? n24715 : n25252;
  assign n25254 = pi16 ? n24712 : n25253;
  assign n25255 = pi20 ? n139 : n12396;
  assign n25256 = pi19 ? n25255 : n32;
  assign n25257 = pi18 ? n139 : n25256;
  assign n25258 = pi17 ? n24722 : n25257;
  assign n25259 = pi16 ? n439 : n25258;
  assign n25260 = pi15 ? n25254 : n25259;
  assign n25261 = pi14 ? n25248 : n25260;
  assign n25262 = pi13 ? n24696 : n25261;
  assign n25263 = pi17 ? n10653 : n25257;
  assign n25264 = pi16 ? n439 : n25263;
  assign n25265 = pi22 ? n6833 : n32;
  assign n25266 = pi21 ? n139 : n25265;
  assign n25267 = pi20 ? n139 : n25266;
  assign n25268 = pi19 ? n25267 : n32;
  assign n25269 = pi18 ? n24730 : n25268;
  assign n25270 = pi17 ? n11568 : n25269;
  assign n25271 = pi16 ? n439 : n25270;
  assign n25272 = pi15 ? n25264 : n25271;
  assign n25273 = pi18 ? n13193 : n25268;
  assign n25274 = pi17 ? n24736 : n25273;
  assign n25275 = pi16 ? n439 : n25274;
  assign n25276 = pi22 ? n3472 : n32;
  assign n25277 = pi21 ? n139 : n25276;
  assign n25278 = pi20 ? n139 : n25277;
  assign n25279 = pi19 ? n25278 : n32;
  assign n25280 = pi18 ? n14115 : n25279;
  assign n25281 = pi17 ? n37 : n25280;
  assign n25282 = pi16 ? n439 : n25281;
  assign n25283 = pi15 ? n25275 : n25282;
  assign n25284 = pi14 ? n25272 : n25283;
  assign n25285 = pi22 ? n13834 : n32;
  assign n25286 = pi21 ? n204 : n25285;
  assign n25287 = pi20 ? n204 : n25286;
  assign n25288 = pi19 ? n25287 : n32;
  assign n25289 = pi18 ? n24752 : n25288;
  assign n25290 = pi17 ? n37 : n25289;
  assign n25291 = pi16 ? n439 : n25290;
  assign n25292 = pi15 ? n24750 : n25291;
  assign n25293 = pi14 ? n25292 : n24768;
  assign n25294 = pi13 ? n25284 : n25293;
  assign n25295 = pi12 ? n25262 : n25294;
  assign n25296 = pi21 ? n233 : n3319;
  assign n25297 = pi20 ? n233 : n25296;
  assign n25298 = pi19 ? n25297 : n32;
  assign n25299 = pi18 ? n24774 : n25298;
  assign n25300 = pi17 ? n37 : n25299;
  assign n25301 = pi16 ? n439 : n25300;
  assign n25302 = pi21 ? n335 : n3339;
  assign n25303 = pi20 ? n335 : n25302;
  assign n25304 = pi19 ? n25303 : n32;
  assign n25305 = pi18 ? n17205 : n25304;
  assign n25306 = pi17 ? n37 : n25305;
  assign n25307 = pi16 ? n439 : n25306;
  assign n25308 = pi15 ? n25301 : n25307;
  assign n25309 = pi14 ? n25308 : n24798;
  assign n25310 = pi13 ? n25309 : n24815;
  assign n25311 = pi20 ? n2091 : n23203;
  assign n25312 = pi19 ? n25311 : n32;
  assign n25313 = pi18 ? n2102 : n25312;
  assign n25314 = pi17 ? n37 : n25313;
  assign n25315 = pi16 ? n439 : n25314;
  assign n25316 = pi15 ? n25315 : n24827;
  assign n25317 = pi20 ? n37 : n21211;
  assign n25318 = pi19 ? n25317 : n32;
  assign n25319 = pi18 ? n37 : n25318;
  assign n25320 = pi17 ? n37 : n25319;
  assign n25321 = pi16 ? n439 : n25320;
  assign n25322 = pi21 ? n24835 : n2700;
  assign n25323 = pi20 ? n37 : n25322;
  assign n25324 = pi19 ? n25323 : n32;
  assign n25325 = pi18 ? n37 : n25324;
  assign n25326 = pi17 ? n37 : n25325;
  assign n25327 = pi16 ? n439 : n25326;
  assign n25328 = pi15 ? n25321 : n25327;
  assign n25329 = pi14 ? n25316 : n25328;
  assign n25330 = pi21 ? n17764 : n32;
  assign n25331 = pi20 ? n37 : n25330;
  assign n25332 = pi19 ? n25331 : n32;
  assign n25333 = pi18 ? n37 : n25332;
  assign n25334 = pi17 ? n37 : n25333;
  assign n25335 = pi16 ? n439 : n25334;
  assign n25336 = pi21 ? n14255 : n32;
  assign n25337 = pi20 ? n363 : n25336;
  assign n25338 = pi19 ? n25337 : n32;
  assign n25339 = pi18 ? n24867 : n25338;
  assign n25340 = pi17 ? n37 : n25339;
  assign n25341 = pi16 ? n439 : n25340;
  assign n25342 = pi15 ? n25335 : n25341;
  assign n25343 = pi14 ? n24856 : n25342;
  assign n25344 = pi13 ? n25329 : n25343;
  assign n25345 = pi12 ? n25310 : n25344;
  assign n25346 = pi11 ? n25295 : n25345;
  assign n25347 = pi22 ? n363 : n2244;
  assign n25348 = pi21 ? n25347 : n32;
  assign n25349 = pi20 ? n7730 : n25348;
  assign n25350 = pi19 ? n25349 : n32;
  assign n25351 = pi18 ? n24881 : n25350;
  assign n25352 = pi17 ? n37 : n25351;
  assign n25353 = pi16 ? n439 : n25352;
  assign n25354 = pi20 ? n37 : n7332;
  assign n25355 = pi19 ? n25354 : n7322;
  assign n25356 = pi21 ? n6401 : n3392;
  assign n25357 = pi21 ? n20460 : n32;
  assign n25358 = pi20 ? n25356 : n25357;
  assign n25359 = pi19 ? n25358 : n32;
  assign n25360 = pi18 ? n25355 : n25359;
  assign n25361 = pi17 ? n37 : n25360;
  assign n25362 = pi16 ? n439 : n25361;
  assign n25363 = pi15 ? n25353 : n25362;
  assign n25364 = pi20 ? n37 : n12501;
  assign n25365 = pi19 ? n25364 : n32;
  assign n25366 = pi18 ? n37 : n25365;
  assign n25367 = pi17 ? n37 : n25366;
  assign n25368 = pi16 ? n439 : n25367;
  assign n25369 = pi20 ? n157 : n12501;
  assign n25370 = pi19 ? n25369 : n32;
  assign n25371 = pi18 ? n24903 : n25370;
  assign n25372 = pi17 ? n37 : n25371;
  assign n25373 = pi16 ? n439 : n25372;
  assign n25374 = pi15 ? n25368 : n25373;
  assign n25375 = pi14 ? n25363 : n25374;
  assign n25376 = pi20 ? n99 : n11674;
  assign n25377 = pi19 ? n25376 : n32;
  assign n25378 = pi18 ? n24914 : n25377;
  assign n25379 = pi17 ? n99 : n25378;
  assign n25380 = pi16 ? n744 : n25379;
  assign n25381 = pi20 ? n4617 : n99;
  assign n25382 = pi19 ? n99 : n25381;
  assign n25383 = pi21 ? n4193 : n32;
  assign n25384 = pi20 ? n99 : n25383;
  assign n25385 = pi19 ? n25384 : n32;
  assign n25386 = pi18 ? n25382 : n25385;
  assign n25387 = pi17 ? n99 : n25386;
  assign n25388 = pi16 ? n744 : n25387;
  assign n25389 = pi15 ? n25380 : n25388;
  assign n25390 = pi20 ? n99 : n13398;
  assign n25391 = pi19 ? n25390 : n32;
  assign n25392 = pi18 ? n99 : n25391;
  assign n25393 = pi17 ? n99 : n25392;
  assign n25394 = pi16 ? n744 : n25393;
  assign n25395 = pi16 ? n744 : n24933;
  assign n25396 = pi15 ? n25394 : n25395;
  assign n25397 = pi14 ? n25389 : n25396;
  assign n25398 = pi13 ? n25375 : n25397;
  assign n25399 = pi21 ? n5145 : n32;
  assign n25400 = pi20 ? n2238 : n25399;
  assign n25401 = pi19 ? n25400 : n32;
  assign n25402 = pi18 ? n99 : n25401;
  assign n25403 = pi17 ? n99 : n25402;
  assign n25404 = pi16 ? n744 : n25403;
  assign n25405 = pi22 ? n157 : n706;
  assign n25406 = pi21 ? n25405 : n32;
  assign n25407 = pi20 ? n2238 : n25406;
  assign n25408 = pi19 ? n25407 : n32;
  assign n25409 = pi18 ? n24944 : n25408;
  assign n25410 = pi17 ? n99 : n25409;
  assign n25411 = pi16 ? n744 : n25410;
  assign n25412 = pi15 ? n25404 : n25411;
  assign n25413 = pi21 ? n739 : n139;
  assign n25414 = pi20 ? n32 : n25413;
  assign n25415 = pi19 ? n32 : n25414;
  assign n25416 = pi18 ? n25415 : n139;
  assign n25417 = pi17 ? n32 : n25416;
  assign n25418 = pi16 ? n25417 : n24961;
  assign n25419 = pi16 ? n915 : n24967;
  assign n25420 = pi15 ? n25418 : n25419;
  assign n25421 = pi14 ? n25412 : n25420;
  assign n25422 = pi13 ? n25421 : n25004;
  assign n25423 = pi12 ? n25398 : n25422;
  assign n25424 = pi20 ? n14953 : n7042;
  assign n25425 = pi19 ? n25424 : n32;
  assign n25426 = pi18 ? n139 : n25425;
  assign n25427 = pi17 ? n139 : n25426;
  assign n25428 = pi16 ? n915 : n25427;
  assign n25429 = pi20 ? n25015 : n7049;
  assign n25430 = pi19 ? n25429 : n32;
  assign n25431 = pi18 ? n25013 : n25430;
  assign n25432 = pi17 ? n139 : n25431;
  assign n25433 = pi16 ? n915 : n25432;
  assign n25434 = pi15 ? n25428 : n25433;
  assign n25435 = pi20 ? n25023 : n5830;
  assign n25436 = pi19 ? n25435 : n32;
  assign n25437 = pi18 ? n25022 : n25436;
  assign n25438 = pi17 ? n139 : n25437;
  assign n25439 = pi16 ? n915 : n25438;
  assign n25440 = pi22 ? n909 : n566;
  assign n25441 = pi21 ? n25440 : n9122;
  assign n25442 = pi20 ? n32 : n25441;
  assign n25443 = pi19 ? n32 : n25442;
  assign n25444 = pi21 ? n580 : n9122;
  assign n25445 = pi20 ? n25444 : n3075;
  assign n25446 = pi21 ? n1531 : n567;
  assign n25447 = pi19 ? n25445 : n25446;
  assign n25448 = pi18 ? n25443 : n25447;
  assign n25449 = pi17 ? n32 : n25448;
  assign n25450 = pi21 ? n3073 : n569;
  assign n25451 = pi20 ? n25450 : n9118;
  assign n25452 = pi19 ? n25450 : n25451;
  assign n25453 = pi21 ? n37 : n9144;
  assign n25454 = pi20 ? n25044 : n25453;
  assign n25455 = pi21 ? n9122 : n3073;
  assign n25456 = pi20 ? n25455 : n9125;
  assign n25457 = pi19 ? n25454 : n25456;
  assign n25458 = pi18 ? n25452 : n25457;
  assign n25459 = pi21 ? n9563 : n567;
  assign n25460 = pi21 ? n9119 : n204;
  assign n25461 = pi20 ? n25459 : n25460;
  assign n25462 = pi19 ? n25461 : n204;
  assign n25463 = pi22 ? n204 : n21511;
  assign n25464 = pi21 ? n204 : n25463;
  assign n25465 = pi20 ? n25464 : n10011;
  assign n25466 = pi19 ? n25465 : n32;
  assign n25467 = pi18 ? n25462 : n25466;
  assign n25468 = pi17 ? n25458 : n25467;
  assign n25469 = pi16 ? n25449 : n25468;
  assign n25470 = pi15 ? n25439 : n25469;
  assign n25471 = pi14 ? n25434 : n25470;
  assign n25472 = pi18 ? n602 : n25066;
  assign n25473 = pi17 ? n32 : n25472;
  assign n25474 = pi21 ? n233 : n12983;
  assign n25475 = pi20 ? n25474 : n2653;
  assign n25476 = pi19 ? n25475 : n32;
  assign n25477 = pi18 ? n25071 : n25476;
  assign n25478 = pi17 ? n335 : n25477;
  assign n25479 = pi16 ? n25473 : n25478;
  assign n25480 = pi18 ? n602 : n25079;
  assign n25481 = pi17 ? n32 : n25480;
  assign n25482 = pi21 ? n233 : n12994;
  assign n25483 = pi20 ? n25482 : n1822;
  assign n25484 = pi19 ? n25483 : n32;
  assign n25485 = pi18 ? n25082 : n25484;
  assign n25486 = pi17 ? n335 : n25485;
  assign n25487 = pi16 ? n25481 : n25486;
  assign n25488 = pi15 ? n25479 : n25487;
  assign n25489 = pi21 ? n6376 : n12994;
  assign n25490 = pi20 ? n25489 : n32;
  assign n25491 = pi19 ? n25490 : n32;
  assign n25492 = pi18 ? n25093 : n25491;
  assign n25493 = pi17 ? n25092 : n25492;
  assign n25494 = pi16 ? n25090 : n25493;
  assign n25495 = pi15 ? n25494 : n25104;
  assign n25496 = pi14 ? n25488 : n25495;
  assign n25497 = pi13 ? n25471 : n25496;
  assign n25498 = pi21 ? n37 : n3404;
  assign n25499 = pi20 ? n25498 : n1921;
  assign n25500 = pi21 ? n25108 : n37;
  assign n25501 = pi20 ? n37 : n25500;
  assign n25502 = pi19 ? n25499 : n25501;
  assign n25503 = pi18 ? n7718 : n25502;
  assign n25504 = pi17 ? n25503 : n25121;
  assign n25505 = pi16 ? n25113 : n25504;
  assign n25506 = pi18 ? n25127 : n25120;
  assign n25507 = pi17 ? n25124 : n25506;
  assign n25508 = pi16 ? n439 : n25507;
  assign n25509 = pi15 ? n25505 : n25508;
  assign n25510 = pi18 ? n25135 : n25120;
  assign n25511 = pi17 ? n25124 : n25510;
  assign n25512 = pi16 ? n439 : n25511;
  assign n25513 = pi21 ? n335 : n19726;
  assign n25514 = pi20 ? n25513 : n32;
  assign n25515 = pi19 ? n25514 : n32;
  assign n25516 = pi18 ? n25154 : n25515;
  assign n25517 = pi17 ? n25152 : n25516;
  assign n25518 = pi16 ? n25143 : n25517;
  assign n25519 = pi15 ? n25512 : n25518;
  assign n25520 = pi14 ? n25509 : n25519;
  assign n25521 = pi18 ? n233 : n23546;
  assign n25522 = pi17 ? n25173 : n25521;
  assign n25523 = pi16 ? n25171 : n25522;
  assign n25524 = pi21 ? n5014 : n20848;
  assign n25525 = pi20 ? n25524 : n32;
  assign n25526 = pi19 ? n25525 : n32;
  assign n25527 = pi18 ? n21243 : n25526;
  assign n25528 = pi17 ? n25191 : n25527;
  assign n25529 = pi16 ? n25185 : n25528;
  assign n25530 = pi15 ? n25523 : n25529;
  assign n25531 = pi21 ? n363 : n2230;
  assign n25532 = pi20 ? n25531 : n32;
  assign n25533 = pi19 ? n25532 : n32;
  assign n25534 = pi18 ? n25201 : n25533;
  assign n25535 = pi17 ? n363 : n25534;
  assign n25536 = pi16 ? n21561 : n25535;
  assign n25537 = pi22 ? n2767 : n706;
  assign n25538 = pi21 ? n363 : n25537;
  assign n25539 = pi20 ? n25538 : n32;
  assign n25540 = pi19 ? n25539 : n32;
  assign n25541 = pi18 ? n25209 : n25540;
  assign n25542 = pi17 ? n363 : n25541;
  assign n25543 = pi16 ? n21561 : n25542;
  assign n25544 = pi15 ? n25536 : n25543;
  assign n25545 = pi14 ? n25530 : n25544;
  assign n25546 = pi13 ? n25520 : n25545;
  assign n25547 = pi12 ? n25497 : n25546;
  assign n25548 = pi11 ? n25423 : n25547;
  assign n25549 = pi10 ? n25346 : n25548;
  assign n25550 = pi09 ? n25234 : n25549;
  assign n25551 = pi08 ? n25222 : n25550;
  assign n25552 = pi19 ? n50 : n32;
  assign n25553 = pi18 ? n37 : n25552;
  assign n25554 = pi17 ? n37 : n25553;
  assign n25555 = pi16 ? n14445 : n25554;
  assign n25556 = pi15 ? n32 : n25555;
  assign n25557 = pi20 ? n37 : n11379;
  assign n25558 = pi19 ? n25557 : n32;
  assign n25559 = pi18 ? n37 : n25558;
  assign n25560 = pi17 ? n37 : n25559;
  assign n25561 = pi16 ? n14445 : n25560;
  assign n25562 = pi20 ? n2974 : n7346;
  assign n25563 = pi19 ? n25562 : n17013;
  assign n25564 = pi20 ? n4202 : n105;
  assign n25565 = pi19 ? n25564 : n32;
  assign n25566 = pi18 ? n25563 : n25565;
  assign n25567 = pi17 ? n37 : n25566;
  assign n25568 = pi16 ? n16595 : n25567;
  assign n25569 = pi15 ? n25561 : n25568;
  assign n25570 = pi14 ? n25556 : n25569;
  assign n25571 = pi13 ? n32 : n25570;
  assign n25572 = pi12 ? n32 : n25571;
  assign n25573 = pi11 ? n32 : n25572;
  assign n25574 = pi10 ? n32 : n25573;
  assign n25575 = pi21 ? n181 : n303;
  assign n25576 = pi20 ? n17960 : n25575;
  assign n25577 = pi19 ? n25576 : n32;
  assign n25578 = pi18 ? n37 : n25577;
  assign n25579 = pi17 ? n37 : n25578;
  assign n25580 = pi16 ? n16595 : n25579;
  assign n25581 = pi21 ? n181 : n588;
  assign n25582 = pi20 ? n37 : n25581;
  assign n25583 = pi19 ? n25582 : n32;
  assign n25584 = pi18 ? n37 : n25583;
  assign n25585 = pi17 ? n37 : n25584;
  assign n25586 = pi16 ? n17010 : n25585;
  assign n25587 = pi15 ? n25580 : n25586;
  assign n25588 = pi20 ? n37 : n11403;
  assign n25589 = pi19 ? n25588 : n32;
  assign n25590 = pi18 ? n37 : n25589;
  assign n25591 = pi17 ? n37 : n25590;
  assign n25592 = pi16 ? n17010 : n25591;
  assign n25593 = pi21 ? n37 : n11427;
  assign n25594 = pi20 ? n37 : n25593;
  assign n25595 = pi19 ? n25594 : n32;
  assign n25596 = pi18 ? n37 : n25595;
  assign n25597 = pi17 ? n37 : n25596;
  assign n25598 = pi16 ? n439 : n25597;
  assign n25599 = pi15 ? n25592 : n25598;
  assign n25600 = pi14 ? n25587 : n25599;
  assign n25601 = pi23 ? n99 : n11910;
  assign n25602 = pi22 ? n25601 : n32;
  assign n25603 = pi21 ? n99 : n25602;
  assign n25604 = pi20 ? n99 : n25603;
  assign n25605 = pi19 ? n25604 : n32;
  assign n25606 = pi18 ? n99 : n25605;
  assign n25607 = pi17 ? n99 : n25606;
  assign n25608 = pi16 ? n24698 : n25607;
  assign n25609 = pi18 ? n199 : n18854;
  assign n25610 = pi17 ? n32 : n25609;
  assign n25611 = pi20 ? n99 : n11459;
  assign n25612 = pi19 ? n25611 : n32;
  assign n25613 = pi18 ? n99 : n25612;
  assign n25614 = pi17 ? n99 : n25613;
  assign n25615 = pi16 ? n25610 : n25614;
  assign n25616 = pi15 ? n25608 : n25615;
  assign n25617 = pi19 ? n99 : n227;
  assign n25618 = pi18 ? n3031 : n25617;
  assign n25619 = pi17 ? n32 : n25618;
  assign n25620 = pi20 ? n219 : n14846;
  assign n25621 = pi19 ? n25620 : n139;
  assign n25622 = pi18 ? n25621 : n139;
  assign n25623 = pi21 ? n139 : n11458;
  assign n25624 = pi20 ? n139 : n25623;
  assign n25625 = pi19 ? n25624 : n32;
  assign n25626 = pi18 ? n139 : n25625;
  assign n25627 = pi17 ? n25622 : n25626;
  assign n25628 = pi16 ? n25619 : n25627;
  assign n25629 = pi23 ? n139 : n16890;
  assign n25630 = pi22 ? n25629 : n32;
  assign n25631 = pi21 ? n139 : n25630;
  assign n25632 = pi20 ? n139 : n25631;
  assign n25633 = pi19 ? n25632 : n32;
  assign n25634 = pi18 ? n139 : n25633;
  assign n25635 = pi17 ? n24722 : n25634;
  assign n25636 = pi16 ? n439 : n25635;
  assign n25637 = pi15 ? n25628 : n25636;
  assign n25638 = pi14 ? n25616 : n25637;
  assign n25639 = pi13 ? n25600 : n25638;
  assign n25640 = pi20 ? n997 : n992;
  assign n25641 = pi19 ? n37 : n25640;
  assign n25642 = pi20 ? n3104 : n942;
  assign n25643 = pi19 ? n25642 : n139;
  assign n25644 = pi18 ? n25641 : n25643;
  assign n25645 = pi17 ? n25644 : n25634;
  assign n25646 = pi16 ? n439 : n25645;
  assign n25647 = pi20 ? n941 : n3083;
  assign n25648 = pi19 ? n25647 : n139;
  assign n25649 = pi18 ? n25648 : n25633;
  assign n25650 = pi17 ? n11568 : n25649;
  assign n25651 = pi16 ? n439 : n25650;
  assign n25652 = pi15 ? n25646 : n25651;
  assign n25653 = pi23 ? n139 : n7393;
  assign n25654 = pi22 ? n25653 : n32;
  assign n25655 = pi21 ? n139 : n25654;
  assign n25656 = pi20 ? n139 : n25655;
  assign n25657 = pi19 ? n25656 : n32;
  assign n25658 = pi18 ? n13193 : n25657;
  assign n25659 = pi17 ? n24736 : n25658;
  assign n25660 = pi16 ? n439 : n25659;
  assign n25661 = pi18 ? n14115 : n25657;
  assign n25662 = pi17 ? n37 : n25661;
  assign n25663 = pi16 ? n439 : n25662;
  assign n25664 = pi15 ? n25660 : n25663;
  assign n25665 = pi14 ? n25652 : n25664;
  assign n25666 = pi23 ? n139 : n10729;
  assign n25667 = pi22 ? n25666 : n32;
  assign n25668 = pi21 ? n37 : n25667;
  assign n25669 = pi20 ? n1583 : n25668;
  assign n25670 = pi19 ? n25669 : n32;
  assign n25671 = pi18 ? n37 : n25670;
  assign n25672 = pi17 ? n37 : n25671;
  assign n25673 = pi16 ? n439 : n25672;
  assign n25674 = pi21 ? n204 : n12404;
  assign n25675 = pi20 ? n204 : n25674;
  assign n25676 = pi19 ? n25675 : n32;
  assign n25677 = pi18 ? n23802 : n25676;
  assign n25678 = pi17 ? n37 : n25677;
  assign n25679 = pi16 ? n439 : n25678;
  assign n25680 = pi15 ? n25673 : n25679;
  assign n25681 = pi19 ? n37 : n18984;
  assign n25682 = pi18 ? n25681 : n25676;
  assign n25683 = pi17 ? n37 : n25682;
  assign n25684 = pi16 ? n439 : n25683;
  assign n25685 = pi21 ? n204 : n7034;
  assign n25686 = pi20 ? n204 : n25685;
  assign n25687 = pi19 ? n25686 : n32;
  assign n25688 = pi18 ? n25681 : n25687;
  assign n25689 = pi17 ? n37 : n25688;
  assign n25690 = pi16 ? n439 : n25689;
  assign n25691 = pi15 ? n25684 : n25690;
  assign n25692 = pi14 ? n25680 : n25691;
  assign n25693 = pi13 ? n25665 : n25692;
  assign n25694 = pi12 ? n25639 : n25693;
  assign n25695 = pi20 ? n233 : n13743;
  assign n25696 = pi19 ? n25695 : n32;
  assign n25697 = pi18 ? n7707 : n25696;
  assign n25698 = pi17 ? n37 : n25697;
  assign n25699 = pi16 ? n439 : n25698;
  assign n25700 = pi21 ? n335 : n4109;
  assign n25701 = pi20 ? n335 : n25700;
  assign n25702 = pi19 ? n25701 : n32;
  assign n25703 = pi18 ? n24789 : n25702;
  assign n25704 = pi17 ? n37 : n25703;
  assign n25705 = pi16 ? n439 : n25704;
  assign n25706 = pi15 ? n25699 : n25705;
  assign n25707 = pi20 ? n569 : n25700;
  assign n25708 = pi19 ? n25707 : n32;
  assign n25709 = pi18 ? n7686 : n25708;
  assign n25710 = pi17 ? n37 : n25709;
  assign n25711 = pi16 ? n439 : n25710;
  assign n25712 = pi15 ? n25705 : n25711;
  assign n25713 = pi14 ? n25706 : n25712;
  assign n25714 = pi18 ? n37 : n25708;
  assign n25715 = pi17 ? n37 : n25714;
  assign n25716 = pi16 ? n439 : n25715;
  assign n25717 = pi20 ? n649 : n25700;
  assign n25718 = pi19 ? n25717 : n32;
  assign n25719 = pi18 ? n37 : n25718;
  assign n25720 = pi17 ? n37 : n25719;
  assign n25721 = pi16 ? n439 : n25720;
  assign n25722 = pi15 ? n25716 : n25721;
  assign n25723 = pi20 ? n37 : n25700;
  assign n25724 = pi19 ? n25723 : n32;
  assign n25725 = pi18 ? n37 : n25724;
  assign n25726 = pi17 ? n37 : n25725;
  assign n25727 = pi16 ? n439 : n25726;
  assign n25728 = pi20 ? n37 : n11602;
  assign n25729 = pi19 ? n25728 : n32;
  assign n25730 = pi18 ? n37 : n25729;
  assign n25731 = pi17 ? n37 : n25730;
  assign n25732 = pi16 ? n439 : n25731;
  assign n25733 = pi15 ? n25727 : n25732;
  assign n25734 = pi14 ? n25722 : n25733;
  assign n25735 = pi13 ? n25713 : n25734;
  assign n25736 = pi20 ? n2094 : n21182;
  assign n25737 = pi19 ? n25736 : n32;
  assign n25738 = pi18 ? n37 : n25737;
  assign n25739 = pi17 ? n37 : n25738;
  assign n25740 = pi16 ? n439 : n25739;
  assign n25741 = pi20 ? n37 : n13322;
  assign n25742 = pi19 ? n25741 : n32;
  assign n25743 = pi18 ? n37 : n25742;
  assign n25744 = pi17 ? n37 : n25743;
  assign n25745 = pi16 ? n439 : n25744;
  assign n25746 = pi15 ? n25740 : n25745;
  assign n25747 = pi21 ? n2106 : n5829;
  assign n25748 = pi20 ? n37 : n25747;
  assign n25749 = pi19 ? n25748 : n32;
  assign n25750 = pi18 ? n37 : n25749;
  assign n25751 = pi17 ? n37 : n25750;
  assign n25752 = pi16 ? n439 : n25751;
  assign n25753 = pi20 ? n37 : n12872;
  assign n25754 = pi19 ? n25753 : n32;
  assign n25755 = pi18 ? n37 : n25754;
  assign n25756 = pi17 ? n37 : n25755;
  assign n25757 = pi16 ? n439 : n25756;
  assign n25758 = pi15 ? n25752 : n25757;
  assign n25759 = pi14 ? n25746 : n25758;
  assign n25760 = pi21 ? n3392 : n928;
  assign n25761 = pi20 ? n37 : n25760;
  assign n25762 = pi19 ? n25761 : n32;
  assign n25763 = pi18 ? n37 : n25762;
  assign n25764 = pi17 ? n37 : n25763;
  assign n25765 = pi16 ? n439 : n25764;
  assign n25766 = pi21 ? n3392 : n1009;
  assign n25767 = pi20 ? n37 : n25766;
  assign n25768 = pi19 ? n25767 : n32;
  assign n25769 = pi18 ? n37 : n25768;
  assign n25770 = pi17 ? n37 : n25769;
  assign n25771 = pi16 ? n439 : n25770;
  assign n25772 = pi15 ? n25765 : n25771;
  assign n25773 = pi23 ? n1432 : n157;
  assign n25774 = pi22 ? n37 : n25773;
  assign n25775 = pi21 ? n25774 : n32;
  assign n25776 = pi20 ? n37 : n25775;
  assign n25777 = pi19 ? n25776 : n32;
  assign n25778 = pi18 ? n37 : n25777;
  assign n25779 = pi17 ? n37 : n25778;
  assign n25780 = pi16 ? n439 : n25779;
  assign n25781 = pi19 ? n5029 : n363;
  assign n25782 = pi21 ? n5054 : n32;
  assign n25783 = pi20 ? n363 : n25782;
  assign n25784 = pi19 ? n25783 : n32;
  assign n25785 = pi18 ? n25781 : n25784;
  assign n25786 = pi17 ? n37 : n25785;
  assign n25787 = pi16 ? n439 : n25786;
  assign n25788 = pi15 ? n25780 : n25787;
  assign n25789 = pi14 ? n25772 : n25788;
  assign n25790 = pi13 ? n25759 : n25789;
  assign n25791 = pi12 ? n25735 : n25790;
  assign n25792 = pi11 ? n25694 : n25791;
  assign n25793 = pi20 ? n7730 : n11665;
  assign n25794 = pi19 ? n25793 : n32;
  assign n25795 = pi18 ? n24881 : n25794;
  assign n25796 = pi17 ? n37 : n25795;
  assign n25797 = pi16 ? n439 : n25796;
  assign n25798 = pi20 ? n37 : n11665;
  assign n25799 = pi19 ? n25798 : n32;
  assign n25800 = pi18 ? n37 : n25799;
  assign n25801 = pi17 ? n37 : n25800;
  assign n25802 = pi16 ? n439 : n25801;
  assign n25803 = pi15 ? n25797 : n25802;
  assign n25804 = pi21 ? n37 : n157;
  assign n25805 = pi20 ? n37 : n25804;
  assign n25806 = pi19 ? n25805 : n157;
  assign n25807 = pi18 ? n25806 : n25370;
  assign n25808 = pi17 ? n37 : n25807;
  assign n25809 = pi16 ? n439 : n25808;
  assign n25810 = pi15 ? n25802 : n25809;
  assign n25811 = pi14 ? n25803 : n25810;
  assign n25812 = pi16 ? n721 : n25379;
  assign n25813 = pi22 ? n745 : n316;
  assign n25814 = pi21 ? n25813 : n32;
  assign n25815 = pi20 ? n99 : n25814;
  assign n25816 = pi19 ? n25815 : n32;
  assign n25817 = pi18 ? n99 : n25816;
  assign n25818 = pi17 ? n99 : n25817;
  assign n25819 = pi16 ? n721 : n25818;
  assign n25820 = pi15 ? n25812 : n25819;
  assign n25821 = pi16 ? n721 : n25393;
  assign n25822 = pi21 ? n6535 : n32;
  assign n25823 = pi20 ? n99 : n25822;
  assign n25824 = pi19 ? n25823 : n32;
  assign n25825 = pi18 ? n99 : n25824;
  assign n25826 = pi17 ? n99 : n25825;
  assign n25827 = pi16 ? n721 : n25826;
  assign n25828 = pi15 ? n25821 : n25827;
  assign n25829 = pi14 ? n25820 : n25828;
  assign n25830 = pi13 ? n25811 : n25829;
  assign n25831 = pi20 ? n776 : n25406;
  assign n25832 = pi19 ? n25831 : n32;
  assign n25833 = pi18 ? n24944 : n25832;
  assign n25834 = pi17 ? n99 : n25833;
  assign n25835 = pi16 ? n721 : n25834;
  assign n25836 = pi15 ? n23968 : n25835;
  assign n25837 = pi20 ? n24957 : n14352;
  assign n25838 = pi19 ? n25837 : n32;
  assign n25839 = pi18 ? n24956 : n25838;
  assign n25840 = pi17 ? n139 : n25839;
  assign n25841 = pi16 ? n24953 : n25840;
  assign n25842 = pi20 ? n18317 : n4008;
  assign n25843 = pi19 ? n25842 : n32;
  assign n25844 = pi18 ? n24963 : n25843;
  assign n25845 = pi17 ? n139 : n25844;
  assign n25846 = pi16 ? n331 : n25845;
  assign n25847 = pi15 ? n25841 : n25846;
  assign n25848 = pi14 ? n25836 : n25847;
  assign n25849 = pi19 ? n204 : n15422;
  assign n25850 = pi21 ? n4056 : n204;
  assign n25851 = pi20 ? n25850 : n37;
  assign n25852 = pi19 ? n25851 : n204;
  assign n25853 = pi18 ? n25849 : n25852;
  assign n25854 = pi20 ? n316 : n4008;
  assign n25855 = pi19 ? n25854 : n32;
  assign n25856 = pi18 ? n24977 : n25855;
  assign n25857 = pi17 ? n25853 : n25856;
  assign n25858 = pi16 ? n11804 : n25857;
  assign n25859 = pi18 ? n24995 : n25855;
  assign n25860 = pi17 ? n204 : n25859;
  assign n25861 = pi16 ? n13493 : n25860;
  assign n25862 = pi15 ? n25858 : n25861;
  assign n25863 = pi20 ? n204 : n1583;
  assign n25864 = pi19 ? n25863 : n204;
  assign n25865 = pi18 ? n204 : n25864;
  assign n25866 = pi17 ? n25865 : n25859;
  assign n25867 = pi16 ? n13846 : n25866;
  assign n25868 = pi21 ? n139 : n4780;
  assign n25869 = pi21 ? n204 : n19311;
  assign n25870 = pi20 ? n25868 : n25869;
  assign n25871 = pi19 ? n15405 : n25870;
  assign n25872 = pi20 ? n1026 : n20391;
  assign n25873 = pi19 ? n25872 : n32;
  assign n25874 = pi18 ? n25871 : n25873;
  assign n25875 = pi17 ? n25865 : n25874;
  assign n25876 = pi16 ? n13846 : n25875;
  assign n25877 = pi15 ? n25867 : n25876;
  assign n25878 = pi14 ? n25862 : n25877;
  assign n25879 = pi13 ? n25848 : n25878;
  assign n25880 = pi12 ? n25830 : n25879;
  assign n25881 = pi20 ? n1026 : n7042;
  assign n25882 = pi19 ? n25881 : n32;
  assign n25883 = pi18 ? n139 : n25882;
  assign n25884 = pi17 ? n139 : n25883;
  assign n25885 = pi16 ? n915 : n25884;
  assign n25886 = pi20 ? n2316 : n6577;
  assign n25887 = pi19 ? n139 : n25886;
  assign n25888 = pi20 ? n6577 : n7049;
  assign n25889 = pi19 ? n25888 : n32;
  assign n25890 = pi18 ? n25887 : n25889;
  assign n25891 = pi17 ? n139 : n25890;
  assign n25892 = pi16 ? n915 : n25891;
  assign n25893 = pi15 ? n25885 : n25892;
  assign n25894 = pi20 ? n1016 : n922;
  assign n25895 = pi19 ? n139 : n25894;
  assign n25896 = pi20 ? n1026 : n5830;
  assign n25897 = pi19 ? n25896 : n32;
  assign n25898 = pi18 ? n25895 : n25897;
  assign n25899 = pi17 ? n139 : n25898;
  assign n25900 = pi16 ? n915 : n25899;
  assign n25901 = pi19 ? n3285 : n649;
  assign n25902 = pi18 ? n9556 : n25901;
  assign n25903 = pi17 ? n32 : n25902;
  assign n25904 = pi19 ? n605 : n4984;
  assign n25905 = pi20 ? n335 : n3335;
  assign n25906 = pi19 ? n25905 : n611;
  assign n25907 = pi18 ? n25904 : n25906;
  assign n25908 = pi19 ? n1090 : n204;
  assign n25909 = pi20 ? n204 : n2653;
  assign n25910 = pi19 ? n25909 : n32;
  assign n25911 = pi18 ? n25908 : n25910;
  assign n25912 = pi17 ? n25907 : n25911;
  assign n25913 = pi16 ? n25903 : n25912;
  assign n25914 = pi15 ? n25900 : n25913;
  assign n25915 = pi14 ? n25893 : n25914;
  assign n25916 = pi19 ? n335 : n233;
  assign n25917 = pi20 ? n233 : n1822;
  assign n25918 = pi19 ? n25917 : n32;
  assign n25919 = pi18 ? n25916 : n25918;
  assign n25920 = pi17 ? n335 : n25919;
  assign n25921 = pi16 ? n7943 : n25920;
  assign n25922 = pi18 ? n7941 : n3352;
  assign n25923 = pi17 ? n32 : n25922;
  assign n25924 = pi20 ? n233 : n32;
  assign n25925 = pi19 ? n25924 : n32;
  assign n25926 = pi18 ? n25082 : n25925;
  assign n25927 = pi17 ? n335 : n25926;
  assign n25928 = pi16 ? n25923 : n25927;
  assign n25929 = pi15 ? n25921 : n25928;
  assign n25930 = pi20 ? n16544 : n32;
  assign n25931 = pi19 ? n25930 : n32;
  assign n25932 = pi18 ? n25093 : n25931;
  assign n25933 = pi17 ? n25092 : n25932;
  assign n25934 = pi16 ? n25090 : n25933;
  assign n25935 = pi19 ? n10681 : n233;
  assign n25936 = pi18 ? n25935 : n25925;
  assign n25937 = pi17 ? n37 : n25936;
  assign n25938 = pi16 ? n439 : n25937;
  assign n25939 = pi15 ? n25934 : n25938;
  assign n25940 = pi14 ? n25929 : n25939;
  assign n25941 = pi13 ? n25915 : n25940;
  assign n25942 = pi23 ? n38 : n233;
  assign n25943 = pi22 ? n25942 : n335;
  assign n25944 = pi21 ? n25943 : n233;
  assign n25945 = pi20 ? n32 : n25944;
  assign n25946 = pi19 ? n32 : n25945;
  assign n25947 = pi21 ? n569 : n233;
  assign n25948 = pi20 ? n25947 : n37;
  assign n25949 = pi20 ? n21148 : n21150;
  assign n25950 = pi19 ? n25948 : n25949;
  assign n25951 = pi18 ? n25946 : n25950;
  assign n25952 = pi17 ? n32 : n25951;
  assign n25953 = pi21 ? n6376 : n2048;
  assign n25954 = pi20 ? n14223 : n25953;
  assign n25955 = pi20 ? n25953 : n16530;
  assign n25956 = pi19 ? n25954 : n25955;
  assign n25957 = pi21 ? n233 : n569;
  assign n25958 = pi20 ? n18431 : n25957;
  assign n25959 = pi21 ? n19386 : n2048;
  assign n25960 = pi20 ? n25959 : n13527;
  assign n25961 = pi19 ? n25958 : n25960;
  assign n25962 = pi18 ? n25956 : n25961;
  assign n25963 = pi20 ? n6362 : n233;
  assign n25964 = pi19 ? n25963 : n233;
  assign n25965 = pi21 ? n233 : n18411;
  assign n25966 = pi20 ? n25965 : n32;
  assign n25967 = pi19 ? n25966 : n32;
  assign n25968 = pi18 ? n25964 : n25967;
  assign n25969 = pi17 ? n25962 : n25968;
  assign n25970 = pi16 ? n25952 : n25969;
  assign n25971 = pi19 ? n21125 : n37;
  assign n25972 = pi18 ? n37 : n25971;
  assign n25973 = pi18 ? n25135 : n25967;
  assign n25974 = pi17 ? n25972 : n25973;
  assign n25975 = pi16 ? n439 : n25974;
  assign n25976 = pi15 ? n25970 : n25975;
  assign n25977 = pi22 ? n233 : n316;
  assign n25978 = pi21 ? n233 : n25977;
  assign n25979 = pi20 ? n25978 : n32;
  assign n25980 = pi19 ? n25979 : n32;
  assign n25981 = pi18 ? n25135 : n25980;
  assign n25982 = pi17 ? n25972 : n25981;
  assign n25983 = pi16 ? n439 : n25982;
  assign n25984 = pi22 ? n25942 : n37;
  assign n25985 = pi21 ? n25984 : n584;
  assign n25986 = pi20 ? n32 : n25985;
  assign n25987 = pi19 ? n32 : n25986;
  assign n25988 = pi21 ? n2007 : n233;
  assign n25989 = pi20 ? n3292 : n25988;
  assign n25990 = pi19 ? n37 : n25989;
  assign n25991 = pi18 ? n25987 : n25990;
  assign n25992 = pi17 ? n32 : n25991;
  assign n25993 = pi21 ? n2048 : n574;
  assign n25994 = pi20 ? n25993 : n9912;
  assign n25995 = pi20 ? n9912 : n233;
  assign n25996 = pi19 ? n25994 : n25995;
  assign n25997 = pi21 ? n584 : n233;
  assign n25998 = pi20 ? n5023 : n25997;
  assign n25999 = pi20 ? n25957 : n7705;
  assign n26000 = pi19 ? n25998 : n25999;
  assign n26001 = pi18 ? n25996 : n26000;
  assign n26002 = pi21 ? n233 : n4912;
  assign n26003 = pi20 ? n18431 : n26002;
  assign n26004 = pi19 ? n233 : n26003;
  assign n26005 = pi21 ? n6361 : n19726;
  assign n26006 = pi20 ? n26005 : n32;
  assign n26007 = pi19 ? n26006 : n32;
  assign n26008 = pi18 ? n26004 : n26007;
  assign n26009 = pi17 ? n26001 : n26008;
  assign n26010 = pi16 ? n25992 : n26009;
  assign n26011 = pi15 ? n25983 : n26010;
  assign n26012 = pi14 ? n25976 : n26011;
  assign n26013 = pi22 ? n8501 : n233;
  assign n26014 = pi21 ? n26013 : n233;
  assign n26015 = pi20 ? n32 : n26014;
  assign n26016 = pi19 ? n32 : n26015;
  assign n26017 = pi20 ? n233 : n25167;
  assign n26018 = pi19 ? n26017 : n19423;
  assign n26019 = pi18 ? n26016 : n26018;
  assign n26020 = pi17 ? n32 : n26019;
  assign n26021 = pi21 ? n233 : n10981;
  assign n26022 = pi20 ? n26021 : n32;
  assign n26023 = pi19 ? n26022 : n32;
  assign n26024 = pi18 ? n233 : n26023;
  assign n26025 = pi17 ? n25173 : n26024;
  assign n26026 = pi16 ? n26020 : n26025;
  assign n26027 = pi23 ? n714 : n363;
  assign n26028 = pi22 ? n26027 : n99;
  assign n26029 = pi21 ? n26028 : n363;
  assign n26030 = pi20 ? n32 : n26029;
  assign n26031 = pi19 ? n32 : n26030;
  assign n26032 = pi18 ? n26031 : n25183;
  assign n26033 = pi17 ? n32 : n26032;
  assign n26034 = pi20 ? n23175 : n363;
  assign n26035 = pi19 ? n26034 : n25186;
  assign n26036 = pi20 ? n233 : n23155;
  assign n26037 = pi20 ? n21222 : n233;
  assign n26038 = pi19 ? n26036 : n26037;
  assign n26039 = pi18 ? n26035 : n26038;
  assign n26040 = pi21 ? n233 : n23157;
  assign n26041 = pi20 ? n233 : n26040;
  assign n26042 = pi19 ? n233 : n26041;
  assign n26043 = pi21 ? n363 : n15889;
  assign n26044 = pi20 ? n26043 : n32;
  assign n26045 = pi19 ? n26044 : n32;
  assign n26046 = pi18 ? n26042 : n26045;
  assign n26047 = pi17 ? n26039 : n26046;
  assign n26048 = pi16 ? n26033 : n26047;
  assign n26049 = pi15 ? n26026 : n26048;
  assign n26050 = pi21 ? n363 : n8486;
  assign n26051 = pi20 ? n26050 : n32;
  assign n26052 = pi19 ? n26051 : n32;
  assign n26053 = pi18 ? n25209 : n26052;
  assign n26054 = pi17 ? n363 : n26053;
  assign n26055 = pi16 ? n21219 : n26054;
  assign n26056 = pi23 ? n1590 : n363;
  assign n26057 = pi22 ? n26056 : n363;
  assign n26058 = pi21 ? n26057 : n363;
  assign n26059 = pi20 ? n32 : n26058;
  assign n26060 = pi19 ? n32 : n26059;
  assign n26061 = pi18 ? n26060 : n363;
  assign n26062 = pi17 ? n32 : n26061;
  assign n26063 = pi16 ? n26062 : n25214;
  assign n26064 = pi15 ? n26055 : n26063;
  assign n26065 = pi14 ? n26049 : n26064;
  assign n26066 = pi13 ? n26012 : n26065;
  assign n26067 = pi12 ? n25941 : n26066;
  assign n26068 = pi11 ? n25880 : n26067;
  assign n26069 = pi10 ? n25792 : n26068;
  assign n26070 = pi09 ? n25574 : n26069;
  assign n26071 = pi21 ? n37 : n5423;
  assign n26072 = pi20 ? n37 : n26071;
  assign n26073 = pi19 ? n26072 : n32;
  assign n26074 = pi18 ? n37 : n26073;
  assign n26075 = pi17 ? n37 : n26074;
  assign n26076 = pi16 ? n14445 : n26075;
  assign n26077 = pi15 ? n26076 : n25568;
  assign n26078 = pi14 ? n25556 : n26077;
  assign n26079 = pi13 ? n32 : n26078;
  assign n26080 = pi12 ? n32 : n26079;
  assign n26081 = pi11 ? n32 : n26080;
  assign n26082 = pi10 ? n32 : n26081;
  assign n26083 = pi20 ? n37 : n11891;
  assign n26084 = pi19 ? n26083 : n32;
  assign n26085 = pi18 ? n37 : n26084;
  assign n26086 = pi17 ? n37 : n26085;
  assign n26087 = pi16 ? n17010 : n26086;
  assign n26088 = pi16 ? n439 : n26086;
  assign n26089 = pi15 ? n26087 : n26088;
  assign n26090 = pi14 ? n25587 : n26089;
  assign n26091 = pi20 ? n99 : n11939;
  assign n26092 = pi19 ? n26091 : n32;
  assign n26093 = pi18 ? n99 : n26092;
  assign n26094 = pi17 ? n99 : n26093;
  assign n26095 = pi16 ? n24698 : n26094;
  assign n26096 = pi16 ? n25610 : n26094;
  assign n26097 = pi15 ? n26095 : n26096;
  assign n26098 = pi21 ? n139 : n11945;
  assign n26099 = pi20 ? n139 : n26098;
  assign n26100 = pi19 ? n26099 : n32;
  assign n26101 = pi18 ? n139 : n26100;
  assign n26102 = pi17 ? n25622 : n26101;
  assign n26103 = pi16 ? n25619 : n26102;
  assign n26104 = pi20 ? n139 : n13184;
  assign n26105 = pi19 ? n26104 : n32;
  assign n26106 = pi18 ? n139 : n26105;
  assign n26107 = pi17 ? n24722 : n26106;
  assign n26108 = pi16 ? n439 : n26107;
  assign n26109 = pi15 ? n26103 : n26108;
  assign n26110 = pi14 ? n26097 : n26109;
  assign n26111 = pi13 ? n26090 : n26110;
  assign n26112 = pi17 ? n25644 : n26106;
  assign n26113 = pi16 ? n439 : n26112;
  assign n26114 = pi18 ? n25648 : n26105;
  assign n26115 = pi17 ? n11568 : n26114;
  assign n26116 = pi16 ? n439 : n26115;
  assign n26117 = pi15 ? n26113 : n26116;
  assign n26118 = pi21 ? n139 : n18905;
  assign n26119 = pi20 ? n139 : n26118;
  assign n26120 = pi19 ? n26119 : n32;
  assign n26121 = pi18 ? n13193 : n26120;
  assign n26122 = pi17 ? n24736 : n26121;
  assign n26123 = pi16 ? n439 : n26122;
  assign n26124 = pi18 ? n14115 : n26120;
  assign n26125 = pi17 ? n37 : n26124;
  assign n26126 = pi16 ? n439 : n26125;
  assign n26127 = pi15 ? n26123 : n26126;
  assign n26128 = pi14 ? n26117 : n26127;
  assign n26129 = pi22 ? n9827 : n688;
  assign n26130 = pi21 ? n37 : n26129;
  assign n26131 = pi20 ? n1583 : n26130;
  assign n26132 = pi19 ? n26131 : n32;
  assign n26133 = pi18 ? n37 : n26132;
  assign n26134 = pi17 ? n37 : n26133;
  assign n26135 = pi16 ? n439 : n26134;
  assign n26136 = pi21 ? n204 : n14351;
  assign n26137 = pi20 ? n204 : n26136;
  assign n26138 = pi19 ? n26137 : n32;
  assign n26139 = pi18 ? n23802 : n26138;
  assign n26140 = pi17 ? n37 : n26139;
  assign n26141 = pi16 ? n439 : n26140;
  assign n26142 = pi15 ? n26135 : n26141;
  assign n26143 = pi18 ? n25681 : n26138;
  assign n26144 = pi17 ? n37 : n26143;
  assign n26145 = pi16 ? n439 : n26144;
  assign n26146 = pi15 ? n26145 : n25690;
  assign n26147 = pi14 ? n26142 : n26146;
  assign n26148 = pi13 ? n26128 : n26147;
  assign n26149 = pi12 ? n26111 : n26148;
  assign n26150 = pi21 ? n233 : n13722;
  assign n26151 = pi20 ? n233 : n26150;
  assign n26152 = pi19 ? n26151 : n32;
  assign n26153 = pi18 ? n7707 : n26152;
  assign n26154 = pi17 ? n37 : n26153;
  assign n26155 = pi16 ? n439 : n26154;
  assign n26156 = pi21 ? n335 : n12825;
  assign n26157 = pi20 ? n335 : n26156;
  assign n26158 = pi19 ? n26157 : n32;
  assign n26159 = pi18 ? n24789 : n26158;
  assign n26160 = pi17 ? n37 : n26159;
  assign n26161 = pi16 ? n439 : n26160;
  assign n26162 = pi15 ? n26155 : n26161;
  assign n26163 = pi22 ? n10768 : n32;
  assign n26164 = pi21 ? n335 : n26163;
  assign n26165 = pi20 ? n569 : n26164;
  assign n26166 = pi19 ? n26165 : n32;
  assign n26167 = pi18 ? n7686 : n26166;
  assign n26168 = pi17 ? n37 : n26167;
  assign n26169 = pi16 ? n439 : n26168;
  assign n26170 = pi15 ? n25705 : n26169;
  assign n26171 = pi14 ? n26162 : n26170;
  assign n26172 = pi21 ? n335 : n5813;
  assign n26173 = pi20 ? n569 : n26172;
  assign n26174 = pi19 ? n26173 : n32;
  assign n26175 = pi18 ? n37 : n26174;
  assign n26176 = pi17 ? n37 : n26175;
  assign n26177 = pi16 ? n439 : n26176;
  assign n26178 = pi20 ? n649 : n26172;
  assign n26179 = pi19 ? n26178 : n32;
  assign n26180 = pi18 ? n37 : n26179;
  assign n26181 = pi17 ? n37 : n26180;
  assign n26182 = pi16 ? n439 : n26181;
  assign n26183 = pi15 ? n26177 : n26182;
  assign n26184 = pi14 ? n26183 : n25733;
  assign n26185 = pi13 ? n26171 : n26184;
  assign n26186 = pi20 ? n37 : n12856;
  assign n26187 = pi19 ? n26186 : n32;
  assign n26188 = pi18 ? n37 : n26187;
  assign n26189 = pi17 ? n37 : n26188;
  assign n26190 = pi16 ? n439 : n26189;
  assign n26191 = pi15 ? n25740 : n26190;
  assign n26192 = pi14 ? n26191 : n25758;
  assign n26193 = pi21 ? n3392 : n2700;
  assign n26194 = pi20 ? n37 : n26193;
  assign n26195 = pi19 ? n26194 : n32;
  assign n26196 = pi18 ? n37 : n26195;
  assign n26197 = pi17 ? n37 : n26196;
  assign n26198 = pi16 ? n439 : n26197;
  assign n26199 = pi15 ? n25765 : n26198;
  assign n26200 = pi22 ? n37 : n3944;
  assign n26201 = pi21 ? n26200 : n2700;
  assign n26202 = pi20 ? n37 : n26201;
  assign n26203 = pi19 ? n26202 : n32;
  assign n26204 = pi18 ? n37 : n26203;
  assign n26205 = pi17 ? n37 : n26204;
  assign n26206 = pi16 ? n439 : n26205;
  assign n26207 = pi21 ? n5054 : n2700;
  assign n26208 = pi20 ? n363 : n26207;
  assign n26209 = pi19 ? n26208 : n32;
  assign n26210 = pi18 ? n25781 : n26209;
  assign n26211 = pi17 ? n37 : n26210;
  assign n26212 = pi16 ? n439 : n26211;
  assign n26213 = pi15 ? n26206 : n26212;
  assign n26214 = pi14 ? n26199 : n26213;
  assign n26215 = pi13 ? n26192 : n26214;
  assign n26216 = pi12 ? n26185 : n26215;
  assign n26217 = pi11 ? n26149 : n26216;
  assign n26218 = pi20 ? n7730 : n12095;
  assign n26219 = pi19 ? n26218 : n32;
  assign n26220 = pi18 ? n24881 : n26219;
  assign n26221 = pi17 ? n37 : n26220;
  assign n26222 = pi16 ? n439 : n26221;
  assign n26223 = pi20 ? n37 : n12095;
  assign n26224 = pi19 ? n26223 : n32;
  assign n26225 = pi18 ? n37 : n26224;
  assign n26226 = pi17 ? n37 : n26225;
  assign n26227 = pi16 ? n439 : n26226;
  assign n26228 = pi15 ? n26222 : n26227;
  assign n26229 = pi20 ? n157 : n12909;
  assign n26230 = pi19 ? n26229 : n32;
  assign n26231 = pi18 ? n25806 : n26230;
  assign n26232 = pi17 ? n37 : n26231;
  assign n26233 = pi16 ? n439 : n26232;
  assign n26234 = pi15 ? n26227 : n26233;
  assign n26235 = pi14 ? n26228 : n26234;
  assign n26236 = pi20 ? n99 : n7407;
  assign n26237 = pi19 ? n26236 : n32;
  assign n26238 = pi18 ? n24914 : n26237;
  assign n26239 = pi17 ? n99 : n26238;
  assign n26240 = pi16 ? n744 : n26239;
  assign n26241 = pi22 ? n745 : n22383;
  assign n26242 = pi21 ? n26241 : n1009;
  assign n26243 = pi20 ? n99 : n26242;
  assign n26244 = pi19 ? n26243 : n32;
  assign n26245 = pi18 ? n99 : n26244;
  assign n26246 = pi17 ? n99 : n26245;
  assign n26247 = pi16 ? n744 : n26246;
  assign n26248 = pi15 ? n26240 : n26247;
  assign n26249 = pi22 ? n316 : n22383;
  assign n26250 = pi21 ? n26249 : n1009;
  assign n26251 = pi20 ? n99 : n26250;
  assign n26252 = pi19 ? n26251 : n32;
  assign n26253 = pi18 ? n99 : n26252;
  assign n26254 = pi17 ? n99 : n26253;
  assign n26255 = pi16 ? n744 : n26254;
  assign n26256 = pi22 ? n157 : n22383;
  assign n26257 = pi21 ? n26256 : n32;
  assign n26258 = pi20 ? n99 : n26257;
  assign n26259 = pi19 ? n26258 : n32;
  assign n26260 = pi18 ? n99 : n26259;
  assign n26261 = pi17 ? n99 : n26260;
  assign n26262 = pi16 ? n744 : n26261;
  assign n26263 = pi15 ? n26255 : n26262;
  assign n26264 = pi14 ? n26248 : n26263;
  assign n26265 = pi13 ? n26235 : n26264;
  assign n26266 = pi20 ? n776 : n25399;
  assign n26267 = pi19 ? n26266 : n32;
  assign n26268 = pi18 ? n24944 : n26267;
  assign n26269 = pi17 ? n99 : n26268;
  assign n26270 = pi16 ? n744 : n26269;
  assign n26271 = pi15 ? n24530 : n26270;
  assign n26272 = pi20 ? n24957 : n4749;
  assign n26273 = pi19 ? n26272 : n32;
  assign n26274 = pi18 ? n24956 : n26273;
  assign n26275 = pi17 ? n139 : n26274;
  assign n26276 = pi16 ? n25417 : n26275;
  assign n26277 = pi20 ? n18317 : n4789;
  assign n26278 = pi19 ? n26277 : n32;
  assign n26279 = pi18 ? n24963 : n26278;
  assign n26280 = pi17 ? n139 : n26279;
  assign n26281 = pi16 ? n331 : n26280;
  assign n26282 = pi15 ? n26276 : n26281;
  assign n26283 = pi14 ? n26271 : n26282;
  assign n26284 = pi20 ? n316 : n4789;
  assign n26285 = pi19 ? n26284 : n32;
  assign n26286 = pi18 ? n24977 : n26285;
  assign n26287 = pi17 ? n25853 : n26286;
  assign n26288 = pi16 ? n11804 : n26287;
  assign n26289 = pi18 ? n24995 : n26285;
  assign n26290 = pi17 ? n204 : n26289;
  assign n26291 = pi16 ? n24565 : n26290;
  assign n26292 = pi15 ? n26288 : n26291;
  assign n26293 = pi21 ? n4208 : n32;
  assign n26294 = pi20 ? n316 : n26293;
  assign n26295 = pi19 ? n26294 : n32;
  assign n26296 = pi18 ? n24995 : n26295;
  assign n26297 = pi17 ? n25865 : n26296;
  assign n26298 = pi16 ? n13477 : n26297;
  assign n26299 = pi22 ? n316 : n1043;
  assign n26300 = pi21 ? n139 : n26299;
  assign n26301 = pi20 ? n26300 : n25869;
  assign n26302 = pi19 ? n15405 : n26301;
  assign n26303 = pi22 ? n4079 : n625;
  assign n26304 = pi21 ? n26303 : n32;
  assign n26305 = pi20 ? n1026 : n26304;
  assign n26306 = pi19 ? n26305 : n32;
  assign n26307 = pi18 ? n26302 : n26306;
  assign n26308 = pi17 ? n25865 : n26307;
  assign n26309 = pi16 ? n21002 : n26308;
  assign n26310 = pi15 ? n26298 : n26309;
  assign n26311 = pi14 ? n26292 : n26310;
  assign n26312 = pi13 ? n26283 : n26311;
  assign n26313 = pi12 ? n26265 : n26312;
  assign n26314 = pi20 ? n1026 : n7003;
  assign n26315 = pi19 ? n26314 : n32;
  assign n26316 = pi18 ? n139 : n26315;
  assign n26317 = pi17 ? n139 : n26316;
  assign n26318 = pi16 ? n2291 : n26317;
  assign n26319 = pi20 ? n6577 : n20391;
  assign n26320 = pi19 ? n26319 : n32;
  assign n26321 = pi18 ? n25887 : n26320;
  assign n26322 = pi17 ? n139 : n26321;
  assign n26323 = pi16 ? n2291 : n26322;
  assign n26324 = pi15 ? n26318 : n26323;
  assign n26325 = pi20 ? n1026 : n7049;
  assign n26326 = pi19 ? n26325 : n32;
  assign n26327 = pi18 ? n25895 : n26326;
  assign n26328 = pi17 ? n139 : n26327;
  assign n26329 = pi16 ? n915 : n26328;
  assign n26330 = pi20 ? n204 : n5830;
  assign n26331 = pi19 ? n26330 : n32;
  assign n26332 = pi18 ? n25908 : n26331;
  assign n26333 = pi17 ? n25907 : n26332;
  assign n26334 = pi16 ? n25903 : n26333;
  assign n26335 = pi15 ? n26329 : n26334;
  assign n26336 = pi14 ? n26324 : n26335;
  assign n26337 = pi20 ? n233 : n2653;
  assign n26338 = pi19 ? n26337 : n32;
  assign n26339 = pi18 ? n25916 : n26338;
  assign n26340 = pi17 ? n335 : n26339;
  assign n26341 = pi16 ? n7943 : n26340;
  assign n26342 = pi18 ? n25082 : n25918;
  assign n26343 = pi17 ? n335 : n26342;
  assign n26344 = pi16 ? n25923 : n26343;
  assign n26345 = pi15 ? n26341 : n26344;
  assign n26346 = pi14 ? n26345 : n25939;
  assign n26347 = pi13 ? n26336 : n26346;
  assign n26348 = pi21 ? n25984 : n37;
  assign n26349 = pi20 ? n32 : n26348;
  assign n26350 = pi19 ? n32 : n26349;
  assign n26351 = pi18 ? n26350 : n8929;
  assign n26352 = pi17 ? n32 : n26351;
  assign n26353 = pi19 ? n21125 : n13337;
  assign n26354 = pi18 ? n26353 : n26000;
  assign n26355 = pi21 ? n233 : n11199;
  assign n26356 = pi22 ? n233 : n2116;
  assign n26357 = pi21 ? n233 : n26356;
  assign n26358 = pi20 ? n26355 : n26357;
  assign n26359 = pi19 ? n233 : n26358;
  assign n26360 = pi22 ? n233 : n583;
  assign n26361 = pi21 ? n26360 : n18411;
  assign n26362 = pi20 ? n26361 : n32;
  assign n26363 = pi19 ? n26362 : n32;
  assign n26364 = pi18 ? n26359 : n26363;
  assign n26365 = pi17 ? n26354 : n26364;
  assign n26366 = pi16 ? n26352 : n26365;
  assign n26367 = pi15 ? n25983 : n26366;
  assign n26368 = pi14 ? n25976 : n26367;
  assign n26369 = pi21 ? n233 : n19438;
  assign n26370 = pi20 ? n26369 : n32;
  assign n26371 = pi19 ? n26370 : n32;
  assign n26372 = pi18 ? n233 : n26371;
  assign n26373 = pi17 ? n25173 : n26372;
  assign n26374 = pi16 ? n26020 : n26373;
  assign n26375 = pi15 ? n26374 : n26048;
  assign n26376 = pi23 ? n13482 : n32;
  assign n26377 = pi22 ? n685 : n26376;
  assign n26378 = pi21 ? n363 : n26377;
  assign n26379 = pi20 ? n26378 : n32;
  assign n26380 = pi19 ? n26379 : n32;
  assign n26381 = pi18 ? n25209 : n26380;
  assign n26382 = pi17 ? n363 : n26381;
  assign n26383 = pi16 ? n21561 : n26382;
  assign n26384 = pi18 ? n25209 : n25204;
  assign n26385 = pi17 ? n363 : n26384;
  assign n26386 = pi16 ? n21561 : n26385;
  assign n26387 = pi15 ? n26383 : n26386;
  assign n26388 = pi14 ? n26375 : n26387;
  assign n26389 = pi13 ? n26368 : n26388;
  assign n26390 = pi12 ? n26347 : n26389;
  assign n26391 = pi11 ? n26313 : n26390;
  assign n26392 = pi10 ? n26217 : n26391;
  assign n26393 = pi09 ? n26082 : n26392;
  assign n26394 = pi08 ? n26070 : n26393;
  assign n26395 = pi07 ? n25551 : n26394;
  assign n26396 = pi06 ? n24646 : n26395;
  assign n26397 = pi19 ? n87 : n32;
  assign n26398 = pi18 ? n37 : n26397;
  assign n26399 = pi17 ? n37 : n26398;
  assign n26400 = pi16 ? n14445 : n26399;
  assign n26401 = pi15 ? n32 : n26400;
  assign n26402 = pi20 ? n37 : n121;
  assign n26403 = pi19 ? n26402 : n32;
  assign n26404 = pi18 ? n37 : n26403;
  assign n26405 = pi17 ? n37 : n26404;
  assign n26406 = pi16 ? n14445 : n26405;
  assign n26407 = pi20 ? n37 : n99;
  assign n26408 = pi19 ? n37 : n26407;
  assign n26409 = pi20 ? n99 : n14887;
  assign n26410 = pi19 ? n26409 : n18853;
  assign n26411 = pi18 ? n26408 : n26410;
  assign n26412 = pi19 ? n122 : n32;
  assign n26413 = pi18 ? n99 : n26412;
  assign n26414 = pi17 ? n26411 : n26413;
  assign n26415 = pi16 ? n16595 : n26414;
  assign n26416 = pi15 ? n26406 : n26415;
  assign n26417 = pi14 ? n26401 : n26416;
  assign n26418 = pi13 ? n32 : n26417;
  assign n26419 = pi12 ? n32 : n26418;
  assign n26420 = pi11 ? n32 : n26419;
  assign n26421 = pi10 ? n32 : n26420;
  assign n26422 = pi19 ? n15951 : n5077;
  assign n26423 = pi18 ? n37 : n26422;
  assign n26424 = pi20 ? n218 : n221;
  assign n26425 = pi19 ? n26424 : n15951;
  assign n26426 = pi20 ? n4202 : n142;
  assign n26427 = pi19 ? n26426 : n32;
  assign n26428 = pi18 ? n26425 : n26427;
  assign n26429 = pi17 ? n26423 : n26428;
  assign n26430 = pi16 ? n16595 : n26429;
  assign n26431 = pi20 ? n2973 : n3039;
  assign n26432 = pi19 ? n26431 : n37;
  assign n26433 = pi20 ? n99 : n13056;
  assign n26434 = pi19 ? n26433 : n32;
  assign n26435 = pi18 ? n26432 : n26434;
  assign n26436 = pi17 ? n37 : n26435;
  assign n26437 = pi16 ? n17010 : n26436;
  assign n26438 = pi15 ? n26430 : n26437;
  assign n26439 = pi20 ? n14887 : n12261;
  assign n26440 = pi19 ? n26439 : n32;
  assign n26441 = pi18 ? n37 : n26440;
  assign n26442 = pi17 ? n37 : n26441;
  assign n26443 = pi16 ? n17010 : n26442;
  assign n26444 = pi16 ? n439 : n26442;
  assign n26445 = pi15 ? n26443 : n26444;
  assign n26446 = pi14 ? n26438 : n26445;
  assign n26447 = pi18 ? n184 : n18854;
  assign n26448 = pi17 ? n32 : n26447;
  assign n26449 = pi16 ? n26448 : n26094;
  assign n26450 = pi15 ? n26449 : n26096;
  assign n26451 = pi22 ? n1504 : n112;
  assign n26452 = pi21 ? n26451 : n2156;
  assign n26453 = pi20 ? n32 : n26452;
  assign n26454 = pi19 ? n32 : n26453;
  assign n26455 = pi22 ? n2160 : n139;
  assign n26456 = pi21 ? n2175 : n26455;
  assign n26457 = pi20 ? n26456 : n139;
  assign n26458 = pi19 ? n5501 : n26457;
  assign n26459 = pi18 ? n26454 : n26458;
  assign n26460 = pi17 ? n32 : n26459;
  assign n26461 = pi17 ? n139 : n26106;
  assign n26462 = pi16 ? n26460 : n26461;
  assign n26463 = pi17 ? n9797 : n26106;
  assign n26464 = pi16 ? n439 : n26463;
  assign n26465 = pi15 ? n26462 : n26464;
  assign n26466 = pi14 ? n26450 : n26465;
  assign n26467 = pi13 ? n26446 : n26466;
  assign n26468 = pi18 ? n13183 : n26105;
  assign n26469 = pi17 ? n9826 : n26468;
  assign n26470 = pi16 ? n439 : n26469;
  assign n26471 = pi20 ? n139 : n3096;
  assign n26472 = pi20 ? n3090 : n139;
  assign n26473 = pi19 ? n26471 : n26472;
  assign n26474 = pi18 ? n26473 : n26105;
  assign n26475 = pi17 ? n18075 : n26474;
  assign n26476 = pi16 ? n439 : n26475;
  assign n26477 = pi15 ? n26470 : n26476;
  assign n26478 = pi19 ? n21712 : n9814;
  assign n26479 = pi18 ? n26478 : n26120;
  assign n26480 = pi17 ? n19830 : n26479;
  assign n26481 = pi16 ? n439 : n26480;
  assign n26482 = pi21 ? n1046 : n139;
  assign n26483 = pi20 ? n26482 : n26118;
  assign n26484 = pi19 ? n26483 : n32;
  assign n26485 = pi18 ? n16093 : n26484;
  assign n26486 = pi17 ? n37 : n26485;
  assign n26487 = pi16 ? n439 : n26486;
  assign n26488 = pi15 ? n26481 : n26487;
  assign n26489 = pi14 ? n26477 : n26488;
  assign n26490 = pi21 ? n916 : n18927;
  assign n26491 = pi20 ? n922 : n26490;
  assign n26492 = pi19 ? n26491 : n32;
  assign n26493 = pi18 ? n16093 : n26492;
  assign n26494 = pi17 ? n37 : n26493;
  assign n26495 = pi16 ? n439 : n26494;
  assign n26496 = pi15 ? n26495 : n26145;
  assign n26497 = pi21 ? n297 : n1056;
  assign n26498 = pi20 ? n37 : n26497;
  assign n26499 = pi19 ? n37 : n26498;
  assign n26500 = pi18 ? n26499 : n26138;
  assign n26501 = pi17 ? n37 : n26500;
  assign n26502 = pi16 ? n439 : n26501;
  assign n26503 = pi19 ? n37 : n20743;
  assign n26504 = pi21 ? n2091 : n11808;
  assign n26505 = pi20 ? n26504 : n25685;
  assign n26506 = pi19 ? n26505 : n32;
  assign n26507 = pi18 ? n26503 : n26506;
  assign n26508 = pi17 ? n37 : n26507;
  assign n26509 = pi16 ? n439 : n26508;
  assign n26510 = pi15 ? n26502 : n26509;
  assign n26511 = pi14 ? n26496 : n26510;
  assign n26512 = pi13 ? n26489 : n26511;
  assign n26513 = pi12 ? n26467 : n26512;
  assign n26514 = pi21 ? n233 : n7041;
  assign n26515 = pi20 ? n7705 : n26514;
  assign n26516 = pi19 ? n26515 : n32;
  assign n26517 = pi18 ? n2102 : n26516;
  assign n26518 = pi17 ? n37 : n26517;
  assign n26519 = pi16 ? n439 : n26518;
  assign n26520 = pi20 ? n605 : n12432;
  assign n26521 = pi19 ? n26520 : n32;
  assign n26522 = pi18 ? n7686 : n26521;
  assign n26523 = pi17 ? n37 : n26522;
  assign n26524 = pi16 ? n439 : n26523;
  assign n26525 = pi15 ? n26519 : n26524;
  assign n26526 = pi20 ? n569 : n12042;
  assign n26527 = pi19 ? n26526 : n32;
  assign n26528 = pi18 ? n37 : n26527;
  assign n26529 = pi17 ? n37 : n26528;
  assign n26530 = pi16 ? n439 : n26529;
  assign n26531 = pi20 ? n577 : n12432;
  assign n26532 = pi19 ? n26531 : n32;
  assign n26533 = pi18 ? n7677 : n26532;
  assign n26534 = pi17 ? n37 : n26533;
  assign n26535 = pi16 ? n439 : n26534;
  assign n26536 = pi15 ? n26530 : n26535;
  assign n26537 = pi14 ? n26525 : n26536;
  assign n26538 = pi21 ? n570 : n7034;
  assign n26539 = pi20 ? n37 : n26538;
  assign n26540 = pi19 ? n26539 : n32;
  assign n26541 = pi18 ? n7686 : n26540;
  assign n26542 = pi17 ? n37 : n26541;
  assign n26543 = pi16 ? n439 : n26542;
  assign n26544 = pi21 ? n569 : n5771;
  assign n26545 = pi20 ? n649 : n26544;
  assign n26546 = pi19 ? n26545 : n32;
  assign n26547 = pi18 ? n24789 : n26546;
  assign n26548 = pi17 ? n37 : n26547;
  assign n26549 = pi16 ? n439 : n26548;
  assign n26550 = pi15 ? n26543 : n26549;
  assign n26551 = pi21 ? n335 : n5771;
  assign n26552 = pi20 ? n37 : n26551;
  assign n26553 = pi19 ? n26552 : n32;
  assign n26554 = pi18 ? n37 : n26553;
  assign n26555 = pi17 ? n37 : n26554;
  assign n26556 = pi16 ? n439 : n26555;
  assign n26557 = pi21 ? n4973 : n7034;
  assign n26558 = pi20 ? n37 : n26557;
  assign n26559 = pi19 ? n26558 : n32;
  assign n26560 = pi18 ? n37 : n26559;
  assign n26561 = pi17 ? n37 : n26560;
  assign n26562 = pi16 ? n439 : n26561;
  assign n26563 = pi15 ? n26556 : n26562;
  assign n26564 = pi14 ? n26550 : n26563;
  assign n26565 = pi13 ? n26537 : n26564;
  assign n26566 = pi21 ? n2091 : n7041;
  assign n26567 = pi20 ? n37 : n26566;
  assign n26568 = pi19 ? n26567 : n32;
  assign n26569 = pi18 ? n37 : n26568;
  assign n26570 = pi17 ? n37 : n26569;
  assign n26571 = pi16 ? n439 : n26570;
  assign n26572 = pi21 ? n3392 : n4101;
  assign n26573 = pi20 ? n37 : n26572;
  assign n26574 = pi19 ? n26573 : n32;
  assign n26575 = pi18 ? n37 : n26574;
  assign n26576 = pi17 ? n37 : n26575;
  assign n26577 = pi16 ? n439 : n26576;
  assign n26578 = pi15 ? n26571 : n26577;
  assign n26579 = pi21 ? n3392 : n7048;
  assign n26580 = pi20 ? n37 : n26579;
  assign n26581 = pi19 ? n26580 : n32;
  assign n26582 = pi18 ? n37 : n26581;
  assign n26583 = pi17 ? n37 : n26582;
  assign n26584 = pi16 ? n439 : n26583;
  assign n26585 = pi21 ? n6401 : n760;
  assign n26586 = pi20 ? n37 : n26585;
  assign n26587 = pi19 ? n26586 : n32;
  assign n26588 = pi18 ? n37 : n26587;
  assign n26589 = pi17 ? n37 : n26588;
  assign n26590 = pi16 ? n439 : n26589;
  assign n26591 = pi15 ? n26584 : n26590;
  assign n26592 = pi14 ? n26578 : n26591;
  assign n26593 = pi21 ? n6401 : n882;
  assign n26594 = pi20 ? n37 : n26593;
  assign n26595 = pi19 ? n26594 : n32;
  assign n26596 = pi18 ? n37 : n26595;
  assign n26597 = pi17 ? n37 : n26596;
  assign n26598 = pi16 ? n439 : n26597;
  assign n26599 = pi21 ? n6401 : n928;
  assign n26600 = pi20 ? n37 : n26599;
  assign n26601 = pi19 ? n26600 : n32;
  assign n26602 = pi18 ? n37 : n26601;
  assign n26603 = pi17 ? n37 : n26602;
  assign n26604 = pi16 ? n439 : n26603;
  assign n26605 = pi15 ? n26598 : n26604;
  assign n26606 = pi20 ? n7730 : n37;
  assign n26607 = pi19 ? n37 : n26606;
  assign n26608 = pi21 ? n6401 : n2469;
  assign n26609 = pi20 ? n37 : n26608;
  assign n26610 = pi19 ? n26609 : n32;
  assign n26611 = pi18 ? n26607 : n26610;
  assign n26612 = pi17 ? n37 : n26611;
  assign n26613 = pi16 ? n439 : n26612;
  assign n26614 = pi19 ? n37 : n24880;
  assign n26615 = pi21 ? n363 : n2469;
  assign n26616 = pi20 ? n363 : n26615;
  assign n26617 = pi19 ? n26616 : n32;
  assign n26618 = pi18 ? n26614 : n26617;
  assign n26619 = pi17 ? n37 : n26618;
  assign n26620 = pi16 ? n439 : n26619;
  assign n26621 = pi15 ? n26613 : n26620;
  assign n26622 = pi14 ? n26605 : n26621;
  assign n26623 = pi13 ? n26592 : n26622;
  assign n26624 = pi12 ? n26565 : n26623;
  assign n26625 = pi11 ? n26513 : n26624;
  assign n26626 = pi21 ? n8567 : n6401;
  assign n26627 = pi20 ? n26626 : n6402;
  assign n26628 = pi19 ? n37 : n26627;
  assign n26629 = pi21 ? n244 : n2553;
  assign n26630 = pi20 ? n37 : n26629;
  assign n26631 = pi19 ? n26630 : n32;
  assign n26632 = pi18 ? n26628 : n26631;
  assign n26633 = pi17 ? n37 : n26632;
  assign n26634 = pi16 ? n439 : n26633;
  assign n26635 = pi20 ? n37 : n7407;
  assign n26636 = pi19 ? n26635 : n32;
  assign n26637 = pi18 ? n37 : n26636;
  assign n26638 = pi17 ? n37 : n26637;
  assign n26639 = pi16 ? n439 : n26638;
  assign n26640 = pi15 ? n26634 : n26639;
  assign n26641 = pi21 ? n6461 : n14277;
  assign n26642 = pi20 ? n157 : n26641;
  assign n26643 = pi19 ? n37 : n26642;
  assign n26644 = pi20 ? n787 : n7407;
  assign n26645 = pi19 ? n26644 : n32;
  assign n26646 = pi18 ? n26643 : n26645;
  assign n26647 = pi17 ? n37 : n26646;
  assign n26648 = pi16 ? n439 : n26647;
  assign n26649 = pi20 ? n157 : n6461;
  assign n26650 = pi19 ? n37 : n26649;
  assign n26651 = pi20 ? n7818 : n12909;
  assign n26652 = pi19 ? n26651 : n32;
  assign n26653 = pi18 ? n26650 : n26652;
  assign n26654 = pi17 ? n37 : n26653;
  assign n26655 = pi16 ? n439 : n26654;
  assign n26656 = pi15 ? n26648 : n26655;
  assign n26657 = pi14 ? n26640 : n26656;
  assign n26658 = pi19 ? n99 : n9715;
  assign n26659 = pi20 ? n99 : n12919;
  assign n26660 = pi19 ? n26659 : n32;
  assign n26661 = pi18 ? n26658 : n26660;
  assign n26662 = pi17 ? n99 : n26661;
  assign n26663 = pi16 ? n721 : n26662;
  assign n26664 = pi18 ? n99 : n26660;
  assign n26665 = pi17 ? n99 : n26664;
  assign n26666 = pi16 ? n721 : n26665;
  assign n26667 = pi15 ? n26663 : n26666;
  assign n26668 = pi19 ? n99 : n20936;
  assign n26669 = pi18 ? n26668 : n26660;
  assign n26670 = pi17 ? n99 : n26669;
  assign n26671 = pi16 ? n721 : n26670;
  assign n26672 = pi20 ? n99 : n12508;
  assign n26673 = pi19 ? n26672 : n32;
  assign n26674 = pi18 ? n26668 : n26673;
  assign n26675 = pi17 ? n99 : n26674;
  assign n26676 = pi16 ? n721 : n26675;
  assign n26677 = pi15 ? n26671 : n26676;
  assign n26678 = pi14 ? n26667 : n26677;
  assign n26679 = pi13 ? n26657 : n26678;
  assign n26680 = pi21 ? n139 : n99;
  assign n26681 = pi20 ? n139 : n26680;
  assign n26682 = pi20 ? n139 : n14846;
  assign n26683 = pi19 ? n26681 : n26682;
  assign n26684 = pi18 ? n139 : n26683;
  assign n26685 = pi20 ? n99 : n6508;
  assign n26686 = pi19 ? n139 : n26685;
  assign n26687 = pi22 ? n157 : n843;
  assign n26688 = pi21 ? n26687 : n32;
  assign n26689 = pi20 ? n157 : n26688;
  assign n26690 = pi19 ? n26689 : n32;
  assign n26691 = pi18 ? n26686 : n26690;
  assign n26692 = pi17 ? n26684 : n26691;
  assign n26693 = pi16 ? n24953 : n26692;
  assign n26694 = pi19 ? n139 : n13371;
  assign n26695 = pi22 ? n157 : n2530;
  assign n26696 = pi21 ? n26695 : n32;
  assign n26697 = pi20 ? n99 : n26696;
  assign n26698 = pi19 ? n26697 : n32;
  assign n26699 = pi18 ? n26694 : n26698;
  assign n26700 = pi17 ? n26684 : n26699;
  assign n26701 = pi16 ? n24953 : n26700;
  assign n26702 = pi15 ? n26693 : n26701;
  assign n26703 = pi20 ? n975 : n6158;
  assign n26704 = pi19 ? n139 : n26703;
  assign n26705 = pi20 ? n1027 : n13429;
  assign n26706 = pi19 ? n26705 : n32;
  assign n26707 = pi18 ? n26704 : n26706;
  assign n26708 = pi17 ? n139 : n26707;
  assign n26709 = pi16 ? n2291 : n26708;
  assign n26710 = pi20 ? n316 : n13429;
  assign n26711 = pi19 ? n26710 : n32;
  assign n26712 = pi18 ? n17418 : n26711;
  assign n26713 = pi17 ? n139 : n26712;
  assign n26714 = pi16 ? n1773 : n26713;
  assign n26715 = pi15 ? n26709 : n26714;
  assign n26716 = pi14 ? n26702 : n26715;
  assign n26717 = pi20 ? n204 : n37;
  assign n26718 = pi19 ? n26717 : n21732;
  assign n26719 = pi18 ? n24984 : n26718;
  assign n26720 = pi19 ? n15421 : n316;
  assign n26721 = pi20 ? n316 : n5667;
  assign n26722 = pi19 ? n26721 : n32;
  assign n26723 = pi18 ? n26720 : n26722;
  assign n26724 = pi17 ? n26719 : n26723;
  assign n26725 = pi16 ? n11804 : n26724;
  assign n26726 = pi19 ? n204 : n3736;
  assign n26727 = pi18 ? n26726 : n26722;
  assign n26728 = pi17 ? n204 : n26727;
  assign n26729 = pi16 ? n13493 : n26728;
  assign n26730 = pi15 ? n26725 : n26729;
  assign n26731 = pi19 ? n204 : n16494;
  assign n26732 = pi18 ? n204 : n26731;
  assign n26733 = pi19 ? n204 : n3732;
  assign n26734 = pi20 ? n2383 : n5667;
  assign n26735 = pi19 ? n26734 : n32;
  assign n26736 = pi18 ? n26733 : n26735;
  assign n26737 = pi17 ? n26732 : n26736;
  assign n26738 = pi16 ? n13846 : n26737;
  assign n26739 = pi20 ? n3087 : n204;
  assign n26740 = pi19 ? n204 : n26739;
  assign n26741 = pi18 ? n204 : n26740;
  assign n26742 = pi20 ? n1016 : n204;
  assign n26743 = pi19 ? n204 : n26742;
  assign n26744 = pi20 ? n204 : n4852;
  assign n26745 = pi19 ? n26744 : n32;
  assign n26746 = pi18 ? n26743 : n26745;
  assign n26747 = pi17 ? n26741 : n26746;
  assign n26748 = pi16 ? n13833 : n26747;
  assign n26749 = pi15 ? n26738 : n26748;
  assign n26750 = pi14 ? n26730 : n26749;
  assign n26751 = pi13 ? n26716 : n26750;
  assign n26752 = pi12 ? n26679 : n26751;
  assign n26753 = pi20 ? n6158 : n8295;
  assign n26754 = pi19 ? n26753 : n32;
  assign n26755 = pi18 ? n25895 : n26754;
  assign n26756 = pi17 ? n139 : n26755;
  assign n26757 = pi16 ? n915 : n26756;
  assign n26758 = pi20 ? n1016 : n4008;
  assign n26759 = pi19 ? n26758 : n32;
  assign n26760 = pi18 ? n23054 : n26759;
  assign n26761 = pi17 ? n139 : n26760;
  assign n26762 = pi16 ? n915 : n26761;
  assign n26763 = pi15 ? n26757 : n26762;
  assign n26764 = pi22 ? n909 : n335;
  assign n26765 = pi21 ? n26764 : n139;
  assign n26766 = pi20 ? n32 : n26765;
  assign n26767 = pi19 ? n32 : n26766;
  assign n26768 = pi21 ? n9126 : n139;
  assign n26769 = pi21 ? n9126 : n1711;
  assign n26770 = pi20 ? n26768 : n26769;
  assign n26771 = pi20 ? n3922 : n10927;
  assign n26772 = pi19 ? n26770 : n26771;
  assign n26773 = pi18 ? n26767 : n26772;
  assign n26774 = pi17 ? n32 : n26773;
  assign n26775 = pi21 ? n9144 : n9146;
  assign n26776 = pi21 ? n295 : n9146;
  assign n26777 = pi20 ? n26775 : n26776;
  assign n26778 = pi19 ? n26777 : n26776;
  assign n26779 = pi21 ? n9119 : n1698;
  assign n26780 = pi20 ? n26779 : n25049;
  assign n26781 = pi21 ? n1711 : n9119;
  assign n26782 = pi20 ? n9127 : n26781;
  assign n26783 = pi19 ? n26780 : n26782;
  assign n26784 = pi18 ? n26778 : n26783;
  assign n26785 = pi21 ? n9144 : n9119;
  assign n26786 = pi20 ? n26785 : n10927;
  assign n26787 = pi21 ? n9122 : n204;
  assign n26788 = pi20 ? n26787 : n5204;
  assign n26789 = pi19 ? n26786 : n26788;
  assign n26790 = pi20 ? n204 : n3210;
  assign n26791 = pi19 ? n26790 : n32;
  assign n26792 = pi18 ? n26789 : n26791;
  assign n26793 = pi17 ? n26784 : n26792;
  assign n26794 = pi16 ? n26774 : n26793;
  assign n26795 = pi19 ? n10957 : n17204;
  assign n26796 = pi18 ? n7941 : n26795;
  assign n26797 = pi17 ? n32 : n26796;
  assign n26798 = pi21 ? n1940 : n233;
  assign n26799 = pi20 ? n26798 : n10011;
  assign n26800 = pi19 ? n26799 : n32;
  assign n26801 = pi18 ? n17534 : n26800;
  assign n26802 = pi17 ? n335 : n26801;
  assign n26803 = pi16 ? n26797 : n26802;
  assign n26804 = pi15 ? n26794 : n26803;
  assign n26805 = pi14 ? n26763 : n26804;
  assign n26806 = pi20 ? n233 : n3398;
  assign n26807 = pi19 ? n26806 : n32;
  assign n26808 = pi18 ? n17540 : n26807;
  assign n26809 = pi17 ? n335 : n26808;
  assign n26810 = pi16 ? n7943 : n26809;
  assign n26811 = pi20 ? n233 : n2679;
  assign n26812 = pi19 ? n26811 : n32;
  assign n26813 = pi18 ? n17540 : n26812;
  assign n26814 = pi17 ? n335 : n26813;
  assign n26815 = pi16 ? n7943 : n26814;
  assign n26816 = pi15 ? n26810 : n26815;
  assign n26817 = pi19 ? n25087 : n37;
  assign n26818 = pi18 ? n37 : n26817;
  assign n26819 = pi20 ? n7705 : n233;
  assign n26820 = pi19 ? n17204 : n26819;
  assign n26821 = pi18 ? n26820 : n26812;
  assign n26822 = pi17 ? n26818 : n26821;
  assign n26823 = pi16 ? n439 : n26822;
  assign n26824 = pi18 ? n3286 : n26817;
  assign n26825 = pi19 ? n18408 : n233;
  assign n26826 = pi20 ? n233 : n2701;
  assign n26827 = pi19 ? n26826 : n32;
  assign n26828 = pi18 ? n26825 : n26827;
  assign n26829 = pi17 ? n26824 : n26828;
  assign n26830 = pi16 ? n439 : n26829;
  assign n26831 = pi15 ? n26823 : n26830;
  assign n26832 = pi14 ? n26816 : n26831;
  assign n26833 = pi13 ? n26805 : n26832;
  assign n26834 = pi22 ? n8880 : n233;
  assign n26835 = pi21 ? n26834 : n233;
  assign n26836 = pi20 ? n32 : n26835;
  assign n26837 = pi19 ? n32 : n26836;
  assign n26838 = pi19 ? n233 : n13337;
  assign n26839 = pi18 ? n26837 : n26838;
  assign n26840 = pi17 ? n32 : n26839;
  assign n26841 = pi19 ? n233 : n13535;
  assign n26842 = pi18 ? n233 : n26841;
  assign n26843 = pi18 ? n233 : n25918;
  assign n26844 = pi17 ? n26842 : n26843;
  assign n26845 = pi16 ? n26840 : n26844;
  assign n26846 = pi21 ? n2091 : n2048;
  assign n26847 = pi20 ? n26846 : n37;
  assign n26848 = pi19 ? n26847 : n37;
  assign n26849 = pi18 ? n37 : n26848;
  assign n26850 = pi18 ? n18113 : n25918;
  assign n26851 = pi17 ? n26849 : n26850;
  assign n26852 = pi16 ? n439 : n26851;
  assign n26853 = pi15 ? n26845 : n26852;
  assign n26854 = pi18 ? n18113 : n25967;
  assign n26855 = pi17 ? n26849 : n26854;
  assign n26856 = pi16 ? n439 : n26855;
  assign n26857 = pi22 ? n55 : n233;
  assign n26858 = pi21 ? n26857 : n233;
  assign n26859 = pi20 ? n32 : n26858;
  assign n26860 = pi19 ? n32 : n26859;
  assign n26861 = pi20 ? n233 : n21124;
  assign n26862 = pi20 ? n14844 : n233;
  assign n26863 = pi19 ? n26861 : n26862;
  assign n26864 = pi18 ? n26860 : n26863;
  assign n26865 = pi17 ? n32 : n26864;
  assign n26866 = pi18 ? n233 : n25980;
  assign n26867 = pi17 ? n233 : n26866;
  assign n26868 = pi16 ? n26865 : n26867;
  assign n26869 = pi15 ? n26856 : n26868;
  assign n26870 = pi14 ? n26853 : n26869;
  assign n26871 = pi21 ? n25162 : n22128;
  assign n26872 = pi20 ? n32 : n26871;
  assign n26873 = pi19 ? n32 : n26872;
  assign n26874 = pi20 ? n363 : n9197;
  assign n26875 = pi19 ? n21222 : n26874;
  assign n26876 = pi18 ? n26873 : n26875;
  assign n26877 = pi17 ? n32 : n26876;
  assign n26878 = pi20 ? n9197 : n233;
  assign n26879 = pi19 ? n26878 : n233;
  assign n26880 = pi21 ? n233 : n9196;
  assign n26881 = pi20 ? n9197 : n26880;
  assign n26882 = pi19 ? n233 : n26881;
  assign n26883 = pi18 ? n26879 : n26882;
  assign n26884 = pi17 ? n26883 : n26866;
  assign n26885 = pi16 ? n26877 : n26884;
  assign n26886 = pi18 ? n23570 : n363;
  assign n26887 = pi17 ? n32 : n26886;
  assign n26888 = pi20 ? n20866 : n363;
  assign n26889 = pi19 ? n26888 : n363;
  assign n26890 = pi21 ? n2721 : n24222;
  assign n26891 = pi21 ? n685 : n363;
  assign n26892 = pi20 ? n26890 : n26891;
  assign n26893 = pi20 ? n26890 : n19084;
  assign n26894 = pi19 ? n26892 : n26893;
  assign n26895 = pi18 ? n26889 : n26894;
  assign n26896 = pi20 ? n24223 : n685;
  assign n26897 = pi21 ? n24222 : n21235;
  assign n26898 = pi21 ? n363 : n24222;
  assign n26899 = pi20 ? n26897 : n26898;
  assign n26900 = pi19 ? n26896 : n26899;
  assign n26901 = pi18 ? n26900 : n25533;
  assign n26902 = pi17 ? n26895 : n26901;
  assign n26903 = pi16 ? n26887 : n26902;
  assign n26904 = pi15 ? n26885 : n26903;
  assign n26905 = pi21 ? n24222 : n363;
  assign n26906 = pi20 ? n19084 : n26905;
  assign n26907 = pi19 ? n363 : n26906;
  assign n26908 = pi22 ? n685 : n21078;
  assign n26909 = pi21 ? n24222 : n26908;
  assign n26910 = pi20 ? n26909 : n32;
  assign n26911 = pi19 ? n26910 : n32;
  assign n26912 = pi18 ? n26907 : n26911;
  assign n26913 = pi17 ? n363 : n26912;
  assign n26914 = pi16 ? n21219 : n26913;
  assign n26915 = pi21 ? n24222 : n3523;
  assign n26916 = pi20 ? n26915 : n32;
  assign n26917 = pi19 ? n26916 : n32;
  assign n26918 = pi18 ? n26907 : n26917;
  assign n26919 = pi17 ? n363 : n26918;
  assign n26920 = pi16 ? n26062 : n26919;
  assign n26921 = pi15 ? n26914 : n26920;
  assign n26922 = pi14 ? n26904 : n26921;
  assign n26923 = pi13 ? n26870 : n26922;
  assign n26924 = pi12 ? n26833 : n26923;
  assign n26925 = pi11 ? n26752 : n26924;
  assign n26926 = pi10 ? n26625 : n26925;
  assign n26927 = pi09 ? n26421 : n26926;
  assign n26928 = pi21 ? n37 : n19793;
  assign n26929 = pi20 ? n14887 : n26928;
  assign n26930 = pi19 ? n26929 : n32;
  assign n26931 = pi18 ? n37 : n26930;
  assign n26932 = pi17 ? n37 : n26931;
  assign n26933 = pi16 ? n17010 : n26932;
  assign n26934 = pi15 ? n26933 : n26444;
  assign n26935 = pi14 ? n26438 : n26934;
  assign n26936 = pi20 ? n99 : n12741;
  assign n26937 = pi19 ? n26936 : n32;
  assign n26938 = pi18 ? n99 : n26937;
  assign n26939 = pi17 ? n99 : n26938;
  assign n26940 = pi16 ? n26448 : n26939;
  assign n26941 = pi16 ? n25610 : n26939;
  assign n26942 = pi15 ? n26940 : n26941;
  assign n26943 = pi21 ? n2175 : n297;
  assign n26944 = pi20 ? n26943 : n139;
  assign n26945 = pi19 ? n14518 : n26944;
  assign n26946 = pi18 ? n14880 : n26945;
  assign n26947 = pi17 ? n32 : n26946;
  assign n26948 = pi20 ? n139 : n14107;
  assign n26949 = pi19 ? n26948 : n32;
  assign n26950 = pi18 ? n139 : n26949;
  assign n26951 = pi17 ? n139 : n26950;
  assign n26952 = pi16 ? n26947 : n26951;
  assign n26953 = pi17 ? n9797 : n26950;
  assign n26954 = pi16 ? n439 : n26953;
  assign n26955 = pi15 ? n26952 : n26954;
  assign n26956 = pi14 ? n26942 : n26955;
  assign n26957 = pi13 ? n26935 : n26956;
  assign n26958 = pi18 ? n13183 : n26949;
  assign n26959 = pi17 ? n9826 : n26958;
  assign n26960 = pi16 ? n439 : n26959;
  assign n26961 = pi18 ? n26473 : n26949;
  assign n26962 = pi17 ? n18075 : n26961;
  assign n26963 = pi16 ? n439 : n26962;
  assign n26964 = pi15 ? n26960 : n26963;
  assign n26965 = pi22 ? n139 : n23369;
  assign n26966 = pi21 ? n139 : n26965;
  assign n26967 = pi20 ? n139 : n26966;
  assign n26968 = pi19 ? n26967 : n32;
  assign n26969 = pi18 ? n26478 : n26968;
  assign n26970 = pi17 ? n19830 : n26969;
  assign n26971 = pi16 ? n439 : n26970;
  assign n26972 = pi22 ? n139 : n23380;
  assign n26973 = pi21 ? n139 : n26972;
  assign n26974 = pi20 ? n26482 : n26973;
  assign n26975 = pi19 ? n26974 : n32;
  assign n26976 = pi18 ? n16093 : n26975;
  assign n26977 = pi17 ? n37 : n26976;
  assign n26978 = pi16 ? n439 : n26977;
  assign n26979 = pi15 ? n26971 : n26978;
  assign n26980 = pi14 ? n26964 : n26979;
  assign n26981 = pi23 ? n10729 : n32;
  assign n26982 = pi22 ? n335 : n26981;
  assign n26983 = pi21 ? n916 : n26982;
  assign n26984 = pi20 ? n922 : n26983;
  assign n26985 = pi19 ? n26984 : n32;
  assign n26986 = pi18 ? n16093 : n26985;
  assign n26987 = pi17 ? n37 : n26986;
  assign n26988 = pi16 ? n439 : n26987;
  assign n26989 = pi21 ? n204 : n20341;
  assign n26990 = pi20 ? n204 : n26989;
  assign n26991 = pi19 ? n26990 : n32;
  assign n26992 = pi18 ? n25681 : n26991;
  assign n26993 = pi17 ? n37 : n26992;
  assign n26994 = pi16 ? n439 : n26993;
  assign n26995 = pi15 ? n26988 : n26994;
  assign n26996 = pi21 ? n204 : n15864;
  assign n26997 = pi20 ? n204 : n26996;
  assign n26998 = pi19 ? n26997 : n32;
  assign n26999 = pi18 ? n26499 : n26998;
  assign n27000 = pi17 ? n37 : n26999;
  assign n27001 = pi16 ? n439 : n27000;
  assign n27002 = pi21 ? n204 : n650;
  assign n27003 = pi20 ? n26504 : n27002;
  assign n27004 = pi19 ? n27003 : n32;
  assign n27005 = pi18 ? n26503 : n27004;
  assign n27006 = pi17 ? n37 : n27005;
  assign n27007 = pi16 ? n439 : n27006;
  assign n27008 = pi15 ? n27001 : n27007;
  assign n27009 = pi14 ? n26995 : n27008;
  assign n27010 = pi13 ? n26980 : n27009;
  assign n27011 = pi12 ? n26957 : n27010;
  assign n27012 = pi20 ? n7705 : n23107;
  assign n27013 = pi19 ? n27012 : n32;
  assign n27014 = pi18 ? n2102 : n27013;
  assign n27015 = pi17 ? n37 : n27014;
  assign n27016 = pi16 ? n439 : n27015;
  assign n27017 = pi21 ? n335 : n5758;
  assign n27018 = pi20 ? n605 : n27017;
  assign n27019 = pi19 ? n27018 : n32;
  assign n27020 = pi18 ? n7686 : n27019;
  assign n27021 = pi17 ? n37 : n27020;
  assign n27022 = pi16 ? n439 : n27021;
  assign n27023 = pi15 ? n27016 : n27022;
  assign n27024 = pi14 ? n27023 : n26536;
  assign n27025 = pi21 ? n574 : n13722;
  assign n27026 = pi20 ? n37 : n27025;
  assign n27027 = pi19 ? n27026 : n32;
  assign n27028 = pi18 ? n37 : n27027;
  assign n27029 = pi17 ? n37 : n27028;
  assign n27030 = pi16 ? n439 : n27029;
  assign n27031 = pi15 ? n26556 : n27030;
  assign n27032 = pi14 ? n26550 : n27031;
  assign n27033 = pi13 ? n27024 : n27032;
  assign n27034 = pi21 ? n3392 : n12825;
  assign n27035 = pi20 ? n37 : n27034;
  assign n27036 = pi19 ? n27035 : n32;
  assign n27037 = pi18 ? n37 : n27036;
  assign n27038 = pi17 ? n37 : n27037;
  assign n27039 = pi16 ? n439 : n27038;
  assign n27040 = pi15 ? n26571 : n27039;
  assign n27041 = pi14 ? n27040 : n26591;
  assign n27042 = pi21 ? n6401 : n5829;
  assign n27043 = pi20 ? n37 : n27042;
  assign n27044 = pi19 ? n27043 : n32;
  assign n27045 = pi18 ? n37 : n27044;
  assign n27046 = pi17 ? n37 : n27045;
  assign n27047 = pi16 ? n439 : n27046;
  assign n27048 = pi21 ? n6401 : n2637;
  assign n27049 = pi20 ? n37 : n27048;
  assign n27050 = pi19 ? n27049 : n32;
  assign n27051 = pi18 ? n37 : n27050;
  assign n27052 = pi17 ? n37 : n27051;
  assign n27053 = pi16 ? n439 : n27052;
  assign n27054 = pi15 ? n27047 : n27053;
  assign n27055 = pi18 ? n26607 : n27050;
  assign n27056 = pi17 ? n37 : n27055;
  assign n27057 = pi16 ? n439 : n27056;
  assign n27058 = pi21 ? n363 : n2637;
  assign n27059 = pi20 ? n363 : n27058;
  assign n27060 = pi19 ? n27059 : n32;
  assign n27061 = pi18 ? n26614 : n27060;
  assign n27062 = pi17 ? n37 : n27061;
  assign n27063 = pi16 ? n439 : n27062;
  assign n27064 = pi15 ? n27057 : n27063;
  assign n27065 = pi14 ? n27054 : n27064;
  assign n27066 = pi13 ? n27041 : n27065;
  assign n27067 = pi12 ? n27033 : n27066;
  assign n27068 = pi11 ? n27011 : n27067;
  assign n27069 = pi19 ? n37 : n6402;
  assign n27070 = pi21 ? n244 : n2637;
  assign n27071 = pi20 ? n37 : n27070;
  assign n27072 = pi19 ? n27071 : n32;
  assign n27073 = pi18 ? n27069 : n27072;
  assign n27074 = pi17 ? n37 : n27073;
  assign n27075 = pi16 ? n439 : n27074;
  assign n27076 = pi21 ? n685 : n2637;
  assign n27077 = pi20 ? n37 : n27076;
  assign n27078 = pi19 ? n27077 : n32;
  assign n27079 = pi18 ? n37 : n27078;
  assign n27080 = pi17 ? n37 : n27079;
  assign n27081 = pi16 ? n439 : n27080;
  assign n27082 = pi15 ? n27075 : n27081;
  assign n27083 = pi20 ? n787 : n27076;
  assign n27084 = pi19 ? n27083 : n32;
  assign n27085 = pi18 ? n26643 : n27084;
  assign n27086 = pi17 ? n37 : n27085;
  assign n27087 = pi16 ? n439 : n27086;
  assign n27088 = pi20 ? n7818 : n13777;
  assign n27089 = pi19 ? n27088 : n32;
  assign n27090 = pi18 ? n26650 : n27089;
  assign n27091 = pi17 ? n37 : n27090;
  assign n27092 = pi16 ? n439 : n27091;
  assign n27093 = pi15 ? n27087 : n27092;
  assign n27094 = pi14 ? n27082 : n27093;
  assign n27095 = pi21 ? n3562 : n928;
  assign n27096 = pi20 ? n99 : n27095;
  assign n27097 = pi19 ? n27096 : n32;
  assign n27098 = pi18 ? n26658 : n27097;
  assign n27099 = pi17 ? n99 : n27098;
  assign n27100 = pi16 ? n744 : n27099;
  assign n27101 = pi18 ? n99 : n27097;
  assign n27102 = pi17 ? n99 : n27101;
  assign n27103 = pi16 ? n744 : n27102;
  assign n27104 = pi15 ? n27100 : n27103;
  assign n27105 = pi18 ? n26668 : n27097;
  assign n27106 = pi17 ? n99 : n27105;
  assign n27107 = pi16 ? n744 : n27106;
  assign n27108 = pi16 ? n744 : n26670;
  assign n27109 = pi15 ? n27107 : n27108;
  assign n27110 = pi14 ? n27104 : n27109;
  assign n27111 = pi13 ? n27094 : n27110;
  assign n27112 = pi20 ? n157 : n6133;
  assign n27113 = pi19 ? n27112 : n32;
  assign n27114 = pi18 ? n26686 : n27113;
  assign n27115 = pi17 ? n26684 : n27114;
  assign n27116 = pi16 ? n25417 : n27115;
  assign n27117 = pi20 ? n99 : n6148;
  assign n27118 = pi19 ? n27117 : n32;
  assign n27119 = pi18 ? n26694 : n27118;
  assign n27120 = pi17 ? n26684 : n27119;
  assign n27121 = pi16 ? n25417 : n27120;
  assign n27122 = pi15 ? n27116 : n27121;
  assign n27123 = pi16 ? n915 : n26708;
  assign n27124 = pi15 ? n27123 : n26714;
  assign n27125 = pi14 ? n27122 : n27124;
  assign n27126 = pi20 ? n204 : n8917;
  assign n27127 = pi19 ? n27126 : n32;
  assign n27128 = pi18 ? n26743 : n27127;
  assign n27129 = pi17 ? n26741 : n27128;
  assign n27130 = pi16 ? n13833 : n27129;
  assign n27131 = pi15 ? n26738 : n27130;
  assign n27132 = pi14 ? n26730 : n27131;
  assign n27133 = pi13 ? n27125 : n27132;
  assign n27134 = pi12 ? n27111 : n27133;
  assign n27135 = pi20 ? n6158 : n9963;
  assign n27136 = pi19 ? n27135 : n32;
  assign n27137 = pi18 ? n25895 : n27136;
  assign n27138 = pi17 ? n139 : n27137;
  assign n27139 = pi16 ? n2291 : n27138;
  assign n27140 = pi16 ? n2291 : n26761;
  assign n27141 = pi15 ? n27139 : n27140;
  assign n27142 = pi21 ? n26764 : n1531;
  assign n27143 = pi20 ? n32 : n27142;
  assign n27144 = pi19 ? n32 : n27143;
  assign n27145 = pi21 ? n567 : n1531;
  assign n27146 = pi21 ? n567 : n820;
  assign n27147 = pi20 ? n27145 : n27146;
  assign n27148 = pi21 ? n10234 : n9122;
  assign n27149 = pi20 ? n3084 : n27148;
  assign n27150 = pi19 ? n27147 : n27149;
  assign n27151 = pi18 ? n27144 : n27150;
  assign n27152 = pi17 ? n32 : n27151;
  assign n27153 = pi21 ? n10234 : n570;
  assign n27154 = pi21 ? n375 : n570;
  assign n27155 = pi20 ? n27153 : n27154;
  assign n27156 = pi19 ? n27155 : n27154;
  assign n27157 = pi20 ? n9120 : n9125;
  assign n27158 = pi20 ? n9127 : n9132;
  assign n27159 = pi19 ? n27157 : n27158;
  assign n27160 = pi18 ? n27156 : n27159;
  assign n27161 = pi21 ? n9144 : n569;
  assign n27162 = pi21 ? n10234 : n9563;
  assign n27163 = pi20 ? n27161 : n27162;
  assign n27164 = pi21 ? n9563 : n204;
  assign n27165 = pi20 ? n27164 : n5204;
  assign n27166 = pi19 ? n27163 : n27165;
  assign n27167 = pi18 ? n27166 : n26791;
  assign n27168 = pi17 ? n27160 : n27167;
  assign n27169 = pi16 ? n27152 : n27168;
  assign n27170 = pi21 ? n567 : n233;
  assign n27171 = pi20 ? n27170 : n3210;
  assign n27172 = pi19 ? n27171 : n32;
  assign n27173 = pi18 ? n17534 : n27172;
  assign n27174 = pi17 ? n335 : n27173;
  assign n27175 = pi16 ? n26797 : n27174;
  assign n27176 = pi15 ? n27169 : n27175;
  assign n27177 = pi14 ? n27141 : n27176;
  assign n27178 = pi20 ? n233 : n10011;
  assign n27179 = pi19 ? n27178 : n32;
  assign n27180 = pi18 ? n17540 : n27179;
  assign n27181 = pi17 ? n335 : n27180;
  assign n27182 = pi16 ? n7943 : n27181;
  assign n27183 = pi18 ? n17540 : n26338;
  assign n27184 = pi17 ? n335 : n27183;
  assign n27185 = pi16 ? n7943 : n27184;
  assign n27186 = pi15 ? n27182 : n27185;
  assign n27187 = pi18 ? n26825 : n26812;
  assign n27188 = pi17 ? n26824 : n27187;
  assign n27189 = pi16 ? n439 : n27188;
  assign n27190 = pi15 ? n26823 : n27189;
  assign n27191 = pi14 ? n27186 : n27190;
  assign n27192 = pi13 ? n27177 : n27191;
  assign n27193 = pi18 ? n26860 : n26838;
  assign n27194 = pi17 ? n32 : n27193;
  assign n27195 = pi18 ? n233 : n26812;
  assign n27196 = pi17 ? n26842 : n27195;
  assign n27197 = pi16 ? n27194 : n27196;
  assign n27198 = pi18 ? n18113 : n26812;
  assign n27199 = pi17 ? n26849 : n27198;
  assign n27200 = pi16 ? n439 : n27199;
  assign n27201 = pi15 ? n27197 : n27200;
  assign n27202 = pi20 ? n25965 : n2701;
  assign n27203 = pi19 ? n27202 : n32;
  assign n27204 = pi18 ? n18113 : n27203;
  assign n27205 = pi17 ? n26849 : n27204;
  assign n27206 = pi16 ? n439 : n27205;
  assign n27207 = pi20 ? n25978 : n1822;
  assign n27208 = pi19 ? n27207 : n32;
  assign n27209 = pi18 ? n233 : n27208;
  assign n27210 = pi17 ? n233 : n27209;
  assign n27211 = pi16 ? n26865 : n27210;
  assign n27212 = pi15 ? n27206 : n27211;
  assign n27213 = pi14 ? n27201 : n27212;
  assign n27214 = pi17 ? n26883 : n27209;
  assign n27215 = pi16 ? n26877 : n27214;
  assign n27216 = pi20 ? n26905 : n26898;
  assign n27217 = pi19 ? n26896 : n27216;
  assign n27218 = pi21 ? n363 : n10325;
  assign n27219 = pi20 ? n27218 : n32;
  assign n27220 = pi19 ? n27219 : n32;
  assign n27221 = pi18 ? n27217 : n27220;
  assign n27222 = pi17 ? n26895 : n27221;
  assign n27223 = pi16 ? n26887 : n27222;
  assign n27224 = pi15 ? n27215 : n27223;
  assign n27225 = pi21 ? n24222 : n2230;
  assign n27226 = pi20 ? n27225 : n32;
  assign n27227 = pi19 ? n27226 : n32;
  assign n27228 = pi18 ? n26907 : n27227;
  assign n27229 = pi17 ? n363 : n27228;
  assign n27230 = pi16 ? n21219 : n27229;
  assign n27231 = pi16 ? n21561 : n26919;
  assign n27232 = pi15 ? n27230 : n27231;
  assign n27233 = pi14 ? n27224 : n27232;
  assign n27234 = pi13 ? n27213 : n27233;
  assign n27235 = pi12 ? n27192 : n27234;
  assign n27236 = pi11 ? n27134 : n27235;
  assign n27237 = pi10 ? n27068 : n27236;
  assign n27238 = pi09 ? n26421 : n27237;
  assign n27239 = pi08 ? n26927 : n27238;
  assign n27240 = pi19 ? n1620 : n32;
  assign n27241 = pi18 ? n37 : n27240;
  assign n27242 = pi17 ? n37 : n27241;
  assign n27243 = pi16 ? n14445 : n27242;
  assign n27244 = pi15 ? n32 : n27243;
  assign n27245 = pi19 ? n37 : n16999;
  assign n27246 = pi20 ? n181 : n37;
  assign n27247 = pi19 ? n27246 : n3039;
  assign n27248 = pi18 ? n27245 : n27247;
  assign n27249 = pi20 ? n181 : n99;
  assign n27250 = pi19 ? n27249 : n99;
  assign n27251 = pi22 ? n99 : n3831;
  assign n27252 = pi21 ? n99 : n27251;
  assign n27253 = pi20 ? n99 : n27252;
  assign n27254 = pi19 ? n27253 : n32;
  assign n27255 = pi18 ? n27250 : n27254;
  assign n27256 = pi17 ? n27248 : n27255;
  assign n27257 = pi16 ? n14445 : n27256;
  assign n27258 = pi18 ? n99 : n27254;
  assign n27259 = pi17 ? n26411 : n27258;
  assign n27260 = pi16 ? n16595 : n27259;
  assign n27261 = pi15 ? n27257 : n27260;
  assign n27262 = pi14 ? n27244 : n27261;
  assign n27263 = pi13 ? n32 : n27262;
  assign n27264 = pi12 ? n32 : n27263;
  assign n27265 = pi11 ? n32 : n27264;
  assign n27266 = pi10 ? n32 : n27265;
  assign n27267 = pi20 ? n14844 : n37;
  assign n27268 = pi19 ? n27267 : n5077;
  assign n27269 = pi18 ? n23649 : n27268;
  assign n27270 = pi22 ? n99 : n18038;
  assign n27271 = pi21 ? n99 : n27270;
  assign n27272 = pi20 ? n99 : n27271;
  assign n27273 = pi19 ? n27272 : n32;
  assign n27274 = pi18 ? n26425 : n27273;
  assign n27275 = pi17 ? n27269 : n27274;
  assign n27276 = pi16 ? n16595 : n27275;
  assign n27277 = pi20 ? n7745 : n3039;
  assign n27278 = pi20 ? n2974 : n37;
  assign n27279 = pi19 ? n27277 : n27278;
  assign n27280 = pi22 ? n99 : n8174;
  assign n27281 = pi21 ? n99 : n27280;
  assign n27282 = pi20 ? n99 : n27281;
  assign n27283 = pi19 ? n27282 : n32;
  assign n27284 = pi18 ? n27279 : n27283;
  assign n27285 = pi17 ? n37 : n27284;
  assign n27286 = pi16 ? n17010 : n27285;
  assign n27287 = pi15 ? n27276 : n27286;
  assign n27288 = pi22 ? n37 : n8198;
  assign n27289 = pi21 ? n37 : n27288;
  assign n27290 = pi20 ? n14887 : n27289;
  assign n27291 = pi19 ? n27290 : n32;
  assign n27292 = pi18 ? n37 : n27291;
  assign n27293 = pi17 ? n37 : n27292;
  assign n27294 = pi16 ? n17010 : n27293;
  assign n27295 = pi22 ? n37 : n17574;
  assign n27296 = pi21 ? n37 : n27295;
  assign n27297 = pi20 ? n14887 : n27296;
  assign n27298 = pi19 ? n27297 : n32;
  assign n27299 = pi18 ? n37 : n27298;
  assign n27300 = pi17 ? n37 : n27299;
  assign n27301 = pi16 ? n439 : n27300;
  assign n27302 = pi15 ? n27294 : n27301;
  assign n27303 = pi14 ? n27287 : n27302;
  assign n27304 = pi16 ? n201 : n26939;
  assign n27305 = pi21 ? n180 : n112;
  assign n27306 = pi20 ? n32 : n27305;
  assign n27307 = pi19 ? n32 : n27306;
  assign n27308 = pi18 ? n27307 : n18854;
  assign n27309 = pi17 ? n32 : n27308;
  assign n27310 = pi16 ? n27309 : n26939;
  assign n27311 = pi15 ? n27304 : n27310;
  assign n27312 = pi18 ? n374 : n14115;
  assign n27313 = pi17 ? n32 : n27312;
  assign n27314 = pi16 ? n27313 : n26951;
  assign n27315 = pi20 ? n37 : n1719;
  assign n27316 = pi19 ? n27315 : n139;
  assign n27317 = pi18 ? n27316 : n139;
  assign n27318 = pi17 ? n27317 : n26950;
  assign n27319 = pi16 ? n439 : n27318;
  assign n27320 = pi15 ? n27314 : n27319;
  assign n27321 = pi14 ? n27311 : n27320;
  assign n27322 = pi13 ? n27303 : n27321;
  assign n27323 = pi20 ? n297 : n5273;
  assign n27324 = pi19 ? n9824 : n27323;
  assign n27325 = pi18 ? n37 : n27324;
  assign n27326 = pi20 ? n9348 : n139;
  assign n27327 = pi19 ? n3578 : n27326;
  assign n27328 = pi18 ? n27327 : n26949;
  assign n27329 = pi17 ? n27325 : n27328;
  assign n27330 = pi16 ? n439 : n27329;
  assign n27331 = pi20 ? n37 : n5273;
  assign n27332 = pi19 ? n37 : n27331;
  assign n27333 = pi18 ? n37 : n27332;
  assign n27334 = pi20 ? n139 : n3086;
  assign n27335 = pi19 ? n27334 : n26472;
  assign n27336 = pi18 ? n27335 : n26949;
  assign n27337 = pi17 ? n27333 : n27336;
  assign n27338 = pi16 ? n439 : n27337;
  assign n27339 = pi15 ? n27330 : n27338;
  assign n27340 = pi20 ? n139 : n13103;
  assign n27341 = pi19 ? n27340 : n32;
  assign n27342 = pi18 ? n16093 : n27341;
  assign n27343 = pi17 ? n19830 : n27342;
  assign n27344 = pi16 ? n439 : n27343;
  assign n27345 = pi21 ? n139 : n19522;
  assign n27346 = pi20 ? n26482 : n27345;
  assign n27347 = pi19 ? n27346 : n32;
  assign n27348 = pi18 ? n16093 : n27347;
  assign n27349 = pi17 ? n37 : n27348;
  assign n27350 = pi16 ? n439 : n27349;
  assign n27351 = pi15 ? n27344 : n27350;
  assign n27352 = pi14 ? n27339 : n27351;
  assign n27353 = pi21 ? n916 : n19522;
  assign n27354 = pi20 ? n922 : n27353;
  assign n27355 = pi19 ? n27354 : n32;
  assign n27356 = pi18 ? n16093 : n27355;
  assign n27357 = pi17 ? n37 : n27356;
  assign n27358 = pi16 ? n439 : n27357;
  assign n27359 = pi20 ? n204 : n22005;
  assign n27360 = pi19 ? n27359 : n32;
  assign n27361 = pi18 ? n26503 : n27360;
  assign n27362 = pi17 ? n37 : n27361;
  assign n27363 = pi16 ? n439 : n27362;
  assign n27364 = pi15 ? n27358 : n27363;
  assign n27365 = pi21 ? n204 : n516;
  assign n27366 = pi20 ? n27365 : n22005;
  assign n27367 = pi19 ? n27366 : n32;
  assign n27368 = pi18 ? n26503 : n27367;
  assign n27369 = pi17 ? n37 : n27368;
  assign n27370 = pi16 ? n439 : n27369;
  assign n27371 = pi21 ? n2091 : n3409;
  assign n27372 = pi21 ? n580 : n650;
  assign n27373 = pi20 ? n27371 : n27372;
  assign n27374 = pi19 ? n27373 : n32;
  assign n27375 = pi18 ? n37 : n27374;
  assign n27376 = pi17 ? n37 : n27375;
  assign n27377 = pi16 ? n439 : n27376;
  assign n27378 = pi15 ? n27370 : n27377;
  assign n27379 = pi14 ? n27364 : n27378;
  assign n27380 = pi13 ? n27352 : n27379;
  assign n27381 = pi12 ? n27322 : n27380;
  assign n27382 = pi21 ? n37 : n22332;
  assign n27383 = pi20 ? n2091 : n27382;
  assign n27384 = pi19 ? n27383 : n32;
  assign n27385 = pi18 ? n37 : n27384;
  assign n27386 = pi17 ? n37 : n27385;
  assign n27387 = pi16 ? n439 : n27386;
  assign n27388 = pi23 ? n37 : n19714;
  assign n27389 = pi22 ? n27388 : n625;
  assign n27390 = pi21 ? n335 : n27389;
  assign n27391 = pi20 ? n605 : n27390;
  assign n27392 = pi19 ? n27391 : n32;
  assign n27393 = pi18 ? n7686 : n27392;
  assign n27394 = pi17 ? n37 : n27393;
  assign n27395 = pi16 ? n439 : n27394;
  assign n27396 = pi15 ? n27387 : n27395;
  assign n27397 = pi24 ? n335 : n157;
  assign n27398 = pi23 ? n37 : n27397;
  assign n27399 = pi22 ? n27398 : n625;
  assign n27400 = pi21 ? n37 : n27399;
  assign n27401 = pi20 ? n647 : n27400;
  assign n27402 = pi19 ? n27401 : n32;
  assign n27403 = pi18 ? n37 : n27402;
  assign n27404 = pi17 ? n37 : n27403;
  assign n27405 = pi16 ? n439 : n27404;
  assign n27406 = pi22 ? n3935 : n625;
  assign n27407 = pi21 ? n335 : n27406;
  assign n27408 = pi20 ? n577 : n27407;
  assign n27409 = pi19 ? n27408 : n32;
  assign n27410 = pi18 ? n7677 : n27409;
  assign n27411 = pi17 ? n37 : n27410;
  assign n27412 = pi16 ? n439 : n27411;
  assign n27413 = pi15 ? n27405 : n27412;
  assign n27414 = pi14 ? n27396 : n27413;
  assign n27415 = pi22 ? n583 : n559;
  assign n27416 = pi21 ? n37 : n27415;
  assign n27417 = pi21 ? n6376 : n6983;
  assign n27418 = pi20 ? n27416 : n27417;
  assign n27419 = pi19 ? n27418 : n32;
  assign n27420 = pi18 ? n7686 : n27419;
  assign n27421 = pi17 ? n37 : n27420;
  assign n27422 = pi16 ? n439 : n27421;
  assign n27423 = pi20 ? n4954 : n13257;
  assign n27424 = pi19 ? n27423 : n32;
  assign n27425 = pi18 ? n24789 : n27424;
  assign n27426 = pi17 ? n37 : n27425;
  assign n27427 = pi16 ? n439 : n27426;
  assign n27428 = pi15 ? n27422 : n27427;
  assign n27429 = pi20 ? n575 : n13257;
  assign n27430 = pi19 ? n27429 : n32;
  assign n27431 = pi18 ? n17225 : n27430;
  assign n27432 = pi17 ? n37 : n27431;
  assign n27433 = pi16 ? n439 : n27432;
  assign n27434 = pi21 ? n2048 : n13280;
  assign n27435 = pi20 ? n37 : n27434;
  assign n27436 = pi19 ? n27435 : n32;
  assign n27437 = pi18 ? n2114 : n27436;
  assign n27438 = pi17 ? n37 : n27437;
  assign n27439 = pi16 ? n439 : n27438;
  assign n27440 = pi15 ? n27433 : n27439;
  assign n27441 = pi14 ? n27428 : n27440;
  assign n27442 = pi13 ? n27414 : n27441;
  assign n27443 = pi20 ? n37 : n15173;
  assign n27444 = pi19 ? n37 : n27443;
  assign n27445 = pi20 ? n37 : n23107;
  assign n27446 = pi19 ? n27445 : n32;
  assign n27447 = pi18 ? n27444 : n27446;
  assign n27448 = pi17 ? n37 : n27447;
  assign n27449 = pi16 ? n439 : n27448;
  assign n27450 = pi21 ? n6401 : n8486;
  assign n27451 = pi20 ? n37 : n27450;
  assign n27452 = pi19 ? n27451 : n32;
  assign n27453 = pi18 ? n37 : n27452;
  assign n27454 = pi17 ? n37 : n27453;
  assign n27455 = pi16 ? n439 : n27454;
  assign n27456 = pi15 ? n27449 : n27455;
  assign n27457 = pi21 ? n3073 : n8486;
  assign n27458 = pi20 ? n37 : n27457;
  assign n27459 = pi19 ? n27458 : n32;
  assign n27460 = pi18 ? n37 : n27459;
  assign n27461 = pi17 ? n37 : n27460;
  assign n27462 = pi16 ? n439 : n27461;
  assign n27463 = pi21 ? n3073 : n7723;
  assign n27464 = pi20 ? n37 : n27463;
  assign n27465 = pi19 ? n27464 : n32;
  assign n27466 = pi18 ? n37 : n27465;
  assign n27467 = pi17 ? n37 : n27466;
  assign n27468 = pi16 ? n439 : n27467;
  assign n27469 = pi15 ? n27462 : n27468;
  assign n27470 = pi14 ? n27456 : n27469;
  assign n27471 = pi21 ? n3392 : n2320;
  assign n27472 = pi20 ? n37 : n27471;
  assign n27473 = pi19 ? n27472 : n32;
  assign n27474 = pi18 ? n37 : n27473;
  assign n27475 = pi17 ? n37 : n27474;
  assign n27476 = pi16 ? n439 : n27475;
  assign n27477 = pi20 ? n8038 : n19091;
  assign n27478 = pi19 ? n15173 : n27477;
  assign n27479 = pi18 ? n374 : n27478;
  assign n27480 = pi17 ? n32 : n27479;
  assign n27481 = pi21 ? n7327 : n5015;
  assign n27482 = pi21 ? n10490 : n5015;
  assign n27483 = pi20 ? n27481 : n27482;
  assign n27484 = pi21 ? n7334 : n5015;
  assign n27485 = pi19 ? n27483 : n27484;
  assign n27486 = pi20 ? n27484 : n22881;
  assign n27487 = pi20 ? n9660 : n13310;
  assign n27488 = pi19 ? n27486 : n27487;
  assign n27489 = pi18 ? n27485 : n27488;
  assign n27490 = pi21 ? n7327 : n363;
  assign n27491 = pi20 ? n7730 : n27490;
  assign n27492 = pi19 ? n27491 : n37;
  assign n27493 = pi21 ? n3392 : n3125;
  assign n27494 = pi20 ? n37 : n27493;
  assign n27495 = pi19 ? n27494 : n32;
  assign n27496 = pi18 ? n27492 : n27495;
  assign n27497 = pi17 ? n27489 : n27496;
  assign n27498 = pi16 ? n27480 : n27497;
  assign n27499 = pi15 ? n27476 : n27498;
  assign n27500 = pi19 ? n23903 : n37;
  assign n27501 = pi21 ? n363 : n3392;
  assign n27502 = pi20 ? n3393 : n27501;
  assign n27503 = pi20 ? n22881 : n15173;
  assign n27504 = pi19 ? n27502 : n27503;
  assign n27505 = pi18 ? n27500 : n27504;
  assign n27506 = pi21 ? n5015 : n3392;
  assign n27507 = pi20 ? n363 : n27506;
  assign n27508 = pi19 ? n7730 : n27507;
  assign n27509 = pi21 ? n3392 : n9246;
  assign n27510 = pi20 ? n15173 : n27509;
  assign n27511 = pi19 ? n27510 : n32;
  assign n27512 = pi18 ? n27508 : n27511;
  assign n27513 = pi17 ? n27505 : n27512;
  assign n27514 = pi16 ? n439 : n27513;
  assign n27515 = pi19 ? n22878 : n37;
  assign n27516 = pi20 ? n3393 : n15173;
  assign n27517 = pi19 ? n27516 : n27503;
  assign n27518 = pi18 ? n27515 : n27517;
  assign n27519 = pi20 ? n7332 : n3393;
  assign n27520 = pi21 ? n5015 : n363;
  assign n27521 = pi20 ? n363 : n27520;
  assign n27522 = pi19 ? n27519 : n27521;
  assign n27523 = pi21 ? n363 : n9246;
  assign n27524 = pi20 ? n363 : n27523;
  assign n27525 = pi19 ? n27524 : n32;
  assign n27526 = pi18 ? n27522 : n27525;
  assign n27527 = pi17 ? n27518 : n27526;
  assign n27528 = pi16 ? n439 : n27527;
  assign n27529 = pi15 ? n27514 : n27528;
  assign n27530 = pi14 ? n27499 : n27529;
  assign n27531 = pi13 ? n27470 : n27530;
  assign n27532 = pi12 ? n27442 : n27531;
  assign n27533 = pi11 ? n27381 : n27532;
  assign n27534 = pi21 ? n2106 : n19958;
  assign n27535 = pi20 ? n37 : n27534;
  assign n27536 = pi19 ? n37 : n27535;
  assign n27537 = pi21 ? n214 : n2637;
  assign n27538 = pi20 ? n37 : n27537;
  assign n27539 = pi19 ? n27538 : n32;
  assign n27540 = pi18 ? n27536 : n27539;
  assign n27541 = pi17 ? n37 : n27540;
  assign n27542 = pi16 ? n439 : n27541;
  assign n27543 = pi22 ? n24834 : n37;
  assign n27544 = pi21 ? n27543 : n37;
  assign n27545 = pi20 ? n27544 : n27076;
  assign n27546 = pi19 ? n27545 : n32;
  assign n27547 = pi18 ? n18193 : n27546;
  assign n27548 = pi17 ? n37 : n27547;
  assign n27549 = pi16 ? n439 : n27548;
  assign n27550 = pi15 ? n27542 : n27549;
  assign n27551 = pi21 ? n6461 : n685;
  assign n27552 = pi20 ? n278 : n27551;
  assign n27553 = pi19 ? n37 : n27552;
  assign n27554 = pi22 ? n7780 : n157;
  assign n27555 = pi21 ? n27554 : n157;
  assign n27556 = pi20 ? n27555 : n27076;
  assign n27557 = pi19 ? n27556 : n32;
  assign n27558 = pi18 ? n27553 : n27557;
  assign n27559 = pi17 ? n37 : n27558;
  assign n27560 = pi16 ? n439 : n27559;
  assign n27561 = pi20 ? n278 : n157;
  assign n27562 = pi19 ? n37 : n27561;
  assign n27563 = pi22 ? n5452 : n2244;
  assign n27564 = pi21 ? n157 : n27563;
  assign n27565 = pi21 ? n20460 : n2637;
  assign n27566 = pi20 ? n27564 : n27565;
  assign n27567 = pi19 ? n27566 : n32;
  assign n27568 = pi18 ? n27562 : n27567;
  assign n27569 = pi17 ? n37 : n27568;
  assign n27570 = pi16 ? n439 : n27569;
  assign n27571 = pi15 ? n27560 : n27570;
  assign n27572 = pi14 ? n27550 : n27571;
  assign n27573 = pi20 ? n2238 : n27095;
  assign n27574 = pi19 ? n27573 : n32;
  assign n27575 = pi18 ? n26658 : n27574;
  assign n27576 = pi17 ? n99 : n27575;
  assign n27577 = pi16 ? n744 : n27576;
  assign n27578 = pi20 ? n99 : n13948;
  assign n27579 = pi19 ? n99 : n27578;
  assign n27580 = pi18 ? n27579 : n27097;
  assign n27581 = pi17 ? n99 : n27580;
  assign n27582 = pi16 ? n744 : n27581;
  assign n27583 = pi15 ? n27577 : n27582;
  assign n27584 = pi20 ? n99 : n7438;
  assign n27585 = pi19 ? n27584 : n32;
  assign n27586 = pi18 ? n27579 : n27585;
  assign n27587 = pi17 ? n99 : n27586;
  assign n27588 = pi16 ? n744 : n27587;
  assign n27589 = pi15 ? n27107 : n27588;
  assign n27590 = pi14 ? n27583 : n27589;
  assign n27591 = pi13 ? n27572 : n27590;
  assign n27592 = pi19 ? n139 : n19134;
  assign n27593 = pi18 ? n27592 : n27113;
  assign n27594 = pi17 ? n26684 : n27593;
  assign n27595 = pi16 ? n25417 : n27594;
  assign n27596 = pi20 ? n99 : n22965;
  assign n27597 = pi19 ? n139 : n27596;
  assign n27598 = pi21 ? n20977 : n99;
  assign n27599 = pi20 ? n27598 : n16506;
  assign n27600 = pi19 ? n27599 : n32;
  assign n27601 = pi18 ? n27597 : n27600;
  assign n27602 = pi17 ? n26684 : n27601;
  assign n27603 = pi16 ? n25417 : n27602;
  assign n27604 = pi15 ? n27595 : n27603;
  assign n27605 = pi20 ? n975 : n204;
  assign n27606 = pi19 ? n139 : n27605;
  assign n27607 = pi20 ? n1027 : n16506;
  assign n27608 = pi19 ? n27607 : n32;
  assign n27609 = pi18 ? n27606 : n27608;
  assign n27610 = pi17 ? n139 : n27609;
  assign n27611 = pi16 ? n915 : n27610;
  assign n27612 = pi20 ? n316 : n16506;
  assign n27613 = pi19 ? n27612 : n32;
  assign n27614 = pi18 ? n17418 : n27613;
  assign n27615 = pi17 ? n139 : n27614;
  assign n27616 = pi16 ? n1773 : n27615;
  assign n27617 = pi15 ? n27611 : n27616;
  assign n27618 = pi14 ? n27604 : n27617;
  assign n27619 = pi21 ? n391 : n204;
  assign n27620 = pi20 ? n204 : n27619;
  assign n27621 = pi19 ? n27620 : n204;
  assign n27622 = pi20 ? n204 : n7900;
  assign n27623 = pi21 ? n3258 : n204;
  assign n27624 = pi21 ? n381 : n204;
  assign n27625 = pi20 ? n27623 : n27624;
  assign n27626 = pi19 ? n27622 : n27625;
  assign n27627 = pi18 ? n27621 : n27626;
  assign n27628 = pi19 ? n24023 : n316;
  assign n27629 = pi20 ? n316 : n6935;
  assign n27630 = pi19 ? n27629 : n32;
  assign n27631 = pi18 ? n27628 : n27630;
  assign n27632 = pi17 ? n27627 : n27631;
  assign n27633 = pi16 ? n11804 : n27632;
  assign n27634 = pi20 ? n7858 : n316;
  assign n27635 = pi19 ? n204 : n27634;
  assign n27636 = pi18 ? n27635 : n27630;
  assign n27637 = pi17 ? n204 : n27636;
  assign n27638 = pi16 ? n24565 : n27637;
  assign n27639 = pi15 ? n27633 : n27638;
  assign n27640 = pi19 ? n204 : n22775;
  assign n27641 = pi18 ? n204 : n27640;
  assign n27642 = pi20 ? n5204 : n1016;
  assign n27643 = pi19 ? n204 : n27642;
  assign n27644 = pi20 ? n6158 : n10335;
  assign n27645 = pi19 ? n27644 : n32;
  assign n27646 = pi18 ? n27643 : n27645;
  assign n27647 = pi17 ? n27641 : n27646;
  assign n27648 = pi16 ? n13493 : n27647;
  assign n27649 = pi18 ? n15397 : n204;
  assign n27650 = pi17 ? n32 : n27649;
  assign n27651 = pi20 ? n3086 : n204;
  assign n27652 = pi19 ? n204 : n27651;
  assign n27653 = pi18 ? n204 : n27652;
  assign n27654 = pi22 ? n4883 : n317;
  assign n27655 = pi21 ? n27654 : n32;
  assign n27656 = pi20 ? n204 : n27655;
  assign n27657 = pi19 ? n27656 : n32;
  assign n27658 = pi18 ? n26743 : n27657;
  assign n27659 = pi17 ? n27653 : n27658;
  assign n27660 = pi16 ? n27650 : n27659;
  assign n27661 = pi15 ? n27648 : n27660;
  assign n27662 = pi14 ? n27639 : n27661;
  assign n27663 = pi13 ? n27618 : n27662;
  assign n27664 = pi12 ? n27591 : n27663;
  assign n27665 = pi20 ? n1016 : n921;
  assign n27666 = pi19 ? n139 : n27665;
  assign n27667 = pi23 ? n204 : n4145;
  assign n27668 = pi22 ? n27667 : n317;
  assign n27669 = pi21 ? n27668 : n32;
  assign n27670 = pi20 ? n6158 : n27669;
  assign n27671 = pi19 ? n27670 : n32;
  assign n27672 = pi18 ? n27666 : n27671;
  assign n27673 = pi17 ? n139 : n27672;
  assign n27674 = pi16 ? n915 : n27673;
  assign n27675 = pi21 ? n9186 : n32;
  assign n27676 = pi20 ? n1016 : n27675;
  assign n27677 = pi19 ? n27676 : n32;
  assign n27678 = pi18 ? n23054 : n27677;
  assign n27679 = pi17 ? n139 : n27678;
  assign n27680 = pi16 ? n915 : n27679;
  assign n27681 = pi15 ? n27674 : n27680;
  assign n27682 = pi19 ? n638 : n6373;
  assign n27683 = pi18 ? n602 : n27682;
  assign n27684 = pi17 ? n32 : n27683;
  assign n27685 = pi20 ? n577 : n604;
  assign n27686 = pi19 ? n27685 : n604;
  assign n27687 = pi20 ? n577 : n605;
  assign n27688 = pi19 ? n335 : n27687;
  assign n27689 = pi18 ? n27686 : n27688;
  assign n27690 = pi20 ? n1089 : n2405;
  assign n27691 = pi19 ? n335 : n27690;
  assign n27692 = pi23 ? n204 : n2766;
  assign n27693 = pi22 ? n27692 : n32;
  assign n27694 = pi21 ? n27693 : n32;
  assign n27695 = pi20 ? n204 : n27694;
  assign n27696 = pi19 ? n27695 : n32;
  assign n27697 = pi18 ? n27691 : n27696;
  assign n27698 = pi17 ? n27689 : n27697;
  assign n27699 = pi16 ? n27684 : n27698;
  assign n27700 = pi18 ? n602 : n26795;
  assign n27701 = pi17 ? n32 : n27700;
  assign n27702 = pi20 ? n13527 : n4102;
  assign n27703 = pi19 ? n27702 : n32;
  assign n27704 = pi18 ? n17534 : n27703;
  assign n27705 = pi17 ? n335 : n27704;
  assign n27706 = pi16 ? n27701 : n27705;
  assign n27707 = pi15 ? n27699 : n27706;
  assign n27708 = pi14 ? n27681 : n27707;
  assign n27709 = pi18 ? n17540 : n19048;
  assign n27710 = pi17 ? n335 : n27709;
  assign n27711 = pi16 ? n7943 : n27710;
  assign n27712 = pi20 ? n16544 : n2579;
  assign n27713 = pi19 ? n27712 : n32;
  assign n27714 = pi18 ? n17540 : n27713;
  assign n27715 = pi17 ? n335 : n27714;
  assign n27716 = pi16 ? n7943 : n27715;
  assign n27717 = pi15 ? n27711 : n27716;
  assign n27718 = pi20 ? n233 : n2638;
  assign n27719 = pi19 ? n27718 : n32;
  assign n27720 = pi18 ? n26820 : n27719;
  assign n27721 = pi17 ? n26818 : n27720;
  assign n27722 = pi16 ? n439 : n27721;
  assign n27723 = pi18 ? n9556 : n27682;
  assign n27724 = pi17 ? n32 : n27723;
  assign n27725 = pi19 ? n17495 : n649;
  assign n27726 = pi20 ? n639 : n581;
  assign n27727 = pi20 ? n649 : n642;
  assign n27728 = pi19 ? n27726 : n27727;
  assign n27729 = pi18 ? n27725 : n27728;
  assign n27730 = pi21 ? n570 : n574;
  assign n27731 = pi20 ? n27730 : n335;
  assign n27732 = pi19 ? n27731 : n233;
  assign n27733 = pi18 ? n27732 : n27719;
  assign n27734 = pi17 ? n27729 : n27733;
  assign n27735 = pi16 ? n27724 : n27734;
  assign n27736 = pi15 ? n27722 : n27735;
  assign n27737 = pi14 ? n27717 : n27736;
  assign n27738 = pi13 ? n27708 : n27737;
  assign n27739 = pi24 ? n32 : n233;
  assign n27740 = pi23 ? n27739 : n37;
  assign n27741 = pi22 ? n27740 : n233;
  assign n27742 = pi21 ? n27741 : n233;
  assign n27743 = pi20 ? n32 : n27742;
  assign n27744 = pi19 ? n32 : n27743;
  assign n27745 = pi18 ? n27744 : n26838;
  assign n27746 = pi17 ? n32 : n27745;
  assign n27747 = pi21 ? n6361 : n2061;
  assign n27748 = pi20 ? n27747 : n233;
  assign n27749 = pi19 ? n233 : n27748;
  assign n27750 = pi18 ? n233 : n27749;
  assign n27751 = pi18 ? n233 : n26338;
  assign n27752 = pi17 ? n27750 : n27751;
  assign n27753 = pi16 ? n27746 : n27752;
  assign n27754 = pi20 ? n2094 : n37;
  assign n27755 = pi19 ? n27754 : n37;
  assign n27756 = pi18 ? n37 : n27755;
  assign n27757 = pi18 ? n18113 : n26338;
  assign n27758 = pi17 ? n27756 : n27757;
  assign n27759 = pi16 ? n439 : n27758;
  assign n27760 = pi15 ? n27753 : n27759;
  assign n27761 = pi17 ? n27756 : n27204;
  assign n27762 = pi16 ? n439 : n27761;
  assign n27763 = pi21 ? n233 : n22128;
  assign n27764 = pi20 ? n233 : n27763;
  assign n27765 = pi20 ? n99 : n233;
  assign n27766 = pi19 ? n27764 : n27765;
  assign n27767 = pi18 ? n26016 : n27766;
  assign n27768 = pi17 ? n32 : n27767;
  assign n27769 = pi16 ? n27768 : n27210;
  assign n27770 = pi15 ? n27762 : n27769;
  assign n27771 = pi14 ? n27760 : n27770;
  assign n27772 = pi22 ? n673 : n99;
  assign n27773 = pi21 ? n25162 : n27772;
  assign n27774 = pi20 ? n32 : n27773;
  assign n27775 = pi19 ? n32 : n27774;
  assign n27776 = pi21 ? n722 : n233;
  assign n27777 = pi20 ? n363 : n27776;
  assign n27778 = pi19 ? n20860 : n27777;
  assign n27779 = pi18 ? n27775 : n27778;
  assign n27780 = pi17 ? n32 : n27779;
  assign n27781 = pi21 ? n233 : n722;
  assign n27782 = pi20 ? n27776 : n27781;
  assign n27783 = pi19 ? n27782 : n27781;
  assign n27784 = pi21 ? n233 : n19920;
  assign n27785 = pi21 ? n23186 : n233;
  assign n27786 = pi20 ? n27784 : n27785;
  assign n27787 = pi21 ? n99 : n2707;
  assign n27788 = pi20 ? n27787 : n26880;
  assign n27789 = pi19 ? n27786 : n27788;
  assign n27790 = pi18 ? n27783 : n27789;
  assign n27791 = pi20 ? n19921 : n15177;
  assign n27792 = pi19 ? n27791 : n233;
  assign n27793 = pi18 ? n27792 : n27208;
  assign n27794 = pi17 ? n27790 : n27793;
  assign n27795 = pi16 ? n27780 : n27794;
  assign n27796 = pi21 ? n363 : n24215;
  assign n27797 = pi20 ? n27796 : n363;
  assign n27798 = pi19 ? n27797 : n363;
  assign n27799 = pi18 ? n363 : n27798;
  assign n27800 = pi20 ? n363 : n26898;
  assign n27801 = pi18 ? n27800 : n27220;
  assign n27802 = pi17 ? n27799 : n27801;
  assign n27803 = pi16 ? n21219 : n27802;
  assign n27804 = pi15 ? n27795 : n27803;
  assign n27805 = pi21 ? n2721 : n2230;
  assign n27806 = pi20 ? n27805 : n32;
  assign n27807 = pi19 ? n27806 : n32;
  assign n27808 = pi18 ? n26907 : n27807;
  assign n27809 = pi17 ? n363 : n27808;
  assign n27810 = pi16 ? n21219 : n27809;
  assign n27811 = pi20 ? n19084 : n363;
  assign n27812 = pi19 ? n363 : n27811;
  assign n27813 = pi22 ? n363 : n15186;
  assign n27814 = pi21 ? n27813 : n3523;
  assign n27815 = pi20 ? n27814 : n32;
  assign n27816 = pi19 ? n27815 : n32;
  assign n27817 = pi18 ? n27812 : n27816;
  assign n27818 = pi17 ? n363 : n27817;
  assign n27819 = pi16 ? n26062 : n27818;
  assign n27820 = pi15 ? n27810 : n27819;
  assign n27821 = pi14 ? n27804 : n27820;
  assign n27822 = pi13 ? n27771 : n27821;
  assign n27823 = pi12 ? n27738 : n27822;
  assign n27824 = pi11 ? n27664 : n27823;
  assign n27825 = pi10 ? n27533 : n27824;
  assign n27826 = pi09 ? n27266 : n27825;
  assign n27827 = pi20 ? n14887 : n13050;
  assign n27828 = pi19 ? n27827 : n32;
  assign n27829 = pi18 ? n37 : n27828;
  assign n27830 = pi17 ? n37 : n27829;
  assign n27831 = pi16 ? n439 : n27830;
  assign n27832 = pi15 ? n27294 : n27831;
  assign n27833 = pi14 ? n27287 : n27832;
  assign n27834 = pi20 ? n99 : n13577;
  assign n27835 = pi19 ? n27834 : n32;
  assign n27836 = pi18 ? n99 : n27835;
  assign n27837 = pi17 ? n99 : n27836;
  assign n27838 = pi16 ? n201 : n27837;
  assign n27839 = pi15 ? n27838 : n27310;
  assign n27840 = pi21 ? n139 : n21725;
  assign n27841 = pi20 ? n139 : n27840;
  assign n27842 = pi19 ? n27841 : n32;
  assign n27843 = pi18 ? n139 : n27842;
  assign n27844 = pi17 ? n139 : n27843;
  assign n27845 = pi16 ? n27313 : n27844;
  assign n27846 = pi17 ? n27317 : n27843;
  assign n27847 = pi16 ? n439 : n27846;
  assign n27848 = pi15 ? n27845 : n27847;
  assign n27849 = pi14 ? n27839 : n27848;
  assign n27850 = pi13 ? n27833 : n27849;
  assign n27851 = pi19 ? n1220 : n32;
  assign n27852 = pi18 ? n27327 : n27851;
  assign n27853 = pi17 ? n27325 : n27852;
  assign n27854 = pi16 ? n439 : n27853;
  assign n27855 = pi22 ? n139 : n3301;
  assign n27856 = pi21 ? n139 : n27855;
  assign n27857 = pi20 ? n139 : n27856;
  assign n27858 = pi19 ? n27857 : n32;
  assign n27859 = pi18 ? n27335 : n27858;
  assign n27860 = pi17 ? n27333 : n27859;
  assign n27861 = pi16 ? n439 : n27860;
  assign n27862 = pi15 ? n27854 : n27861;
  assign n27863 = pi20 ? n139 : n13603;
  assign n27864 = pi19 ? n27863 : n32;
  assign n27865 = pi18 ? n16093 : n27864;
  assign n27866 = pi17 ? n19830 : n27865;
  assign n27867 = pi16 ? n439 : n27866;
  assign n27868 = pi22 ? n139 : n759;
  assign n27869 = pi21 ? n139 : n27868;
  assign n27870 = pi20 ? n26482 : n27869;
  assign n27871 = pi19 ? n27870 : n32;
  assign n27872 = pi18 ? n16093 : n27871;
  assign n27873 = pi17 ? n37 : n27872;
  assign n27874 = pi16 ? n439 : n27873;
  assign n27875 = pi15 ? n27867 : n27874;
  assign n27876 = pi14 ? n27862 : n27875;
  assign n27877 = pi21 ? n916 : n27868;
  assign n27878 = pi20 ? n922 : n27877;
  assign n27879 = pi19 ? n27878 : n32;
  assign n27880 = pi18 ? n16093 : n27879;
  assign n27881 = pi17 ? n37 : n27880;
  assign n27882 = pi16 ? n439 : n27881;
  assign n27883 = pi20 ? n204 : n21474;
  assign n27884 = pi19 ? n27883 : n32;
  assign n27885 = pi18 ? n26503 : n27884;
  assign n27886 = pi17 ? n37 : n27885;
  assign n27887 = pi16 ? n439 : n27886;
  assign n27888 = pi15 ? n27882 : n27887;
  assign n27889 = pi20 ? n27365 : n21474;
  assign n27890 = pi19 ? n27889 : n32;
  assign n27891 = pi18 ? n26503 : n27890;
  assign n27892 = pi17 ? n37 : n27891;
  assign n27893 = pi16 ? n439 : n27892;
  assign n27894 = pi21 ? n580 : n665;
  assign n27895 = pi20 ? n27371 : n27894;
  assign n27896 = pi19 ? n27895 : n32;
  assign n27897 = pi18 ? n37 : n27896;
  assign n27898 = pi17 ? n37 : n27897;
  assign n27899 = pi16 ? n439 : n27898;
  assign n27900 = pi15 ? n27893 : n27899;
  assign n27901 = pi14 ? n27888 : n27900;
  assign n27902 = pi13 ? n27876 : n27901;
  assign n27903 = pi12 ? n27850 : n27902;
  assign n27904 = pi20 ? n2091 : n1409;
  assign n27905 = pi19 ? n27904 : n32;
  assign n27906 = pi18 ? n37 : n27905;
  assign n27907 = pi17 ? n37 : n27906;
  assign n27908 = pi16 ? n439 : n27907;
  assign n27909 = pi22 ? n583 : n317;
  assign n27910 = pi21 ? n335 : n27909;
  assign n27911 = pi20 ? n605 : n27910;
  assign n27912 = pi19 ? n27911 : n32;
  assign n27913 = pi18 ? n7686 : n27912;
  assign n27914 = pi17 ? n37 : n27913;
  assign n27915 = pi16 ? n439 : n27914;
  assign n27916 = pi15 ? n27908 : n27915;
  assign n27917 = pi22 ? n583 : n2468;
  assign n27918 = pi21 ? n37 : n27917;
  assign n27919 = pi20 ? n647 : n27918;
  assign n27920 = pi19 ? n27919 : n32;
  assign n27921 = pi18 ? n37 : n27920;
  assign n27922 = pi17 ? n37 : n27921;
  assign n27923 = pi16 ? n439 : n27922;
  assign n27924 = pi22 ? n3935 : n2468;
  assign n27925 = pi21 ? n335 : n27924;
  assign n27926 = pi20 ? n577 : n27925;
  assign n27927 = pi19 ? n27926 : n32;
  assign n27928 = pi18 ? n7677 : n27927;
  assign n27929 = pi17 ? n37 : n27928;
  assign n27930 = pi16 ? n439 : n27929;
  assign n27931 = pi15 ? n27923 : n27930;
  assign n27932 = pi14 ? n27916 : n27931;
  assign n27933 = pi20 ? n561 : n27434;
  assign n27934 = pi19 ? n27933 : n32;
  assign n27935 = pi18 ? n2114 : n27934;
  assign n27936 = pi17 ? n37 : n27935;
  assign n27937 = pi16 ? n439 : n27936;
  assign n27938 = pi15 ? n27433 : n27937;
  assign n27939 = pi14 ? n27428 : n27938;
  assign n27940 = pi13 ? n27932 : n27939;
  assign n27941 = pi21 ? n20629 : n8486;
  assign n27942 = pi20 ? n37 : n27941;
  assign n27943 = pi19 ? n27942 : n32;
  assign n27944 = pi18 ? n37 : n27943;
  assign n27945 = pi17 ? n37 : n27944;
  assign n27946 = pi16 ? n439 : n27945;
  assign n27947 = pi21 ? n7025 : n7723;
  assign n27948 = pi20 ? n37 : n27947;
  assign n27949 = pi19 ? n27948 : n32;
  assign n27950 = pi18 ? n37 : n27949;
  assign n27951 = pi17 ? n37 : n27950;
  assign n27952 = pi16 ? n439 : n27951;
  assign n27953 = pi15 ? n27946 : n27952;
  assign n27954 = pi14 ? n27456 : n27953;
  assign n27955 = pi21 ? n3392 : n7327;
  assign n27956 = pi20 ? n15173 : n27955;
  assign n27957 = pi19 ? n27956 : n27477;
  assign n27958 = pi18 ? n374 : n27957;
  assign n27959 = pi17 ? n32 : n27958;
  assign n27960 = pi21 ? n7326 : n5015;
  assign n27961 = pi20 ? n27960 : n27482;
  assign n27962 = pi21 ? n8567 : n5015;
  assign n27963 = pi19 ? n27961 : n27962;
  assign n27964 = pi20 ? n27962 : n22881;
  assign n27965 = pi21 ? n5015 : n6401;
  assign n27966 = pi20 ? n27965 : n8568;
  assign n27967 = pi19 ? n27964 : n27966;
  assign n27968 = pi18 ? n27963 : n27967;
  assign n27969 = pi19 ? n27490 : n37;
  assign n27970 = pi21 ? n3392 : n20889;
  assign n27971 = pi20 ? n37 : n27970;
  assign n27972 = pi19 ? n27971 : n32;
  assign n27973 = pi18 ? n27969 : n27972;
  assign n27974 = pi17 ? n27968 : n27973;
  assign n27975 = pi16 ? n27959 : n27974;
  assign n27976 = pi15 ? n27476 : n27975;
  assign n27977 = pi21 ? n3392 : n1512;
  assign n27978 = pi20 ? n15173 : n27977;
  assign n27979 = pi19 ? n27978 : n32;
  assign n27980 = pi18 ? n27508 : n27979;
  assign n27981 = pi17 ? n27505 : n27980;
  assign n27982 = pi16 ? n439 : n27981;
  assign n27983 = pi21 ? n363 : n1512;
  assign n27984 = pi20 ? n363 : n27983;
  assign n27985 = pi19 ? n27984 : n32;
  assign n27986 = pi18 ? n27522 : n27985;
  assign n27987 = pi17 ? n27518 : n27986;
  assign n27988 = pi16 ? n439 : n27987;
  assign n27989 = pi15 ? n27982 : n27988;
  assign n27990 = pi14 ? n27976 : n27989;
  assign n27991 = pi13 ? n27954 : n27990;
  assign n27992 = pi12 ? n27940 : n27991;
  assign n27993 = pi11 ? n27903 : n27992;
  assign n27994 = pi23 ? n20627 : n157;
  assign n27995 = pi22 ? n37 : n27994;
  assign n27996 = pi21 ? n27995 : n760;
  assign n27997 = pi20 ? n37 : n27996;
  assign n27998 = pi19 ? n27997 : n32;
  assign n27999 = pi18 ? n27536 : n27998;
  assign n28000 = pi17 ? n37 : n27999;
  assign n28001 = pi16 ? n439 : n28000;
  assign n28002 = pi21 ? n685 : n760;
  assign n28003 = pi20 ? n27544 : n28002;
  assign n28004 = pi19 ? n28003 : n32;
  assign n28005 = pi18 ? n18193 : n28004;
  assign n28006 = pi17 ? n37 : n28005;
  assign n28007 = pi16 ? n439 : n28006;
  assign n28008 = pi15 ? n28001 : n28007;
  assign n28009 = pi20 ? n27555 : n28002;
  assign n28010 = pi19 ? n28009 : n32;
  assign n28011 = pi18 ? n27553 : n28010;
  assign n28012 = pi17 ? n37 : n28011;
  assign n28013 = pi16 ? n439 : n28012;
  assign n28014 = pi22 ? n112 : n164;
  assign n28015 = pi21 ? n157 : n28014;
  assign n28016 = pi21 ? n20460 : n5829;
  assign n28017 = pi20 ? n28015 : n28016;
  assign n28018 = pi19 ? n28017 : n32;
  assign n28019 = pi18 ? n27562 : n28018;
  assign n28020 = pi17 ? n37 : n28019;
  assign n28021 = pi16 ? n439 : n28020;
  assign n28022 = pi15 ? n28013 : n28021;
  assign n28023 = pi14 ? n28008 : n28022;
  assign n28024 = pi21 ? n3562 : n882;
  assign n28025 = pi20 ? n2238 : n28024;
  assign n28026 = pi19 ? n28025 : n32;
  assign n28027 = pi18 ? n26658 : n28026;
  assign n28028 = pi17 ? n99 : n28027;
  assign n28029 = pi16 ? n721 : n28028;
  assign n28030 = pi16 ? n721 : n27581;
  assign n28031 = pi15 ? n28029 : n28030;
  assign n28032 = pi16 ? n721 : n27106;
  assign n28033 = pi21 ? n6132 : n928;
  assign n28034 = pi20 ? n99 : n28033;
  assign n28035 = pi19 ? n28034 : n32;
  assign n28036 = pi18 ? n27579 : n28035;
  assign n28037 = pi17 ? n99 : n28036;
  assign n28038 = pi16 ? n721 : n28037;
  assign n28039 = pi15 ? n28032 : n28038;
  assign n28040 = pi14 ? n28031 : n28039;
  assign n28041 = pi13 ? n28023 : n28040;
  assign n28042 = pi20 ? n157 : n7438;
  assign n28043 = pi19 ? n28042 : n32;
  assign n28044 = pi18 ? n27592 : n28043;
  assign n28045 = pi17 ? n26684 : n28044;
  assign n28046 = pi16 ? n24953 : n28045;
  assign n28047 = pi20 ? n27598 : n16476;
  assign n28048 = pi19 ? n28047 : n32;
  assign n28049 = pi18 ? n27597 : n28048;
  assign n28050 = pi17 ? n26684 : n28049;
  assign n28051 = pi16 ? n24953 : n28050;
  assign n28052 = pi15 ? n28046 : n28051;
  assign n28053 = pi20 ? n1027 : n7622;
  assign n28054 = pi19 ? n28053 : n32;
  assign n28055 = pi18 ? n27606 : n28054;
  assign n28056 = pi17 ? n139 : n28055;
  assign n28057 = pi16 ? n2291 : n28056;
  assign n28058 = pi15 ? n28057 : n27616;
  assign n28059 = pi14 ? n28052 : n28058;
  assign n28060 = pi16 ? n13493 : n27637;
  assign n28061 = pi15 ? n27633 : n28060;
  assign n28062 = pi21 ? n21980 : n32;
  assign n28063 = pi20 ? n6158 : n28062;
  assign n28064 = pi19 ? n28063 : n32;
  assign n28065 = pi18 ? n27643 : n28064;
  assign n28066 = pi17 ? n27641 : n28065;
  assign n28067 = pi16 ? n13493 : n28066;
  assign n28068 = pi22 ? n4079 : n2192;
  assign n28069 = pi21 ? n28068 : n32;
  assign n28070 = pi20 ? n204 : n28069;
  assign n28071 = pi19 ? n28070 : n32;
  assign n28072 = pi18 ? n26743 : n28071;
  assign n28073 = pi17 ? n27653 : n28072;
  assign n28074 = pi16 ? n27650 : n28073;
  assign n28075 = pi15 ? n28067 : n28074;
  assign n28076 = pi14 ? n28061 : n28075;
  assign n28077 = pi13 ? n28059 : n28076;
  assign n28078 = pi12 ? n28041 : n28077;
  assign n28079 = pi20 ? n6158 : n28069;
  assign n28080 = pi19 ? n28079 : n32;
  assign n28081 = pi18 ? n27666 : n28080;
  assign n28082 = pi17 ? n139 : n28081;
  assign n28083 = pi16 ? n2291 : n28082;
  assign n28084 = pi21 ? n20524 : n32;
  assign n28085 = pi20 ? n1016 : n28084;
  assign n28086 = pi19 ? n28085 : n32;
  assign n28087 = pi18 ? n23054 : n28086;
  assign n28088 = pi17 ? n139 : n28087;
  assign n28089 = pi16 ? n2291 : n28088;
  assign n28090 = pi15 ? n28083 : n28089;
  assign n28091 = pi18 ? n10397 : n27682;
  assign n28092 = pi17 ? n32 : n28091;
  assign n28093 = pi20 ? n204 : n27675;
  assign n28094 = pi19 ? n28093 : n32;
  assign n28095 = pi18 ? n27691 : n28094;
  assign n28096 = pi17 ? n27689 : n28095;
  assign n28097 = pi16 ? n28092 : n28096;
  assign n28098 = pi18 ? n10397 : n26795;
  assign n28099 = pi17 ? n32 : n28098;
  assign n28100 = pi16 ? n28099 : n27705;
  assign n28101 = pi15 ? n28097 : n28100;
  assign n28102 = pi14 ? n28090 : n28101;
  assign n28103 = pi18 ? n17540 : n19584;
  assign n28104 = pi17 ? n335 : n28103;
  assign n28105 = pi16 ? n2425 : n28104;
  assign n28106 = pi20 ? n16544 : n3340;
  assign n28107 = pi19 ? n28106 : n32;
  assign n28108 = pi18 ? n17540 : n28107;
  assign n28109 = pi17 ? n335 : n28108;
  assign n28110 = pi16 ? n7943 : n28109;
  assign n28111 = pi15 ? n28105 : n28110;
  assign n28112 = pi14 ? n28111 : n27736;
  assign n28113 = pi13 ? n28102 : n28112;
  assign n28114 = pi16 ? n27194 : n27752;
  assign n28115 = pi15 ? n28114 : n27759;
  assign n28116 = pi20 ? n25965 : n2653;
  assign n28117 = pi19 ? n28116 : n32;
  assign n28118 = pi18 ? n18113 : n28117;
  assign n28119 = pi17 ? n27756 : n28118;
  assign n28120 = pi16 ? n439 : n28119;
  assign n28121 = pi20 ? n25978 : n2653;
  assign n28122 = pi19 ? n28121 : n32;
  assign n28123 = pi18 ? n233 : n28122;
  assign n28124 = pi17 ? n233 : n28123;
  assign n28125 = pi16 ? n27768 : n28124;
  assign n28126 = pi15 ? n28120 : n28125;
  assign n28127 = pi14 ? n28115 : n28126;
  assign n28128 = pi21 ? n363 : n3445;
  assign n28129 = pi20 ? n28128 : n32;
  assign n28130 = pi19 ? n28129 : n32;
  assign n28131 = pi18 ? n27800 : n28130;
  assign n28132 = pi17 ? n27799 : n28131;
  assign n28133 = pi16 ? n21219 : n28132;
  assign n28134 = pi15 ? n27795 : n28133;
  assign n28135 = pi21 ? n2721 : n10325;
  assign n28136 = pi20 ? n28135 : n32;
  assign n28137 = pi19 ? n28136 : n32;
  assign n28138 = pi18 ? n26907 : n28137;
  assign n28139 = pi17 ? n363 : n28138;
  assign n28140 = pi16 ? n21219 : n28139;
  assign n28141 = pi21 ? n27813 : n5178;
  assign n28142 = pi20 ? n28141 : n32;
  assign n28143 = pi19 ? n28142 : n32;
  assign n28144 = pi18 ? n27812 : n28143;
  assign n28145 = pi17 ? n363 : n28144;
  assign n28146 = pi16 ? n21561 : n28145;
  assign n28147 = pi15 ? n28140 : n28146;
  assign n28148 = pi14 ? n28134 : n28147;
  assign n28149 = pi13 ? n28127 : n28148;
  assign n28150 = pi12 ? n28113 : n28149;
  assign n28151 = pi11 ? n28078 : n28150;
  assign n28152 = pi10 ? n27993 : n28151;
  assign n28153 = pi09 ? n27266 : n28152;
  assign n28154 = pi08 ? n27826 : n28153;
  assign n28155 = pi07 ? n27239 : n28154;
  assign n28156 = pi22 ? n32 : n20563;
  assign n28157 = pi21 ? n28156 : n20563;
  assign n28158 = pi20 ? n32 : n28157;
  assign n28159 = pi19 ? n32 : n28158;
  assign n28160 = pi18 ? n28159 : n37;
  assign n28161 = pi17 ? n32 : n28160;
  assign n28162 = pi19 ? n23648 : n20657;
  assign n28163 = pi19 ? n16999 : n32;
  assign n28164 = pi18 ? n28162 : n28163;
  assign n28165 = pi17 ? n37 : n28164;
  assign n28166 = pi16 ? n28161 : n28165;
  assign n28167 = pi15 ? n32 : n28166;
  assign n28168 = pi18 ? n14443 : n26408;
  assign n28169 = pi17 ? n32 : n28168;
  assign n28170 = pi19 ? n99 : n32;
  assign n28171 = pi18 ? n99 : n28170;
  assign n28172 = pi17 ? n99 : n28171;
  assign n28173 = pi16 ? n28169 : n28172;
  assign n28174 = pi18 ? n16593 : n14842;
  assign n28175 = pi17 ? n32 : n28174;
  assign n28176 = pi16 ? n28175 : n28172;
  assign n28177 = pi15 ? n28173 : n28176;
  assign n28178 = pi14 ? n28167 : n28177;
  assign n28179 = pi13 ? n32 : n28178;
  assign n28180 = pi12 ? n32 : n28179;
  assign n28181 = pi11 ? n32 : n28180;
  assign n28182 = pi10 ? n32 : n28181;
  assign n28183 = pi19 ? n37 : n3050;
  assign n28184 = pi19 ? n4583 : n220;
  assign n28185 = pi18 ? n28183 : n28184;
  assign n28186 = pi19 ? n22702 : n32;
  assign n28187 = pi18 ? n14845 : n28186;
  assign n28188 = pi17 ? n28185 : n28187;
  assign n28189 = pi16 ? n16595 : n28188;
  assign n28190 = pi20 ? n2973 : n99;
  assign n28191 = pi19 ? n37 : n28190;
  assign n28192 = pi18 ? n17008 : n28191;
  assign n28193 = pi17 ? n32 : n28192;
  assign n28194 = pi20 ? n99 : n14844;
  assign n28195 = pi19 ? n99 : n28194;
  assign n28196 = pi20 ? n99 : n1658;
  assign n28197 = pi19 ? n28196 : n32;
  assign n28198 = pi18 ? n28195 : n28197;
  assign n28199 = pi17 ? n99 : n28198;
  assign n28200 = pi16 ? n28193 : n28199;
  assign n28201 = pi15 ? n28189 : n28200;
  assign n28202 = pi19 ? n37 : n23645;
  assign n28203 = pi18 ? n17008 : n28202;
  assign n28204 = pi17 ? n32 : n28203;
  assign n28205 = pi20 ? n14887 : n2973;
  assign n28206 = pi19 ? n28205 : n3038;
  assign n28207 = pi19 ? n2973 : n21640;
  assign n28208 = pi18 ? n28206 : n28207;
  assign n28209 = pi20 ? n23290 : n7745;
  assign n28210 = pi20 ? n21643 : n219;
  assign n28211 = pi19 ? n28209 : n28210;
  assign n28212 = pi20 ? n99 : n4549;
  assign n28213 = pi19 ? n28212 : n32;
  assign n28214 = pi18 ? n28211 : n28213;
  assign n28215 = pi17 ? n28208 : n28214;
  assign n28216 = pi16 ? n28204 : n28215;
  assign n28217 = pi20 ? n14887 : n37;
  assign n28218 = pi19 ? n37 : n28217;
  assign n28219 = pi20 ? n2176 : n37;
  assign n28220 = pi19 ? n28219 : n3039;
  assign n28221 = pi18 ? n28218 : n28220;
  assign n28222 = pi20 ? n218 : n2976;
  assign n28223 = pi20 ? n2973 : n7747;
  assign n28224 = pi19 ? n28222 : n28223;
  assign n28225 = pi20 ? n218 : n13920;
  assign n28226 = pi19 ? n28225 : n32;
  assign n28227 = pi18 ? n28224 : n28226;
  assign n28228 = pi17 ? n28221 : n28227;
  assign n28229 = pi16 ? n439 : n28228;
  assign n28230 = pi15 ? n28216 : n28229;
  assign n28231 = pi14 ? n28201 : n28230;
  assign n28232 = pi21 ? n180 : n2164;
  assign n28233 = pi20 ? n32 : n28232;
  assign n28234 = pi19 ? n32 : n28233;
  assign n28235 = pi20 ? n4202 : n99;
  assign n28236 = pi19 ? n28235 : n99;
  assign n28237 = pi18 ? n28234 : n28236;
  assign n28238 = pi17 ? n32 : n28237;
  assign n28239 = pi22 ? n99 : n10510;
  assign n28240 = pi21 ? n99 : n28239;
  assign n28241 = pi20 ? n99 : n28240;
  assign n28242 = pi19 ? n28241 : n32;
  assign n28243 = pi18 ? n99 : n28242;
  assign n28244 = pi17 ? n99 : n28243;
  assign n28245 = pi16 ? n28238 : n28244;
  assign n28246 = pi21 ? n99 : n4247;
  assign n28247 = pi19 ? n99 : n28246;
  assign n28248 = pi18 ? n99 : n28247;
  assign n28249 = pi21 ? n4237 : n28239;
  assign n28250 = pi20 ? n4247 : n28249;
  assign n28251 = pi19 ? n28250 : n32;
  assign n28252 = pi18 ? n99 : n28251;
  assign n28253 = pi17 ? n28248 : n28252;
  assign n28254 = pi16 ? n25610 : n28253;
  assign n28255 = pi15 ? n28245 : n28254;
  assign n28256 = pi19 ? n9824 : n8765;
  assign n28257 = pi19 ? n13093 : n139;
  assign n28258 = pi18 ? n28256 : n28257;
  assign n28259 = pi22 ? n139 : n1196;
  assign n28260 = pi21 ? n139 : n28259;
  assign n28261 = pi20 ? n139 : n28260;
  assign n28262 = pi19 ? n28261 : n32;
  assign n28263 = pi18 ? n139 : n28262;
  assign n28264 = pi17 ? n28258 : n28263;
  assign n28265 = pi16 ? n439 : n28264;
  assign n28266 = pi18 ? n15029 : n28257;
  assign n28267 = pi22 ? n139 : n13969;
  assign n28268 = pi21 ? n916 : n28267;
  assign n28269 = pi20 ? n139 : n28268;
  assign n28270 = pi19 ? n28269 : n32;
  assign n28271 = pi18 ? n139 : n28270;
  assign n28272 = pi17 ? n28266 : n28271;
  assign n28273 = pi16 ? n439 : n28272;
  assign n28274 = pi15 ? n28265 : n28273;
  assign n28275 = pi14 ? n28255 : n28274;
  assign n28276 = pi13 ? n28231 : n28275;
  assign n28277 = pi19 ? n37 : n15033;
  assign n28278 = pi18 ? n37 : n28277;
  assign n28279 = pi20 ? n3092 : n3086;
  assign n28280 = pi20 ? n13613 : n3096;
  assign n28281 = pi19 ? n28279 : n28280;
  assign n28282 = pi23 ? n37 : n531;
  assign n28283 = pi22 ? n139 : n28282;
  assign n28284 = pi21 ? n139 : n28283;
  assign n28285 = pi20 ? n139 : n28284;
  assign n28286 = pi19 ? n28285 : n32;
  assign n28287 = pi18 ? n28281 : n28286;
  assign n28288 = pi17 ? n28278 : n28287;
  assign n28289 = pi16 ? n439 : n28288;
  assign n28290 = pi20 ? n1003 : n37;
  assign n28291 = pi19 ? n28290 : n9824;
  assign n28292 = pi23 ? n37 : n624;
  assign n28293 = pi22 ? n139 : n28292;
  assign n28294 = pi21 ? n139 : n28293;
  assign n28295 = pi20 ? n139 : n28294;
  assign n28296 = pi19 ? n28295 : n32;
  assign n28297 = pi18 ? n28291 : n28296;
  assign n28298 = pi17 ? n16094 : n28297;
  assign n28299 = pi16 ? n439 : n28298;
  assign n28300 = pi15 ? n28289 : n28299;
  assign n28301 = pi21 ? n139 : n20300;
  assign n28302 = pi20 ? n139 : n28301;
  assign n28303 = pi19 ? n28302 : n32;
  assign n28304 = pi18 ? n17061 : n28303;
  assign n28305 = pi17 ? n12372 : n28304;
  assign n28306 = pi16 ? n439 : n28305;
  assign n28307 = pi19 ? n9824 : n13168;
  assign n28308 = pi18 ? n37 : n28307;
  assign n28309 = pi19 ? n3083 : n18934;
  assign n28310 = pi21 ? n139 : n20308;
  assign n28311 = pi20 ? n139 : n28310;
  assign n28312 = pi19 ? n28311 : n32;
  assign n28313 = pi18 ? n28309 : n28312;
  assign n28314 = pi17 ? n28308 : n28313;
  assign n28315 = pi16 ? n439 : n28314;
  assign n28316 = pi15 ? n28306 : n28315;
  assign n28317 = pi14 ? n28300 : n28316;
  assign n28318 = pi18 ? n37 : n20760;
  assign n28319 = pi22 ? n139 : n20317;
  assign n28320 = pi21 ? n139 : n28319;
  assign n28321 = pi20 ? n139 : n28320;
  assign n28322 = pi19 ? n28321 : n32;
  assign n28323 = pi18 ? n16093 : n28322;
  assign n28324 = pi17 ? n28318 : n28323;
  assign n28325 = pi16 ? n439 : n28324;
  assign n28326 = pi20 ? n139 : n14086;
  assign n28327 = pi19 ? n28326 : n32;
  assign n28328 = pi18 ? n14115 : n28327;
  assign n28329 = pi17 ? n19830 : n28328;
  assign n28330 = pi16 ? n439 : n28329;
  assign n28331 = pi15 ? n28325 : n28330;
  assign n28332 = pi21 ? n335 : n21355;
  assign n28333 = pi20 ? n335 : n28332;
  assign n28334 = pi19 ? n28333 : n32;
  assign n28335 = pi18 ? n7677 : n28334;
  assign n28336 = pi17 ? n37 : n28335;
  assign n28337 = pi16 ? n439 : n28336;
  assign n28338 = pi21 ? n2007 : n20800;
  assign n28339 = pi20 ? n3335 : n28338;
  assign n28340 = pi19 ? n28339 : n32;
  assign n28341 = pi18 ? n14149 : n28340;
  assign n28342 = pi17 ? n37 : n28341;
  assign n28343 = pi16 ? n439 : n28342;
  assign n28344 = pi15 ? n28337 : n28343;
  assign n28345 = pi14 ? n28331 : n28344;
  assign n28346 = pi13 ? n28317 : n28345;
  assign n28347 = pi12 ? n28276 : n28346;
  assign n28348 = pi22 ? n335 : n13626;
  assign n28349 = pi21 ? n2007 : n28348;
  assign n28350 = pi20 ? n649 : n28349;
  assign n28351 = pi19 ? n28350 : n32;
  assign n28352 = pi18 ? n37 : n28351;
  assign n28353 = pi17 ? n37 : n28352;
  assign n28354 = pi16 ? n439 : n28353;
  assign n28355 = pi21 ? n335 : n20800;
  assign n28356 = pi20 ? n335 : n28355;
  assign n28357 = pi19 ? n28356 : n32;
  assign n28358 = pi18 ? n37 : n28357;
  assign n28359 = pi17 ? n37 : n28358;
  assign n28360 = pi16 ? n439 : n28359;
  assign n28361 = pi15 ? n28354 : n28360;
  assign n28362 = pi18 ? n7686 : n28357;
  assign n28363 = pi17 ? n37 : n28362;
  assign n28364 = pi16 ? n439 : n28363;
  assign n28365 = pi19 ? n37 : n643;
  assign n28366 = pi18 ? n37 : n28365;
  assign n28367 = pi20 ? n577 : n603;
  assign n28368 = pi19 ? n37 : n28367;
  assign n28369 = pi21 ? n570 : n20800;
  assign n28370 = pi20 ? n335 : n28369;
  assign n28371 = pi19 ? n28370 : n32;
  assign n28372 = pi18 ? n28368 : n28371;
  assign n28373 = pi17 ? n28366 : n28372;
  assign n28374 = pi16 ? n439 : n28373;
  assign n28375 = pi15 ? n28364 : n28374;
  assign n28376 = pi14 ? n28361 : n28375;
  assign n28377 = pi21 ? n335 : n567;
  assign n28378 = pi20 ? n28377 : n570;
  assign n28379 = pi19 ? n37 : n28378;
  assign n28380 = pi18 ? n22068 : n28379;
  assign n28381 = pi20 ? n639 : n603;
  assign n28382 = pi19 ? n28381 : n16516;
  assign n28383 = pi18 ? n28382 : n28357;
  assign n28384 = pi17 ? n28380 : n28383;
  assign n28385 = pi16 ? n439 : n28384;
  assign n28386 = pi21 ? n569 : n20800;
  assign n28387 = pi20 ? n335 : n28386;
  assign n28388 = pi19 ? n28387 : n32;
  assign n28389 = pi18 ? n17205 : n28388;
  assign n28390 = pi17 ? n37 : n28389;
  assign n28391 = pi16 ? n439 : n28390;
  assign n28392 = pi15 ? n28385 : n28391;
  assign n28393 = pi21 ? n2007 : n6376;
  assign n28394 = pi20 ? n37 : n28393;
  assign n28395 = pi19 ? n37 : n28394;
  assign n28396 = pi22 ? n2060 : n4899;
  assign n28397 = pi21 ? n11199 : n28396;
  assign n28398 = pi21 ? n5014 : n665;
  assign n28399 = pi20 ? n28397 : n28398;
  assign n28400 = pi19 ? n28399 : n32;
  assign n28401 = pi18 ? n28395 : n28400;
  assign n28402 = pi17 ? n37 : n28401;
  assign n28403 = pi16 ? n439 : n28402;
  assign n28404 = pi21 ? n5015 : n4920;
  assign n28405 = pi21 ? n2048 : n14168;
  assign n28406 = pi20 ? n28404 : n28405;
  assign n28407 = pi19 ? n28406 : n32;
  assign n28408 = pi18 ? n19093 : n28407;
  assign n28409 = pi17 ? n37 : n28408;
  assign n28410 = pi16 ? n439 : n28409;
  assign n28411 = pi15 ? n28403 : n28410;
  assign n28412 = pi14 ? n28392 : n28411;
  assign n28413 = pi13 ? n28376 : n28412;
  assign n28414 = pi21 ? n19958 : n1423;
  assign n28415 = pi20 ? n37 : n28414;
  assign n28416 = pi19 ? n28415 : n32;
  assign n28417 = pi18 ? n37 : n28416;
  assign n28418 = pi17 ? n37 : n28417;
  assign n28419 = pi16 ? n439 : n28418;
  assign n28420 = pi21 ? n37 : n2230;
  assign n28421 = pi20 ? n9660 : n28420;
  assign n28422 = pi19 ? n28421 : n32;
  assign n28423 = pi18 ? n37 : n28422;
  assign n28424 = pi17 ? n37 : n28423;
  assign n28425 = pi16 ? n439 : n28424;
  assign n28426 = pi15 ? n28419 : n28425;
  assign n28427 = pi20 ? n37 : n28420;
  assign n28428 = pi19 ? n28427 : n32;
  assign n28429 = pi18 ? n37 : n28428;
  assign n28430 = pi17 ? n37 : n28429;
  assign n28431 = pi16 ? n439 : n28430;
  assign n28432 = pi19 ? n691 : n32;
  assign n28433 = pi18 ? n37 : n28432;
  assign n28434 = pi17 ? n37 : n28433;
  assign n28435 = pi16 ? n439 : n28434;
  assign n28436 = pi15 ? n28431 : n28435;
  assign n28437 = pi14 ? n28426 : n28436;
  assign n28438 = pi22 ? n24857 : n706;
  assign n28439 = pi21 ? n3392 : n28438;
  assign n28440 = pi20 ? n37 : n28439;
  assign n28441 = pi19 ? n28440 : n32;
  assign n28442 = pi18 ? n37 : n28441;
  assign n28443 = pi17 ? n37 : n28442;
  assign n28444 = pi16 ? n439 : n28443;
  assign n28445 = pi20 ? n13310 : n37;
  assign n28446 = pi19 ? n37 : n28445;
  assign n28447 = pi23 ? n363 : n842;
  assign n28448 = pi22 ? n28447 : n32;
  assign n28449 = pi21 ? n3392 : n28448;
  assign n28450 = pi20 ? n37 : n28449;
  assign n28451 = pi19 ? n28450 : n32;
  assign n28452 = pi18 ? n28446 : n28451;
  assign n28453 = pi17 ? n37 : n28452;
  assign n28454 = pi16 ? n439 : n28453;
  assign n28455 = pi15 ? n28444 : n28454;
  assign n28456 = pi20 ? n19091 : n7730;
  assign n28457 = pi20 ? n22881 : n3393;
  assign n28458 = pi19 ? n28456 : n28457;
  assign n28459 = pi18 ? n374 : n28458;
  assign n28460 = pi17 ? n32 : n28459;
  assign n28461 = pi19 ? n363 : n27520;
  assign n28462 = pi19 ? n27520 : n363;
  assign n28463 = pi18 ? n28461 : n28462;
  assign n28464 = pi20 ? n10496 : n363;
  assign n28465 = pi19 ? n28464 : n363;
  assign n28466 = pi23 ? n363 : n531;
  assign n28467 = pi22 ? n28466 : n32;
  assign n28468 = pi21 ? n37 : n28467;
  assign n28469 = pi20 ? n22881 : n28468;
  assign n28470 = pi19 ? n28469 : n32;
  assign n28471 = pi18 ? n28465 : n28470;
  assign n28472 = pi17 ? n28463 : n28471;
  assign n28473 = pi16 ? n28460 : n28472;
  assign n28474 = pi21 ? n2957 : n1512;
  assign n28475 = pi20 ? n37 : n28474;
  assign n28476 = pi19 ? n28475 : n32;
  assign n28477 = pi18 ? n37 : n28476;
  assign n28478 = pi17 ? n37 : n28477;
  assign n28479 = pi16 ? n439 : n28478;
  assign n28480 = pi15 ? n28473 : n28479;
  assign n28481 = pi14 ? n28455 : n28480;
  assign n28482 = pi13 ? n28437 : n28481;
  assign n28483 = pi12 ? n28413 : n28482;
  assign n28484 = pi11 ? n28347 : n28483;
  assign n28485 = pi21 ? n19933 : n685;
  assign n28486 = pi20 ? n37 : n28485;
  assign n28487 = pi19 ? n37 : n28486;
  assign n28488 = pi21 ? n2106 : n748;
  assign n28489 = pi20 ? n37 : n28488;
  assign n28490 = pi19 ? n28489 : n32;
  assign n28491 = pi18 ? n28487 : n28490;
  assign n28492 = pi17 ? n37 : n28491;
  assign n28493 = pi16 ? n439 : n28492;
  assign n28494 = pi20 ? n24493 : n244;
  assign n28495 = pi19 ? n28494 : n37;
  assign n28496 = pi20 ? n37 : n273;
  assign n28497 = pi22 ? n157 : n889;
  assign n28498 = pi21 ? n37 : n28497;
  assign n28499 = pi20 ? n273 : n28498;
  assign n28500 = pi19 ? n28496 : n28499;
  assign n28501 = pi18 ? n28495 : n28500;
  assign n28502 = pi21 ? n272 : n23932;
  assign n28503 = pi20 ? n24493 : n28502;
  assign n28504 = pi20 ? n278 : n7829;
  assign n28505 = pi19 ? n28503 : n28504;
  assign n28506 = pi22 ? n112 : n685;
  assign n28507 = pi21 ? n28506 : n3319;
  assign n28508 = pi20 ? n685 : n28507;
  assign n28509 = pi19 ? n28508 : n32;
  assign n28510 = pi18 ? n28505 : n28509;
  assign n28511 = pi17 ? n28501 : n28510;
  assign n28512 = pi16 ? n439 : n28511;
  assign n28513 = pi15 ? n28493 : n28512;
  assign n28514 = pi20 ? n25804 : n16279;
  assign n28515 = pi19 ? n37 : n28514;
  assign n28516 = pi21 ? n3445 : n685;
  assign n28517 = pi20 ? n28516 : n28002;
  assign n28518 = pi19 ? n28517 : n32;
  assign n28519 = pi18 ? n28515 : n28518;
  assign n28520 = pi17 ? n37 : n28519;
  assign n28521 = pi16 ? n439 : n28520;
  assign n28522 = pi20 ? n25804 : n157;
  assign n28523 = pi19 ? n37 : n28522;
  assign n28524 = pi21 ? n3562 : n157;
  assign n28525 = pi21 ? n19178 : n882;
  assign n28526 = pi20 ? n28524 : n28525;
  assign n28527 = pi19 ? n28526 : n32;
  assign n28528 = pi18 ? n28523 : n28527;
  assign n28529 = pi17 ? n37 : n28528;
  assign n28530 = pi16 ? n439 : n28529;
  assign n28531 = pi15 ? n28521 : n28530;
  assign n28532 = pi14 ? n28513 : n28531;
  assign n28533 = pi20 ? n99 : n2330;
  assign n28534 = pi19 ? n28533 : n32;
  assign n28535 = pi18 ? n99 : n28534;
  assign n28536 = pi17 ? n99 : n28535;
  assign n28537 = pi16 ? n744 : n28536;
  assign n28538 = pi20 ? n776 : n27095;
  assign n28539 = pi19 ? n28538 : n32;
  assign n28540 = pi18 ? n10010 : n28539;
  assign n28541 = pi17 ? n99 : n28540;
  assign n28542 = pi16 ? n744 : n28541;
  assign n28543 = pi15 ? n28537 : n28542;
  assign n28544 = pi20 ? n99 : n27598;
  assign n28545 = pi19 ? n99 : n28544;
  assign n28546 = pi18 ? n28545 : n28035;
  assign n28547 = pi17 ? n99 : n28546;
  assign n28548 = pi16 ? n744 : n28547;
  assign n28549 = pi15 ? n27103 : n28548;
  assign n28550 = pi14 ? n28543 : n28549;
  assign n28551 = pi13 ? n28532 : n28550;
  assign n28552 = pi22 ? n316 : n158;
  assign n28553 = pi21 ? n159 : n28552;
  assign n28554 = pi20 ? n26680 : n28553;
  assign n28555 = pi19 ? n139 : n28554;
  assign n28556 = pi21 ? n8632 : n1009;
  assign n28557 = pi20 ? n2238 : n28556;
  assign n28558 = pi19 ? n28557 : n32;
  assign n28559 = pi18 ? n28555 : n28558;
  assign n28560 = pi17 ? n26684 : n28559;
  assign n28561 = pi16 ? n25417 : n28560;
  assign n28562 = pi20 ? n18317 : n16476;
  assign n28563 = pi19 ? n28562 : n32;
  assign n28564 = pi18 ? n9111 : n28563;
  assign n28565 = pi17 ? n139 : n28564;
  assign n28566 = pi16 ? n915 : n28565;
  assign n28567 = pi15 ? n28561 : n28566;
  assign n28568 = pi20 ? n3731 : n16476;
  assign n28569 = pi19 ? n28568 : n32;
  assign n28570 = pi18 ? n18328 : n28569;
  assign n28571 = pi17 ? n139 : n28570;
  assign n28572 = pi16 ? n915 : n28571;
  assign n28573 = pi18 ? n990 : n11552;
  assign n28574 = pi17 ? n32 : n28573;
  assign n28575 = pi21 ? n1056 : n37;
  assign n28576 = pi20 ? n37 : n28575;
  assign n28577 = pi19 ? n28576 : n37;
  assign n28578 = pi21 ? n139 : n1056;
  assign n28579 = pi20 ? n37 : n28578;
  assign n28580 = pi19 ? n18934 : n28579;
  assign n28581 = pi18 ? n28577 : n28580;
  assign n28582 = pi20 ? n3096 : n37;
  assign n28583 = pi21 ? n1056 : n316;
  assign n28584 = pi20 ? n28583 : n316;
  assign n28585 = pi19 ? n28582 : n28584;
  assign n28586 = pi20 ? n4437 : n16476;
  assign n28587 = pi19 ? n28586 : n32;
  assign n28588 = pi18 ? n28585 : n28587;
  assign n28589 = pi17 ? n28581 : n28588;
  assign n28590 = pi16 ? n28574 : n28589;
  assign n28591 = pi15 ? n28572 : n28590;
  assign n28592 = pi14 ? n28567 : n28591;
  assign n28593 = pi20 ? n1068 : n204;
  assign n28594 = pi19 ? n204 : n28593;
  assign n28595 = pi18 ? n13844 : n28594;
  assign n28596 = pi17 ? n32 : n28595;
  assign n28597 = pi20 ? n1059 : n2383;
  assign n28598 = pi19 ? n28597 : n7858;
  assign n28599 = pi20 ? n7858 : n1059;
  assign n28600 = pi21 ? n1027 : n391;
  assign n28601 = pi20 ? n28600 : n7909;
  assign n28602 = pi19 ? n28599 : n28601;
  assign n28603 = pi18 ? n28598 : n28602;
  assign n28604 = pi20 ? n1060 : n1018;
  assign n28605 = pi19 ? n28604 : n316;
  assign n28606 = pi20 ? n316 : n13398;
  assign n28607 = pi19 ? n28606 : n32;
  assign n28608 = pi18 ? n28605 : n28607;
  assign n28609 = pi17 ? n28603 : n28608;
  assign n28610 = pi16 ? n28596 : n28609;
  assign n28611 = pi21 ? n20102 : n2319;
  assign n28612 = pi20 ? n204 : n28611;
  assign n28613 = pi19 ? n204 : n28612;
  assign n28614 = pi20 ? n1059 : n14748;
  assign n28615 = pi19 ? n28614 : n32;
  assign n28616 = pi18 ? n28613 : n28615;
  assign n28617 = pi17 ? n204 : n28616;
  assign n28618 = pi16 ? n24565 : n28617;
  assign n28619 = pi15 ? n28610 : n28618;
  assign n28620 = pi19 ? n204 : n13494;
  assign n28621 = pi18 ? n204 : n28620;
  assign n28622 = pi20 ? n204 : n28062;
  assign n28623 = pi19 ? n28622 : n32;
  assign n28624 = pi18 ? n204 : n28623;
  assign n28625 = pi17 ? n28621 : n28624;
  assign n28626 = pi16 ? n13846 : n28625;
  assign n28627 = pi21 ? n204 : n820;
  assign n28628 = pi20 ? n28627 : n21011;
  assign n28629 = pi19 ? n204 : n28628;
  assign n28630 = pi18 ? n204 : n28629;
  assign n28631 = pi20 ? n204 : n16944;
  assign n28632 = pi19 ? n28631 : n32;
  assign n28633 = pi18 ? n204 : n28632;
  assign n28634 = pi17 ? n28630 : n28633;
  assign n28635 = pi16 ? n13833 : n28634;
  assign n28636 = pi15 ? n28626 : n28635;
  assign n28637 = pi14 ? n28619 : n28636;
  assign n28638 = pi13 ? n28592 : n28637;
  assign n28639 = pi12 ? n28551 : n28638;
  assign n28640 = pi20 ? n1016 : n28069;
  assign n28641 = pi19 ? n28640 : n32;
  assign n28642 = pi18 ? n11765 : n28641;
  assign n28643 = pi17 ? n139 : n28642;
  assign n28644 = pi16 ? n915 : n28643;
  assign n28645 = pi19 ? n335 : n2068;
  assign n28646 = pi18 ? n602 : n28645;
  assign n28647 = pi17 ? n32 : n28646;
  assign n28648 = pi19 ? n335 : n11815;
  assign n28649 = pi22 ? n139 : n233;
  assign n28650 = pi21 ? n335 : n28649;
  assign n28651 = pi20 ? n28650 : n28084;
  assign n28652 = pi19 ? n28651 : n32;
  assign n28653 = pi18 ? n28648 : n28652;
  assign n28654 = pi17 ? n335 : n28653;
  assign n28655 = pi16 ? n28647 : n28654;
  assign n28656 = pi15 ? n28644 : n28655;
  assign n28657 = pi20 ? n6377 : n8958;
  assign n28658 = pi19 ? n28657 : n32;
  assign n28659 = pi18 ? n335 : n28658;
  assign n28660 = pi17 ? n335 : n28659;
  assign n28661 = pi16 ? n2035 : n28660;
  assign n28662 = pi20 ? n6377 : n7733;
  assign n28663 = pi19 ? n28662 : n32;
  assign n28664 = pi18 ? n335 : n28663;
  assign n28665 = pi17 ? n335 : n28664;
  assign n28666 = pi16 ? n7943 : n28665;
  assign n28667 = pi15 ? n28661 : n28666;
  assign n28668 = pi14 ? n28656 : n28667;
  assign n28669 = pi21 ? n2061 : n233;
  assign n28670 = pi20 ? n28669 : n4102;
  assign n28671 = pi19 ? n28670 : n32;
  assign n28672 = pi18 ? n15438 : n28671;
  assign n28673 = pi17 ? n335 : n28672;
  assign n28674 = pi16 ? n7943 : n28673;
  assign n28675 = pi20 ? n233 : n6417;
  assign n28676 = pi19 ? n28675 : n32;
  assign n28677 = pi18 ? n15438 : n28676;
  assign n28678 = pi17 ? n335 : n28677;
  assign n28679 = pi16 ? n7943 : n28678;
  assign n28680 = pi15 ? n28674 : n28679;
  assign n28681 = pi19 ? n17486 : n335;
  assign n28682 = pi18 ? n335 : n28681;
  assign n28683 = pi21 ? n16562 : n233;
  assign n28684 = pi20 ? n28683 : n6417;
  assign n28685 = pi19 ? n28684 : n32;
  assign n28686 = pi18 ? n15438 : n28685;
  assign n28687 = pi17 ? n28682 : n28686;
  assign n28688 = pi16 ? n2035 : n28687;
  assign n28689 = pi21 ? n19386 : n335;
  assign n28690 = pi20 ? n335 : n28689;
  assign n28691 = pi19 ? n28690 : n335;
  assign n28692 = pi18 ? n335 : n28691;
  assign n28693 = pi17 ? n28692 : n27709;
  assign n28694 = pi16 ? n7943 : n28693;
  assign n28695 = pi15 ? n28688 : n28694;
  assign n28696 = pi14 ? n28680 : n28695;
  assign n28697 = pi13 ? n28668 : n28696;
  assign n28698 = pi21 ? n26857 : n6361;
  assign n28699 = pi20 ? n32 : n28698;
  assign n28700 = pi19 ? n32 : n28699;
  assign n28701 = pi21 ? n6361 : n6376;
  assign n28702 = pi20 ? n18431 : n28701;
  assign n28703 = pi19 ? n28702 : n15470;
  assign n28704 = pi18 ? n28700 : n28703;
  assign n28705 = pi17 ? n32 : n28704;
  assign n28706 = pi20 ? n15465 : n16544;
  assign n28707 = pi19 ? n233 : n28706;
  assign n28708 = pi18 ? n233 : n28707;
  assign n28709 = pi20 ? n233 : n5830;
  assign n28710 = pi19 ? n28709 : n32;
  assign n28711 = pi18 ? n233 : n28710;
  assign n28712 = pi17 ? n28708 : n28711;
  assign n28713 = pi16 ? n28705 : n28712;
  assign n28714 = pi19 ? n6355 : n37;
  assign n28715 = pi20 ? n37 : n6358;
  assign n28716 = pi19 ? n28715 : n6359;
  assign n28717 = pi18 ? n28714 : n28716;
  assign n28718 = pi20 ? n37 : n21124;
  assign n28719 = pi19 ? n28718 : n233;
  assign n28720 = pi18 ? n28719 : n27719;
  assign n28721 = pi17 ? n28717 : n28720;
  assign n28722 = pi16 ? n439 : n28721;
  assign n28723 = pi15 ? n28713 : n28722;
  assign n28724 = pi19 ? n37 : n233;
  assign n28725 = pi18 ? n28724 : n26338;
  assign n28726 = pi17 ? n37 : n28725;
  assign n28727 = pi16 ? n439 : n28726;
  assign n28728 = pi21 ? n25162 : n5014;
  assign n28729 = pi20 ? n32 : n28728;
  assign n28730 = pi19 ? n32 : n28729;
  assign n28731 = pi20 ? n26880 : n23155;
  assign n28732 = pi21 ? n722 : n99;
  assign n28733 = pi20 ? n28732 : n99;
  assign n28734 = pi19 ? n28731 : n28733;
  assign n28735 = pi18 ? n28730 : n28734;
  assign n28736 = pi17 ? n32 : n28735;
  assign n28737 = pi21 ? n22128 : n99;
  assign n28738 = pi20 ? n28737 : n233;
  assign n28739 = pi19 ? n28738 : n9197;
  assign n28740 = pi20 ? n25166 : n233;
  assign n28741 = pi19 ? n26881 : n28740;
  assign n28742 = pi18 ? n28739 : n28741;
  assign n28743 = pi21 ? n99 : n233;
  assign n28744 = pi21 ? n22128 : n233;
  assign n28745 = pi20 ? n28743 : n28744;
  assign n28746 = pi22 ? n685 : n233;
  assign n28747 = pi21 ? n233 : n28746;
  assign n28748 = pi20 ? n233 : n28747;
  assign n28749 = pi19 ? n28745 : n28748;
  assign n28750 = pi21 ? n233 : n12635;
  assign n28751 = pi20 ? n28750 : n2653;
  assign n28752 = pi19 ? n28751 : n32;
  assign n28753 = pi18 ? n28749 : n28752;
  assign n28754 = pi17 ? n28742 : n28753;
  assign n28755 = pi16 ? n28736 : n28754;
  assign n28756 = pi15 ? n28727 : n28755;
  assign n28757 = pi14 ? n28723 : n28756;
  assign n28758 = pi22 ? n26027 : n363;
  assign n28759 = pi21 ? n28758 : n363;
  assign n28760 = pi20 ? n32 : n28759;
  assign n28761 = pi19 ? n32 : n28760;
  assign n28762 = pi18 ? n28761 : n363;
  assign n28763 = pi17 ? n32 : n28762;
  assign n28764 = pi20 ? n23162 : n363;
  assign n28765 = pi19 ? n363 : n28764;
  assign n28766 = pi18 ? n363 : n28765;
  assign n28767 = pi20 ? n363 : n685;
  assign n28768 = pi19 ? n363 : n28767;
  assign n28769 = pi21 ? n363 : n5113;
  assign n28770 = pi20 ? n28769 : n1822;
  assign n28771 = pi19 ? n28770 : n32;
  assign n28772 = pi18 ? n28768 : n28771;
  assign n28773 = pi17 ? n28766 : n28772;
  assign n28774 = pi16 ? n28763 : n28773;
  assign n28775 = pi20 ? n19084 : n18194;
  assign n28776 = pi19 ? n363 : n28775;
  assign n28777 = pi20 ? n28769 : n32;
  assign n28778 = pi19 ? n28777 : n32;
  assign n28779 = pi18 ? n28776 : n28778;
  assign n28780 = pi17 ? n363 : n28779;
  assign n28781 = pi16 ? n21219 : n28780;
  assign n28782 = pi15 ? n28774 : n28781;
  assign n28783 = pi21 ? n363 : n2200;
  assign n28784 = pi20 ? n28783 : n32;
  assign n28785 = pi19 ? n28784 : n32;
  assign n28786 = pi18 ? n363 : n28785;
  assign n28787 = pi17 ? n363 : n28786;
  assign n28788 = pi16 ? n21219 : n28787;
  assign n28789 = pi18 ? n363 : n25533;
  assign n28790 = pi17 ? n363 : n28789;
  assign n28791 = pi16 ? n26062 : n28790;
  assign n28792 = pi15 ? n28788 : n28791;
  assign n28793 = pi14 ? n28782 : n28792;
  assign n28794 = pi13 ? n28757 : n28793;
  assign n28795 = pi12 ? n28697 : n28794;
  assign n28796 = pi11 ? n28639 : n28795;
  assign n28797 = pi10 ? n28484 : n28796;
  assign n28798 = pi09 ? n28182 : n28797;
  assign n28799 = pi19 ? n1666 : n32;
  assign n28800 = pi18 ? n99 : n28799;
  assign n28801 = pi17 ? n99 : n28800;
  assign n28802 = pi16 ? n28238 : n28801;
  assign n28803 = pi15 ? n28802 : n28254;
  assign n28804 = pi19 ? n1795 : n32;
  assign n28805 = pi18 ? n139 : n28804;
  assign n28806 = pi17 ? n28258 : n28805;
  assign n28807 = pi16 ? n439 : n28806;
  assign n28808 = pi20 ? n139 : n4366;
  assign n28809 = pi19 ? n28808 : n32;
  assign n28810 = pi18 ? n139 : n28809;
  assign n28811 = pi17 ? n28266 : n28810;
  assign n28812 = pi16 ? n439 : n28811;
  assign n28813 = pi15 ? n28807 : n28812;
  assign n28814 = pi14 ? n28803 : n28813;
  assign n28815 = pi13 ? n28231 : n28814;
  assign n28816 = pi20 ? n139 : n1811;
  assign n28817 = pi19 ? n28816 : n32;
  assign n28818 = pi18 ? n28281 : n28817;
  assign n28819 = pi17 ? n28278 : n28818;
  assign n28820 = pi16 ? n439 : n28819;
  assign n28821 = pi22 ? n139 : n559;
  assign n28822 = pi21 ? n139 : n28821;
  assign n28823 = pi20 ? n139 : n28822;
  assign n28824 = pi19 ? n28823 : n32;
  assign n28825 = pi18 ? n28291 : n28824;
  assign n28826 = pi17 ? n16094 : n28825;
  assign n28827 = pi16 ? n439 : n28826;
  assign n28828 = pi15 ? n28820 : n28827;
  assign n28829 = pi20 ? n139 : n14953;
  assign n28830 = pi19 ? n28829 : n32;
  assign n28831 = pi18 ? n17061 : n28830;
  assign n28832 = pi17 ? n12372 : n28831;
  assign n28833 = pi16 ? n439 : n28832;
  assign n28834 = pi20 ? n139 : n14542;
  assign n28835 = pi19 ? n28834 : n32;
  assign n28836 = pi18 ? n28309 : n28835;
  assign n28837 = pi17 ? n28308 : n28836;
  assign n28838 = pi16 ? n439 : n28837;
  assign n28839 = pi15 ? n28833 : n28838;
  assign n28840 = pi14 ? n28828 : n28839;
  assign n28841 = pi22 ? n139 : n5782;
  assign n28842 = pi21 ? n139 : n28841;
  assign n28843 = pi20 ? n139 : n28842;
  assign n28844 = pi19 ? n28843 : n32;
  assign n28845 = pi18 ? n16093 : n28844;
  assign n28846 = pi17 ? n28318 : n28845;
  assign n28847 = pi16 ? n439 : n28846;
  assign n28848 = pi21 ? n139 : n5235;
  assign n28849 = pi20 ? n139 : n28848;
  assign n28850 = pi19 ? n28849 : n32;
  assign n28851 = pi18 ? n14115 : n28850;
  assign n28852 = pi17 ? n19830 : n28851;
  assign n28853 = pi16 ? n439 : n28852;
  assign n28854 = pi15 ? n28847 : n28853;
  assign n28855 = pi22 ? n335 : n2299;
  assign n28856 = pi21 ? n335 : n28855;
  assign n28857 = pi20 ? n335 : n28856;
  assign n28858 = pi19 ? n28857 : n32;
  assign n28859 = pi18 ? n7677 : n28858;
  assign n28860 = pi17 ? n37 : n28859;
  assign n28861 = pi16 ? n439 : n28860;
  assign n28862 = pi21 ? n2007 : n15100;
  assign n28863 = pi20 ? n3335 : n28862;
  assign n28864 = pi19 ? n28863 : n32;
  assign n28865 = pi18 ? n14149 : n28864;
  assign n28866 = pi17 ? n37 : n28865;
  assign n28867 = pi16 ? n439 : n28866;
  assign n28868 = pi15 ? n28861 : n28867;
  assign n28869 = pi14 ? n28854 : n28868;
  assign n28870 = pi13 ? n28840 : n28869;
  assign n28871 = pi12 ? n28815 : n28870;
  assign n28872 = pi22 ? n335 : n16771;
  assign n28873 = pi21 ? n2007 : n28872;
  assign n28874 = pi20 ? n649 : n28873;
  assign n28875 = pi19 ? n28874 : n32;
  assign n28876 = pi18 ? n37 : n28875;
  assign n28877 = pi17 ? n37 : n28876;
  assign n28878 = pi16 ? n439 : n28877;
  assign n28879 = pi22 ? n335 : n3338;
  assign n28880 = pi21 ? n335 : n28879;
  assign n28881 = pi20 ? n335 : n28880;
  assign n28882 = pi19 ? n28881 : n32;
  assign n28883 = pi18 ? n37 : n28882;
  assign n28884 = pi17 ? n37 : n28883;
  assign n28885 = pi16 ? n439 : n28884;
  assign n28886 = pi15 ? n28878 : n28885;
  assign n28887 = pi14 ? n28886 : n28375;
  assign n28888 = pi21 ? n2007 : n11199;
  assign n28889 = pi20 ? n37 : n28888;
  assign n28890 = pi19 ? n37 : n28889;
  assign n28891 = pi21 ? n11199 : n13349;
  assign n28892 = pi20 ? n28891 : n28398;
  assign n28893 = pi19 ? n28892 : n32;
  assign n28894 = pi18 ? n28890 : n28893;
  assign n28895 = pi17 ? n37 : n28894;
  assign n28896 = pi16 ? n439 : n28895;
  assign n28897 = pi15 ? n28896 : n28410;
  assign n28898 = pi14 ? n28392 : n28897;
  assign n28899 = pi13 ? n28887 : n28898;
  assign n28900 = pi21 ? n3392 : n8957;
  assign n28901 = pi20 ? n37 : n28900;
  assign n28902 = pi19 ? n28901 : n32;
  assign n28903 = pi18 ? n37 : n28902;
  assign n28904 = pi17 ? n37 : n28903;
  assign n28905 = pi16 ? n439 : n28904;
  assign n28906 = pi21 ? n3392 : n21387;
  assign n28907 = pi20 ? n37 : n28906;
  assign n28908 = pi19 ? n28907 : n32;
  assign n28909 = pi18 ? n28446 : n28908;
  assign n28910 = pi17 ? n37 : n28909;
  assign n28911 = pi16 ? n439 : n28910;
  assign n28912 = pi15 ? n28905 : n28911;
  assign n28913 = pi21 ? n37 : n21387;
  assign n28914 = pi20 ? n22881 : n28913;
  assign n28915 = pi19 ? n28914 : n32;
  assign n28916 = pi18 ? n28465 : n28915;
  assign n28917 = pi17 ? n28463 : n28916;
  assign n28918 = pi16 ? n28460 : n28917;
  assign n28919 = pi21 ? n2957 : n2256;
  assign n28920 = pi20 ? n37 : n28919;
  assign n28921 = pi19 ? n28920 : n32;
  assign n28922 = pi18 ? n37 : n28921;
  assign n28923 = pi17 ? n37 : n28922;
  assign n28924 = pi16 ? n439 : n28923;
  assign n28925 = pi15 ? n28918 : n28924;
  assign n28926 = pi14 ? n28912 : n28925;
  assign n28927 = pi13 ? n28437 : n28926;
  assign n28928 = pi12 ? n28899 : n28927;
  assign n28929 = pi11 ? n28871 : n28928;
  assign n28930 = pi21 ? n2106 : n2256;
  assign n28931 = pi20 ? n37 : n28930;
  assign n28932 = pi19 ? n28931 : n32;
  assign n28933 = pi18 ? n28487 : n28932;
  assign n28934 = pi17 ? n37 : n28933;
  assign n28935 = pi16 ? n439 : n28934;
  assign n28936 = pi21 ? n244 : n8658;
  assign n28937 = pi20 ? n24493 : n28936;
  assign n28938 = pi19 ? n28937 : n37;
  assign n28939 = pi21 ? n157 : n22379;
  assign n28940 = pi20 ? n37 : n28939;
  assign n28941 = pi21 ? n157 : n28497;
  assign n28942 = pi20 ? n28941 : n28498;
  assign n28943 = pi19 ? n28940 : n28942;
  assign n28944 = pi18 ? n28938 : n28943;
  assign n28945 = pi21 ? n28506 : n4094;
  assign n28946 = pi20 ? n685 : n28945;
  assign n28947 = pi19 ? n28946 : n32;
  assign n28948 = pi18 ? n28505 : n28947;
  assign n28949 = pi17 ? n28944 : n28948;
  assign n28950 = pi16 ? n439 : n28949;
  assign n28951 = pi15 ? n28935 : n28950;
  assign n28952 = pi20 ? n28516 : n15197;
  assign n28953 = pi19 ? n28952 : n32;
  assign n28954 = pi18 ? n28515 : n28953;
  assign n28955 = pi17 ? n37 : n28954;
  assign n28956 = pi16 ? n439 : n28955;
  assign n28957 = pi21 ? n19178 : n2320;
  assign n28958 = pi20 ? n28524 : n28957;
  assign n28959 = pi19 ? n28958 : n32;
  assign n28960 = pi18 ? n28523 : n28959;
  assign n28961 = pi17 ? n37 : n28960;
  assign n28962 = pi16 ? n439 : n28961;
  assign n28963 = pi15 ? n28956 : n28962;
  assign n28964 = pi14 ? n28951 : n28963;
  assign n28965 = pi20 ? n99 : n3619;
  assign n28966 = pi19 ? n28965 : n32;
  assign n28967 = pi18 ? n99 : n28966;
  assign n28968 = pi17 ? n99 : n28967;
  assign n28969 = pi16 ? n721 : n28968;
  assign n28970 = pi20 ? n776 : n28024;
  assign n28971 = pi19 ? n28970 : n32;
  assign n28972 = pi18 ? n10010 : n28971;
  assign n28973 = pi17 ? n99 : n28972;
  assign n28974 = pi16 ? n721 : n28973;
  assign n28975 = pi15 ? n28969 : n28974;
  assign n28976 = pi20 ? n99 : n28024;
  assign n28977 = pi19 ? n28976 : n32;
  assign n28978 = pi18 ? n99 : n28977;
  assign n28979 = pi17 ? n99 : n28978;
  assign n28980 = pi16 ? n721 : n28979;
  assign n28981 = pi20 ? n99 : n883;
  assign n28982 = pi19 ? n28981 : n32;
  assign n28983 = pi18 ? n28545 : n28982;
  assign n28984 = pi17 ? n99 : n28983;
  assign n28985 = pi16 ? n721 : n28984;
  assign n28986 = pi15 ? n28980 : n28985;
  assign n28987 = pi14 ? n28975 : n28986;
  assign n28988 = pi13 ? n28964 : n28987;
  assign n28989 = pi22 ? n316 : n2160;
  assign n28990 = pi21 ? n159 : n28989;
  assign n28991 = pi20 ? n26680 : n28990;
  assign n28992 = pi19 ? n139 : n28991;
  assign n28993 = pi21 ? n8632 : n928;
  assign n28994 = pi20 ? n2238 : n28993;
  assign n28995 = pi19 ? n28994 : n32;
  assign n28996 = pi18 ? n28992 : n28995;
  assign n28997 = pi17 ? n26684 : n28996;
  assign n28998 = pi16 ? n24953 : n28997;
  assign n28999 = pi20 ? n18317 : n18386;
  assign n29000 = pi19 ? n28999 : n32;
  assign n29001 = pi18 ? n9111 : n29000;
  assign n29002 = pi17 ? n139 : n29001;
  assign n29003 = pi16 ? n2291 : n29002;
  assign n29004 = pi15 ? n28998 : n29003;
  assign n29005 = pi16 ? n2291 : n28571;
  assign n29006 = pi15 ? n29005 : n28590;
  assign n29007 = pi14 ? n29004 : n29006;
  assign n29008 = pi21 ? n2876 : n346;
  assign n29009 = pi20 ? n204 : n29008;
  assign n29010 = pi19 ? n204 : n29009;
  assign n29011 = pi21 ? n204 : n19302;
  assign n29012 = pi22 ? n316 : n6365;
  assign n29013 = pi21 ? n29012 : n32;
  assign n29014 = pi20 ? n29011 : n29013;
  assign n29015 = pi19 ? n29014 : n32;
  assign n29016 = pi18 ? n29010 : n29015;
  assign n29017 = pi17 ? n204 : n29016;
  assign n29018 = pi16 ? n13493 : n29017;
  assign n29019 = pi15 ? n28610 : n29018;
  assign n29020 = pi20 ? n204 : n1072;
  assign n29021 = pi19 ? n29020 : n32;
  assign n29022 = pi18 ? n204 : n29021;
  assign n29023 = pi17 ? n28621 : n29022;
  assign n29024 = pi16 ? n13846 : n29023;
  assign n29025 = pi20 ? n204 : n19439;
  assign n29026 = pi19 ? n29025 : n32;
  assign n29027 = pi18 ? n204 : n29026;
  assign n29028 = pi17 ? n28630 : n29027;
  assign n29029 = pi16 ? n13833 : n29028;
  assign n29030 = pi15 ? n29024 : n29029;
  assign n29031 = pi14 ? n29019 : n29030;
  assign n29032 = pi13 ? n29007 : n29031;
  assign n29033 = pi12 ? n28988 : n29032;
  assign n29034 = pi22 ? n4079 : n759;
  assign n29035 = pi21 ? n29034 : n32;
  assign n29036 = pi20 ? n1016 : n29035;
  assign n29037 = pi19 ? n29036 : n32;
  assign n29038 = pi18 ? n11765 : n29037;
  assign n29039 = pi17 ? n139 : n29038;
  assign n29040 = pi16 ? n915 : n29039;
  assign n29041 = pi22 ? n3762 : n396;
  assign n29042 = pi21 ? n29041 : n32;
  assign n29043 = pi20 ? n28650 : n29042;
  assign n29044 = pi19 ? n29043 : n32;
  assign n29045 = pi18 ? n28648 : n29044;
  assign n29046 = pi17 ? n335 : n29045;
  assign n29047 = pi16 ? n28647 : n29046;
  assign n29048 = pi15 ? n29040 : n29047;
  assign n29049 = pi20 ? n6377 : n9463;
  assign n29050 = pi19 ? n29049 : n32;
  assign n29051 = pi18 ? n335 : n29050;
  assign n29052 = pi17 ? n335 : n29051;
  assign n29053 = pi16 ? n2035 : n29052;
  assign n29054 = pi20 ? n6377 : n24937;
  assign n29055 = pi19 ? n29054 : n32;
  assign n29056 = pi18 ? n335 : n29055;
  assign n29057 = pi17 ? n335 : n29056;
  assign n29058 = pi16 ? n2425 : n29057;
  assign n29059 = pi15 ? n29053 : n29058;
  assign n29060 = pi14 ? n29048 : n29059;
  assign n29061 = pi22 ? n2121 : n706;
  assign n29062 = pi21 ? n29061 : n32;
  assign n29063 = pi20 ? n28669 : n29062;
  assign n29064 = pi19 ? n29063 : n32;
  assign n29065 = pi18 ? n15438 : n29064;
  assign n29066 = pi17 ? n335 : n29065;
  assign n29067 = pi16 ? n7943 : n29066;
  assign n29068 = pi18 ? n15438 : n18115;
  assign n29069 = pi17 ? n335 : n29068;
  assign n29070 = pi16 ? n7943 : n29069;
  assign n29071 = pi15 ? n29067 : n29070;
  assign n29072 = pi20 ? n28683 : n4110;
  assign n29073 = pi19 ? n29072 : n32;
  assign n29074 = pi18 ? n15438 : n29073;
  assign n29075 = pi17 ? n28682 : n29074;
  assign n29076 = pi16 ? n2035 : n29075;
  assign n29077 = pi18 ? n17540 : n28676;
  assign n29078 = pi17 ? n28692 : n29077;
  assign n29079 = pi16 ? n7943 : n29078;
  assign n29080 = pi15 ? n29076 : n29079;
  assign n29081 = pi14 ? n29071 : n29080;
  assign n29082 = pi13 ? n29060 : n29081;
  assign n29083 = pi20 ? n233 : n4116;
  assign n29084 = pi19 ? n29083 : n32;
  assign n29085 = pi18 ? n233 : n29084;
  assign n29086 = pi17 ? n28708 : n29085;
  assign n29087 = pi16 ? n28705 : n29086;
  assign n29088 = pi18 ? n28719 : n28710;
  assign n29089 = pi17 ? n28717 : n29088;
  assign n29090 = pi16 ? n439 : n29089;
  assign n29091 = pi15 ? n29087 : n29090;
  assign n29092 = pi18 ? n28724 : n27179;
  assign n29093 = pi17 ? n37 : n29092;
  assign n29094 = pi16 ? n439 : n29093;
  assign n29095 = pi15 ? n29094 : n28755;
  assign n29096 = pi14 ? n29091 : n29095;
  assign n29097 = pi20 ? n28769 : n2653;
  assign n29098 = pi19 ? n29097 : n32;
  assign n29099 = pi18 ? n28768 : n29098;
  assign n29100 = pi17 ? n28766 : n29099;
  assign n29101 = pi16 ? n28763 : n29100;
  assign n29102 = pi18 ? n28776 : n28771;
  assign n29103 = pi17 ? n363 : n29102;
  assign n29104 = pi16 ? n21219 : n29103;
  assign n29105 = pi15 ? n29101 : n29104;
  assign n29106 = pi18 ? n363 : n28778;
  assign n29107 = pi17 ? n363 : n29106;
  assign n29108 = pi16 ? n21219 : n29107;
  assign n29109 = pi18 ? n363 : n27220;
  assign n29110 = pi17 ? n363 : n29109;
  assign n29111 = pi16 ? n26062 : n29110;
  assign n29112 = pi15 ? n29108 : n29111;
  assign n29113 = pi14 ? n29105 : n29112;
  assign n29114 = pi13 ? n29096 : n29113;
  assign n29115 = pi12 ? n29082 : n29114;
  assign n29116 = pi11 ? n29033 : n29115;
  assign n29117 = pi10 ? n28929 : n29116;
  assign n29118 = pi09 ? n28182 : n29117;
  assign n29119 = pi08 ? n28798 : n29118;
  assign n29120 = pi20 ? n2974 : n3888;
  assign n29121 = pi19 ? n29120 : n9972;
  assign n29122 = pi19 ? n21611 : n2935;
  assign n29123 = pi18 ? n29121 : n29122;
  assign n29124 = pi17 ? n37 : n29123;
  assign n29125 = pi16 ? n28161 : n29124;
  assign n29126 = pi15 ? n32 : n29125;
  assign n29127 = pi20 ? n14829 : n32;
  assign n29128 = pi19 ? n99 : n29127;
  assign n29129 = pi18 ? n99 : n29128;
  assign n29130 = pi17 ? n99 : n29129;
  assign n29131 = pi16 ? n28169 : n29130;
  assign n29132 = pi22 ? n39 : n20563;
  assign n29133 = pi22 ? n20563 : n37;
  assign n29134 = pi21 ? n29132 : n29133;
  assign n29135 = pi20 ? n32 : n29134;
  assign n29136 = pi19 ? n32 : n29135;
  assign n29137 = pi21 ? n37 : n2168;
  assign n29138 = pi20 ? n37 : n29137;
  assign n29139 = pi19 ? n29138 : n99;
  assign n29140 = pi18 ? n29136 : n29139;
  assign n29141 = pi17 ? n32 : n29140;
  assign n29142 = pi16 ? n29141 : n29130;
  assign n29143 = pi15 ? n29131 : n29142;
  assign n29144 = pi14 ? n29126 : n29143;
  assign n29145 = pi13 ? n32 : n29144;
  assign n29146 = pi12 ? n32 : n29145;
  assign n29147 = pi11 ? n32 : n29146;
  assign n29148 = pi10 ? n32 : n29147;
  assign n29149 = pi19 ? n37 : n14525;
  assign n29150 = pi18 ? n16593 : n29149;
  assign n29151 = pi17 ? n32 : n29150;
  assign n29152 = pi19 ? n23706 : n3806;
  assign n29153 = pi20 ? n3888 : n2755;
  assign n29154 = pi19 ? n29153 : n6043;
  assign n29155 = pi18 ? n29152 : n29154;
  assign n29156 = pi19 ? n18512 : n3825;
  assign n29157 = pi20 ? n14835 : n32;
  assign n29158 = pi19 ? n22702 : n29157;
  assign n29159 = pi18 ? n29156 : n29158;
  assign n29160 = pi17 ? n29155 : n29159;
  assign n29161 = pi16 ? n29151 : n29160;
  assign n29162 = pi19 ? n37 : n18853;
  assign n29163 = pi18 ? n17008 : n29162;
  assign n29164 = pi17 ? n32 : n29163;
  assign n29165 = pi20 ? n99 : n3042;
  assign n29166 = pi19 ? n99 : n29165;
  assign n29167 = pi20 ? n14847 : n32;
  assign n29168 = pi19 ? n10837 : n29167;
  assign n29169 = pi18 ? n29166 : n29168;
  assign n29170 = pi17 ? n99 : n29169;
  assign n29171 = pi16 ? n29164 : n29170;
  assign n29172 = pi15 ? n29161 : n29171;
  assign n29173 = pi20 ? n2983 : n3814;
  assign n29174 = pi19 ? n37 : n29173;
  assign n29175 = pi18 ? n17008 : n29174;
  assign n29176 = pi17 ? n32 : n29175;
  assign n29177 = pi19 ? n21634 : n226;
  assign n29178 = pi19 ? n226 : n99;
  assign n29179 = pi18 ? n29177 : n29178;
  assign n29180 = pi19 ? n17016 : n17972;
  assign n29181 = pi20 ? n15978 : n32;
  assign n29182 = pi19 ? n28196 : n29181;
  assign n29183 = pi18 ? n29180 : n29182;
  assign n29184 = pi17 ? n29179 : n29183;
  assign n29185 = pi16 ? n29176 : n29184;
  assign n29186 = pi19 ? n37 : n3046;
  assign n29187 = pi20 ? n218 : n219;
  assign n29188 = pi19 ? n9972 : n29187;
  assign n29189 = pi18 ? n29186 : n29188;
  assign n29190 = pi20 ? n4617 : n7745;
  assign n29191 = pi20 ? n221 : n23624;
  assign n29192 = pi19 ? n29190 : n29191;
  assign n29193 = pi20 ? n221 : n1658;
  assign n29194 = pi19 ? n29193 : n32;
  assign n29195 = pi18 ? n29192 : n29194;
  assign n29196 = pi17 ? n29189 : n29195;
  assign n29197 = pi16 ? n439 : n29196;
  assign n29198 = pi15 ? n29185 : n29197;
  assign n29199 = pi14 ? n29172 : n29198;
  assign n29200 = pi18 ? n374 : n18854;
  assign n29201 = pi17 ? n32 : n29200;
  assign n29202 = pi16 ? n29201 : n28801;
  assign n29203 = pi20 ? n13612 : n15594;
  assign n29204 = pi20 ? n1743 : n942;
  assign n29205 = pi19 ? n29203 : n29204;
  assign n29206 = pi18 ? n374 : n29205;
  assign n29207 = pi17 ? n32 : n29206;
  assign n29208 = pi19 ? n1804 : n1806;
  assign n29209 = pi18 ? n29208 : n967;
  assign n29210 = pi21 ? n139 : n862;
  assign n29211 = pi20 ? n139 : n29210;
  assign n29212 = pi19 ? n29211 : n32;
  assign n29213 = pi18 ? n139 : n29212;
  assign n29214 = pi17 ? n29209 : n29213;
  assign n29215 = pi16 ? n29207 : n29214;
  assign n29216 = pi15 ? n29202 : n29215;
  assign n29217 = pi20 ? n5257 : n139;
  assign n29218 = pi19 ? n29217 : n139;
  assign n29219 = pi18 ? n28256 : n29218;
  assign n29220 = pi19 ? n3578 : n3626;
  assign n29221 = pi19 ? n12589 : n32;
  assign n29222 = pi18 ? n29220 : n29221;
  assign n29223 = pi17 ? n29219 : n29222;
  assign n29224 = pi16 ? n439 : n29223;
  assign n29225 = pi18 ? n14963 : n28257;
  assign n29226 = pi20 ? n139 : n916;
  assign n29227 = pi19 ? n29226 : n32;
  assign n29228 = pi18 ? n139 : n29227;
  assign n29229 = pi17 ? n29225 : n29228;
  assign n29230 = pi16 ? n439 : n29229;
  assign n29231 = pi15 ? n29224 : n29230;
  assign n29232 = pi14 ? n29216 : n29231;
  assign n29233 = pi13 ? n29199 : n29232;
  assign n29234 = pi19 ? n9824 : n942;
  assign n29235 = pi19 ? n942 : n139;
  assign n29236 = pi18 ? n29234 : n29235;
  assign n29237 = pi20 ? n139 : n3090;
  assign n29238 = pi20 ? n939 : n3096;
  assign n29239 = pi19 ? n29237 : n29238;
  assign n29240 = pi18 ? n29239 : n28804;
  assign n29241 = pi17 ? n29236 : n29240;
  assign n29242 = pi16 ? n439 : n29241;
  assign n29243 = pi19 ? n23761 : n9824;
  assign n29244 = pi18 ? n29243 : n28830;
  assign n29245 = pi17 ? n16094 : n29244;
  assign n29246 = pi16 ? n439 : n29245;
  assign n29247 = pi15 ? n29242 : n29246;
  assign n29248 = pi20 ? n3086 : n947;
  assign n29249 = pi19 ? n37 : n29248;
  assign n29250 = pi18 ? n37 : n29249;
  assign n29251 = pi20 ? n1003 : n3671;
  assign n29252 = pi20 ? n3083 : n3090;
  assign n29253 = pi19 ? n29251 : n29252;
  assign n29254 = pi18 ? n29253 : n28830;
  assign n29255 = pi17 ? n29250 : n29254;
  assign n29256 = pi16 ? n439 : n29255;
  assign n29257 = pi19 ? n37 : n377;
  assign n29258 = pi18 ? n374 : n29257;
  assign n29259 = pi17 ? n32 : n29258;
  assign n29260 = pi20 ? n13147 : n942;
  assign n29261 = pi19 ? n29260 : n942;
  assign n29262 = pi18 ? n18083 : n29261;
  assign n29263 = pi18 ? n7927 : n28835;
  assign n29264 = pi17 ? n29262 : n29263;
  assign n29265 = pi16 ? n29259 : n29264;
  assign n29266 = pi15 ? n29256 : n29265;
  assign n29267 = pi14 ? n29247 : n29266;
  assign n29268 = pi20 ? n3104 : n3083;
  assign n29269 = pi19 ? n29268 : n27331;
  assign n29270 = pi18 ? n29269 : n28835;
  assign n29271 = pi17 ? n18075 : n29270;
  assign n29272 = pi16 ? n439 : n29271;
  assign n29273 = pi20 ? n37 : n13613;
  assign n29274 = pi19 ? n29273 : n17110;
  assign n29275 = pi21 ? n10930 : n14978;
  assign n29276 = pi20 ? n10927 : n29275;
  assign n29277 = pi19 ? n29276 : n32;
  assign n29278 = pi18 ? n29274 : n29277;
  assign n29279 = pi17 ? n37 : n29278;
  assign n29280 = pi16 ? n439 : n29279;
  assign n29281 = pi15 ? n29272 : n29280;
  assign n29282 = pi21 ? n335 : n9900;
  assign n29283 = pi20 ? n335 : n29282;
  assign n29284 = pi19 ? n29283 : n32;
  assign n29285 = pi18 ? n7677 : n29284;
  assign n29286 = pi17 ? n37 : n29285;
  assign n29287 = pi16 ? n439 : n29286;
  assign n29288 = pi21 ? n335 : n22278;
  assign n29289 = pi20 ? n649 : n29288;
  assign n29290 = pi19 ? n29289 : n32;
  assign n29291 = pi18 ? n37 : n29290;
  assign n29292 = pi17 ? n37 : n29291;
  assign n29293 = pi16 ? n439 : n29292;
  assign n29294 = pi15 ? n29287 : n29293;
  assign n29295 = pi14 ? n29281 : n29294;
  assign n29296 = pi13 ? n29267 : n29295;
  assign n29297 = pi12 ? n29233 : n29296;
  assign n29298 = pi21 ? n570 : n28872;
  assign n29299 = pi20 ? n649 : n29298;
  assign n29300 = pi19 ? n29299 : n32;
  assign n29301 = pi18 ? n37 : n29300;
  assign n29302 = pi17 ? n37 : n29301;
  assign n29303 = pi16 ? n439 : n29302;
  assign n29304 = pi20 ? n335 : n15648;
  assign n29305 = pi19 ? n29304 : n32;
  assign n29306 = pi18 ? n37 : n29305;
  assign n29307 = pi17 ? n37 : n29306;
  assign n29308 = pi16 ? n439 : n29307;
  assign n29309 = pi15 ? n29303 : n29308;
  assign n29310 = pi22 ? n335 : n747;
  assign n29311 = pi21 ? n335 : n29310;
  assign n29312 = pi20 ? n335 : n29311;
  assign n29313 = pi19 ? n29312 : n32;
  assign n29314 = pi18 ? n7686 : n29313;
  assign n29315 = pi17 ? n37 : n29314;
  assign n29316 = pi16 ? n439 : n29315;
  assign n29317 = pi20 ? n649 : n4939;
  assign n29318 = pi19 ? n37 : n29317;
  assign n29319 = pi22 ? n37 : n3301;
  assign n29320 = pi21 ? n37 : n29319;
  assign n29321 = pi20 ? n335 : n29320;
  assign n29322 = pi19 ? n29321 : n32;
  assign n29323 = pi18 ? n29318 : n29322;
  assign n29324 = pi17 ? n15129 : n29323;
  assign n29325 = pi16 ? n439 : n29324;
  assign n29326 = pi15 ? n29316 : n29325;
  assign n29327 = pi14 ? n29309 : n29326;
  assign n29328 = pi20 ? n581 : n4971;
  assign n29329 = pi19 ? n3332 : n29328;
  assign n29330 = pi19 ? n4971 : n335;
  assign n29331 = pi18 ? n29329 : n29330;
  assign n29332 = pi19 ? n28367 : n16516;
  assign n29333 = pi22 ? n335 : n3301;
  assign n29334 = pi21 ? n335 : n29333;
  assign n29335 = pi20 ? n335 : n29334;
  assign n29336 = pi19 ? n29335 : n32;
  assign n29337 = pi18 ? n29332 : n29336;
  assign n29338 = pi17 ? n29331 : n29337;
  assign n29339 = pi16 ? n3360 : n29338;
  assign n29340 = pi20 ? n639 : n638;
  assign n29341 = pi19 ? n37 : n29340;
  assign n29342 = pi18 ? n37 : n29341;
  assign n29343 = pi21 ? n6361 : n7658;
  assign n29344 = pi20 ? n335 : n29343;
  assign n29345 = pi19 ? n29344 : n32;
  assign n29346 = pi18 ? n21770 : n29345;
  assign n29347 = pi17 ? n29342 : n29346;
  assign n29348 = pi16 ? n439 : n29347;
  assign n29349 = pi15 ? n29339 : n29348;
  assign n29350 = pi18 ? n37 : n27444;
  assign n29351 = pi20 ? n19422 : n25128;
  assign n29352 = pi19 ? n29351 : n32;
  assign n29353 = pi18 ? n19093 : n29352;
  assign n29354 = pi17 ? n29350 : n29353;
  assign n29355 = pi16 ? n439 : n29354;
  assign n29356 = pi21 ? n3392 : n5015;
  assign n29357 = pi20 ? n37 : n29356;
  assign n29358 = pi19 ? n37 : n29357;
  assign n29359 = pi21 ? n363 : n2091;
  assign n29360 = pi20 ? n29359 : n24081;
  assign n29361 = pi19 ? n29360 : n32;
  assign n29362 = pi18 ? n29358 : n29361;
  assign n29363 = pi17 ? n37 : n29362;
  assign n29364 = pi16 ? n439 : n29363;
  assign n29365 = pi15 ? n29355 : n29364;
  assign n29366 = pi14 ? n29349 : n29365;
  assign n29367 = pi13 ? n29327 : n29366;
  assign n29368 = pi20 ? n37 : n2782;
  assign n29369 = pi19 ? n29368 : n32;
  assign n29370 = pi18 ? n37 : n29369;
  assign n29371 = pi17 ? n37 : n29370;
  assign n29372 = pi16 ? n439 : n29371;
  assign n29373 = pi21 ? n3392 : n1423;
  assign n29374 = pi20 ? n37 : n29373;
  assign n29375 = pi19 ? n29374 : n32;
  assign n29376 = pi18 ? n37 : n29375;
  assign n29377 = pi17 ? n37 : n29376;
  assign n29378 = pi16 ? n439 : n29377;
  assign n29379 = pi15 ? n29372 : n29378;
  assign n29380 = pi19 ? n1410 : n32;
  assign n29381 = pi18 ? n37 : n29380;
  assign n29382 = pi17 ? n37 : n29381;
  assign n29383 = pi16 ? n439 : n29382;
  assign n29384 = pi19 ? n1418 : n32;
  assign n29385 = pi18 ? n37 : n29384;
  assign n29386 = pi17 ? n37 : n29385;
  assign n29387 = pi16 ? n439 : n29386;
  assign n29388 = pi15 ? n29383 : n29387;
  assign n29389 = pi14 ? n29379 : n29388;
  assign n29390 = pi22 ? n3944 : n317;
  assign n29391 = pi21 ? n3392 : n29390;
  assign n29392 = pi20 ? n37 : n29391;
  assign n29393 = pi19 ? n29392 : n32;
  assign n29394 = pi18 ? n37 : n29393;
  assign n29395 = pi17 ? n37 : n29394;
  assign n29396 = pi16 ? n439 : n29395;
  assign n29397 = pi15 ? n29396 : n28905;
  assign n29398 = pi20 ? n9660 : n37;
  assign n29399 = pi19 ? n37 : n29398;
  assign n29400 = pi20 ? n363 : n22881;
  assign n29401 = pi19 ? n5029 : n29400;
  assign n29402 = pi18 ? n29399 : n29401;
  assign n29403 = pi20 ? n24865 : n363;
  assign n29404 = pi19 ? n15173 : n29403;
  assign n29405 = pi20 ? n15173 : n28913;
  assign n29406 = pi19 ? n29405 : n32;
  assign n29407 = pi18 ? n29404 : n29406;
  assign n29408 = pi17 ? n29402 : n29407;
  assign n29409 = pi16 ? n439 : n29408;
  assign n29410 = pi21 ? n20629 : n7723;
  assign n29411 = pi20 ? n37 : n29410;
  assign n29412 = pi19 ? n29411 : n32;
  assign n29413 = pi18 ? n37 : n29412;
  assign n29414 = pi17 ? n37 : n29413;
  assign n29415 = pi16 ? n439 : n29414;
  assign n29416 = pi15 ? n29409 : n29415;
  assign n29417 = pi14 ? n29397 : n29416;
  assign n29418 = pi13 ? n29389 : n29417;
  assign n29419 = pi12 ? n29367 : n29418;
  assign n29420 = pi11 ? n29297 : n29419;
  assign n29421 = pi21 ? n2106 : n14246;
  assign n29422 = pi21 ? n6089 : n7723;
  assign n29423 = pi20 ? n29421 : n29422;
  assign n29424 = pi19 ? n29423 : n32;
  assign n29425 = pi18 ? n2731 : n29424;
  assign n29426 = pi17 ? n37 : n29425;
  assign n29427 = pi16 ? n439 : n29426;
  assign n29428 = pi20 ? n221 : n99;
  assign n29429 = pi19 ? n21611 : n29428;
  assign n29430 = pi18 ? n374 : n29429;
  assign n29431 = pi17 ? n32 : n29430;
  assign n29432 = pi19 ? n2238 : n99;
  assign n29433 = pi21 ? n272 : n99;
  assign n29434 = pi20 ? n7818 : n29433;
  assign n29435 = pi19 ? n20936 : n29434;
  assign n29436 = pi18 ? n29432 : n29435;
  assign n29437 = pi20 ? n219 : n2238;
  assign n29438 = pi20 ? n787 : n7829;
  assign n29439 = pi19 ? n29437 : n29438;
  assign n29440 = pi20 ? n685 : n15197;
  assign n29441 = pi19 ? n29440 : n32;
  assign n29442 = pi18 ? n29439 : n29441;
  assign n29443 = pi17 ? n29436 : n29442;
  assign n29444 = pi16 ? n29431 : n29443;
  assign n29445 = pi15 ? n29427 : n29444;
  assign n29446 = pi20 ? n22666 : n37;
  assign n29447 = pi19 ? n37 : n29446;
  assign n29448 = pi18 ? n374 : n29447;
  assign n29449 = pi17 ? n32 : n29448;
  assign n29450 = pi20 ? n2982 : n14844;
  assign n29451 = pi19 ? n29450 : n5077;
  assign n29452 = pi20 ? n5077 : n7747;
  assign n29453 = pi20 ? n7747 : n15960;
  assign n29454 = pi19 ? n29452 : n29453;
  assign n29455 = pi18 ? n29451 : n29454;
  assign n29456 = pi20 ? n14887 : n7745;
  assign n29457 = pi20 ? n219 : n157;
  assign n29458 = pi19 ? n29456 : n29457;
  assign n29459 = pi20 ? n9747 : n3619;
  assign n29460 = pi19 ? n29459 : n32;
  assign n29461 = pi18 ? n29458 : n29460;
  assign n29462 = pi17 ? n29455 : n29461;
  assign n29463 = pi16 ? n29449 : n29462;
  assign n29464 = pi20 ? n2982 : n14887;
  assign n29465 = pi19 ? n29464 : n28217;
  assign n29466 = pi18 ? n184 : n29465;
  assign n29467 = pi17 ? n32 : n29466;
  assign n29468 = pi20 ? n2973 : n181;
  assign n29469 = pi19 ? n29468 : n5077;
  assign n29470 = pi18 ? n29469 : n29454;
  assign n29471 = pi20 ? n14530 : n7745;
  assign n29472 = pi20 ? n220 : n157;
  assign n29473 = pi19 ? n29471 : n29472;
  assign n29474 = pi21 ? n3562 : n777;
  assign n29475 = pi20 ? n29474 : n17369;
  assign n29476 = pi19 ? n29475 : n32;
  assign n29477 = pi18 ? n29473 : n29476;
  assign n29478 = pi17 ? n29470 : n29477;
  assign n29479 = pi16 ? n29467 : n29478;
  assign n29480 = pi15 ? n29463 : n29479;
  assign n29481 = pi14 ? n29445 : n29480;
  assign n29482 = pi16 ? n744 : n28968;
  assign n29483 = pi21 ? n3562 : n2835;
  assign n29484 = pi20 ? n99 : n29483;
  assign n29485 = pi19 ? n29484 : n32;
  assign n29486 = pi18 ? n10010 : n29485;
  assign n29487 = pi17 ? n99 : n29486;
  assign n29488 = pi16 ? n744 : n29487;
  assign n29489 = pi15 ? n29482 : n29488;
  assign n29490 = pi21 ? n20977 : n2835;
  assign n29491 = pi20 ? n99 : n29490;
  assign n29492 = pi19 ? n29491 : n32;
  assign n29493 = pi18 ? n99 : n29492;
  assign n29494 = pi17 ? n99 : n29493;
  assign n29495 = pi16 ? n744 : n29494;
  assign n29496 = pi20 ? n99 : n15287;
  assign n29497 = pi19 ? n29496 : n32;
  assign n29498 = pi18 ? n28545 : n29497;
  assign n29499 = pi17 ? n99 : n29498;
  assign n29500 = pi16 ? n744 : n29499;
  assign n29501 = pi15 ? n29495 : n29500;
  assign n29502 = pi14 ? n29489 : n29501;
  assign n29503 = pi13 ? n29481 : n29502;
  assign n29504 = pi20 ? n26680 : n22965;
  assign n29505 = pi19 ? n139 : n29504;
  assign n29506 = pi21 ? n20977 : n928;
  assign n29507 = pi20 ? n99 : n29506;
  assign n29508 = pi19 ? n29507 : n32;
  assign n29509 = pi18 ? n29505 : n29508;
  assign n29510 = pi17 ? n26684 : n29509;
  assign n29511 = pi16 ? n25417 : n29510;
  assign n29512 = pi21 ? n139 : n4712;
  assign n29513 = pi20 ? n139 : n29512;
  assign n29514 = pi20 ? n139 : n9773;
  assign n29515 = pi19 ? n29513 : n29514;
  assign n29516 = pi18 ? n139 : n29515;
  assign n29517 = pi17 ? n29516 : n29001;
  assign n29518 = pi16 ? n915 : n29517;
  assign n29519 = pi15 ? n29511 : n29518;
  assign n29520 = pi21 ? n139 : n919;
  assign n29521 = pi20 ? n139 : n29520;
  assign n29522 = pi20 ? n139 : n6208;
  assign n29523 = pi19 ? n29521 : n29522;
  assign n29524 = pi18 ? n139 : n29523;
  assign n29525 = pi21 ? n316 : n1039;
  assign n29526 = pi20 ? n29525 : n1030;
  assign n29527 = pi19 ? n29526 : n32;
  assign n29528 = pi18 ? n11798 : n29527;
  assign n29529 = pi17 ? n29524 : n29528;
  assign n29530 = pi16 ? n915 : n29529;
  assign n29531 = pi19 ? n139 : n13462;
  assign n29532 = pi18 ? n990 : n29531;
  assign n29533 = pi17 ? n32 : n29532;
  assign n29534 = pi20 ? n1906 : n1057;
  assign n29535 = pi19 ? n29534 : n7634;
  assign n29536 = pi20 ? n7634 : n921;
  assign n29537 = pi21 ? n139 : n1578;
  assign n29538 = pi20 ? n1057 : n29537;
  assign n29539 = pi19 ? n29536 : n29538;
  assign n29540 = pi18 ? n29535 : n29539;
  assign n29541 = pi20 ? n26482 : n1063;
  assign n29542 = pi20 ? n2318 : n2353;
  assign n29543 = pi19 ? n29541 : n29542;
  assign n29544 = pi20 ? n316 : n1030;
  assign n29545 = pi19 ? n29544 : n32;
  assign n29546 = pi18 ? n29543 : n29545;
  assign n29547 = pi17 ? n29540 : n29546;
  assign n29548 = pi16 ? n29533 : n29547;
  assign n29549 = pi15 ? n29530 : n29548;
  assign n29550 = pi14 ? n29519 : n29549;
  assign n29551 = pi21 ? n916 : n19302;
  assign n29552 = pi20 ? n204 : n29551;
  assign n29553 = pi19 ? n204 : n29552;
  assign n29554 = pi21 ? n19302 : n921;
  assign n29555 = pi20 ? n29554 : n15370;
  assign n29556 = pi19 ? n29555 : n32;
  assign n29557 = pi18 ? n29553 : n29556;
  assign n29558 = pi17 ? n204 : n29557;
  assign n29559 = pi16 ? n13493 : n29558;
  assign n29560 = pi18 ? n204 : n22273;
  assign n29561 = pi17 ? n204 : n29560;
  assign n29562 = pi16 ? n24565 : n29561;
  assign n29563 = pi15 ? n29559 : n29562;
  assign n29564 = pi20 ? n1063 : n21732;
  assign n29565 = pi19 ? n204 : n29564;
  assign n29566 = pi18 ? n204 : n29565;
  assign n29567 = pi20 ? n204 : n16476;
  assign n29568 = pi19 ? n29567 : n32;
  assign n29569 = pi18 ? n204 : n29568;
  assign n29570 = pi17 ? n29566 : n29569;
  assign n29571 = pi16 ? n13846 : n29570;
  assign n29572 = pi21 ? n297 : n204;
  assign n29573 = pi20 ? n28627 : n29572;
  assign n29574 = pi19 ? n204 : n29573;
  assign n29575 = pi18 ? n204 : n29574;
  assign n29576 = pi17 ? n29575 : n29022;
  assign n29577 = pi16 ? n27650 : n29576;
  assign n29578 = pi15 ? n29571 : n29577;
  assign n29579 = pi14 ? n29563 : n29578;
  assign n29580 = pi13 ? n29550 : n29579;
  assign n29581 = pi12 ? n29503 : n29580;
  assign n29582 = pi20 ? n6577 : n11236;
  assign n29583 = pi19 ? n29582 : n32;
  assign n29584 = pi18 ? n12556 : n29583;
  assign n29585 = pi17 ? n139 : n29584;
  assign n29586 = pi16 ? n915 : n29585;
  assign n29587 = pi18 ? n7941 : n28645;
  assign n29588 = pi17 ? n32 : n29587;
  assign n29589 = pi21 ? n6376 : n1083;
  assign n29590 = pi20 ? n335 : n29589;
  assign n29591 = pi19 ? n335 : n29590;
  assign n29592 = pi21 ? n1929 : n6376;
  assign n29593 = pi20 ? n29592 : n14327;
  assign n29594 = pi19 ? n29593 : n32;
  assign n29595 = pi18 ? n29591 : n29594;
  assign n29596 = pi17 ? n335 : n29595;
  assign n29597 = pi16 ? n29588 : n29596;
  assign n29598 = pi15 ? n29586 : n29597;
  assign n29599 = pi20 ? n28701 : n8917;
  assign n29600 = pi19 ? n29599 : n32;
  assign n29601 = pi18 ? n335 : n29600;
  assign n29602 = pi17 ? n335 : n29601;
  assign n29603 = pi16 ? n7943 : n29602;
  assign n29604 = pi19 ? n335 : n25069;
  assign n29605 = pi20 ? n6377 : n5759;
  assign n29606 = pi19 ? n29605 : n32;
  assign n29607 = pi18 ? n29604 : n29606;
  assign n29608 = pi17 ? n335 : n29607;
  assign n29609 = pi16 ? n2035 : n29608;
  assign n29610 = pi15 ? n29603 : n29609;
  assign n29611 = pi14 ? n29598 : n29610;
  assign n29612 = pi20 ? n2062 : n233;
  assign n29613 = pi19 ? n335 : n29612;
  assign n29614 = pi20 ? n6362 : n6367;
  assign n29615 = pi19 ? n29614 : n32;
  assign n29616 = pi18 ? n29613 : n29615;
  assign n29617 = pi17 ? n335 : n29616;
  assign n29618 = pi16 ? n2035 : n29617;
  assign n29619 = pi20 ? n233 : n7042;
  assign n29620 = pi19 ? n29619 : n32;
  assign n29621 = pi18 ? n15438 : n29620;
  assign n29622 = pi17 ? n335 : n29621;
  assign n29623 = pi16 ? n2035 : n29622;
  assign n29624 = pi15 ? n29618 : n29623;
  assign n29625 = pi21 ? n570 : n4902;
  assign n29626 = pi20 ? n335 : n29625;
  assign n29627 = pi19 ? n29626 : n335;
  assign n29628 = pi18 ? n335 : n29627;
  assign n29629 = pi20 ? n6362 : n4102;
  assign n29630 = pi19 ? n29629 : n32;
  assign n29631 = pi18 ? n15438 : n29630;
  assign n29632 = pi17 ? n29628 : n29631;
  assign n29633 = pi16 ? n2035 : n29632;
  assign n29634 = pi21 ? n335 : n4912;
  assign n29635 = pi20 ? n335 : n29634;
  assign n29636 = pi19 ? n29635 : n612;
  assign n29637 = pi18 ? n335 : n29636;
  assign n29638 = pi20 ? n13527 : n15465;
  assign n29639 = pi19 ? n335 : n29638;
  assign n29640 = pi18 ? n29639 : n19584;
  assign n29641 = pi17 ? n29637 : n29640;
  assign n29642 = pi16 ? n2035 : n29641;
  assign n29643 = pi15 ? n29633 : n29642;
  assign n29644 = pi14 ? n29624 : n29643;
  assign n29645 = pi13 ? n29611 : n29644;
  assign n29646 = pi20 ? n13251 : n335;
  assign n29647 = pi19 ? n8914 : n29646;
  assign n29648 = pi18 ? n7941 : n29647;
  assign n29649 = pi17 ? n32 : n29648;
  assign n29650 = pi21 ? n335 : n19386;
  assign n29651 = pi20 ? n233 : n29650;
  assign n29652 = pi19 ? n233 : n29651;
  assign n29653 = pi18 ? n233 : n29652;
  assign n29654 = pi18 ? n233 : n28676;
  assign n29655 = pi17 ? n29653 : n29654;
  assign n29656 = pi16 ? n29649 : n29655;
  assign n29657 = pi21 ? n8881 : n580;
  assign n29658 = pi20 ? n32 : n29657;
  assign n29659 = pi19 ? n32 : n29658;
  assign n29660 = pi20 ? n3289 : n3292;
  assign n29661 = pi19 ? n29660 : n37;
  assign n29662 = pi18 ? n29659 : n29661;
  assign n29663 = pi17 ? n32 : n29662;
  assign n29664 = pi19 ? n2049 : n3405;
  assign n29665 = pi21 ? n3409 : n26356;
  assign n29666 = pi20 ? n3405 : n29665;
  assign n29667 = pi21 ? n233 : n4891;
  assign n29668 = pi20 ? n29667 : n2094;
  assign n29669 = pi19 ? n29666 : n29668;
  assign n29670 = pi18 ? n29664 : n29669;
  assign n29671 = pi21 ? n2048 : n3404;
  assign n29672 = pi20 ? n21124 : n29671;
  assign n29673 = pi19 ? n29672 : n233;
  assign n29674 = pi18 ? n29673 : n19048;
  assign n29675 = pi17 ? n29670 : n29674;
  assign n29676 = pi16 ? n29663 : n29675;
  assign n29677 = pi15 ? n29656 : n29676;
  assign n29678 = pi18 ? n28724 : n28710;
  assign n29679 = pi17 ? n37 : n29678;
  assign n29680 = pi16 ? n439 : n29679;
  assign n29681 = pi23 ? n21554 : n99;
  assign n29682 = pi22 ? n29681 : n99;
  assign n29683 = pi21 ? n29682 : n363;
  assign n29684 = pi20 ? n32 : n29683;
  assign n29685 = pi19 ? n32 : n29684;
  assign n29686 = pi21 ? n363 : n22549;
  assign n29687 = pi20 ? n722 : n29686;
  assign n29688 = pi22 ? n11047 : n363;
  assign n29689 = pi21 ? n29688 : n99;
  assign n29690 = pi22 ? n4543 : n99;
  assign n29691 = pi21 ? n29690 : n99;
  assign n29692 = pi20 ? n29689 : n29691;
  assign n29693 = pi19 ? n29687 : n29692;
  assign n29694 = pi18 ? n29685 : n29693;
  assign n29695 = pi17 ? n32 : n29694;
  assign n29696 = pi21 ? n14936 : n6089;
  assign n29697 = pi21 ? n14936 : n28746;
  assign n29698 = pi20 ? n29696 : n29697;
  assign n29699 = pi21 ? n5458 : n9196;
  assign n29700 = pi19 ? n29698 : n29699;
  assign n29701 = pi22 ? n5452 : n11047;
  assign n29702 = pi22 ? n685 : n4543;
  assign n29703 = pi21 ? n29701 : n29702;
  assign n29704 = pi20 ? n29699 : n29703;
  assign n29705 = pi22 ? n11047 : n685;
  assign n29706 = pi22 ? n24606 : n5452;
  assign n29707 = pi21 ? n29705 : n29706;
  assign n29708 = pi23 ? n685 : n233;
  assign n29709 = pi22 ? n24606 : n29708;
  assign n29710 = pi21 ? n99 : n29709;
  assign n29711 = pi20 ? n29707 : n29710;
  assign n29712 = pi19 ? n29704 : n29711;
  assign n29713 = pi18 ? n29700 : n29712;
  assign n29714 = pi21 ? n6089 : n14936;
  assign n29715 = pi22 ? n685 : n24606;
  assign n29716 = pi21 ? n29715 : n5458;
  assign n29717 = pi20 ? n29714 : n29716;
  assign n29718 = pi22 ? n233 : n29708;
  assign n29719 = pi21 ? n29718 : n28746;
  assign n29720 = pi22 ? n29708 : n233;
  assign n29721 = pi21 ? n29720 : n28746;
  assign n29722 = pi20 ? n29719 : n29721;
  assign n29723 = pi19 ? n29717 : n29722;
  assign n29724 = pi21 ? n28746 : n685;
  assign n29725 = pi20 ? n29724 : n2638;
  assign n29726 = pi19 ? n29725 : n32;
  assign n29727 = pi18 ? n29723 : n29726;
  assign n29728 = pi17 ? n29713 : n29727;
  assign n29729 = pi16 ? n29695 : n29728;
  assign n29730 = pi15 ? n29680 : n29729;
  assign n29731 = pi14 ? n29677 : n29730;
  assign n29732 = pi22 ? n715 : n363;
  assign n29733 = pi21 ? n29732 : n363;
  assign n29734 = pi20 ? n32 : n29733;
  assign n29735 = pi19 ? n32 : n29734;
  assign n29736 = pi18 ? n29735 : n363;
  assign n29737 = pi17 ? n32 : n29736;
  assign n29738 = pi20 ? n25181 : n363;
  assign n29739 = pi19 ? n363 : n29738;
  assign n29740 = pi18 ? n363 : n29739;
  assign n29741 = pi21 ? n24222 : n685;
  assign n29742 = pi20 ? n29741 : n2653;
  assign n29743 = pi19 ? n29742 : n32;
  assign n29744 = pi18 ? n28768 : n29743;
  assign n29745 = pi17 ? n29740 : n29744;
  assign n29746 = pi16 ? n29737 : n29745;
  assign n29747 = pi18 ? n23174 : n363;
  assign n29748 = pi17 ? n32 : n29747;
  assign n29749 = pi20 ? n363 : n18194;
  assign n29750 = pi19 ? n363 : n29749;
  assign n29751 = pi20 ? n28128 : n1822;
  assign n29752 = pi19 ? n29751 : n32;
  assign n29753 = pi18 ? n29750 : n29752;
  assign n29754 = pi17 ? n363 : n29753;
  assign n29755 = pi16 ? n29748 : n29754;
  assign n29756 = pi15 ? n29746 : n29755;
  assign n29757 = pi21 ? n363 : n3436;
  assign n29758 = pi20 ? n29757 : n32;
  assign n29759 = pi19 ? n29758 : n32;
  assign n29760 = pi18 ? n363 : n29759;
  assign n29761 = pi17 ? n363 : n29760;
  assign n29762 = pi16 ? n26887 : n29761;
  assign n29763 = pi22 ? n2419 : n363;
  assign n29764 = pi21 ? n29763 : n363;
  assign n29765 = pi20 ? n32 : n29764;
  assign n29766 = pi19 ? n32 : n29765;
  assign n29767 = pi18 ? n29766 : n363;
  assign n29768 = pi17 ? n32 : n29767;
  assign n29769 = pi16 ? n29768 : n28787;
  assign n29770 = pi15 ? n29762 : n29769;
  assign n29771 = pi14 ? n29756 : n29770;
  assign n29772 = pi13 ? n29731 : n29771;
  assign n29773 = pi12 ? n29645 : n29772;
  assign n29774 = pi11 ? n29581 : n29773;
  assign n29775 = pi10 ? n29420 : n29774;
  assign n29776 = pi09 ? n29148 : n29775;
  assign n29777 = pi20 ? n5077 : n3888;
  assign n29778 = pi20 ? n99 : n22666;
  assign n29779 = pi19 ? n29777 : n29778;
  assign n29780 = pi19 ? n22685 : n29127;
  assign n29781 = pi18 ? n29779 : n29780;
  assign n29782 = pi17 ? n37 : n29781;
  assign n29783 = pi16 ? n28161 : n29782;
  assign n29784 = pi15 ? n32 : n29783;
  assign n29785 = pi20 ? n37 : n21635;
  assign n29786 = pi19 ? n29785 : n99;
  assign n29787 = pi18 ? n29136 : n29786;
  assign n29788 = pi17 ? n32 : n29787;
  assign n29789 = pi16 ? n29788 : n29130;
  assign n29790 = pi15 ? n29131 : n29789;
  assign n29791 = pi14 ? n29784 : n29790;
  assign n29792 = pi13 ? n32 : n29791;
  assign n29793 = pi12 ? n32 : n29792;
  assign n29794 = pi11 ? n32 : n29793;
  assign n29795 = pi10 ? n32 : n29794;
  assign n29796 = pi20 ? n3814 : n2185;
  assign n29797 = pi19 ? n23706 : n29796;
  assign n29798 = pi20 ? n4619 : n2185;
  assign n29799 = pi19 ? n29798 : n5509;
  assign n29800 = pi18 ? n29797 : n29799;
  assign n29801 = pi17 ? n29800 : n29159;
  assign n29802 = pi16 ? n29151 : n29801;
  assign n29803 = pi15 ? n29802 : n29171;
  assign n29804 = pi14 ? n29803 : n29198;
  assign n29805 = pi18 ? n99 : n28213;
  assign n29806 = pi17 ? n99 : n29805;
  assign n29807 = pi16 ? n29201 : n29806;
  assign n29808 = pi15 ? n29807 : n29215;
  assign n29809 = pi19 ? n12589 : n2555;
  assign n29810 = pi18 ? n29220 : n29809;
  assign n29811 = pi17 ? n29219 : n29810;
  assign n29812 = pi16 ? n439 : n29811;
  assign n29813 = pi19 ? n29226 : n2555;
  assign n29814 = pi18 ? n139 : n29813;
  assign n29815 = pi17 ? n29225 : n29814;
  assign n29816 = pi16 ? n439 : n29815;
  assign n29817 = pi15 ? n29812 : n29816;
  assign n29818 = pi14 ? n29808 : n29817;
  assign n29819 = pi13 ? n29804 : n29818;
  assign n29820 = pi19 ? n139 : n2555;
  assign n29821 = pi18 ? n29239 : n29820;
  assign n29822 = pi17 ? n29236 : n29821;
  assign n29823 = pi16 ? n439 : n29822;
  assign n29824 = pi19 ? n139 : n2680;
  assign n29825 = pi18 ? n29243 : n29824;
  assign n29826 = pi17 ? n16094 : n29825;
  assign n29827 = pi16 ? n439 : n29826;
  assign n29828 = pi15 ? n29823 : n29827;
  assign n29829 = pi18 ? n29253 : n29824;
  assign n29830 = pi17 ? n29250 : n29829;
  assign n29831 = pi16 ? n439 : n29830;
  assign n29832 = pi19 ? n139 : n2702;
  assign n29833 = pi18 ? n7927 : n29832;
  assign n29834 = pi17 ? n29262 : n29833;
  assign n29835 = pi16 ? n29259 : n29834;
  assign n29836 = pi15 ? n29831 : n29835;
  assign n29837 = pi14 ? n29828 : n29836;
  assign n29838 = pi22 ? n139 : n364;
  assign n29839 = pi21 ? n139 : n29838;
  assign n29840 = pi20 ? n139 : n29839;
  assign n29841 = pi19 ? n29840 : n1823;
  assign n29842 = pi18 ? n29269 : n29841;
  assign n29843 = pi17 ? n18075 : n29842;
  assign n29844 = pi16 ? n439 : n29843;
  assign n29845 = pi19 ? n29273 : n12370;
  assign n29846 = pi21 ? n9133 : n9122;
  assign n29847 = pi22 ? n295 : n448;
  assign n29848 = pi21 ? n10930 : n29847;
  assign n29849 = pi20 ? n29846 : n29848;
  assign n29850 = pi19 ? n29849 : n1823;
  assign n29851 = pi18 ? n29845 : n29850;
  assign n29852 = pi17 ? n37 : n29851;
  assign n29853 = pi16 ? n439 : n29852;
  assign n29854 = pi15 ? n29844 : n29853;
  assign n29855 = pi19 ? n29283 : n1823;
  assign n29856 = pi18 ? n7677 : n29855;
  assign n29857 = pi17 ? n37 : n29856;
  assign n29858 = pi16 ? n439 : n29857;
  assign n29859 = pi20 ? n649 : n2062;
  assign n29860 = pi19 ? n29859 : n32;
  assign n29861 = pi18 ? n37 : n29860;
  assign n29862 = pi17 ? n37 : n29861;
  assign n29863 = pi16 ? n439 : n29862;
  assign n29864 = pi15 ? n29858 : n29863;
  assign n29865 = pi14 ? n29854 : n29864;
  assign n29866 = pi13 ? n29837 : n29865;
  assign n29867 = pi12 ? n29819 : n29866;
  assign n29868 = pi22 ? n335 : n686;
  assign n29869 = pi21 ? n570 : n29868;
  assign n29870 = pi20 ? n649 : n29869;
  assign n29871 = pi19 ? n29870 : n32;
  assign n29872 = pi18 ? n37 : n29871;
  assign n29873 = pi17 ? n37 : n29872;
  assign n29874 = pi16 ? n439 : n29873;
  assign n29875 = pi22 ? n335 : n6393;
  assign n29876 = pi21 ? n335 : n29875;
  assign n29877 = pi20 ? n335 : n29876;
  assign n29878 = pi19 ? n29877 : n32;
  assign n29879 = pi18 ? n37 : n29878;
  assign n29880 = pi17 ? n37 : n29879;
  assign n29881 = pi16 ? n439 : n29880;
  assign n29882 = pi15 ? n29874 : n29881;
  assign n29883 = pi14 ? n29882 : n29326;
  assign n29884 = pi13 ? n29883 : n29366;
  assign n29885 = pi21 ? n3392 : n689;
  assign n29886 = pi20 ? n37 : n29885;
  assign n29887 = pi19 ? n29886 : n32;
  assign n29888 = pi18 ? n37 : n29887;
  assign n29889 = pi17 ? n37 : n29888;
  assign n29890 = pi16 ? n439 : n29889;
  assign n29891 = pi15 ? n29396 : n29890;
  assign n29892 = pi20 ? n15173 : n690;
  assign n29893 = pi19 ? n29892 : n32;
  assign n29894 = pi18 ? n29404 : n29893;
  assign n29895 = pi17 ? n29402 : n29894;
  assign n29896 = pi16 ? n439 : n29895;
  assign n29897 = pi21 ? n2957 : n696;
  assign n29898 = pi20 ? n37 : n29897;
  assign n29899 = pi19 ? n29898 : n32;
  assign n29900 = pi18 ? n37 : n29899;
  assign n29901 = pi17 ? n37 : n29900;
  assign n29902 = pi16 ? n439 : n29901;
  assign n29903 = pi15 ? n29896 : n29902;
  assign n29904 = pi14 ? n29891 : n29903;
  assign n29905 = pi13 ? n29389 : n29904;
  assign n29906 = pi12 ? n29884 : n29905;
  assign n29907 = pi11 ? n29867 : n29906;
  assign n29908 = pi21 ? n6089 : n696;
  assign n29909 = pi20 ? n29421 : n29908;
  assign n29910 = pi19 ? n29909 : n32;
  assign n29911 = pi18 ? n2731 : n29910;
  assign n29912 = pi17 ? n37 : n29911;
  assign n29913 = pi16 ? n439 : n29912;
  assign n29914 = pi20 ? n685 : n15729;
  assign n29915 = pi19 ? n29914 : n32;
  assign n29916 = pi18 ? n29439 : n29915;
  assign n29917 = pi17 ? n29436 : n29916;
  assign n29918 = pi16 ? n29431 : n29917;
  assign n29919 = pi15 ? n29913 : n29918;
  assign n29920 = pi20 ? n9747 : n5245;
  assign n29921 = pi19 ? n29920 : n32;
  assign n29922 = pi18 ? n29458 : n29921;
  assign n29923 = pi17 ? n29455 : n29922;
  assign n29924 = pi16 ? n29449 : n29923;
  assign n29925 = pi20 ? n29474 : n3563;
  assign n29926 = pi19 ? n29925 : n32;
  assign n29927 = pi18 ? n29473 : n29926;
  assign n29928 = pi17 ? n29470 : n29927;
  assign n29929 = pi16 ? n29467 : n29928;
  assign n29930 = pi15 ? n29924 : n29929;
  assign n29931 = pi14 ? n29919 : n29930;
  assign n29932 = pi20 ? n99 : n17369;
  assign n29933 = pi19 ? n29932 : n32;
  assign n29934 = pi18 ? n10010 : n29933;
  assign n29935 = pi17 ? n99 : n29934;
  assign n29936 = pi16 ? n721 : n29935;
  assign n29937 = pi15 ? n28969 : n29936;
  assign n29938 = pi21 ? n20977 : n2320;
  assign n29939 = pi20 ? n99 : n29938;
  assign n29940 = pi19 ? n29939 : n32;
  assign n29941 = pi18 ? n99 : n29940;
  assign n29942 = pi17 ? n99 : n29941;
  assign n29943 = pi16 ? n721 : n29942;
  assign n29944 = pi15 ? n29943 : n28985;
  assign n29945 = pi14 ? n29937 : n29944;
  assign n29946 = pi13 ? n29931 : n29945;
  assign n29947 = pi21 ? n20977 : n882;
  assign n29948 = pi20 ? n99 : n29947;
  assign n29949 = pi19 ? n29948 : n32;
  assign n29950 = pi18 ? n29505 : n29949;
  assign n29951 = pi17 ? n26684 : n29950;
  assign n29952 = pi16 ? n24953 : n29951;
  assign n29953 = pi21 ? n204 : n2678;
  assign n29954 = pi20 ? n18317 : n29953;
  assign n29955 = pi19 ? n29954 : n32;
  assign n29956 = pi18 ? n9111 : n29955;
  assign n29957 = pi17 ? n29516 : n29956;
  assign n29958 = pi16 ? n2291 : n29957;
  assign n29959 = pi15 ? n29952 : n29958;
  assign n29960 = pi21 ? n1027 : n2678;
  assign n29961 = pi20 ? n29525 : n29960;
  assign n29962 = pi19 ? n29961 : n32;
  assign n29963 = pi18 ? n11798 : n29962;
  assign n29964 = pi17 ? n29524 : n29963;
  assign n29965 = pi16 ? n2291 : n29964;
  assign n29966 = pi20 ? n316 : n2889;
  assign n29967 = pi19 ? n29966 : n32;
  assign n29968 = pi18 ? n29543 : n29967;
  assign n29969 = pi17 ? n29540 : n29968;
  assign n29970 = pi16 ? n29533 : n29969;
  assign n29971 = pi15 ? n29965 : n29970;
  assign n29972 = pi14 ? n29959 : n29971;
  assign n29973 = pi21 ? n1018 : n2700;
  assign n29974 = pi20 ? n7466 : n29973;
  assign n29975 = pi19 ? n29974 : n32;
  assign n29976 = pi18 ? n29553 : n29975;
  assign n29977 = pi17 ? n204 : n29976;
  assign n29978 = pi16 ? n13493 : n29977;
  assign n29979 = pi20 ? n204 : n17892;
  assign n29980 = pi19 ? n29979 : n32;
  assign n29981 = pi18 ? n204 : n29980;
  assign n29982 = pi17 ? n204 : n29981;
  assign n29983 = pi16 ? n13493 : n29982;
  assign n29984 = pi15 ? n29978 : n29983;
  assign n29985 = pi18 ? n204 : n21695;
  assign n29986 = pi17 ? n29566 : n29985;
  assign n29987 = pi16 ? n13846 : n29986;
  assign n29988 = pi15 ? n29987 : n29577;
  assign n29989 = pi14 ? n29984 : n29988;
  assign n29990 = pi13 ? n29972 : n29989;
  assign n29991 = pi12 ? n29946 : n29990;
  assign n29992 = pi22 ? n204 : n685;
  assign n29993 = pi21 ? n29992 : n32;
  assign n29994 = pi20 ? n6577 : n29993;
  assign n29995 = pi19 ? n29994 : n32;
  assign n29996 = pi18 ? n12556 : n29995;
  assign n29997 = pi17 ? n139 : n29996;
  assign n29998 = pi16 ? n915 : n29997;
  assign n29999 = pi21 ? n4938 : n6376;
  assign n30000 = pi20 ? n29999 : n1101;
  assign n30001 = pi19 ? n30000 : n32;
  assign n30002 = pi18 ? n29591 : n30001;
  assign n30003 = pi17 ? n335 : n30002;
  assign n30004 = pi16 ? n29588 : n30003;
  assign n30005 = pi15 ? n29998 : n30004;
  assign n30006 = pi21 ? n23543 : n32;
  assign n30007 = pi20 ? n28701 : n30006;
  assign n30008 = pi19 ? n30007 : n32;
  assign n30009 = pi18 ? n335 : n30008;
  assign n30010 = pi17 ? n335 : n30009;
  assign n30011 = pi16 ? n7943 : n30010;
  assign n30012 = pi20 ? n6377 : n8917;
  assign n30013 = pi19 ? n30012 : n32;
  assign n30014 = pi18 ? n29604 : n30013;
  assign n30015 = pi17 ? n335 : n30014;
  assign n30016 = pi16 ? n10399 : n30015;
  assign n30017 = pi15 ? n30011 : n30016;
  assign n30018 = pi14 ? n30005 : n30017;
  assign n30019 = pi13 ? n30018 : n29644;
  assign n30020 = pi18 ? n233 : n29620;
  assign n30021 = pi17 ? n29653 : n30020;
  assign n30022 = pi16 ? n29649 : n30021;
  assign n30023 = pi21 ? n180 : n580;
  assign n30024 = pi20 ? n32 : n30023;
  assign n30025 = pi19 ? n32 : n30024;
  assign n30026 = pi19 ? n11632 : n37;
  assign n30027 = pi18 ? n30025 : n30026;
  assign n30028 = pi17 ? n32 : n30027;
  assign n30029 = pi18 ? n29673 : n19584;
  assign n30030 = pi17 ? n29670 : n30029;
  assign n30031 = pi16 ? n30028 : n30030;
  assign n30032 = pi15 ? n30022 : n30031;
  assign n30033 = pi20 ? n233 : n7049;
  assign n30034 = pi19 ? n30033 : n32;
  assign n30035 = pi18 ? n28724 : n30034;
  assign n30036 = pi17 ? n37 : n30035;
  assign n30037 = pi16 ? n439 : n30036;
  assign n30038 = pi18 ? n23149 : n29693;
  assign n30039 = pi17 ? n32 : n30038;
  assign n30040 = pi21 ? n5458 : n29702;
  assign n30041 = pi20 ? n29699 : n30040;
  assign n30042 = pi21 ? n767 : n5453;
  assign n30043 = pi20 ? n30042 : n5454;
  assign n30044 = pi19 ? n30041 : n30043;
  assign n30045 = pi18 ? n29700 : n30044;
  assign n30046 = pi21 ? n6089 : n5458;
  assign n30047 = pi20 ? n14295 : n30046;
  assign n30048 = pi22 ? n15186 : n233;
  assign n30049 = pi21 ? n30048 : n28746;
  assign n30050 = pi20 ? n29719 : n30049;
  assign n30051 = pi19 ? n30047 : n30050;
  assign n30052 = pi20 ? n29724 : n4116;
  assign n30053 = pi19 ? n30052 : n32;
  assign n30054 = pi18 ? n30051 : n30053;
  assign n30055 = pi17 ? n30045 : n30054;
  assign n30056 = pi16 ? n30039 : n30055;
  assign n30057 = pi15 ? n30037 : n30056;
  assign n30058 = pi14 ? n30032 : n30057;
  assign n30059 = pi22 ? n29681 : n363;
  assign n30060 = pi21 ? n30059 : n363;
  assign n30061 = pi20 ? n32 : n30060;
  assign n30062 = pi19 ? n32 : n30061;
  assign n30063 = pi18 ? n30062 : n363;
  assign n30064 = pi17 ? n32 : n30063;
  assign n30065 = pi20 ? n29741 : n10011;
  assign n30066 = pi19 ? n30065 : n32;
  assign n30067 = pi18 ? n28768 : n30066;
  assign n30068 = pi17 ? n29740 : n30067;
  assign n30069 = pi16 ? n30064 : n30068;
  assign n30070 = pi20 ? n28128 : n2653;
  assign n30071 = pi19 ? n30070 : n32;
  assign n30072 = pi18 ? n29750 : n30071;
  assign n30073 = pi17 ? n363 : n30072;
  assign n30074 = pi16 ? n29748 : n30073;
  assign n30075 = pi15 ? n30069 : n30074;
  assign n30076 = pi16 ? n29748 : n29761;
  assign n30077 = pi23 ? n21554 : n335;
  assign n30078 = pi22 ? n30077 : n363;
  assign n30079 = pi21 ? n30078 : n363;
  assign n30080 = pi20 ? n32 : n30079;
  assign n30081 = pi19 ? n32 : n30080;
  assign n30082 = pi18 ? n30081 : n363;
  assign n30083 = pi17 ? n32 : n30082;
  assign n30084 = pi16 ? n30083 : n28787;
  assign n30085 = pi15 ? n30076 : n30084;
  assign n30086 = pi14 ? n30075 : n30085;
  assign n30087 = pi13 ? n30058 : n30086;
  assign n30088 = pi12 ? n30019 : n30087;
  assign n30089 = pi11 ? n29991 : n30088;
  assign n30090 = pi10 ? n29907 : n30089;
  assign n30091 = pi09 ? n29795 : n30090;
  assign n30092 = pi08 ? n29776 : n30091;
  assign n30093 = pi07 ? n29119 : n30092;
  assign n30094 = pi06 ? n28155 : n30093;
  assign n30095 = pi05 ? n26396 : n30094;
  assign n30096 = pi21 ? n29133 : n37;
  assign n30097 = pi20 ? n30096 : n37;
  assign n30098 = pi19 ? n30097 : n222;
  assign n30099 = pi18 ? n28159 : n30098;
  assign n30100 = pi17 ? n32 : n30099;
  assign n30101 = pi19 ? n227 : n3050;
  assign n30102 = pi18 ? n30101 : n4584;
  assign n30103 = pi19 ? n99 : n2991;
  assign n30104 = pi18 ? n99 : n30103;
  assign n30105 = pi17 ? n30102 : n30104;
  assign n30106 = pi16 ? n30100 : n30105;
  assign n30107 = pi15 ? n32 : n30106;
  assign n30108 = pi21 ? n37 : n112;
  assign n30109 = pi20 ? n30096 : n30108;
  assign n30110 = pi19 ? n30109 : n99;
  assign n30111 = pi18 ? n28159 : n30110;
  assign n30112 = pi17 ? n32 : n30111;
  assign n30113 = pi17 ? n99 : n30104;
  assign n30114 = pi16 ? n30112 : n30113;
  assign n30115 = pi23 ? n32 : n20564;
  assign n30116 = pi22 ? n30115 : n20563;
  assign n30117 = pi21 ? n30116 : n20563;
  assign n30118 = pi20 ? n32 : n30117;
  assign n30119 = pi19 ? n32 : n30118;
  assign n30120 = pi21 ? n37 : n29133;
  assign n30121 = pi20 ? n30120 : n14844;
  assign n30122 = pi19 ? n30121 : n99;
  assign n30123 = pi18 ? n30119 : n30122;
  assign n30124 = pi17 ? n32 : n30123;
  assign n30125 = pi19 ? n99 : n3024;
  assign n30126 = pi18 ? n99 : n30125;
  assign n30127 = pi17 ? n99 : n30126;
  assign n30128 = pi16 ? n30124 : n30127;
  assign n30129 = pi15 ? n30114 : n30128;
  assign n30130 = pi14 ? n30107 : n30129;
  assign n30131 = pi13 ? n32 : n30130;
  assign n30132 = pi12 ? n32 : n30131;
  assign n30133 = pi11 ? n32 : n30132;
  assign n30134 = pi10 ? n32 : n30133;
  assign n30135 = pi21 ? n29132 : n20563;
  assign n30136 = pi20 ? n32 : n30135;
  assign n30137 = pi19 ? n32 : n30136;
  assign n30138 = pi20 ? n30096 : n5077;
  assign n30139 = pi19 ? n30138 : n99;
  assign n30140 = pi18 ? n30137 : n30139;
  assign n30141 = pi17 ? n32 : n30140;
  assign n30142 = pi16 ? n30141 : n30127;
  assign n30143 = pi22 ? n64 : n20563;
  assign n30144 = pi21 ? n30143 : n29133;
  assign n30145 = pi20 ? n32 : n30144;
  assign n30146 = pi19 ? n32 : n30145;
  assign n30147 = pi18 ? n30146 : n29162;
  assign n30148 = pi17 ? n32 : n30147;
  assign n30149 = pi19 ? n99 : n3068;
  assign n30150 = pi18 ? n99 : n30149;
  assign n30151 = pi17 ? n99 : n30150;
  assign n30152 = pi16 ? n30148 : n30151;
  assign n30153 = pi15 ? n30142 : n30152;
  assign n30154 = pi23 ? n32 : n20563;
  assign n30155 = pi22 ? n30154 : n20563;
  assign n30156 = pi21 ? n30155 : n29133;
  assign n30157 = pi20 ? n32 : n30156;
  assign n30158 = pi19 ? n32 : n30157;
  assign n30159 = pi20 ? n21635 : n99;
  assign n30160 = pi19 ? n30159 : n99;
  assign n30161 = pi18 ? n30158 : n30160;
  assign n30162 = pi17 ? n32 : n30161;
  assign n30163 = pi20 ? n17032 : n32;
  assign n30164 = pi19 ? n99 : n30163;
  assign n30165 = pi18 ? n99 : n30164;
  assign n30166 = pi17 ? n99 : n30165;
  assign n30167 = pi16 ? n30162 : n30166;
  assign n30168 = pi22 ? n55 : n20563;
  assign n30169 = pi21 ? n30168 : n37;
  assign n30170 = pi20 ? n32 : n30169;
  assign n30171 = pi19 ? n32 : n30170;
  assign n30172 = pi20 ? n21635 : n2968;
  assign n30173 = pi20 ? n3884 : n221;
  assign n30174 = pi19 ? n30172 : n30173;
  assign n30175 = pi18 ? n30171 : n30174;
  assign n30176 = pi17 ? n32 : n30175;
  assign n30177 = pi20 ? n3042 : n219;
  assign n30178 = pi19 ? n227 : n30177;
  assign n30179 = pi18 ? n30178 : n4584;
  assign n30180 = pi19 ? n99 : n29167;
  assign n30181 = pi18 ? n99 : n30180;
  assign n30182 = pi17 ? n30179 : n30181;
  assign n30183 = pi16 ? n30176 : n30182;
  assign n30184 = pi15 ? n30167 : n30183;
  assign n30185 = pi14 ? n30153 : n30184;
  assign n30186 = pi21 ? n2957 : n1143;
  assign n30187 = pi20 ? n30186 : n99;
  assign n30188 = pi19 ? n30187 : n99;
  assign n30189 = pi18 ? n374 : n30188;
  assign n30190 = pi17 ? n32 : n30189;
  assign n30191 = pi19 ? n99 : n29181;
  assign n30192 = pi18 ? n99 : n30191;
  assign n30193 = pi17 ? n99 : n30192;
  assign n30194 = pi16 ? n30190 : n30193;
  assign n30195 = pi23 ? n20563 : n37;
  assign n30196 = pi22 ? n55 : n30195;
  assign n30197 = pi21 ? n30196 : n37;
  assign n30198 = pi20 ? n32 : n30197;
  assign n30199 = pi19 ? n32 : n30198;
  assign n30200 = pi18 ? n30199 : n37;
  assign n30201 = pi17 ? n32 : n30200;
  assign n30202 = pi19 ? n13094 : n15033;
  assign n30203 = pi18 ? n15003 : n30202;
  assign n30204 = pi20 ? n3092 : n3104;
  assign n30205 = pi21 ? n820 : n1531;
  assign n30206 = pi20 ? n30205 : n3645;
  assign n30207 = pi19 ? n30204 : n30206;
  assign n30208 = pi24 ? n139 : n37;
  assign n30209 = pi23 ? n37 : n30208;
  assign n30210 = pi22 ? n139 : n30209;
  assign n30211 = pi21 ? n139 : n30210;
  assign n30212 = pi20 ? n942 : n30211;
  assign n30213 = pi19 ? n30212 : n2471;
  assign n30214 = pi18 ? n30207 : n30213;
  assign n30215 = pi17 ? n30203 : n30214;
  assign n30216 = pi16 ? n30201 : n30215;
  assign n30217 = pi15 ? n30194 : n30216;
  assign n30218 = pi20 ? n8729 : n1704;
  assign n30219 = pi20 ? n13119 : n1694;
  assign n30220 = pi19 ? n30218 : n30219;
  assign n30221 = pi18 ? n374 : n30220;
  assign n30222 = pi17 ? n32 : n30221;
  assign n30223 = pi20 ? n12014 : n15594;
  assign n30224 = pi19 ? n30223 : n1800;
  assign n30225 = pi20 ? n939 : n992;
  assign n30226 = pi19 ? n30225 : n1800;
  assign n30227 = pi18 ? n30224 : n30226;
  assign n30228 = pi20 ? n139 : n1757;
  assign n30229 = pi19 ? n30228 : n139;
  assign n30230 = pi18 ? n30229 : n29820;
  assign n30231 = pi17 ? n30227 : n30230;
  assign n30232 = pi16 ? n30222 : n30231;
  assign n30233 = pi19 ? n8743 : n942;
  assign n30234 = pi18 ? n30233 : n29235;
  assign n30235 = pi20 ? n939 : n3086;
  assign n30236 = pi19 ? n940 : n30235;
  assign n30237 = pi18 ? n30236 : n29820;
  assign n30238 = pi17 ? n30234 : n30237;
  assign n30239 = pi16 ? n439 : n30238;
  assign n30240 = pi15 ? n30232 : n30239;
  assign n30241 = pi14 ? n30217 : n30240;
  assign n30242 = pi13 ? n30185 : n30241;
  assign n30243 = pi18 ? n29243 : n29820;
  assign n30244 = pi17 ? n12372 : n30243;
  assign n30245 = pi16 ? n439 : n30244;
  assign n30246 = pi20 ? n37 : n1743;
  assign n30247 = pi19 ? n37 : n30246;
  assign n30248 = pi18 ? n374 : n30247;
  assign n30249 = pi17 ? n32 : n30248;
  assign n30250 = pi20 ? n13119 : n1693;
  assign n30251 = pi19 ? n30250 : n3604;
  assign n30252 = pi20 ? n1693 : n3645;
  assign n30253 = pi19 ? n30252 : n947;
  assign n30254 = pi18 ? n30251 : n30253;
  assign n30255 = pi21 ? n1211 : n820;
  assign n30256 = pi20 ? n997 : n30255;
  assign n30257 = pi21 ? n139 : n375;
  assign n30258 = pi20 ? n30257 : n3086;
  assign n30259 = pi19 ? n30256 : n30258;
  assign n30260 = pi19 ? n9769 : n2680;
  assign n30261 = pi18 ? n30259 : n30260;
  assign n30262 = pi17 ? n30254 : n30261;
  assign n30263 = pi16 ? n30249 : n30262;
  assign n30264 = pi15 ? n30245 : n30263;
  assign n30265 = pi20 ? n3104 : n939;
  assign n30266 = pi19 ? n37 : n30265;
  assign n30267 = pi18 ? n17061 : n30266;
  assign n30268 = pi20 ? n3086 : n13147;
  assign n30269 = pi19 ? n30268 : n18912;
  assign n30270 = pi18 ? n30269 : n29824;
  assign n30271 = pi17 ? n30267 : n30270;
  assign n30272 = pi16 ? n439 : n30271;
  assign n30273 = pi18 ? n37 : n17061;
  assign n30274 = pi18 ? n17061 : n29832;
  assign n30275 = pi17 ? n30273 : n30274;
  assign n30276 = pi16 ? n439 : n30275;
  assign n30277 = pi15 ? n30272 : n30276;
  assign n30278 = pi14 ? n30264 : n30277;
  assign n30279 = pi20 ? n8707 : n37;
  assign n30280 = pi19 ? n37 : n30279;
  assign n30281 = pi18 ? n374 : n30280;
  assign n30282 = pi17 ? n32 : n30281;
  assign n30283 = pi19 ? n15002 : n10641;
  assign n30284 = pi19 ? n1795 : n2702;
  assign n30285 = pi18 ? n30283 : n30284;
  assign n30286 = pi17 ? n12372 : n30285;
  assign n30287 = pi16 ? n30282 : n30286;
  assign n30288 = pi21 ? n567 : n335;
  assign n30289 = pi20 ? n30288 : n2062;
  assign n30290 = pi19 ? n30289 : n1823;
  assign n30291 = pi18 ? n7677 : n30290;
  assign n30292 = pi17 ? n37 : n30291;
  assign n30293 = pi16 ? n439 : n30292;
  assign n30294 = pi15 ? n30287 : n30293;
  assign n30295 = pi20 ? n577 : n2062;
  assign n30296 = pi19 ? n30295 : n1823;
  assign n30297 = pi18 ? n37 : n30296;
  assign n30298 = pi17 ? n37 : n30297;
  assign n30299 = pi16 ? n439 : n30298;
  assign n30300 = pi21 ? n570 : n2061;
  assign n30301 = pi20 ? n37 : n30300;
  assign n30302 = pi19 ? n30301 : n32;
  assign n30303 = pi18 ? n37 : n30302;
  assign n30304 = pi17 ? n37 : n30303;
  assign n30305 = pi16 ? n439 : n30304;
  assign n30306 = pi15 ? n30299 : n30305;
  assign n30307 = pi14 ? n30294 : n30306;
  assign n30308 = pi13 ? n30278 : n30307;
  assign n30309 = pi12 ? n30242 : n30308;
  assign n30310 = pi19 ? n2095 : n32;
  assign n30311 = pi18 ? n37 : n30310;
  assign n30312 = pi17 ? n37 : n30311;
  assign n30313 = pi16 ? n439 : n30312;
  assign n30314 = pi20 ? n7646 : n4974;
  assign n30315 = pi19 ? n37 : n30314;
  assign n30316 = pi18 ? n37 : n30315;
  assign n30317 = pi20 ? n642 : n9912;
  assign n30318 = pi20 ? n9912 : n639;
  assign n30319 = pi19 ? n30317 : n30318;
  assign n30320 = pi21 ? n569 : n2091;
  assign n30321 = pi20 ? n335 : n30320;
  assign n30322 = pi19 ? n30321 : n32;
  assign n30323 = pi18 ? n30319 : n30322;
  assign n30324 = pi17 ? n30316 : n30323;
  assign n30325 = pi16 ? n439 : n30324;
  assign n30326 = pi15 ? n30313 : n30325;
  assign n30327 = pi20 ? n577 : n6324;
  assign n30328 = pi19 ? n37 : n30327;
  assign n30329 = pi18 ? n37 : n30328;
  assign n30330 = pi19 ? n3330 : n12628;
  assign n30331 = pi20 ? n610 : n2094;
  assign n30332 = pi19 ? n30331 : n32;
  assign n30333 = pi18 ? n30330 : n30332;
  assign n30334 = pi17 ? n30329 : n30333;
  assign n30335 = pi16 ? n439 : n30334;
  assign n30336 = pi20 ? n577 : n610;
  assign n30337 = pi19 ? n37 : n30336;
  assign n30338 = pi18 ? n37 : n30337;
  assign n30339 = pi19 ? n3330 : n23838;
  assign n30340 = pi20 ? n647 : n25125;
  assign n30341 = pi19 ? n30340 : n32;
  assign n30342 = pi18 ? n30339 : n30341;
  assign n30343 = pi17 ? n30338 : n30342;
  assign n30344 = pi16 ? n439 : n30343;
  assign n30345 = pi15 ? n30335 : n30344;
  assign n30346 = pi14 ? n30326 : n30345;
  assign n30347 = pi22 ? n233 : n566;
  assign n30348 = pi21 ? n30347 : n233;
  assign n30349 = pi20 ? n335 : n30348;
  assign n30350 = pi19 ? n30349 : n32;
  assign n30351 = pi18 ? n6374 : n30350;
  assign n30352 = pi17 ? n6339 : n30351;
  assign n30353 = pi16 ? n439 : n30352;
  assign n30354 = pi21 ? n1943 : n233;
  assign n30355 = pi20 ? n30354 : n25965;
  assign n30356 = pi19 ? n30355 : n32;
  assign n30357 = pi18 ? n14149 : n30356;
  assign n30358 = pi17 ? n37 : n30357;
  assign n30359 = pi16 ? n439 : n30358;
  assign n30360 = pi15 ? n30353 : n30359;
  assign n30361 = pi21 ? n233 : n685;
  assign n30362 = pi20 ? n2722 : n30361;
  assign n30363 = pi19 ? n30362 : n32;
  assign n30364 = pi18 ? n37 : n30363;
  assign n30365 = pi17 ? n37 : n30364;
  assign n30366 = pi16 ? n439 : n30365;
  assign n30367 = pi21 ? n2106 : n3445;
  assign n30368 = pi20 ? n15173 : n30367;
  assign n30369 = pi19 ? n30368 : n32;
  assign n30370 = pi18 ? n19093 : n30369;
  assign n30371 = pi17 ? n37 : n30370;
  assign n30372 = pi16 ? n439 : n30371;
  assign n30373 = pi15 ? n30366 : n30372;
  assign n30374 = pi14 ? n30360 : n30373;
  assign n30375 = pi13 ? n30346 : n30374;
  assign n30376 = pi21 ? n3392 : n3436;
  assign n30377 = pi20 ? n15173 : n30376;
  assign n30378 = pi19 ? n30377 : n32;
  assign n30379 = pi18 ? n5030 : n30378;
  assign n30380 = pi17 ? n37 : n30379;
  assign n30381 = pi16 ? n439 : n30380;
  assign n30382 = pi19 ? n2141 : n32;
  assign n30383 = pi18 ? n37 : n30382;
  assign n30384 = pi17 ? n37 : n30383;
  assign n30385 = pi16 ? n439 : n30384;
  assign n30386 = pi15 ? n30381 : n30385;
  assign n30387 = pi14 ? n30386 : n30385;
  assign n30388 = pi20 ? n3393 : n27520;
  assign n30389 = pi19 ? n37 : n30388;
  assign n30390 = pi22 ? n363 : n396;
  assign n30391 = pi21 ? n37 : n30390;
  assign n30392 = pi20 ? n22881 : n30391;
  assign n30393 = pi19 ? n30392 : n32;
  assign n30394 = pi18 ? n30389 : n30393;
  assign n30395 = pi17 ? n37 : n30394;
  assign n30396 = pi16 ? n439 : n30395;
  assign n30397 = pi20 ? n15173 : n9660;
  assign n30398 = pi19 ? n37 : n30397;
  assign n30399 = pi18 ? n37 : n30398;
  assign n30400 = pi20 ? n7730 : n27520;
  assign n30401 = pi19 ? n37 : n30400;
  assign n30402 = pi20 ? n363 : n25531;
  assign n30403 = pi19 ? n30402 : n32;
  assign n30404 = pi18 ? n30401 : n30403;
  assign n30405 = pi17 ? n30399 : n30404;
  assign n30406 = pi16 ? n439 : n30405;
  assign n30407 = pi15 ? n30396 : n30406;
  assign n30408 = pi21 ? n37 : n22919;
  assign n30409 = pi20 ? n37 : n30408;
  assign n30410 = pi19 ? n30409 : n32;
  assign n30411 = pi18 ? n37 : n30410;
  assign n30412 = pi17 ? n37 : n30411;
  assign n30413 = pi16 ? n439 : n30412;
  assign n30414 = pi21 ? n157 : n37;
  assign n30415 = pi20 ? n30414 : n30408;
  assign n30416 = pi19 ? n30415 : n32;
  assign n30417 = pi18 ? n37 : n30416;
  assign n30418 = pi17 ? n37 : n30417;
  assign n30419 = pi16 ? n439 : n30418;
  assign n30420 = pi15 ? n30413 : n30419;
  assign n30421 = pi14 ? n30407 : n30420;
  assign n30422 = pi13 ? n30387 : n30421;
  assign n30423 = pi12 ? n30375 : n30422;
  assign n30424 = pi11 ? n30309 : n30423;
  assign n30425 = pi20 ? n37 : n16279;
  assign n30426 = pi19 ? n37 : n30425;
  assign n30427 = pi18 ? n30426 : n29915;
  assign n30428 = pi17 ? n37 : n30427;
  assign n30429 = pi16 ? n439 : n30428;
  assign n30430 = pi21 ? n796 : n218;
  assign n30431 = pi20 ? n32 : n30430;
  assign n30432 = pi19 ? n32 : n30431;
  assign n30433 = pi18 ? n30432 : n99;
  assign n30434 = pi17 ? n32 : n30433;
  assign n30435 = pi20 ? n99 : n21852;
  assign n30436 = pi19 ? n99 : n30435;
  assign n30437 = pi21 ? n6089 : n8341;
  assign n30438 = pi21 ? n19153 : n3494;
  assign n30439 = pi20 ? n30437 : n30438;
  assign n30440 = pi19 ? n30439 : n32;
  assign n30441 = pi18 ? n30436 : n30440;
  assign n30442 = pi17 ? n99 : n30441;
  assign n30443 = pi16 ? n30434 : n30442;
  assign n30444 = pi15 ? n30429 : n30443;
  assign n30445 = pi21 ? n157 : n20977;
  assign n30446 = pi20 ? n30445 : n3563;
  assign n30447 = pi19 ? n30446 : n32;
  assign n30448 = pi18 ? n9985 : n30447;
  assign n30449 = pi17 ? n99 : n30448;
  assign n30450 = pi16 ? n201 : n30449;
  assign n30451 = pi19 ? n99 : n27596;
  assign n30452 = pi21 ? n20977 : n3523;
  assign n30453 = pi20 ? n99 : n30452;
  assign n30454 = pi19 ? n30453 : n32;
  assign n30455 = pi18 ? n30451 : n30454;
  assign n30456 = pi17 ? n99 : n30455;
  assign n30457 = pi16 ? n801 : n30456;
  assign n30458 = pi15 ? n30450 : n30457;
  assign n30459 = pi14 ? n30444 : n30458;
  assign n30460 = pi16 ? n744 : n29942;
  assign n30461 = pi21 ? n777 : n2320;
  assign n30462 = pi20 ? n99 : n30461;
  assign n30463 = pi19 ? n30462 : n32;
  assign n30464 = pi18 ? n99 : n30463;
  assign n30465 = pi17 ? n99 : n30464;
  assign n30466 = pi16 ? n744 : n30465;
  assign n30467 = pi15 ? n30460 : n30466;
  assign n30468 = pi19 ? n99 : n22704;
  assign n30469 = pi18 ? n742 : n30468;
  assign n30470 = pi17 ? n32 : n30469;
  assign n30471 = pi19 ? n139 : n26682;
  assign n30472 = pi18 ? n139 : n30471;
  assign n30473 = pi20 ? n139 : n99;
  assign n30474 = pi19 ? n139 : n30473;
  assign n30475 = pi21 ? n316 : n99;
  assign n30476 = pi20 ? n30475 : n30461;
  assign n30477 = pi19 ? n30476 : n32;
  assign n30478 = pi18 ? n30474 : n30477;
  assign n30479 = pi17 ? n30472 : n30478;
  assign n30480 = pi16 ? n30470 : n30479;
  assign n30481 = pi20 ? n139 : n19208;
  assign n30482 = pi19 ? n139 : n30481;
  assign n30483 = pi20 ? n316 : n2330;
  assign n30484 = pi19 ? n30483 : n32;
  assign n30485 = pi18 ? n30482 : n30484;
  assign n30486 = pi17 ? n30472 : n30485;
  assign n30487 = pi16 ? n30470 : n30486;
  assign n30488 = pi15 ? n30480 : n30487;
  assign n30489 = pi14 ? n30467 : n30488;
  assign n30490 = pi13 ? n30459 : n30489;
  assign n30491 = pi18 ? n10078 : n30484;
  assign n30492 = pi17 ? n139 : n30491;
  assign n30493 = pi16 ? n915 : n30492;
  assign n30494 = pi20 ? n347 : n4437;
  assign n30495 = pi19 ? n139 : n30494;
  assign n30496 = pi20 ? n316 : n980;
  assign n30497 = pi19 ? n30496 : n32;
  assign n30498 = pi18 ? n30495 : n30497;
  assign n30499 = pi17 ? n139 : n30498;
  assign n30500 = pi16 ? n915 : n30499;
  assign n30501 = pi15 ? n30493 : n30500;
  assign n30502 = pi20 ? n922 : n976;
  assign n30503 = pi19 ? n1795 : n30502;
  assign n30504 = pi18 ? n29531 : n30503;
  assign n30505 = pi20 ? n6568 : n1016;
  assign n30506 = pi19 ? n30505 : n18327;
  assign n30507 = pi18 ? n30506 : n30497;
  assign n30508 = pi17 ? n30504 : n30507;
  assign n30509 = pi16 ? n331 : n30508;
  assign n30510 = pi20 ? n942 : n297;
  assign n30511 = pi19 ? n30510 : n24974;
  assign n30512 = pi18 ? n913 : n30511;
  assign n30513 = pi17 ? n32 : n30512;
  assign n30514 = pi19 ? n26742 : n2318;
  assign n30515 = pi21 ? n346 : n1860;
  assign n30516 = pi20 ? n204 : n30515;
  assign n30517 = pi19 ? n15398 : n30516;
  assign n30518 = pi18 ? n30514 : n30517;
  assign n30519 = pi20 ? n6158 : n2353;
  assign n30520 = pi19 ? n204 : n30519;
  assign n30521 = pi19 ? n2378 : n32;
  assign n30522 = pi18 ? n30520 : n30521;
  assign n30523 = pi17 ? n30518 : n30522;
  assign n30524 = pi16 ? n30513 : n30523;
  assign n30525 = pi15 ? n30509 : n30524;
  assign n30526 = pi14 ? n30501 : n30525;
  assign n30527 = pi20 ? n1026 : n5199;
  assign n30528 = pi19 ? n30527 : n204;
  assign n30529 = pi18 ? n3597 : n30528;
  assign n30530 = pi17 ? n32 : n30529;
  assign n30531 = pi21 ? n204 : n2700;
  assign n30532 = pi20 ? n204 : n30531;
  assign n30533 = pi19 ? n30532 : n32;
  assign n30534 = pi18 ? n204 : n30533;
  assign n30535 = pi17 ? n204 : n30534;
  assign n30536 = pi16 ? n30530 : n30535;
  assign n30537 = pi20 ? n8154 : n5229;
  assign n30538 = pi19 ? n30537 : n204;
  assign n30539 = pi18 ? n913 : n30538;
  assign n30540 = pi17 ? n32 : n30539;
  assign n30541 = pi20 ? n204 : n23406;
  assign n30542 = pi19 ? n30541 : n32;
  assign n30543 = pi18 ? n204 : n30542;
  assign n30544 = pi17 ? n204 : n30543;
  assign n30545 = pi16 ? n30540 : n30544;
  assign n30546 = pi15 ? n30536 : n30545;
  assign n30547 = pi21 ? n326 : n37;
  assign n30548 = pi20 ? n32 : n30547;
  assign n30549 = pi19 ? n32 : n30548;
  assign n30550 = pi20 ? n939 : n1003;
  assign n30551 = pi19 ? n30550 : n998;
  assign n30552 = pi18 ? n30549 : n30551;
  assign n30553 = pi17 ? n32 : n30552;
  assign n30554 = pi19 ? n139 : n940;
  assign n30555 = pi18 ? n139 : n30554;
  assign n30556 = pi19 ? n139 : n16473;
  assign n30557 = pi18 ? n30556 : n30542;
  assign n30558 = pi17 ? n30555 : n30557;
  assign n30559 = pi16 ? n30553 : n30558;
  assign n30560 = pi18 ? n329 : n22746;
  assign n30561 = pi17 ? n32 : n30560;
  assign n30562 = pi21 ? n139 : n3073;
  assign n30563 = pi20 ? n139 : n30562;
  assign n30564 = pi19 ? n139 : n30563;
  assign n30565 = pi18 ? n139 : n30564;
  assign n30566 = pi20 ? n204 : n29993;
  assign n30567 = pi19 ? n30566 : n32;
  assign n30568 = pi18 ? n30556 : n30567;
  assign n30569 = pi17 ? n30565 : n30568;
  assign n30570 = pi16 ? n30561 : n30569;
  assign n30571 = pi15 ? n30559 : n30570;
  assign n30572 = pi14 ? n30546 : n30571;
  assign n30573 = pi13 ? n30526 : n30572;
  assign n30574 = pi12 ? n30490 : n30573;
  assign n30575 = pi21 ? n326 : n295;
  assign n30576 = pi20 ? n32 : n30575;
  assign n30577 = pi19 ? n32 : n30576;
  assign n30578 = pi21 ? n1043 : n375;
  assign n30579 = pi20 ? n30578 : n15594;
  assign n30580 = pi20 ? n12014 : n1699;
  assign n30581 = pi19 ? n30579 : n30580;
  assign n30582 = pi18 ? n30577 : n30581;
  assign n30583 = pi17 ? n32 : n30582;
  assign n30584 = pi21 ? n9144 : n375;
  assign n30585 = pi19 ? n26781 : n30584;
  assign n30586 = pi20 ? n30584 : n26785;
  assign n30587 = pi21 ? n25048 : n9122;
  assign n30588 = pi20 ? n30587 : n26768;
  assign n30589 = pi19 ? n30586 : n30588;
  assign n30590 = pi18 ? n30585 : n30589;
  assign n30591 = pi21 ? n9126 : n1698;
  assign n30592 = pi20 ? n30591 : n25044;
  assign n30593 = pi21 ? n916 : n11808;
  assign n30594 = pi20 ? n9141 : n30593;
  assign n30595 = pi19 ? n30592 : n30594;
  assign n30596 = pi21 ? n28649 : n9144;
  assign n30597 = pi20 ? n30596 : n29993;
  assign n30598 = pi19 ? n30597 : n32;
  assign n30599 = pi18 ? n30595 : n30598;
  assign n30600 = pi17 ? n30590 : n30599;
  assign n30601 = pi16 ? n30583 : n30600;
  assign n30602 = pi20 ? n604 : n571;
  assign n30603 = pi19 ? n30602 : n335;
  assign n30604 = pi18 ? n602 : n30603;
  assign n30605 = pi17 ? n32 : n30604;
  assign n30606 = pi21 ? n25977 : n32;
  assign n30607 = pi20 ? n7980 : n30606;
  assign n30608 = pi19 ? n30607 : n32;
  assign n30609 = pi18 ? n17487 : n30608;
  assign n30610 = pi17 ? n335 : n30609;
  assign n30611 = pi16 ? n30605 : n30610;
  assign n30612 = pi15 ? n30601 : n30611;
  assign n30613 = pi19 ? n28367 : n10957;
  assign n30614 = pi18 ? n602 : n30613;
  assign n30615 = pi17 ? n32 : n30614;
  assign n30616 = pi19 ? n335 : n647;
  assign n30617 = pi19 ? n2073 : n335;
  assign n30618 = pi18 ? n30616 : n30617;
  assign n30619 = pi20 ? n15457 : n30006;
  assign n30620 = pi19 ? n30619 : n32;
  assign n30621 = pi18 ? n17487 : n30620;
  assign n30622 = pi17 ? n30618 : n30621;
  assign n30623 = pi16 ? n30615 : n30622;
  assign n30624 = pi19 ? n14166 : n10957;
  assign n30625 = pi18 ? n3349 : n30624;
  assign n30626 = pi17 ? n32 : n30625;
  assign n30627 = pi20 ? n642 : n647;
  assign n30628 = pi19 ? n612 : n30627;
  assign n30629 = pi20 ? n603 : n604;
  assign n30630 = pi19 ? n2073 : n30629;
  assign n30631 = pi18 ? n30628 : n30630;
  assign n30632 = pi20 ? n603 : n18121;
  assign n30633 = pi19 ? n4984 : n30632;
  assign n30634 = pi20 ? n7980 : n8917;
  assign n30635 = pi19 ? n30634 : n32;
  assign n30636 = pi18 ? n30633 : n30635;
  assign n30637 = pi17 ? n30631 : n30636;
  assign n30638 = pi16 ? n30626 : n30637;
  assign n30639 = pi15 ? n30623 : n30638;
  assign n30640 = pi14 ? n30612 : n30639;
  assign n30641 = pi20 ? n569 : n603;
  assign n30642 = pi19 ? n335 : n30641;
  assign n30643 = pi18 ? n12625 : n30642;
  assign n30644 = pi17 ? n32 : n30643;
  assign n30645 = pi19 ? n603 : n335;
  assign n30646 = pi18 ? n30645 : n335;
  assign n30647 = pi20 ? n233 : n15446;
  assign n30648 = pi19 ? n30647 : n32;
  assign n30649 = pi18 ? n19406 : n30648;
  assign n30650 = pi17 ? n30646 : n30649;
  assign n30651 = pi16 ? n30644 : n30650;
  assign n30652 = pi19 ? n7685 : n19379;
  assign n30653 = pi18 ? n374 : n30652;
  assign n30654 = pi17 ? n32 : n30653;
  assign n30655 = pi20 ? n604 : n577;
  assign n30656 = pi19 ? n30655 : n6341;
  assign n30657 = pi21 ? n2048 : n569;
  assign n30658 = pi20 ? n15469 : n30657;
  assign n30659 = pi19 ? n4984 : n30658;
  assign n30660 = pi18 ? n30656 : n30659;
  assign n30661 = pi20 ? n642 : n610;
  assign n30662 = pi19 ? n30661 : n13532;
  assign n30663 = pi20 ? n233 : n5759;
  assign n30664 = pi19 ? n30663 : n32;
  assign n30665 = pi18 ? n30662 : n30664;
  assign n30666 = pi17 ? n30660 : n30665;
  assign n30667 = pi16 ? n30654 : n30666;
  assign n30668 = pi15 ? n30651 : n30667;
  assign n30669 = pi18 ? n9556 : n4985;
  assign n30670 = pi17 ? n32 : n30669;
  assign n30671 = pi20 ? n21124 : n605;
  assign n30672 = pi19 ? n612 : n30671;
  assign n30673 = pi20 ? n605 : n647;
  assign n30674 = pi21 ? n2048 : n335;
  assign n30675 = pi20 ? n30657 : n30674;
  assign n30676 = pi19 ? n30673 : n30675;
  assign n30677 = pi18 ? n30672 : n30676;
  assign n30678 = pi20 ? n3335 : n13527;
  assign n30679 = pi19 ? n30678 : n19358;
  assign n30680 = pi18 ? n30679 : n30664;
  assign n30681 = pi17 ? n30677 : n30680;
  assign n30682 = pi16 ? n30670 : n30681;
  assign n30683 = pi21 ? n10394 : n569;
  assign n30684 = pi20 ? n32 : n30683;
  assign n30685 = pi19 ? n32 : n30684;
  assign n30686 = pi20 ? n604 : n3335;
  assign n30687 = pi19 ? n605 : n30686;
  assign n30688 = pi18 ? n30685 : n30687;
  assign n30689 = pi17 ? n32 : n30688;
  assign n30690 = pi21 ? n30347 : n567;
  assign n30691 = pi20 ? n30690 : n2004;
  assign n30692 = pi19 ? n7591 : n30691;
  assign n30693 = pi21 ? n569 : n2061;
  assign n30694 = pi20 ? n2004 : n30693;
  assign n30695 = pi20 ? n610 : n30288;
  assign n30696 = pi19 ? n30694 : n30695;
  assign n30697 = pi18 ? n30692 : n30696;
  assign n30698 = pi20 ? n6377 : n233;
  assign n30699 = pi19 ? n24115 : n30698;
  assign n30700 = pi22 ? n233 : n3935;
  assign n30701 = pi21 ? n233 : n30700;
  assign n30702 = pi20 ? n30701 : n7724;
  assign n30703 = pi19 ? n30702 : n32;
  assign n30704 = pi18 ? n30699 : n30703;
  assign n30705 = pi17 ? n30697 : n30704;
  assign n30706 = pi16 ? n30689 : n30705;
  assign n30707 = pi15 ? n30682 : n30706;
  assign n30708 = pi14 ? n30668 : n30707;
  assign n30709 = pi13 ? n30640 : n30708;
  assign n30710 = pi21 ? n574 : n580;
  assign n30711 = pi20 ? n30710 : n638;
  assign n30712 = pi20 ? n604 : n27730;
  assign n30713 = pi19 ? n30711 : n30712;
  assign n30714 = pi18 ? n558 : n30713;
  assign n30715 = pi17 ? n32 : n30714;
  assign n30716 = pi21 ? n570 : n6376;
  assign n30717 = pi20 ? n30716 : n21150;
  assign n30718 = pi21 ? n233 : n567;
  assign n30719 = pi21 ? n560 : n567;
  assign n30720 = pi20 ? n30718 : n30719;
  assign n30721 = pi19 ? n30717 : n30720;
  assign n30722 = pi21 ? n2048 : n567;
  assign n30723 = pi20 ? n30722 : n233;
  assign n30724 = pi21 ? n233 : n2007;
  assign n30725 = pi20 ? n233 : n30724;
  assign n30726 = pi19 ? n30723 : n30725;
  assign n30727 = pi18 ? n30721 : n30726;
  assign n30728 = pi21 ? n233 : n30347;
  assign n30729 = pi20 ? n30728 : n16544;
  assign n30730 = pi19 ? n30729 : n233;
  assign n30731 = pi20 ? n233 : n7724;
  assign n30732 = pi19 ? n30731 : n32;
  assign n30733 = pi18 ? n30730 : n30732;
  assign n30734 = pi17 ? n30727 : n30733;
  assign n30735 = pi16 ? n30715 : n30734;
  assign n30736 = pi19 ? n7717 : n37;
  assign n30737 = pi21 ? n560 : n2091;
  assign n30738 = pi20 ? n37 : n30737;
  assign n30739 = pi19 ? n30738 : n2050;
  assign n30740 = pi18 ? n30736 : n30739;
  assign n30741 = pi21 ? n2091 : n4891;
  assign n30742 = pi20 ? n21124 : n30741;
  assign n30743 = pi20 ? n17777 : n233;
  assign n30744 = pi19 ? n30742 : n30743;
  assign n30745 = pi20 ? n233 : n3210;
  assign n30746 = pi19 ? n30745 : n32;
  assign n30747 = pi18 ? n30744 : n30746;
  assign n30748 = pi17 ? n30740 : n30747;
  assign n30749 = pi16 ? n439 : n30748;
  assign n30750 = pi15 ? n30735 : n30749;
  assign n30751 = pi21 ? n685 : n28746;
  assign n30752 = pi20 ? n2094 : n30751;
  assign n30753 = pi19 ? n37 : n30752;
  assign n30754 = pi20 ? n30361 : n3210;
  assign n30755 = pi19 ? n30754 : n32;
  assign n30756 = pi18 ? n30753 : n30755;
  assign n30757 = pi17 ? n37 : n30756;
  assign n30758 = pi16 ? n439 : n30757;
  assign n30759 = pi22 ? n715 : n4543;
  assign n30760 = pi21 ? n30759 : n99;
  assign n30761 = pi20 ? n32 : n30760;
  assign n30762 = pi19 ? n32 : n30761;
  assign n30763 = pi21 ? n29690 : n22549;
  assign n30764 = pi20 ? n30763 : n28732;
  assign n30765 = pi21 ? n22557 : n99;
  assign n30766 = pi21 ? n22549 : n99;
  assign n30767 = pi20 ? n30765 : n30766;
  assign n30768 = pi19 ? n30764 : n30767;
  assign n30769 = pi18 ? n30762 : n30768;
  assign n30770 = pi17 ? n32 : n30769;
  assign n30771 = pi21 ? n22549 : n5453;
  assign n30772 = pi20 ? n30766 : n30771;
  assign n30773 = pi21 ? n99 : n29690;
  assign n30774 = pi19 ? n30772 : n30773;
  assign n30775 = pi21 ? n22549 : n767;
  assign n30776 = pi20 ? n30773 : n30775;
  assign n30777 = pi21 ? n22549 : n6089;
  assign n30778 = pi21 ? n4551 : n99;
  assign n30779 = pi20 ? n30777 : n30778;
  assign n30780 = pi19 ? n30776 : n30779;
  assign n30781 = pi18 ? n30774 : n30780;
  assign n30782 = pi21 ? n5458 : n22549;
  assign n30783 = pi20 ? n30782 : n30042;
  assign n30784 = pi22 ? n99 : n15186;
  assign n30785 = pi21 ? n3444 : n30784;
  assign n30786 = pi20 ? n30785 : n685;
  assign n30787 = pi19 ? n30783 : n30786;
  assign n30788 = pi22 ? n685 : n15186;
  assign n30789 = pi21 ? n30788 : n685;
  assign n30790 = pi20 ? n30789 : n4116;
  assign n30791 = pi19 ? n30790 : n32;
  assign n30792 = pi18 ? n30787 : n30791;
  assign n30793 = pi17 ? n30781 : n30792;
  assign n30794 = pi16 ? n30770 : n30793;
  assign n30795 = pi15 ? n30758 : n30794;
  assign n30796 = pi14 ? n30750 : n30795;
  assign n30797 = pi18 ? n23149 : n363;
  assign n30798 = pi17 ? n32 : n30797;
  assign n30799 = pi19 ? n363 : n27800;
  assign n30800 = pi20 ? n24223 : n10011;
  assign n30801 = pi19 ? n30800 : n32;
  assign n30802 = pi18 ? n30799 : n30801;
  assign n30803 = pi17 ? n363 : n30802;
  assign n30804 = pi16 ? n30798 : n30803;
  assign n30805 = pi20 ? n363 : n26905;
  assign n30806 = pi19 ? n363 : n30805;
  assign n30807 = pi22 ? n363 : n2299;
  assign n30808 = pi21 ? n363 : n30807;
  assign n30809 = pi20 ? n30808 : n2653;
  assign n30810 = pi19 ? n30809 : n32;
  assign n30811 = pi18 ? n30806 : n30810;
  assign n30812 = pi17 ? n363 : n30811;
  assign n30813 = pi16 ? n21219 : n30812;
  assign n30814 = pi15 ? n30804 : n30813;
  assign n30815 = pi20 ? n30808 : n32;
  assign n30816 = pi19 ? n30815 : n32;
  assign n30817 = pi18 ? n363 : n30816;
  assign n30818 = pi17 ? n363 : n30817;
  assign n30819 = pi16 ? n21219 : n30818;
  assign n30820 = pi22 ? n363 : n6415;
  assign n30821 = pi21 ? n685 : n30820;
  assign n30822 = pi20 ? n30821 : n32;
  assign n30823 = pi19 ? n30822 : n32;
  assign n30824 = pi18 ? n363 : n30823;
  assign n30825 = pi17 ? n363 : n30824;
  assign n30826 = pi16 ? n26062 : n30825;
  assign n30827 = pi15 ? n30819 : n30826;
  assign n30828 = pi14 ? n30814 : n30827;
  assign n30829 = pi13 ? n30796 : n30828;
  assign n30830 = pi12 ? n30709 : n30829;
  assign n30831 = pi11 ? n30574 : n30830;
  assign n30832 = pi10 ? n30424 : n30831;
  assign n30833 = pi09 ? n30134 : n30832;
  assign n30834 = pi18 ? n30137 : n30110;
  assign n30835 = pi17 ? n32 : n30834;
  assign n30836 = pi16 ? n30835 : n30113;
  assign n30837 = pi15 ? n30836 : n30128;
  assign n30838 = pi14 ? n30107 : n30837;
  assign n30839 = pi13 ? n32 : n30838;
  assign n30840 = pi12 ? n32 : n30839;
  assign n30841 = pi11 ? n32 : n30840;
  assign n30842 = pi10 ? n32 : n30841;
  assign n30843 = pi22 ? n30195 : n37;
  assign n30844 = pi21 ? n29133 : n30843;
  assign n30845 = pi20 ? n30844 : n5077;
  assign n30846 = pi19 ? n30845 : n99;
  assign n30847 = pi18 ? n30137 : n30846;
  assign n30848 = pi17 ? n32 : n30847;
  assign n30849 = pi16 ? n30848 : n30127;
  assign n30850 = pi15 ? n30849 : n30152;
  assign n30851 = pi19 ? n26407 : n99;
  assign n30852 = pi18 ? n30158 : n30851;
  assign n30853 = pi17 ? n32 : n30852;
  assign n30854 = pi16 ? n30853 : n30166;
  assign n30855 = pi17 ? n30179 : n30192;
  assign n30856 = pi16 ? n30176 : n30855;
  assign n30857 = pi15 ? n30854 : n30856;
  assign n30858 = pi14 ? n30850 : n30857;
  assign n30859 = pi21 ? n2957 : n181;
  assign n30860 = pi20 ? n30859 : n99;
  assign n30861 = pi19 ? n30860 : n99;
  assign n30862 = pi18 ? n374 : n30861;
  assign n30863 = pi17 ? n32 : n30862;
  assign n30864 = pi16 ? n30863 : n29130;
  assign n30865 = pi23 ? n20564 : n20563;
  assign n30866 = pi22 ? n30865 : n20563;
  assign n30867 = pi23 ? n37 : n20563;
  assign n30868 = pi25 ? n98 : n32;
  assign n30869 = pi23 ? n37 : n30868;
  assign n30870 = pi22 ? n30867 : n30869;
  assign n30871 = pi21 ? n30866 : n30870;
  assign n30872 = pi20 ? n32 : n30871;
  assign n30873 = pi19 ? n32 : n30872;
  assign n30874 = pi18 ? n30873 : n37;
  assign n30875 = pi17 ? n32 : n30874;
  assign n30876 = pi20 ? n942 : n992;
  assign n30877 = pi19 ? n30876 : n2471;
  assign n30878 = pi18 ? n30207 : n30877;
  assign n30879 = pi17 ? n30203 : n30878;
  assign n30880 = pi16 ? n30875 : n30879;
  assign n30881 = pi15 ? n30864 : n30880;
  assign n30882 = pi20 ? n3075 : n1704;
  assign n30883 = pi19 ? n30882 : n30219;
  assign n30884 = pi18 ? n374 : n30883;
  assign n30885 = pi17 ? n32 : n30884;
  assign n30886 = pi19 ? n139 : n2567;
  assign n30887 = pi18 ? n30229 : n30886;
  assign n30888 = pi17 ? n30227 : n30887;
  assign n30889 = pi16 ? n30885 : n30888;
  assign n30890 = pi21 ? n23362 : n32;
  assign n30891 = pi20 ? n30890 : n32;
  assign n30892 = pi19 ? n139 : n30891;
  assign n30893 = pi18 ? n30236 : n30892;
  assign n30894 = pi17 ? n30234 : n30893;
  assign n30895 = pi16 ? n439 : n30894;
  assign n30896 = pi15 ? n30889 : n30895;
  assign n30897 = pi14 ? n30881 : n30896;
  assign n30898 = pi13 ? n30858 : n30897;
  assign n30899 = pi21 ? n23370 : n32;
  assign n30900 = pi20 ? n30899 : n32;
  assign n30901 = pi19 ? n139 : n30900;
  assign n30902 = pi18 ? n29243 : n30901;
  assign n30903 = pi17 ? n12372 : n30902;
  assign n30904 = pi16 ? n439 : n30903;
  assign n30905 = pi19 ? n9769 : n2580;
  assign n30906 = pi18 ? n30259 : n30905;
  assign n30907 = pi17 ? n30254 : n30906;
  assign n30908 = pi16 ? n30249 : n30907;
  assign n30909 = pi15 ? n30904 : n30908;
  assign n30910 = pi19 ? n139 : n2639;
  assign n30911 = pi18 ? n30269 : n30910;
  assign n30912 = pi17 ? n30267 : n30911;
  assign n30913 = pi16 ? n439 : n30912;
  assign n30914 = pi18 ? n17061 : n30910;
  assign n30915 = pi17 ? n30273 : n30914;
  assign n30916 = pi16 ? n439 : n30915;
  assign n30917 = pi15 ? n30913 : n30916;
  assign n30918 = pi14 ? n30909 : n30917;
  assign n30919 = pi19 ? n1795 : n2654;
  assign n30920 = pi18 ? n30283 : n30919;
  assign n30921 = pi17 ? n12372 : n30920;
  assign n30922 = pi16 ? n30282 : n30921;
  assign n30923 = pi19 ? n30289 : n2471;
  assign n30924 = pi18 ? n7677 : n30923;
  assign n30925 = pi17 ? n37 : n30924;
  assign n30926 = pi16 ? n439 : n30925;
  assign n30927 = pi15 ? n30922 : n30926;
  assign n30928 = pi19 ? n30295 : n2680;
  assign n30929 = pi18 ? n37 : n30928;
  assign n30930 = pi17 ? n37 : n30929;
  assign n30931 = pi16 ? n439 : n30930;
  assign n30932 = pi19 ? n30301 : n2680;
  assign n30933 = pi18 ? n37 : n30932;
  assign n30934 = pi17 ? n37 : n30933;
  assign n30935 = pi16 ? n439 : n30934;
  assign n30936 = pi15 ? n30931 : n30935;
  assign n30937 = pi14 ? n30927 : n30936;
  assign n30938 = pi13 ? n30918 : n30937;
  assign n30939 = pi12 ? n30898 : n30938;
  assign n30940 = pi19 ? n2095 : n2702;
  assign n30941 = pi18 ? n37 : n30940;
  assign n30942 = pi17 ? n37 : n30941;
  assign n30943 = pi16 ? n439 : n30942;
  assign n30944 = pi19 ? n30321 : n1823;
  assign n30945 = pi18 ? n30319 : n30944;
  assign n30946 = pi17 ? n30316 : n30945;
  assign n30947 = pi16 ? n439 : n30946;
  assign n30948 = pi15 ? n30943 : n30947;
  assign n30949 = pi14 ? n30948 : n30345;
  assign n30950 = pi21 ? n4900 : n233;
  assign n30951 = pi20 ? n335 : n30950;
  assign n30952 = pi19 ? n30951 : n32;
  assign n30953 = pi18 ? n6374 : n30952;
  assign n30954 = pi17 ? n6339 : n30953;
  assign n30955 = pi16 ? n439 : n30954;
  assign n30956 = pi20 ? n25146 : n25965;
  assign n30957 = pi19 ? n30956 : n32;
  assign n30958 = pi18 ? n37 : n30957;
  assign n30959 = pi17 ? n37 : n30958;
  assign n30960 = pi16 ? n439 : n30959;
  assign n30961 = pi15 ? n30955 : n30960;
  assign n30962 = pi14 ? n30961 : n30373;
  assign n30963 = pi13 ? n30949 : n30962;
  assign n30964 = pi21 ? n37 : n10785;
  assign n30965 = pi20 ? n37 : n30964;
  assign n30966 = pi19 ? n30965 : n32;
  assign n30967 = pi18 ? n37 : n30966;
  assign n30968 = pi17 ? n37 : n30967;
  assign n30969 = pi16 ? n439 : n30968;
  assign n30970 = pi15 ? n30381 : n30969;
  assign n30971 = pi14 ? n30970 : n30385;
  assign n30972 = pi21 ? n37 : n2193;
  assign n30973 = pi20 ? n22881 : n30972;
  assign n30974 = pi19 ? n30973 : n32;
  assign n30975 = pi18 ? n30389 : n30974;
  assign n30976 = pi17 ? n37 : n30975;
  assign n30977 = pi16 ? n439 : n30976;
  assign n30978 = pi15 ? n30977 : n30406;
  assign n30979 = pi19 ? n1425 : n32;
  assign n30980 = pi18 ? n37 : n30979;
  assign n30981 = pi17 ? n37 : n30980;
  assign n30982 = pi16 ? n439 : n30981;
  assign n30983 = pi20 ? n30414 : n1424;
  assign n30984 = pi19 ? n30983 : n32;
  assign n30985 = pi18 ? n37 : n30984;
  assign n30986 = pi17 ? n37 : n30985;
  assign n30987 = pi16 ? n439 : n30986;
  assign n30988 = pi15 ? n30982 : n30987;
  assign n30989 = pi14 ? n30978 : n30988;
  assign n30990 = pi13 ? n30971 : n30989;
  assign n30991 = pi12 ? n30963 : n30990;
  assign n30992 = pi11 ? n30939 : n30991;
  assign n30993 = pi20 ? n685 : n2214;
  assign n30994 = pi19 ? n30993 : n32;
  assign n30995 = pi18 ? n30426 : n30994;
  assign n30996 = pi17 ? n37 : n30995;
  assign n30997 = pi16 ? n439 : n30996;
  assign n30998 = pi21 ? n1505 : n218;
  assign n30999 = pi20 ? n32 : n30998;
  assign n31000 = pi19 ? n32 : n30999;
  assign n31001 = pi18 ? n31000 : n99;
  assign n31002 = pi17 ? n32 : n31001;
  assign n31003 = pi21 ? n775 : n5178;
  assign n31004 = pi20 ? n30437 : n31003;
  assign n31005 = pi19 ? n31004 : n32;
  assign n31006 = pi18 ? n19124 : n31005;
  assign n31007 = pi17 ? n99 : n31006;
  assign n31008 = pi16 ? n31002 : n31007;
  assign n31009 = pi15 ? n30997 : n31008;
  assign n31010 = pi21 ? n3562 : n5178;
  assign n31011 = pi20 ? n30445 : n31010;
  assign n31012 = pi19 ? n31011 : n32;
  assign n31013 = pi18 ? n9985 : n31012;
  assign n31014 = pi17 ? n99 : n31013;
  assign n31015 = pi16 ? n201 : n31014;
  assign n31016 = pi21 ? n20977 : n5178;
  assign n31017 = pi20 ? n99 : n31016;
  assign n31018 = pi19 ? n31017 : n32;
  assign n31019 = pi18 ? n30451 : n31018;
  assign n31020 = pi17 ? n99 : n31019;
  assign n31021 = pi16 ? n801 : n31020;
  assign n31022 = pi15 ? n31015 : n31021;
  assign n31023 = pi14 ? n31009 : n31022;
  assign n31024 = pi18 ? n99 : n30454;
  assign n31025 = pi17 ? n99 : n31024;
  assign n31026 = pi16 ? n744 : n31025;
  assign n31027 = pi21 ? n777 : n3523;
  assign n31028 = pi20 ? n99 : n31027;
  assign n31029 = pi19 ? n31028 : n32;
  assign n31030 = pi18 ? n99 : n31029;
  assign n31031 = pi17 ? n99 : n31030;
  assign n31032 = pi16 ? n721 : n31031;
  assign n31033 = pi15 ? n31026 : n31032;
  assign n31034 = pi18 ? n719 : n30468;
  assign n31035 = pi17 ? n32 : n31034;
  assign n31036 = pi20 ? n30475 : n31027;
  assign n31037 = pi19 ? n31036 : n32;
  assign n31038 = pi18 ? n30474 : n31037;
  assign n31039 = pi17 ? n30472 : n31038;
  assign n31040 = pi16 ? n31035 : n31039;
  assign n31041 = pi19 ? n3630 : n32;
  assign n31042 = pi18 ? n30482 : n31041;
  assign n31043 = pi17 ? n30472 : n31042;
  assign n31044 = pi16 ? n31035 : n31043;
  assign n31045 = pi15 ? n31040 : n31044;
  assign n31046 = pi14 ? n31033 : n31045;
  assign n31047 = pi13 ? n31023 : n31046;
  assign n31048 = pi18 ? n10078 : n31041;
  assign n31049 = pi17 ? n139 : n31048;
  assign n31050 = pi16 ? n2291 : n31049;
  assign n31051 = pi16 ? n2291 : n30499;
  assign n31052 = pi15 ? n31050 : n31051;
  assign n31053 = pi16 ? n1575 : n30508;
  assign n31054 = pi15 ? n31053 : n30524;
  assign n31055 = pi14 ? n31052 : n31054;
  assign n31056 = pi18 ? n204 : n24370;
  assign n31057 = pi17 ? n204 : n31056;
  assign n31058 = pi16 ? n30530 : n31057;
  assign n31059 = pi21 ? n11808 : n928;
  assign n31060 = pi20 ? n204 : n31059;
  assign n31061 = pi19 ? n31060 : n32;
  assign n31062 = pi18 ? n204 : n31061;
  assign n31063 = pi17 ? n204 : n31062;
  assign n31064 = pi16 ? n30540 : n31063;
  assign n31065 = pi15 ? n31058 : n31064;
  assign n31066 = pi18 ? n30556 : n31061;
  assign n31067 = pi17 ? n30555 : n31066;
  assign n31068 = pi16 ? n30553 : n31067;
  assign n31069 = pi21 ? n29992 : n2700;
  assign n31070 = pi20 ? n204 : n31069;
  assign n31071 = pi19 ? n31070 : n32;
  assign n31072 = pi18 ? n30556 : n31071;
  assign n31073 = pi17 ? n30565 : n31072;
  assign n31074 = pi16 ? n30561 : n31073;
  assign n31075 = pi15 ? n31068 : n31074;
  assign n31076 = pi14 ? n31065 : n31075;
  assign n31077 = pi13 ? n31055 : n31076;
  assign n31078 = pi12 ? n31047 : n31077;
  assign n31079 = pi21 ? n326 : n375;
  assign n31080 = pi20 ? n32 : n31079;
  assign n31081 = pi19 ? n32 : n31080;
  assign n31082 = pi21 ? n3668 : n375;
  assign n31083 = pi20 ? n31082 : n5255;
  assign n31084 = pi20 ? n12014 : n3075;
  assign n31085 = pi19 ? n31083 : n31084;
  assign n31086 = pi18 ? n31081 : n31085;
  assign n31087 = pi17 ? n32 : n31086;
  assign n31088 = pi21 ? n9144 : n37;
  assign n31089 = pi19 ? n9132 : n31088;
  assign n31090 = pi20 ? n31088 : n27161;
  assign n31091 = pi21 ? n9124 : n9563;
  assign n31092 = pi20 ? n31091 : n27145;
  assign n31093 = pi19 ? n31090 : n31092;
  assign n31094 = pi18 ? n31089 : n31093;
  assign n31095 = pi21 ? n567 : n3073;
  assign n31096 = pi21 ? n569 : n10234;
  assign n31097 = pi20 ? n31095 : n31096;
  assign n31098 = pi19 ? n31097 : n30594;
  assign n31099 = pi20 ? n30596 : n31069;
  assign n31100 = pi19 ? n31099 : n32;
  assign n31101 = pi18 ? n31098 : n31100;
  assign n31102 = pi17 ? n31094 : n31101;
  assign n31103 = pi16 ? n31087 : n31102;
  assign n31104 = pi21 ? n25977 : n1009;
  assign n31105 = pi20 ? n7980 : n31104;
  assign n31106 = pi19 ? n31105 : n32;
  assign n31107 = pi18 ? n17487 : n31106;
  assign n31108 = pi17 ? n335 : n31107;
  assign n31109 = pi16 ? n30605 : n31108;
  assign n31110 = pi15 ? n31103 : n31109;
  assign n31111 = pi20 ? n15457 : n30606;
  assign n31112 = pi19 ? n31111 : n32;
  assign n31113 = pi18 ? n17487 : n31112;
  assign n31114 = pi17 ? n30618 : n31113;
  assign n31115 = pi16 ? n30615 : n31114;
  assign n31116 = pi20 ? n7980 : n30006;
  assign n31117 = pi19 ? n31116 : n32;
  assign n31118 = pi18 ? n30633 : n31117;
  assign n31119 = pi17 ? n30631 : n31118;
  assign n31120 = pi16 ? n30626 : n31119;
  assign n31121 = pi15 ? n31115 : n31120;
  assign n31122 = pi14 ? n31110 : n31121;
  assign n31123 = pi18 ? n19406 : n20844;
  assign n31124 = pi17 ? n30646 : n31123;
  assign n31125 = pi16 ? n30644 : n31124;
  assign n31126 = pi20 ? n233 : n4852;
  assign n31127 = pi19 ? n31126 : n32;
  assign n31128 = pi18 ? n30662 : n31127;
  assign n31129 = pi17 ? n30660 : n31128;
  assign n31130 = pi16 ? n30654 : n31129;
  assign n31131 = pi15 ? n31125 : n31130;
  assign n31132 = pi18 ? n30679 : n30648;
  assign n31133 = pi17 ? n30677 : n31132;
  assign n31134 = pi16 ? n30670 : n31133;
  assign n31135 = pi21 ? n555 : n569;
  assign n31136 = pi20 ? n32 : n31135;
  assign n31137 = pi19 ? n32 : n31136;
  assign n31138 = pi18 ? n31137 : n30687;
  assign n31139 = pi17 ? n32 : n31138;
  assign n31140 = pi20 ? n30701 : n8295;
  assign n31141 = pi19 ? n31140 : n32;
  assign n31142 = pi18 ? n30699 : n31141;
  assign n31143 = pi17 ? n30697 : n31142;
  assign n31144 = pi16 ? n31139 : n31143;
  assign n31145 = pi15 ? n31134 : n31144;
  assign n31146 = pi14 ? n31131 : n31145;
  assign n31147 = pi13 ? n31122 : n31146;
  assign n31148 = pi20 ? n233 : n9482;
  assign n31149 = pi19 ? n31148 : n32;
  assign n31150 = pi18 ? n30730 : n31149;
  assign n31151 = pi17 ? n30727 : n31150;
  assign n31152 = pi16 ? n30715 : n31151;
  assign n31153 = pi20 ? n233 : n4008;
  assign n31154 = pi19 ? n31153 : n32;
  assign n31155 = pi18 ? n30744 : n31154;
  assign n31156 = pi17 ? n30740 : n31155;
  assign n31157 = pi16 ? n439 : n31156;
  assign n31158 = pi15 ? n31152 : n31157;
  assign n31159 = pi20 ? n30789 : n7724;
  assign n31160 = pi19 ? n31159 : n32;
  assign n31161 = pi18 ? n30787 : n31160;
  assign n31162 = pi17 ? n30781 : n31161;
  assign n31163 = pi16 ? n30770 : n31162;
  assign n31164 = pi15 ? n30758 : n31163;
  assign n31165 = pi14 ? n31158 : n31164;
  assign n31166 = pi20 ? n24223 : n3210;
  assign n31167 = pi19 ? n31166 : n32;
  assign n31168 = pi18 ? n30799 : n31167;
  assign n31169 = pi17 ? n363 : n31168;
  assign n31170 = pi16 ? n30798 : n31169;
  assign n31171 = pi23 ? n7420 : n316;
  assign n31172 = pi22 ? n363 : n31171;
  assign n31173 = pi21 ? n363 : n31172;
  assign n31174 = pi20 ? n31173 : n10011;
  assign n31175 = pi19 ? n31174 : n32;
  assign n31176 = pi18 ? n30806 : n31175;
  assign n31177 = pi17 ? n363 : n31176;
  assign n31178 = pi16 ? n21219 : n31177;
  assign n31179 = pi15 ? n31170 : n31178;
  assign n31180 = pi20 ? n31173 : n1822;
  assign n31181 = pi19 ? n31180 : n32;
  assign n31182 = pi18 ? n363 : n31181;
  assign n31183 = pi17 ? n363 : n31182;
  assign n31184 = pi16 ? n21219 : n31183;
  assign n31185 = pi22 ? n363 : n8328;
  assign n31186 = pi21 ? n685 : n31185;
  assign n31187 = pi20 ? n31186 : n32;
  assign n31188 = pi19 ? n31187 : n32;
  assign n31189 = pi18 ? n363 : n31188;
  assign n31190 = pi17 ? n363 : n31189;
  assign n31191 = pi16 ? n26062 : n31190;
  assign n31192 = pi15 ? n31184 : n31191;
  assign n31193 = pi14 ? n31179 : n31192;
  assign n31194 = pi13 ? n31165 : n31193;
  assign n31195 = pi12 ? n31147 : n31194;
  assign n31196 = pi11 ? n31078 : n31195;
  assign n31197 = pi10 ? n30992 : n31196;
  assign n31198 = pi09 ? n30842 : n31197;
  assign n31199 = pi08 ? n30833 : n31198;
  assign n31200 = pi22 ? n30867 : n37;
  assign n31201 = pi21 ? n29132 : n31200;
  assign n31202 = pi20 ? n32 : n31201;
  assign n31203 = pi19 ? n32 : n31202;
  assign n31204 = pi22 ? n30195 : n30867;
  assign n31205 = pi21 ? n31204 : n37;
  assign n31206 = pi20 ? n31205 : n37;
  assign n31207 = pi19 ? n31206 : n16999;
  assign n31208 = pi18 ? n31203 : n31207;
  assign n31209 = pi17 ? n32 : n31208;
  assign n31210 = pi20 ? n3039 : n5077;
  assign n31211 = pi19 ? n31210 : n16999;
  assign n31212 = pi20 ? n226 : n37;
  assign n31213 = pi19 ? n31212 : n21611;
  assign n31214 = pi18 ? n31211 : n31213;
  assign n31215 = pi19 ? n99 : n3834;
  assign n31216 = pi18 ? n99 : n31215;
  assign n31217 = pi17 ? n31214 : n31216;
  assign n31218 = pi16 ? n31209 : n31217;
  assign n31219 = pi15 ? n32 : n31218;
  assign n31220 = pi21 ? n20563 : n37;
  assign n31221 = pi20 ? n20563 : n31220;
  assign n31222 = pi19 ? n31221 : n26407;
  assign n31223 = pi18 ? n30119 : n31222;
  assign n31224 = pi17 ? n32 : n31223;
  assign n31225 = pi17 ? n99 : n31216;
  assign n31226 = pi16 ? n31224 : n31225;
  assign n31227 = pi22 ? n39 : n30195;
  assign n31228 = pi21 ? n31227 : n37;
  assign n31229 = pi20 ? n32 : n31228;
  assign n31230 = pi19 ? n32 : n31229;
  assign n31231 = pi19 ? n37 : n19773;
  assign n31232 = pi18 ? n31230 : n31231;
  assign n31233 = pi17 ? n32 : n31232;
  assign n31234 = pi20 ? n16991 : n32;
  assign n31235 = pi19 ? n99 : n31234;
  assign n31236 = pi18 ? n99 : n31235;
  assign n31237 = pi17 ? n99 : n31236;
  assign n31238 = pi16 ? n31233 : n31237;
  assign n31239 = pi15 ? n31226 : n31238;
  assign n31240 = pi14 ? n31219 : n31239;
  assign n31241 = pi13 ? n32 : n31240;
  assign n31242 = pi12 ? n32 : n31241;
  assign n31243 = pi11 ? n32 : n31242;
  assign n31244 = pi10 ? n32 : n31243;
  assign n31245 = pi22 ? n64 : n30195;
  assign n31246 = pi21 ? n31245 : n31200;
  assign n31247 = pi20 ? n32 : n31246;
  assign n31248 = pi19 ? n32 : n31247;
  assign n31249 = pi18 ? n31248 : n23649;
  assign n31250 = pi17 ? n32 : n31249;
  assign n31251 = pi19 ? n23645 : n29456;
  assign n31252 = pi20 ? n5420 : n14887;
  assign n31253 = pi19 ? n31252 : n7747;
  assign n31254 = pi18 ? n31251 : n31253;
  assign n31255 = pi21 ? n2160 : n37;
  assign n31256 = pi20 ? n99 : n31255;
  assign n31257 = pi19 ? n99 : n31256;
  assign n31258 = pi20 ? n18040 : n32;
  assign n31259 = pi19 ? n99 : n31258;
  assign n31260 = pi18 ? n31257 : n31259;
  assign n31261 = pi17 ? n31254 : n31260;
  assign n31262 = pi16 ? n31250 : n31261;
  assign n31263 = pi21 ? n30155 : n20563;
  assign n31264 = pi20 ? n32 : n31263;
  assign n31265 = pi19 ? n32 : n31264;
  assign n31266 = pi21 ? n20563 : n29133;
  assign n31267 = pi20 ? n31266 : n37;
  assign n31268 = pi19 ? n31267 : n27249;
  assign n31269 = pi18 ? n31265 : n31268;
  assign n31270 = pi17 ? n32 : n31269;
  assign n31271 = pi23 ? n11962 : n586;
  assign n31272 = pi22 ? n31271 : n32;
  assign n31273 = pi21 ? n31272 : n32;
  assign n31274 = pi20 ? n31273 : n32;
  assign n31275 = pi19 ? n99 : n31274;
  assign n31276 = pi18 ? n99 : n31275;
  assign n31277 = pi17 ? n99 : n31276;
  assign n31278 = pi16 ? n31270 : n31277;
  assign n31279 = pi15 ? n31262 : n31278;
  assign n31280 = pi20 ? n31220 : n37;
  assign n31281 = pi19 ? n31280 : n99;
  assign n31282 = pi18 ? n30158 : n31281;
  assign n31283 = pi17 ? n32 : n31282;
  assign n31284 = pi23 ? n11910 : n5630;
  assign n31285 = pi22 ? n31284 : n32;
  assign n31286 = pi21 ? n31285 : n32;
  assign n31287 = pi20 ? n31286 : n32;
  assign n31288 = pi19 ? n99 : n31287;
  assign n31289 = pi18 ? n99 : n31288;
  assign n31290 = pi17 ? n99 : n31289;
  assign n31291 = pi16 ? n31283 : n31290;
  assign n31292 = pi23 ? n38 : n20563;
  assign n31293 = pi22 ? n31292 : n20563;
  assign n31294 = pi22 ? n20563 : n30867;
  assign n31295 = pi21 ? n31293 : n31294;
  assign n31296 = pi20 ? n32 : n31295;
  assign n31297 = pi19 ? n32 : n31296;
  assign n31298 = pi21 ? n31200 : n37;
  assign n31299 = pi20 ? n31298 : n37;
  assign n31300 = pi19 ? n31299 : n37;
  assign n31301 = pi18 ? n31297 : n31300;
  assign n31302 = pi17 ? n32 : n31301;
  assign n31303 = pi19 ? n20657 : n3039;
  assign n31304 = pi18 ? n37 : n31303;
  assign n31305 = pi20 ? n7747 : n3046;
  assign n31306 = pi20 ? n17584 : n32;
  assign n31307 = pi19 ? n31305 : n31306;
  assign n31308 = pi18 ? n28217 : n31307;
  assign n31309 = pi17 ? n31304 : n31308;
  assign n31310 = pi16 ? n31302 : n31309;
  assign n31311 = pi15 ? n31291 : n31310;
  assign n31312 = pi14 ? n31279 : n31311;
  assign n31313 = pi21 ? n30866 : n20563;
  assign n31314 = pi20 ? n32 : n31313;
  assign n31315 = pi19 ? n32 : n31314;
  assign n31316 = pi18 ? n31315 : n37;
  assign n31317 = pi17 ? n32 : n31316;
  assign n31318 = pi20 ? n37 : n14530;
  assign n31319 = pi19 ? n37 : n31318;
  assign n31320 = pi20 ? n17024 : n37;
  assign n31321 = pi19 ? n31320 : n2970;
  assign n31322 = pi18 ? n31319 : n31321;
  assign n31323 = pi20 ? n2185 : n14512;
  assign n31324 = pi20 ? n3822 : n22651;
  assign n31325 = pi19 ? n31323 : n31324;
  assign n31326 = pi21 ? n2981 : n181;
  assign n31327 = pi20 ? n21638 : n31326;
  assign n31328 = pi24 ? n37 : n157;
  assign n31329 = pi23 ? n31328 : n32;
  assign n31330 = pi22 ? n31329 : n32;
  assign n31331 = pi21 ? n31330 : n32;
  assign n31332 = pi20 ? n31331 : n32;
  assign n31333 = pi19 ? n31327 : n31332;
  assign n31334 = pi18 ? n31325 : n31333;
  assign n31335 = pi17 ? n31322 : n31334;
  assign n31336 = pi16 ? n31317 : n31335;
  assign n31337 = pi19 ? n18070 : n37;
  assign n31338 = pi19 ? n9769 : n31332;
  assign n31339 = pi18 ? n31337 : n31338;
  assign n31340 = pi17 ? n37 : n31339;
  assign n31341 = pi16 ? n439 : n31340;
  assign n31342 = pi15 ? n31336 : n31341;
  assign n31343 = pi19 ? n8765 : n2567;
  assign n31344 = pi18 ? n37 : n31343;
  assign n31345 = pi17 ? n37 : n31344;
  assign n31346 = pi16 ? n439 : n31345;
  assign n31347 = pi21 ? n31293 : n31200;
  assign n31348 = pi20 ? n32 : n31347;
  assign n31349 = pi19 ? n32 : n31348;
  assign n31350 = pi18 ? n31349 : n37;
  assign n31351 = pi17 ? n32 : n31350;
  assign n31352 = pi19 ? n3104 : n37;
  assign n31353 = pi18 ? n31352 : n30886;
  assign n31354 = pi17 ? n37 : n31353;
  assign n31355 = pi16 ? n31351 : n31354;
  assign n31356 = pi15 ? n31346 : n31355;
  assign n31357 = pi14 ? n31342 : n31356;
  assign n31358 = pi13 ? n31312 : n31357;
  assign n31359 = pi19 ? n139 : n2580;
  assign n31360 = pi18 ? n37 : n31359;
  assign n31361 = pi17 ? n37 : n31360;
  assign n31362 = pi16 ? n439 : n31361;
  assign n31363 = pi20 ? n3083 : n37;
  assign n31364 = pi19 ? n31363 : n37;
  assign n31365 = pi19 ? n8765 : n2580;
  assign n31366 = pi18 ? n31364 : n31365;
  assign n31367 = pi17 ? n30273 : n31366;
  assign n31368 = pi16 ? n439 : n31367;
  assign n31369 = pi15 ? n31362 : n31368;
  assign n31370 = pi20 ? n3104 : n3090;
  assign n31371 = pi19 ? n37 : n31370;
  assign n31372 = pi18 ? n37 : n31371;
  assign n31373 = pi20 ? n13121 : n8742;
  assign n31374 = pi19 ? n31373 : n29260;
  assign n31375 = pi18 ? n31374 : n30910;
  assign n31376 = pi17 ? n31372 : n31375;
  assign n31377 = pi16 ? n439 : n31376;
  assign n31378 = pi15 ? n31377 : n30916;
  assign n31379 = pi14 ? n31369 : n31378;
  assign n31380 = pi21 ? n1696 : n569;
  assign n31381 = pi21 ? n335 : n20218;
  assign n31382 = pi20 ? n31380 : n31381;
  assign n31383 = pi19 ? n31382 : n2654;
  assign n31384 = pi18 ? n37 : n31383;
  assign n31385 = pi17 ? n37 : n31384;
  assign n31386 = pi16 ? n439 : n31385;
  assign n31387 = pi20 ? n577 : n14383;
  assign n31388 = pi19 ? n31387 : n2471;
  assign n31389 = pi18 ? n37 : n31388;
  assign n31390 = pi17 ? n37 : n31389;
  assign n31391 = pi16 ? n439 : n31390;
  assign n31392 = pi15 ? n31386 : n31391;
  assign n31393 = pi20 ? n649 : n21199;
  assign n31394 = pi19 ? n31393 : n2555;
  assign n31395 = pi18 ? n37 : n31394;
  assign n31396 = pi17 ? n37 : n31395;
  assign n31397 = pi16 ? n439 : n31396;
  assign n31398 = pi19 ? n2095 : n2580;
  assign n31399 = pi18 ? n37 : n31398;
  assign n31400 = pi17 ? n37 : n31399;
  assign n31401 = pi16 ? n439 : n31400;
  assign n31402 = pi15 ? n31397 : n31401;
  assign n31403 = pi14 ? n31392 : n31402;
  assign n31404 = pi13 ? n31379 : n31403;
  assign n31405 = pi12 ? n31358 : n31404;
  assign n31406 = pi19 ? n2095 : n2680;
  assign n31407 = pi18 ? n37 : n31406;
  assign n31408 = pi17 ? n37 : n31407;
  assign n31409 = pi16 ? n439 : n31408;
  assign n31410 = pi21 ? n37 : n2074;
  assign n31411 = pi20 ? n610 : n31410;
  assign n31412 = pi19 ? n31411 : n2680;
  assign n31413 = pi18 ? n37 : n31412;
  assign n31414 = pi17 ? n37 : n31413;
  assign n31415 = pi16 ? n439 : n31414;
  assign n31416 = pi15 ? n31409 : n31415;
  assign n31417 = pi20 ? n37 : n7587;
  assign n31418 = pi19 ? n37 : n31417;
  assign n31419 = pi18 ? n31418 : n31412;
  assign n31420 = pi17 ? n37 : n31419;
  assign n31421 = pi16 ? n439 : n31420;
  assign n31422 = pi20 ? n647 : n8927;
  assign n31423 = pi19 ? n31422 : n2680;
  assign n31424 = pi18 ? n37 : n31423;
  assign n31425 = pi17 ? n37 : n31424;
  assign n31426 = pi16 ? n439 : n31425;
  assign n31427 = pi15 ? n31421 : n31426;
  assign n31428 = pi14 ? n31416 : n31427;
  assign n31429 = pi19 ? n30698 : n2680;
  assign n31430 = pi18 ? n37 : n31429;
  assign n31431 = pi17 ? n37 : n31430;
  assign n31432 = pi16 ? n439 : n31431;
  assign n31433 = pi20 ? n8927 : n25965;
  assign n31434 = pi19 ? n31433 : n2702;
  assign n31435 = pi18 ? n37 : n31434;
  assign n31436 = pi17 ? n37 : n31435;
  assign n31437 = pi16 ? n439 : n31436;
  assign n31438 = pi15 ? n31432 : n31437;
  assign n31439 = pi20 ? n2107 : n2729;
  assign n31440 = pi19 ? n31439 : n2702;
  assign n31441 = pi18 ? n37 : n31440;
  assign n31442 = pi17 ? n37 : n31441;
  assign n31443 = pi16 ? n439 : n31442;
  assign n31444 = pi22 ? n685 : n686;
  assign n31445 = pi21 ? n37 : n31444;
  assign n31446 = pi20 ? n37 : n31445;
  assign n31447 = pi19 ? n31446 : n1823;
  assign n31448 = pi18 ? n37 : n31447;
  assign n31449 = pi17 ? n37 : n31448;
  assign n31450 = pi16 ? n439 : n31449;
  assign n31451 = pi15 ? n31443 : n31450;
  assign n31452 = pi14 ? n31438 : n31451;
  assign n31453 = pi13 ? n31428 : n31452;
  assign n31454 = pi21 ? n37 : n14255;
  assign n31455 = pi20 ? n37 : n31454;
  assign n31456 = pi19 ? n31455 : n32;
  assign n31457 = pi18 ? n37 : n31456;
  assign n31458 = pi17 ? n37 : n31457;
  assign n31459 = pi16 ? n439 : n31458;
  assign n31460 = pi19 ? n2723 : n32;
  assign n31461 = pi18 ? n37 : n31460;
  assign n31462 = pi17 ? n37 : n31461;
  assign n31463 = pi16 ? n439 : n31462;
  assign n31464 = pi22 ? n295 : n685;
  assign n31465 = pi21 ? n37 : n31464;
  assign n31466 = pi20 ? n37 : n31465;
  assign n31467 = pi19 ? n31466 : n32;
  assign n31468 = pi18 ? n37 : n31467;
  assign n31469 = pi17 ? n37 : n31468;
  assign n31470 = pi16 ? n439 : n31469;
  assign n31471 = pi15 ? n31463 : n31470;
  assign n31472 = pi14 ? n31459 : n31471;
  assign n31473 = pi21 ? n37 : n3436;
  assign n31474 = pi20 ? n22881 : n31473;
  assign n31475 = pi19 ? n31474 : n32;
  assign n31476 = pi18 ? n7732 : n31475;
  assign n31477 = pi17 ? n37 : n31476;
  assign n31478 = pi16 ? n439 : n31477;
  assign n31479 = pi20 ? n3393 : n10494;
  assign n31480 = pi19 ? n37 : n31479;
  assign n31481 = pi18 ? n37 : n31480;
  assign n31482 = pi20 ? n7322 : n19091;
  assign n31483 = pi20 ? n19091 : n21826;
  assign n31484 = pi19 ? n31482 : n31483;
  assign n31485 = pi21 ? n363 : n1423;
  assign n31486 = pi20 ? n363 : n31485;
  assign n31487 = pi19 ? n31486 : n32;
  assign n31488 = pi18 ? n31484 : n31487;
  assign n31489 = pi17 ? n31481 : n31488;
  assign n31490 = pi16 ? n439 : n31489;
  assign n31491 = pi15 ? n31478 : n31490;
  assign n31492 = pi20 ? n19959 : n1424;
  assign n31493 = pi19 ? n31492 : n32;
  assign n31494 = pi18 ? n37 : n31493;
  assign n31495 = pi17 ? n37 : n31494;
  assign n31496 = pi16 ? n439 : n31495;
  assign n31497 = pi21 ? n157 : n19958;
  assign n31498 = pi20 ? n31497 : n1424;
  assign n31499 = pi19 ? n31498 : n32;
  assign n31500 = pi18 ? n37 : n31499;
  assign n31501 = pi17 ? n37 : n31500;
  assign n31502 = pi16 ? n439 : n31501;
  assign n31503 = pi15 ? n31496 : n31502;
  assign n31504 = pi14 ? n31491 : n31503;
  assign n31505 = pi13 ? n31472 : n31504;
  assign n31506 = pi12 ? n31453 : n31505;
  assign n31507 = pi11 ? n31405 : n31506;
  assign n31508 = pi19 ? n226 : n18853;
  assign n31509 = pi18 ? n15526 : n31508;
  assign n31510 = pi17 ? n32 : n31509;
  assign n31511 = pi19 ? n3050 : n4583;
  assign n31512 = pi20 ? n776 : n13948;
  assign n31513 = pi19 ? n219 : n31512;
  assign n31514 = pi18 ? n31511 : n31513;
  assign n31515 = pi21 ? n99 : n244;
  assign n31516 = pi20 ? n31515 : n157;
  assign n31517 = pi19 ? n99 : n31516;
  assign n31518 = pi18 ? n31517 : n30994;
  assign n31519 = pi17 ? n31514 : n31518;
  assign n31520 = pi16 ? n31510 : n31519;
  assign n31521 = pi18 ? n3031 : n18854;
  assign n31522 = pi17 ? n32 : n31521;
  assign n31523 = pi19 ? n18853 : n2255;
  assign n31524 = pi20 ? n776 : n5179;
  assign n31525 = pi19 ? n31524 : n32;
  assign n31526 = pi18 ? n31523 : n31525;
  assign n31527 = pi17 ? n99 : n31526;
  assign n31528 = pi16 ? n31522 : n31527;
  assign n31529 = pi15 ? n31520 : n31528;
  assign n31530 = pi16 ? n1676 : n31014;
  assign n31531 = pi18 ? n374 : n15541;
  assign n31532 = pi17 ? n32 : n31531;
  assign n31533 = pi20 ? n18291 : n31027;
  assign n31534 = pi19 ? n31533 : n32;
  assign n31535 = pi18 ? n99 : n31534;
  assign n31536 = pi17 ? n99 : n31535;
  assign n31537 = pi16 ? n31532 : n31536;
  assign n31538 = pi15 ? n31530 : n31537;
  assign n31539 = pi14 ? n31529 : n31538;
  assign n31540 = pi16 ? n801 : n31025;
  assign n31541 = pi21 ? n746 : n3523;
  assign n31542 = pi20 ? n99 : n31541;
  assign n31543 = pi19 ? n31542 : n32;
  assign n31544 = pi18 ? n99 : n31543;
  assign n31545 = pi17 ? n99 : n31544;
  assign n31546 = pi16 ? n744 : n31545;
  assign n31547 = pi15 ? n31540 : n31546;
  assign n31548 = pi20 ? n139 : n22965;
  assign n31549 = pi19 ? n139 : n31548;
  assign n31550 = pi21 ? n159 : n3523;
  assign n31551 = pi20 ? n30475 : n31550;
  assign n31552 = pi19 ? n31551 : n32;
  assign n31553 = pi18 ? n31549 : n31552;
  assign n31554 = pi17 ? n30472 : n31553;
  assign n31555 = pi16 ? n30470 : n31554;
  assign n31556 = pi16 ? n30470 : n31043;
  assign n31557 = pi15 ? n31555 : n31556;
  assign n31558 = pi14 ? n31547 : n31557;
  assign n31559 = pi13 ? n31539 : n31558;
  assign n31560 = pi21 ? n8143 : n1531;
  assign n31561 = pi20 ? n32 : n31560;
  assign n31562 = pi19 ? n32 : n31561;
  assign n31563 = pi18 ? n31562 : n139;
  assign n31564 = pi17 ? n32 : n31563;
  assign n31565 = pi19 ? n139 : n14318;
  assign n31566 = pi18 ? n139 : n31565;
  assign n31567 = pi17 ? n31566 : n30491;
  assign n31568 = pi16 ? n31564 : n31567;
  assign n31569 = pi21 ? n326 : n1531;
  assign n31570 = pi20 ? n32 : n31569;
  assign n31571 = pi19 ? n32 : n31570;
  assign n31572 = pi18 ? n31571 : n139;
  assign n31573 = pi17 ? n32 : n31572;
  assign n31574 = pi20 ? n6650 : n1008;
  assign n31575 = pi19 ? n139 : n31574;
  assign n31576 = pi18 ? n139 : n31575;
  assign n31577 = pi20 ? n139 : n7909;
  assign n31578 = pi19 ? n139 : n31577;
  assign n31579 = pi18 ? n31578 : n30484;
  assign n31580 = pi17 ? n31576 : n31579;
  assign n31581 = pi16 ? n31573 : n31580;
  assign n31582 = pi15 ? n31568 : n31581;
  assign n31583 = pi20 ? n3083 : n997;
  assign n31584 = pi20 ? n947 : n922;
  assign n31585 = pi19 ? n31583 : n31584;
  assign n31586 = pi18 ? n374 : n31585;
  assign n31587 = pi17 ? n32 : n31586;
  assign n31588 = pi21 ? n204 : n919;
  assign n31589 = pi20 ? n31588 : n29520;
  assign n31590 = pi19 ? n18361 : n31589;
  assign n31591 = pi20 ? n2318 : n1068;
  assign n31592 = pi19 ? n29520 : n31591;
  assign n31593 = pi18 ? n31590 : n31592;
  assign n31594 = pi20 ? n927 : n975;
  assign n31595 = pi19 ? n1016 : n31594;
  assign n31596 = pi18 ? n31595 : n30484;
  assign n31597 = pi17 ? n31593 : n31596;
  assign n31598 = pi16 ? n31587 : n31597;
  assign n31599 = pi21 ? n935 : n1698;
  assign n31600 = pi20 ? n32 : n31599;
  assign n31601 = pi19 ? n32 : n31600;
  assign n31602 = pi20 ? n1693 : n13119;
  assign n31603 = pi21 ? n1696 : n297;
  assign n31604 = pi20 ? n31603 : n37;
  assign n31605 = pi19 ? n31602 : n31604;
  assign n31606 = pi18 ? n31601 : n31605;
  assign n31607 = pi17 ? n32 : n31606;
  assign n31608 = pi20 ? n204 : n139;
  assign n31609 = pi19 ? n15398 : n31608;
  assign n31610 = pi18 ? n30514 : n31609;
  assign n31611 = pi20 ? n29572 : n204;
  assign n31612 = pi20 ? n2318 : n6568;
  assign n31613 = pi19 ? n31611 : n31612;
  assign n31614 = pi21 ? n916 : n2637;
  assign n31615 = pi20 ? n922 : n31614;
  assign n31616 = pi19 ? n31615 : n32;
  assign n31617 = pi18 ? n31613 : n31616;
  assign n31618 = pi17 ? n31610 : n31617;
  assign n31619 = pi16 ? n31607 : n31618;
  assign n31620 = pi15 ? n31598 : n31619;
  assign n31621 = pi14 ? n31582 : n31620;
  assign n31622 = pi21 ? n910 : n1711;
  assign n31623 = pi20 ? n32 : n31622;
  assign n31624 = pi19 ? n32 : n31623;
  assign n31625 = pi21 ? n820 : n916;
  assign n31626 = pi20 ? n31625 : n5199;
  assign n31627 = pi19 ? n139 : n31626;
  assign n31628 = pi18 ? n31624 : n31627;
  assign n31629 = pi17 ? n32 : n31628;
  assign n31630 = pi23 ? n1598 : n32;
  assign n31631 = pi22 ? n31630 : n32;
  assign n31632 = pi21 ? n204 : n31631;
  assign n31633 = pi20 ? n204 : n31632;
  assign n31634 = pi19 ? n31633 : n32;
  assign n31635 = pi18 ? n204 : n31634;
  assign n31636 = pi17 ? n204 : n31635;
  assign n31637 = pi16 ? n31629 : n31636;
  assign n31638 = pi20 ? n3075 : n14066;
  assign n31639 = pi21 ? n37 : n1049;
  assign n31640 = pi20 ? n31639 : n204;
  assign n31641 = pi19 ? n31638 : n31640;
  assign n31642 = pi18 ? n8706 : n31641;
  assign n31643 = pi17 ? n32 : n31642;
  assign n31644 = pi21 ? n204 : n3397;
  assign n31645 = pi20 ? n204 : n31644;
  assign n31646 = pi19 ? n31645 : n32;
  assign n31647 = pi18 ? n204 : n31646;
  assign n31648 = pi17 ? n204 : n31647;
  assign n31649 = pi16 ? n31643 : n31648;
  assign n31650 = pi15 ? n31637 : n31649;
  assign n31651 = pi20 ? n1003 : n14039;
  assign n31652 = pi20 ? n1003 : n14068;
  assign n31653 = pi19 ? n31651 : n31652;
  assign n31654 = pi18 ? n31081 : n31653;
  assign n31655 = pi17 ? n32 : n31654;
  assign n31656 = pi19 ? n9769 : n16473;
  assign n31657 = pi23 ? n21112 : n32;
  assign n31658 = pi22 ? n31657 : n32;
  assign n31659 = pi21 ? n11808 : n31658;
  assign n31660 = pi20 ? n204 : n31659;
  assign n31661 = pi19 ? n31660 : n32;
  assign n31662 = pi18 ? n31656 : n31661;
  assign n31663 = pi17 ? n139 : n31662;
  assign n31664 = pi16 ? n31655 : n31663;
  assign n31665 = pi18 ? n329 : n8766;
  assign n31666 = pi17 ? n32 : n31665;
  assign n31667 = pi19 ? n139 : n13100;
  assign n31668 = pi18 ? n139 : n31667;
  assign n31669 = pi21 ? n11808 : n2700;
  assign n31670 = pi20 ? n204 : n31669;
  assign n31671 = pi19 ? n31670 : n32;
  assign n31672 = pi18 ? n30556 : n31671;
  assign n31673 = pi17 ? n31668 : n31672;
  assign n31674 = pi16 ? n31666 : n31673;
  assign n31675 = pi15 ? n31664 : n31674;
  assign n31676 = pi14 ? n31650 : n31675;
  assign n31677 = pi13 ? n31621 : n31676;
  assign n31678 = pi12 ? n31559 : n31677;
  assign n31679 = pi20 ? n647 : n3289;
  assign n31680 = pi19 ? n644 : n31679;
  assign n31681 = pi20 ? n605 : n638;
  assign n31682 = pi19 ? n3289 : n31681;
  assign n31683 = pi18 ? n31680 : n31682;
  assign n31684 = pi20 ? n571 : n639;
  assign n31685 = pi20 ? n604 : n16544;
  assign n31686 = pi19 ? n31684 : n31685;
  assign n31687 = pi21 ? n233 : n11808;
  assign n31688 = pi22 ? n233 : n3762;
  assign n31689 = pi21 ? n31688 : n2700;
  assign n31690 = pi20 ? n31687 : n31689;
  assign n31691 = pi19 ? n31690 : n32;
  assign n31692 = pi18 ? n31686 : n31691;
  assign n31693 = pi17 ? n31683 : n31692;
  assign n31694 = pi16 ? n439 : n31693;
  assign n31695 = pi21 ? n569 : n1943;
  assign n31696 = pi20 ? n577 : n31695;
  assign n31697 = pi20 ? n604 : n30288;
  assign n31698 = pi19 ? n31696 : n31697;
  assign n31699 = pi18 ? n3349 : n31698;
  assign n31700 = pi17 ? n32 : n31699;
  assign n31701 = pi19 ? n16516 : n335;
  assign n31702 = pi18 ? n31701 : n335;
  assign n31703 = pi21 ? n8869 : n1009;
  assign n31704 = pi20 ? n7980 : n31703;
  assign n31705 = pi19 ? n31704 : n32;
  assign n31706 = pi18 ? n335 : n31705;
  assign n31707 = pi17 ? n31702 : n31706;
  assign n31708 = pi16 ? n31700 : n31707;
  assign n31709 = pi15 ? n31694 : n31708;
  assign n31710 = pi18 ? n3349 : n30613;
  assign n31711 = pi17 ? n32 : n31710;
  assign n31712 = pi22 ? n10400 : n3338;
  assign n31713 = pi21 ? n31712 : n32;
  assign n31714 = pi20 ? n15457 : n31713;
  assign n31715 = pi19 ? n31714 : n32;
  assign n31716 = pi18 ? n335 : n31715;
  assign n31717 = pi17 ? n30618 : n31716;
  assign n31718 = pi16 ? n31711 : n31717;
  assign n31719 = pi20 ? n335 : n610;
  assign n31720 = pi19 ? n14166 : n31719;
  assign n31721 = pi18 ? n3349 : n31720;
  assign n31722 = pi17 ? n32 : n31721;
  assign n31723 = pi21 ? n335 : n2007;
  assign n31724 = pi20 ? n7646 : n31723;
  assign n31725 = pi19 ? n612 : n31724;
  assign n31726 = pi20 ? n31723 : n10093;
  assign n31727 = pi20 ? n571 : n604;
  assign n31728 = pi19 ? n31726 : n31727;
  assign n31729 = pi18 ? n31725 : n31728;
  assign n31730 = pi20 ? n3335 : n605;
  assign n31731 = pi19 ? n31730 : n28367;
  assign n31732 = pi20 ? n15465 : n16519;
  assign n31733 = pi19 ? n31732 : n32;
  assign n31734 = pi18 ? n31731 : n31733;
  assign n31735 = pi17 ? n31729 : n31734;
  assign n31736 = pi16 ? n31722 : n31735;
  assign n31737 = pi15 ? n31718 : n31736;
  assign n31738 = pi14 ? n31709 : n31737;
  assign n31739 = pi21 ? n12608 : n569;
  assign n31740 = pi20 ? n32 : n31739;
  assign n31741 = pi19 ? n32 : n31740;
  assign n31742 = pi20 ? n3335 : n604;
  assign n31743 = pi21 ? n4938 : n569;
  assign n31744 = pi20 ? n31743 : n2004;
  assign n31745 = pi19 ? n31742 : n31744;
  assign n31746 = pi18 ? n31741 : n31745;
  assign n31747 = pi17 ? n32 : n31746;
  assign n31748 = pi19 ? n577 : n610;
  assign n31749 = pi21 ? n13253 : n335;
  assign n31750 = pi20 ? n31749 : n605;
  assign n31751 = pi19 ? n611 : n31750;
  assign n31752 = pi18 ? n31748 : n31751;
  assign n31753 = pi19 ? n612 : n19405;
  assign n31754 = pi21 ? n15689 : n32;
  assign n31755 = pi20 ? n233 : n31754;
  assign n31756 = pi19 ? n31755 : n32;
  assign n31757 = pi18 ? n31753 : n31756;
  assign n31758 = pi17 ? n31752 : n31757;
  assign n31759 = pi16 ? n31747 : n31758;
  assign n31760 = pi21 ? n2091 : n335;
  assign n31761 = pi20 ? n604 : n31760;
  assign n31762 = pi20 ? n2092 : n647;
  assign n31763 = pi19 ? n31761 : n31762;
  assign n31764 = pi21 ? n335 : n2048;
  assign n31765 = pi20 ? n31764 : n13527;
  assign n31766 = pi20 ? n15465 : n25957;
  assign n31767 = pi19 ? n31765 : n31766;
  assign n31768 = pi18 ? n31763 : n31767;
  assign n31769 = pi21 ? n13253 : n233;
  assign n31770 = pi21 ? n569 : n6376;
  assign n31771 = pi20 ? n31769 : n31770;
  assign n31772 = pi19 ? n31771 : n7981;
  assign n31773 = pi20 ? n233 : n8273;
  assign n31774 = pi19 ? n31773 : n32;
  assign n31775 = pi18 ? n31772 : n31774;
  assign n31776 = pi17 ? n31768 : n31775;
  assign n31777 = pi16 ? n30654 : n31776;
  assign n31778 = pi15 ? n31759 : n31777;
  assign n31779 = pi18 ? n8884 : n4985;
  assign n31780 = pi17 ? n32 : n31779;
  assign n31781 = pi20 ? n335 : n30674;
  assign n31782 = pi20 ? n14223 : n31764;
  assign n31783 = pi19 ? n31781 : n31782;
  assign n31784 = pi19 ? n13527 : n31766;
  assign n31785 = pi18 ? n31783 : n31784;
  assign n31786 = pi20 ? n28669 : n13527;
  assign n31787 = pi19 ? n31786 : n233;
  assign n31788 = pi18 ? n31787 : n30648;
  assign n31789 = pi17 ? n31785 : n31788;
  assign n31790 = pi16 ? n31780 : n31789;
  assign n31791 = pi20 ? n570 : n3335;
  assign n31792 = pi19 ? n648 : n31791;
  assign n31793 = pi18 ? n374 : n31792;
  assign n31794 = pi17 ? n32 : n31793;
  assign n31795 = pi20 ? n6358 : n639;
  assign n31796 = pi19 ? n649 : n31795;
  assign n31797 = pi20 ? n639 : n25947;
  assign n31798 = pi21 ? n6361 : n37;
  assign n31799 = pi20 ? n21160 : n31798;
  assign n31800 = pi19 ? n31797 : n31799;
  assign n31801 = pi18 ? n31796 : n31800;
  assign n31802 = pi21 ? n13253 : n2048;
  assign n31803 = pi20 ? n31802 : n30354;
  assign n31804 = pi19 ? n31803 : n233;
  assign n31805 = pi18 ? n31804 : n30648;
  assign n31806 = pi17 ? n31801 : n31805;
  assign n31807 = pi16 ? n31794 : n31806;
  assign n31808 = pi15 ? n31790 : n31807;
  assign n31809 = pi14 ? n31778 : n31808;
  assign n31810 = pi13 ? n31738 : n31809;
  assign n31811 = pi21 ? n2048 : n2091;
  assign n31812 = pi20 ? n37 : n31811;
  assign n31813 = pi19 ? n31812 : n6359;
  assign n31814 = pi20 ? n233 : n6358;
  assign n31815 = pi19 ? n7706 : n31814;
  assign n31816 = pi18 ? n31813 : n31815;
  assign n31817 = pi20 ? n14223 : n8927;
  assign n31818 = pi19 ? n31817 : n233;
  assign n31819 = pi18 ? n31818 : n30664;
  assign n31820 = pi17 ? n31816 : n31819;
  assign n31821 = pi16 ? n439 : n31820;
  assign n31822 = pi20 ? n233 : n7035;
  assign n31823 = pi19 ? n31822 : n32;
  assign n31824 = pi18 ? n19910 : n31823;
  assign n31825 = pi17 ? n37 : n31824;
  assign n31826 = pi16 ? n439 : n31825;
  assign n31827 = pi15 ? n31821 : n31826;
  assign n31828 = pi20 ? n685 : n7724;
  assign n31829 = pi19 ? n31828 : n32;
  assign n31830 = pi18 ? n16239 : n31829;
  assign n31831 = pi17 ? n37 : n31830;
  assign n31832 = pi16 ? n439 : n31831;
  assign n31833 = pi22 ? n4537 : n363;
  assign n31834 = pi21 ? n31833 : n99;
  assign n31835 = pi20 ? n31834 : n99;
  assign n31836 = pi19 ? n99 : n31835;
  assign n31837 = pi18 ? n99 : n31836;
  assign n31838 = pi20 ? n99 : n25199;
  assign n31839 = pi19 ? n99 : n31838;
  assign n31840 = pi18 ? n31839 : n31829;
  assign n31841 = pi17 ? n31837 : n31840;
  assign n31842 = pi16 ? n721 : n31841;
  assign n31843 = pi15 ? n31832 : n31842;
  assign n31844 = pi14 ? n31827 : n31843;
  assign n31845 = pi18 ? n26031 : n363;
  assign n31846 = pi17 ? n32 : n31845;
  assign n31847 = pi20 ? n19084 : n3210;
  assign n31848 = pi19 ? n31847 : n32;
  assign n31849 = pi18 ? n30799 : n31848;
  assign n31850 = pi17 ? n363 : n31849;
  assign n31851 = pi16 ? n31846 : n31850;
  assign n31852 = pi20 ? n19084 : n10011;
  assign n31853 = pi19 ? n31852 : n32;
  assign n31854 = pi18 ? n363 : n31853;
  assign n31855 = pi17 ? n363 : n31854;
  assign n31856 = pi16 ? n21219 : n31855;
  assign n31857 = pi15 ? n31851 : n31856;
  assign n31858 = pi20 ? n2721 : n1822;
  assign n31859 = pi19 ? n31858 : n32;
  assign n31860 = pi18 ? n363 : n31859;
  assign n31861 = pi17 ? n363 : n31860;
  assign n31862 = pi16 ? n21219 : n31861;
  assign n31863 = pi22 ? n157 : n1475;
  assign n31864 = pi21 ? n685 : n31863;
  assign n31865 = pi20 ? n31864 : n32;
  assign n31866 = pi19 ? n31865 : n32;
  assign n31867 = pi18 ? n30799 : n31866;
  assign n31868 = pi17 ? n363 : n31867;
  assign n31869 = pi16 ? n26062 : n31868;
  assign n31870 = pi15 ? n31862 : n31869;
  assign n31871 = pi14 ? n31857 : n31870;
  assign n31872 = pi13 ? n31844 : n31871;
  assign n31873 = pi12 ? n31810 : n31872;
  assign n31874 = pi11 ? n31678 : n31873;
  assign n31875 = pi10 ? n31507 : n31874;
  assign n31876 = pi09 ? n31244 : n31875;
  assign n31877 = pi22 ? n30867 : n20563;
  assign n31878 = pi21 ? n31877 : n30195;
  assign n31879 = pi20 ? n20563 : n31878;
  assign n31880 = pi19 ? n31879 : n16999;
  assign n31881 = pi18 ? n30119 : n31880;
  assign n31882 = pi17 ? n32 : n31881;
  assign n31883 = pi16 ? n31882 : n31217;
  assign n31884 = pi15 ? n32 : n31883;
  assign n31885 = pi22 ? n30195 : n20563;
  assign n31886 = pi21 ? n30116 : n31885;
  assign n31887 = pi20 ? n32 : n31886;
  assign n31888 = pi19 ? n32 : n31887;
  assign n31889 = pi22 ? n30867 : n30195;
  assign n31890 = pi22 ? n37 : n30867;
  assign n31891 = pi21 ? n31889 : n31890;
  assign n31892 = pi20 ? n31891 : n31298;
  assign n31893 = pi19 ? n31892 : n19773;
  assign n31894 = pi18 ? n31888 : n31893;
  assign n31895 = pi17 ? n32 : n31894;
  assign n31896 = pi16 ? n31895 : n31237;
  assign n31897 = pi15 ? n31226 : n31896;
  assign n31898 = pi14 ? n31884 : n31897;
  assign n31899 = pi13 ? n32 : n31898;
  assign n31900 = pi12 ? n32 : n31899;
  assign n31901 = pi11 ? n32 : n31900;
  assign n31902 = pi10 ? n32 : n31901;
  assign n31903 = pi21 ? n30843 : n37;
  assign n31904 = pi20 ? n20563 : n31903;
  assign n31905 = pi19 ? n31904 : n23648;
  assign n31906 = pi18 ? n31265 : n31905;
  assign n31907 = pi17 ? n32 : n31906;
  assign n31908 = pi20 ? n17001 : n32;
  assign n31909 = pi19 ? n99 : n31908;
  assign n31910 = pi18 ? n31257 : n31909;
  assign n31911 = pi17 ? n31254 : n31910;
  assign n31912 = pi16 ? n31907 : n31911;
  assign n31913 = pi21 ? n20563 : n31294;
  assign n31914 = pi20 ? n31913 : n37;
  assign n31915 = pi19 ? n31914 : n27249;
  assign n31916 = pi18 ? n31265 : n31915;
  assign n31917 = pi17 ? n32 : n31916;
  assign n31918 = pi20 ? n18052 : n32;
  assign n31919 = pi19 ? n99 : n31918;
  assign n31920 = pi18 ? n99 : n31919;
  assign n31921 = pi17 ? n99 : n31920;
  assign n31922 = pi16 ? n31917 : n31921;
  assign n31923 = pi15 ? n31912 : n31922;
  assign n31924 = pi22 ? n20563 : n30195;
  assign n31925 = pi21 ? n20563 : n31924;
  assign n31926 = pi20 ? n31925 : n37;
  assign n31927 = pi19 ? n31926 : n99;
  assign n31928 = pi18 ? n31265 : n31927;
  assign n31929 = pi17 ? n32 : n31928;
  assign n31930 = pi21 ? n10165 : n32;
  assign n31931 = pi20 ? n31930 : n32;
  assign n31932 = pi19 ? n99 : n31931;
  assign n31933 = pi18 ? n99 : n31932;
  assign n31934 = pi17 ? n99 : n31933;
  assign n31935 = pi16 ? n31929 : n31934;
  assign n31936 = pi21 ? n31293 : n20563;
  assign n31937 = pi20 ? n32 : n31936;
  assign n31938 = pi19 ? n32 : n31937;
  assign n31939 = pi19 ? n31280 : n37;
  assign n31940 = pi18 ? n31938 : n31939;
  assign n31941 = pi17 ? n32 : n31940;
  assign n31942 = pi19 ? n31305 : n30163;
  assign n31943 = pi18 ? n28217 : n31942;
  assign n31944 = pi17 ? n31304 : n31943;
  assign n31945 = pi16 ? n31941 : n31944;
  assign n31946 = pi15 ? n31935 : n31945;
  assign n31947 = pi14 ? n31923 : n31946;
  assign n31948 = pi21 ? n31889 : n37;
  assign n31949 = pi20 ? n31948 : n37;
  assign n31950 = pi19 ? n31949 : n37;
  assign n31951 = pi18 ? n31938 : n31950;
  assign n31952 = pi17 ? n32 : n31951;
  assign n31953 = pi18 ? n37 : n14883;
  assign n31954 = pi20 ? n21635 : n7346;
  assign n31955 = pi19 ? n23302 : n31954;
  assign n31956 = pi20 ? n2970 : n21635;
  assign n31957 = pi20 ? n16621 : n32;
  assign n31958 = pi19 ? n31956 : n31957;
  assign n31959 = pi18 ? n31955 : n31958;
  assign n31960 = pi17 ? n31953 : n31959;
  assign n31961 = pi16 ? n31952 : n31960;
  assign n31962 = pi23 ? n157 : n531;
  assign n31963 = pi22 ? n31962 : n32;
  assign n31964 = pi21 ? n31963 : n32;
  assign n31965 = pi20 ? n31964 : n32;
  assign n31966 = pi19 ? n9769 : n31965;
  assign n31967 = pi18 ? n31337 : n31966;
  assign n31968 = pi17 ? n37 : n31967;
  assign n31969 = pi16 ? n31317 : n31968;
  assign n31970 = pi15 ? n31961 : n31969;
  assign n31971 = pi19 ? n8765 : n3158;
  assign n31972 = pi18 ? n37 : n31971;
  assign n31973 = pi17 ? n37 : n31972;
  assign n31974 = pi16 ? n31317 : n31973;
  assign n31975 = pi19 ? n139 : n3177;
  assign n31976 = pi18 ? n31352 : n31975;
  assign n31977 = pi17 ? n37 : n31976;
  assign n31978 = pi16 ? n31317 : n31977;
  assign n31979 = pi15 ? n31974 : n31978;
  assign n31980 = pi14 ? n31970 : n31979;
  assign n31981 = pi13 ? n31947 : n31980;
  assign n31982 = pi22 ? n31292 : n30867;
  assign n31983 = pi21 ? n31982 : n37;
  assign n31984 = pi20 ? n32 : n31983;
  assign n31985 = pi19 ? n32 : n31984;
  assign n31986 = pi18 ? n31985 : n37;
  assign n31987 = pi17 ? n32 : n31986;
  assign n31988 = pi20 ? n17619 : n32;
  assign n31989 = pi19 ? n139 : n31988;
  assign n31990 = pi18 ? n37 : n31989;
  assign n31991 = pi17 ? n37 : n31990;
  assign n31992 = pi16 ? n31987 : n31991;
  assign n31993 = pi23 ? n20564 : n37;
  assign n31994 = pi22 ? n31993 : n30195;
  assign n31995 = pi21 ? n31994 : n37;
  assign n31996 = pi20 ? n32 : n31995;
  assign n31997 = pi19 ? n32 : n31996;
  assign n31998 = pi18 ? n31997 : n37;
  assign n31999 = pi17 ? n32 : n31998;
  assign n32000 = pi19 ? n8765 : n4111;
  assign n32001 = pi18 ? n31364 : n32000;
  assign n32002 = pi17 ? n30273 : n32001;
  assign n32003 = pi16 ? n31999 : n32002;
  assign n32004 = pi15 ? n31992 : n32003;
  assign n32005 = pi19 ? n139 : n4117;
  assign n32006 = pi18 ? n31374 : n32005;
  assign n32007 = pi17 ? n31372 : n32006;
  assign n32008 = pi16 ? n31999 : n32007;
  assign n32009 = pi22 ? n31292 : n37;
  assign n32010 = pi21 ? n32009 : n37;
  assign n32011 = pi20 ? n32 : n32010;
  assign n32012 = pi19 ? n32 : n32011;
  assign n32013 = pi18 ? n32012 : n37;
  assign n32014 = pi17 ? n32 : n32013;
  assign n32015 = pi19 ? n139 : n5831;
  assign n32016 = pi18 ? n17061 : n32015;
  assign n32017 = pi17 ? n30273 : n32016;
  assign n32018 = pi16 ? n32014 : n32017;
  assign n32019 = pi15 ? n32008 : n32018;
  assign n32020 = pi14 ? n32004 : n32019;
  assign n32021 = pi20 ? n649 : n31381;
  assign n32022 = pi19 ? n32021 : n10012;
  assign n32023 = pi18 ? n37 : n32022;
  assign n32024 = pi17 ? n37 : n32023;
  assign n32025 = pi16 ? n439 : n32024;
  assign n32026 = pi19 ? n31387 : n31957;
  assign n32027 = pi18 ? n37 : n32026;
  assign n32028 = pi17 ? n37 : n32027;
  assign n32029 = pi16 ? n439 : n32028;
  assign n32030 = pi15 ? n32025 : n32029;
  assign n32031 = pi19 ? n31393 : n2567;
  assign n32032 = pi18 ? n37 : n32031;
  assign n32033 = pi17 ? n37 : n32032;
  assign n32034 = pi16 ? n439 : n32033;
  assign n32035 = pi15 ? n32034 : n31401;
  assign n32036 = pi14 ? n32030 : n32035;
  assign n32037 = pi13 ? n32020 : n32036;
  assign n32038 = pi12 ? n31981 : n32037;
  assign n32039 = pi19 ? n2095 : n2639;
  assign n32040 = pi18 ? n37 : n32039;
  assign n32041 = pi17 ? n37 : n32040;
  assign n32042 = pi16 ? n439 : n32041;
  assign n32043 = pi19 ? n31411 : n2654;
  assign n32044 = pi18 ? n37 : n32043;
  assign n32045 = pi17 ? n37 : n32044;
  assign n32046 = pi16 ? n439 : n32045;
  assign n32047 = pi15 ? n32042 : n32046;
  assign n32048 = pi19 ? n31411 : n2555;
  assign n32049 = pi18 ? n31418 : n32048;
  assign n32050 = pi17 ? n37 : n32049;
  assign n32051 = pi16 ? n439 : n32050;
  assign n32052 = pi15 ? n32051 : n31426;
  assign n32053 = pi14 ? n32047 : n32052;
  assign n32054 = pi13 ? n32053 : n31452;
  assign n32055 = pi21 ? n363 : n2147;
  assign n32056 = pi20 ? n363 : n32055;
  assign n32057 = pi19 ? n32056 : n32;
  assign n32058 = pi18 ? n31484 : n32057;
  assign n32059 = pi17 ? n31481 : n32058;
  assign n32060 = pi16 ? n439 : n32059;
  assign n32061 = pi15 ? n31478 : n32060;
  assign n32062 = pi20 ? n19959 : n2148;
  assign n32063 = pi19 ? n32062 : n32;
  assign n32064 = pi18 ? n37 : n32063;
  assign n32065 = pi17 ? n37 : n32064;
  assign n32066 = pi16 ? n439 : n32065;
  assign n32067 = pi20 ? n31497 : n2148;
  assign n32068 = pi19 ? n32067 : n32;
  assign n32069 = pi18 ? n37 : n32068;
  assign n32070 = pi17 ? n37 : n32069;
  assign n32071 = pi16 ? n439 : n32070;
  assign n32072 = pi15 ? n32066 : n32071;
  assign n32073 = pi14 ? n32061 : n32072;
  assign n32074 = pi13 ? n31472 : n32073;
  assign n32075 = pi12 ? n32054 : n32074;
  assign n32076 = pi11 ? n32038 : n32075;
  assign n32077 = pi20 ? n685 : n16787;
  assign n32078 = pi19 ? n32077 : n32;
  assign n32079 = pi18 ? n31517 : n32078;
  assign n32080 = pi17 ? n31514 : n32079;
  assign n32081 = pi16 ? n31510 : n32080;
  assign n32082 = pi21 ? n157 : n397;
  assign n32083 = pi20 ? n776 : n32082;
  assign n32084 = pi19 ? n32083 : n32;
  assign n32085 = pi18 ? n31523 : n32084;
  assign n32086 = pi17 ? n99 : n32085;
  assign n32087 = pi16 ? n31522 : n32086;
  assign n32088 = pi15 ? n32081 : n32087;
  assign n32089 = pi21 ? n3562 : n397;
  assign n32090 = pi20 ? n30445 : n32089;
  assign n32091 = pi19 ? n32090 : n32;
  assign n32092 = pi18 ? n9985 : n32091;
  assign n32093 = pi17 ? n99 : n32092;
  assign n32094 = pi16 ? n1676 : n32093;
  assign n32095 = pi21 ? n777 : n5178;
  assign n32096 = pi20 ? n18291 : n32095;
  assign n32097 = pi19 ? n32096 : n32;
  assign n32098 = pi18 ? n99 : n32097;
  assign n32099 = pi17 ? n99 : n32098;
  assign n32100 = pi16 ? n31532 : n32099;
  assign n32101 = pi15 ? n32094 : n32100;
  assign n32102 = pi14 ? n32088 : n32101;
  assign n32103 = pi18 ? n99 : n31018;
  assign n32104 = pi17 ? n99 : n32103;
  assign n32105 = pi16 ? n801 : n32104;
  assign n32106 = pi21 ? n3493 : n5178;
  assign n32107 = pi20 ? n99 : n32106;
  assign n32108 = pi19 ? n32107 : n32;
  assign n32109 = pi18 ? n99 : n32108;
  assign n32110 = pi17 ? n99 : n32109;
  assign n32111 = pi16 ? n744 : n32110;
  assign n32112 = pi15 ? n32105 : n32111;
  assign n32113 = pi21 ? n159 : n5178;
  assign n32114 = pi20 ? n30475 : n32113;
  assign n32115 = pi19 ? n32114 : n32;
  assign n32116 = pi18 ? n31549 : n32115;
  assign n32117 = pi17 ? n30472 : n32116;
  assign n32118 = pi16 ? n30470 : n32117;
  assign n32119 = pi19 ? n5276 : n32;
  assign n32120 = pi18 ? n30482 : n32119;
  assign n32121 = pi17 ? n30472 : n32120;
  assign n32122 = pi16 ? n30470 : n32121;
  assign n32123 = pi15 ? n32118 : n32122;
  assign n32124 = pi14 ? n32112 : n32123;
  assign n32125 = pi13 ? n32102 : n32124;
  assign n32126 = pi24 ? n204 : n13481;
  assign n32127 = pi23 ? n316 : n32126;
  assign n32128 = pi22 ? n32127 : n32;
  assign n32129 = pi21 ? n316 : n32128;
  assign n32130 = pi20 ? n316 : n32129;
  assign n32131 = pi19 ? n32130 : n32;
  assign n32132 = pi18 ? n10078 : n32131;
  assign n32133 = pi17 ? n31566 : n32132;
  assign n32134 = pi16 ? n31564 : n32133;
  assign n32135 = pi20 ? n316 : n2816;
  assign n32136 = pi19 ? n32135 : n32;
  assign n32137 = pi18 ? n31578 : n32136;
  assign n32138 = pi17 ? n31576 : n32137;
  assign n32139 = pi16 ? n31573 : n32138;
  assign n32140 = pi15 ? n32134 : n32139;
  assign n32141 = pi18 ? n31595 : n32136;
  assign n32142 = pi17 ? n31593 : n32141;
  assign n32143 = pi16 ? n31587 : n32142;
  assign n32144 = pi21 ? n935 : n3668;
  assign n32145 = pi20 ? n32 : n32144;
  assign n32146 = pi19 ? n32 : n32145;
  assign n32147 = pi20 ? n1693 : n13121;
  assign n32148 = pi19 ? n32147 : n31604;
  assign n32149 = pi18 ? n32146 : n32148;
  assign n32150 = pi17 ? n32 : n32149;
  assign n32151 = pi21 ? n916 : n760;
  assign n32152 = pi20 ? n922 : n32151;
  assign n32153 = pi19 ? n32152 : n32;
  assign n32154 = pi18 ? n31613 : n32153;
  assign n32155 = pi17 ? n31610 : n32154;
  assign n32156 = pi16 ? n32150 : n32155;
  assign n32157 = pi15 ? n32143 : n32156;
  assign n32158 = pi14 ? n32140 : n32157;
  assign n32159 = pi21 ? n204 : n3319;
  assign n32160 = pi20 ? n204 : n32159;
  assign n32161 = pi19 ? n32160 : n32;
  assign n32162 = pi18 ? n204 : n32161;
  assign n32163 = pi17 ? n204 : n32162;
  assign n32164 = pi16 ? n31629 : n32163;
  assign n32165 = pi21 ? n204 : n3339;
  assign n32166 = pi20 ? n204 : n32165;
  assign n32167 = pi19 ? n32166 : n32;
  assign n32168 = pi18 ? n204 : n32167;
  assign n32169 = pi17 ? n204 : n32168;
  assign n32170 = pi16 ? n31643 : n32169;
  assign n32171 = pi15 ? n32164 : n32170;
  assign n32172 = pi21 ? n11808 : n2578;
  assign n32173 = pi20 ? n204 : n32172;
  assign n32174 = pi19 ? n32173 : n32;
  assign n32175 = pi18 ? n31656 : n32174;
  assign n32176 = pi17 ? n139 : n32175;
  assign n32177 = pi16 ? n31655 : n32176;
  assign n32178 = pi21 ? n11808 : n2637;
  assign n32179 = pi20 ? n204 : n32178;
  assign n32180 = pi19 ? n32179 : n32;
  assign n32181 = pi18 ? n30556 : n32180;
  assign n32182 = pi17 ? n31668 : n32181;
  assign n32183 = pi16 ? n31666 : n32182;
  assign n32184 = pi15 ? n32177 : n32183;
  assign n32185 = pi14 ? n32171 : n32184;
  assign n32186 = pi13 ? n32158 : n32185;
  assign n32187 = pi12 ? n32125 : n32186;
  assign n32188 = pi20 ? n31687 : n22582;
  assign n32189 = pi19 ? n32188 : n32;
  assign n32190 = pi18 ? n31686 : n32189;
  assign n32191 = pi17 ? n31683 : n32190;
  assign n32192 = pi16 ? n439 : n32191;
  assign n32193 = pi21 ? n8869 : n928;
  assign n32194 = pi20 ? n7980 : n32193;
  assign n32195 = pi19 ? n32194 : n32;
  assign n32196 = pi18 ? n335 : n32195;
  assign n32197 = pi17 ? n31702 : n32196;
  assign n32198 = pi16 ? n31700 : n32197;
  assign n32199 = pi15 ? n32192 : n32198;
  assign n32200 = pi21 ? n11837 : n32;
  assign n32201 = pi20 ? n15457 : n32200;
  assign n32202 = pi19 ? n32201 : n32;
  assign n32203 = pi18 ? n335 : n32202;
  assign n32204 = pi17 ? n30618 : n32203;
  assign n32205 = pi16 ? n31711 : n32204;
  assign n32206 = pi20 ? n15465 : n16944;
  assign n32207 = pi19 ? n32206 : n32;
  assign n32208 = pi18 ? n31731 : n32207;
  assign n32209 = pi17 ? n31729 : n32208;
  assign n32210 = pi16 ? n31722 : n32209;
  assign n32211 = pi15 ? n32205 : n32210;
  assign n32212 = pi14 ? n32199 : n32211;
  assign n32213 = pi20 ? n233 : n9441;
  assign n32214 = pi19 ? n32213 : n32;
  assign n32215 = pi18 ? n31753 : n32214;
  assign n32216 = pi17 ? n31752 : n32215;
  assign n32217 = pi16 ? n31747 : n32216;
  assign n32218 = pi20 ? n233 : n16519;
  assign n32219 = pi19 ? n32218 : n32;
  assign n32220 = pi18 ? n31772 : n32219;
  assign n32221 = pi17 ? n31768 : n32220;
  assign n32222 = pi16 ? n30654 : n32221;
  assign n32223 = pi15 ? n32217 : n32222;
  assign n32224 = pi18 ? n374 : n4985;
  assign n32225 = pi17 ? n32 : n32224;
  assign n32226 = pi18 ? n31787 : n32219;
  assign n32227 = pi17 ? n31785 : n32226;
  assign n32228 = pi16 ? n32225 : n32227;
  assign n32229 = pi18 ? n31804 : n20844;
  assign n32230 = pi17 ? n31801 : n32229;
  assign n32231 = pi16 ? n31794 : n32230;
  assign n32232 = pi15 ? n32228 : n32231;
  assign n32233 = pi14 ? n32223 : n32232;
  assign n32234 = pi13 ? n32212 : n32233;
  assign n32235 = pi18 ? n31818 : n31127;
  assign n32236 = pi17 ? n31816 : n32235;
  assign n32237 = pi16 ? n439 : n32236;
  assign n32238 = pi18 ? n19910 : n31127;
  assign n32239 = pi17 ? n37 : n32238;
  assign n32240 = pi16 ? n439 : n32239;
  assign n32241 = pi15 ? n32237 : n32240;
  assign n32242 = pi20 ? n685 : n8295;
  assign n32243 = pi19 ? n32242 : n32;
  assign n32244 = pi18 ? n16239 : n32243;
  assign n32245 = pi17 ? n37 : n32244;
  assign n32246 = pi16 ? n439 : n32245;
  assign n32247 = pi18 ? n31839 : n32243;
  assign n32248 = pi17 ? n31837 : n32247;
  assign n32249 = pi16 ? n721 : n32248;
  assign n32250 = pi15 ? n32246 : n32249;
  assign n32251 = pi14 ? n32241 : n32250;
  assign n32252 = pi20 ? n19084 : n4008;
  assign n32253 = pi19 ? n32252 : n32;
  assign n32254 = pi18 ? n30799 : n32253;
  assign n32255 = pi17 ? n363 : n32254;
  assign n32256 = pi16 ? n31846 : n32255;
  assign n32257 = pi21 ? n19697 : n32;
  assign n32258 = pi20 ? n19084 : n32257;
  assign n32259 = pi19 ? n32258 : n32;
  assign n32260 = pi18 ? n363 : n32259;
  assign n32261 = pi17 ? n363 : n32260;
  assign n32262 = pi16 ? n21219 : n32261;
  assign n32263 = pi15 ? n32256 : n32262;
  assign n32264 = pi16 ? n21561 : n31861;
  assign n32265 = pi16 ? n21561 : n31868;
  assign n32266 = pi15 ? n32264 : n32265;
  assign n32267 = pi14 ? n32263 : n32266;
  assign n32268 = pi13 ? n32251 : n32267;
  assign n32269 = pi12 ? n32234 : n32268;
  assign n32270 = pi11 ? n32187 : n32269;
  assign n32271 = pi10 ? n32076 : n32270;
  assign n32272 = pi09 ? n31902 : n32271;
  assign n32273 = pi08 ? n31876 : n32272;
  assign n32274 = pi07 ? n31199 : n32273;
  assign n32275 = pi19 ? n20563 : n31280;
  assign n32276 = pi18 ? n30119 : n32275;
  assign n32277 = pi17 ? n32 : n32276;
  assign n32278 = pi20 ? n3046 : n220;
  assign n32279 = pi19 ? n37 : n32278;
  assign n32280 = pi18 ? n37 : n32279;
  assign n32281 = pi19 ? n99 : n4561;
  assign n32282 = pi18 ? n99 : n32281;
  assign n32283 = pi17 ? n32280 : n32282;
  assign n32284 = pi16 ? n32277 : n32283;
  assign n32285 = pi15 ? n32 : n32284;
  assign n32286 = pi21 ? n31294 : n37;
  assign n32287 = pi20 ? n32286 : n37;
  assign n32288 = pi19 ? n20563 : n32287;
  assign n32289 = pi18 ? n30137 : n32288;
  assign n32290 = pi17 ? n32 : n32289;
  assign n32291 = pi18 ? n37 : n30851;
  assign n32292 = pi17 ? n32291 : n32282;
  assign n32293 = pi16 ? n32290 : n32292;
  assign n32294 = pi20 ? n20563 : n31266;
  assign n32295 = pi19 ? n32294 : n37;
  assign n32296 = pi18 ? n30119 : n32295;
  assign n32297 = pi17 ? n32 : n32296;
  assign n32298 = pi19 ? n26407 : n19773;
  assign n32299 = pi18 ? n37 : n32298;
  assign n32300 = pi22 ? n745 : n32;
  assign n32301 = pi21 ? n32300 : n32;
  assign n32302 = pi20 ? n32301 : n32;
  assign n32303 = pi19 ? n99 : n32302;
  assign n32304 = pi18 ? n99 : n32303;
  assign n32305 = pi17 ? n32299 : n32304;
  assign n32306 = pi16 ? n32297 : n32305;
  assign n32307 = pi15 ? n32293 : n32306;
  assign n32308 = pi14 ? n32285 : n32307;
  assign n32309 = pi13 ? n32 : n32308;
  assign n32310 = pi12 ? n32 : n32309;
  assign n32311 = pi11 ? n32 : n32310;
  assign n32312 = pi10 ? n32 : n32311;
  assign n32313 = pi21 ? n20563 : n30843;
  assign n32314 = pi20 ? n20563 : n32313;
  assign n32315 = pi19 ? n32314 : n37;
  assign n32316 = pi18 ? n31265 : n32315;
  assign n32317 = pi17 ? n32 : n32316;
  assign n32318 = pi22 ? n1656 : n32;
  assign n32319 = pi21 ? n32318 : n32;
  assign n32320 = pi20 ? n32319 : n32;
  assign n32321 = pi19 ? n99 : n32320;
  assign n32322 = pi18 ? n18854 : n32321;
  assign n32323 = pi17 ? n37 : n32322;
  assign n32324 = pi16 ? n32317 : n32323;
  assign n32325 = pi18 ? n31265 : n32295;
  assign n32326 = pi17 ? n32 : n32325;
  assign n32327 = pi20 ? n7747 : n7745;
  assign n32328 = pi20 ? n2181 : n2191;
  assign n32329 = pi19 ? n32327 : n32328;
  assign n32330 = pi18 ? n27245 : n32329;
  assign n32331 = pi18 ? n99 : n32321;
  assign n32332 = pi17 ? n32330 : n32331;
  assign n32333 = pi16 ? n32326 : n32332;
  assign n32334 = pi15 ? n32324 : n32333;
  assign n32335 = pi20 ? n2974 : n220;
  assign n32336 = pi19 ? n31221 : n32335;
  assign n32337 = pi18 ? n31265 : n32336;
  assign n32338 = pi17 ? n32 : n32337;
  assign n32339 = pi19 ? n29428 : n18853;
  assign n32340 = pi19 ? n99 : n219;
  assign n32341 = pi18 ? n32339 : n32340;
  assign n32342 = pi21 ? n11427 : n32;
  assign n32343 = pi20 ? n32342 : n32;
  assign n32344 = pi19 ? n99 : n32343;
  assign n32345 = pi18 ? n28236 : n32344;
  assign n32346 = pi17 ? n32341 : n32345;
  assign n32347 = pi16 ? n32338 : n32346;
  assign n32348 = pi20 ? n20563 : n37;
  assign n32349 = pi19 ? n32348 : n37;
  assign n32350 = pi18 ? n31315 : n32349;
  assign n32351 = pi17 ? n32 : n32350;
  assign n32352 = pi20 ? n2973 : n2958;
  assign n32353 = pi20 ? n2973 : n5077;
  assign n32354 = pi19 ? n32352 : n32353;
  assign n32355 = pi20 ? n181 : n2191;
  assign n32356 = pi21 ? n10511 : n32;
  assign n32357 = pi20 ? n32356 : n32;
  assign n32358 = pi19 ? n32355 : n32357;
  assign n32359 = pi18 ? n32354 : n32358;
  assign n32360 = pi17 ? n37 : n32359;
  assign n32361 = pi16 ? n32351 : n32360;
  assign n32362 = pi15 ? n32347 : n32361;
  assign n32363 = pi14 ? n32334 : n32362;
  assign n32364 = pi20 ? n18017 : n32;
  assign n32365 = pi19 ? n9824 : n32364;
  assign n32366 = pi18 ? n37 : n32365;
  assign n32367 = pi17 ? n37 : n32366;
  assign n32368 = pi16 ? n32351 : n32367;
  assign n32369 = pi19 ? n31926 : n37;
  assign n32370 = pi18 ? n31315 : n32369;
  assign n32371 = pi17 ? n32 : n32370;
  assign n32372 = pi19 ? n37 : n32364;
  assign n32373 = pi18 ? n37 : n32372;
  assign n32374 = pi17 ? n37 : n32373;
  assign n32375 = pi16 ? n32371 : n32374;
  assign n32376 = pi15 ? n32368 : n32375;
  assign n32377 = pi19 ? n31267 : n37;
  assign n32378 = pi18 ? n31315 : n32377;
  assign n32379 = pi17 ? n32 : n32378;
  assign n32380 = pi16 ? n32379 : n31973;
  assign n32381 = pi18 ? n31315 : n31939;
  assign n32382 = pi17 ? n32 : n32381;
  assign n32383 = pi16 ? n32382 : n31973;
  assign n32384 = pi15 ? n32380 : n32383;
  assign n32385 = pi14 ? n32376 : n32384;
  assign n32386 = pi13 ? n32363 : n32385;
  assign n32387 = pi18 ? n31938 : n37;
  assign n32388 = pi17 ? n32 : n32387;
  assign n32389 = pi19 ? n8765 : n31988;
  assign n32390 = pi18 ? n37 : n32389;
  assign n32391 = pi17 ? n37 : n32390;
  assign n32392 = pi16 ? n32388 : n32391;
  assign n32393 = pi18 ? n31297 : n37;
  assign n32394 = pi17 ? n32 : n32393;
  assign n32395 = pi19 ? n9769 : n31988;
  assign n32396 = pi18 ? n37 : n32395;
  assign n32397 = pi17 ? n37 : n32396;
  assign n32398 = pi16 ? n32394 : n32397;
  assign n32399 = pi15 ? n32392 : n32398;
  assign n32400 = pi21 ? n30866 : n31294;
  assign n32401 = pi20 ? n32 : n32400;
  assign n32402 = pi19 ? n32 : n32401;
  assign n32403 = pi18 ? n32402 : n37;
  assign n32404 = pi17 ? n32 : n32403;
  assign n32405 = pi21 ? n24338 : n32;
  assign n32406 = pi20 ? n32405 : n32;
  assign n32407 = pi19 ? n139 : n32406;
  assign n32408 = pi18 ? n37 : n32407;
  assign n32409 = pi17 ? n37 : n32408;
  assign n32410 = pi16 ? n32404 : n32409;
  assign n32411 = pi21 ? n30866 : n37;
  assign n32412 = pi20 ? n32 : n32411;
  assign n32413 = pi19 ? n32 : n32412;
  assign n32414 = pi18 ? n32413 : n37;
  assign n32415 = pi17 ? n32 : n32414;
  assign n32416 = pi20 ? n3096 : n9143;
  assign n32417 = pi19 ? n32416 : n5005;
  assign n32418 = pi18 ? n37 : n32417;
  assign n32419 = pi17 ? n37 : n32418;
  assign n32420 = pi16 ? n32415 : n32419;
  assign n32421 = pi15 ? n32410 : n32420;
  assign n32422 = pi14 ? n32399 : n32421;
  assign n32423 = pi19 ? n10681 : n3127;
  assign n32424 = pi18 ? n37 : n32423;
  assign n32425 = pi17 ? n37 : n32424;
  assign n32426 = pi16 ? n32415 : n32425;
  assign n32427 = pi22 ? n31292 : n30195;
  assign n32428 = pi21 ? n32427 : n37;
  assign n32429 = pi20 ? n32 : n32428;
  assign n32430 = pi19 ? n32 : n32429;
  assign n32431 = pi18 ? n32430 : n37;
  assign n32432 = pi17 ? n32 : n32431;
  assign n32433 = pi19 ? n12628 : n31957;
  assign n32434 = pi18 ? n37 : n32433;
  assign n32435 = pi17 ? n37 : n32434;
  assign n32436 = pi16 ? n32432 : n32435;
  assign n32437 = pi15 ? n32426 : n32436;
  assign n32438 = pi20 ? n37 : n20377;
  assign n32439 = pi19 ? n32438 : n2580;
  assign n32440 = pi18 ? n37 : n32439;
  assign n32441 = pi17 ? n37 : n32440;
  assign n32442 = pi16 ? n32014 : n32441;
  assign n32443 = pi19 ? n32438 : n4111;
  assign n32444 = pi18 ? n37 : n32443;
  assign n32445 = pi17 ? n37 : n32444;
  assign n32446 = pi16 ? n439 : n32445;
  assign n32447 = pi15 ? n32442 : n32446;
  assign n32448 = pi14 ? n32437 : n32447;
  assign n32449 = pi13 ? n32422 : n32448;
  assign n32450 = pi12 ? n32386 : n32449;
  assign n32451 = pi16 ? n439 : n32441;
  assign n32452 = pi19 ? n8802 : n37;
  assign n32453 = pi20 ? n571 : n17715;
  assign n32454 = pi19 ? n32453 : n2580;
  assign n32455 = pi18 ? n32452 : n32454;
  assign n32456 = pi17 ? n15070 : n32455;
  assign n32457 = pi16 ? n439 : n32456;
  assign n32458 = pi15 ? n32451 : n32457;
  assign n32459 = pi20 ? n649 : n15465;
  assign n32460 = pi19 ? n32459 : n2580;
  assign n32461 = pi18 ? n7677 : n32460;
  assign n32462 = pi17 ? n37 : n32461;
  assign n32463 = pi16 ? n439 : n32462;
  assign n32464 = pi20 ? n21148 : n18121;
  assign n32465 = pi19 ? n32464 : n2580;
  assign n32466 = pi18 ? n37 : n32465;
  assign n32467 = pi17 ? n15070 : n32466;
  assign n32468 = pi16 ? n439 : n32467;
  assign n32469 = pi15 ? n32463 : n32468;
  assign n32470 = pi14 ? n32458 : n32469;
  assign n32471 = pi21 ? n580 : n2091;
  assign n32472 = pi20 ? n32471 : n233;
  assign n32473 = pi19 ? n32472 : n2580;
  assign n32474 = pi18 ? n37 : n32473;
  assign n32475 = pi17 ? n37 : n32474;
  assign n32476 = pi16 ? n439 : n32475;
  assign n32477 = pi21 ? n37 : n24222;
  assign n32478 = pi20 ? n37 : n32477;
  assign n32479 = pi19 ? n32478 : n2639;
  assign n32480 = pi18 ? n37 : n32479;
  assign n32481 = pi17 ? n37 : n32480;
  assign n32482 = pi16 ? n439 : n32481;
  assign n32483 = pi15 ? n32476 : n32482;
  assign n32484 = pi19 ? n5029 : n7833;
  assign n32485 = pi18 ? n37 : n32484;
  assign n32486 = pi17 ? n37 : n32485;
  assign n32487 = pi16 ? n439 : n32486;
  assign n32488 = pi19 ? n5029 : n2654;
  assign n32489 = pi18 ? n37 : n32488;
  assign n32490 = pi17 ? n37 : n32489;
  assign n32491 = pi16 ? n439 : n32490;
  assign n32492 = pi15 ? n32487 : n32491;
  assign n32493 = pi14 ? n32483 : n32492;
  assign n32494 = pi13 ? n32470 : n32493;
  assign n32495 = pi19 ? n24494 : n2702;
  assign n32496 = pi18 ? n37 : n32495;
  assign n32497 = pi17 ? n37 : n32496;
  assign n32498 = pi16 ? n439 : n32497;
  assign n32499 = pi19 ? n5072 : n2702;
  assign n32500 = pi18 ? n37 : n32499;
  assign n32501 = pi17 ? n37 : n32500;
  assign n32502 = pi16 ? n439 : n32501;
  assign n32503 = pi15 ? n32498 : n32502;
  assign n32504 = pi19 ? n2108 : n2702;
  assign n32505 = pi18 ? n37 : n32504;
  assign n32506 = pi17 ? n37 : n32505;
  assign n32507 = pi16 ? n439 : n32506;
  assign n32508 = pi19 ? n2108 : n1823;
  assign n32509 = pi18 ? n37 : n32508;
  assign n32510 = pi17 ? n37 : n32509;
  assign n32511 = pi16 ? n439 : n32510;
  assign n32512 = pi15 ? n32507 : n32511;
  assign n32513 = pi14 ? n32503 : n32512;
  assign n32514 = pi21 ? n37 : n24858;
  assign n32515 = pi20 ? n37 : n32514;
  assign n32516 = pi19 ? n32515 : n1823;
  assign n32517 = pi18 ? n37 : n32516;
  assign n32518 = pi17 ? n37 : n32517;
  assign n32519 = pi16 ? n439 : n32518;
  assign n32520 = pi22 ? n37 : n759;
  assign n32521 = pi21 ? n37 : n32520;
  assign n32522 = pi20 ? n37 : n32521;
  assign n32523 = pi19 ? n32522 : n32;
  assign n32524 = pi18 ? n37 : n32523;
  assign n32525 = pi17 ? n37 : n32524;
  assign n32526 = pi16 ? n439 : n32525;
  assign n32527 = pi15 ? n32519 : n32526;
  assign n32528 = pi21 ? n37 : n6897;
  assign n32529 = pi20 ? n37 : n32528;
  assign n32530 = pi19 ? n32529 : n32;
  assign n32531 = pi18 ? n37 : n32530;
  assign n32532 = pi17 ? n37 : n32531;
  assign n32533 = pi16 ? n439 : n32532;
  assign n32534 = pi20 ? n37 : n30414;
  assign n32535 = pi19 ? n37 : n32534;
  assign n32536 = pi21 ? n272 : n6897;
  assign n32537 = pi20 ? n157 : n32536;
  assign n32538 = pi19 ? n32537 : n32;
  assign n32539 = pi18 ? n32535 : n32538;
  assign n32540 = pi17 ? n37 : n32539;
  assign n32541 = pi16 ? n439 : n32540;
  assign n32542 = pi15 ? n32533 : n32541;
  assign n32543 = pi14 ? n32527 : n32542;
  assign n32544 = pi13 ? n32513 : n32543;
  assign n32545 = pi12 ? n32494 : n32544;
  assign n32546 = pi11 ? n32450 : n32545;
  assign n32547 = pi18 ? n30851 : n19135;
  assign n32548 = pi20 ? n15263 : n221;
  assign n32549 = pi19 ? n32548 : n11445;
  assign n32550 = pi20 ? n157 : n20013;
  assign n32551 = pi19 ? n32550 : n32;
  assign n32552 = pi18 ? n32549 : n32551;
  assign n32553 = pi17 ? n32547 : n32552;
  assign n32554 = pi16 ? n439 : n32553;
  assign n32555 = pi20 ? n37 : n16008;
  assign n32556 = pi19 ? n37 : n32555;
  assign n32557 = pi18 ? n374 : n32556;
  assign n32558 = pi17 ? n32 : n32557;
  assign n32559 = pi20 ? n2238 : n6523;
  assign n32560 = pi19 ? n99 : n32559;
  assign n32561 = pi18 ? n30851 : n32560;
  assign n32562 = pi21 ? n777 : n1143;
  assign n32563 = pi20 ? n32562 : n99;
  assign n32564 = pi19 ? n32563 : n19134;
  assign n32565 = pi19 ? n6544 : n32;
  assign n32566 = pi18 ? n32564 : n32565;
  assign n32567 = pi17 ? n32561 : n32566;
  assign n32568 = pi16 ? n32558 : n32567;
  assign n32569 = pi15 ? n32554 : n32568;
  assign n32570 = pi20 ? n99 : n6503;
  assign n32571 = pi19 ? n99 : n32570;
  assign n32572 = pi22 ? n157 : n430;
  assign n32573 = pi21 ? n157 : n32572;
  assign n32574 = pi20 ? n157 : n32573;
  assign n32575 = pi19 ? n32574 : n32;
  assign n32576 = pi18 ? n32571 : n32575;
  assign n32577 = pi17 ? n99 : n32576;
  assign n32578 = pi16 ? n23698 : n32577;
  assign n32579 = pi22 ? n99 : n1484;
  assign n32580 = pi21 ? n99 : n32579;
  assign n32581 = pi20 ? n99 : n32580;
  assign n32582 = pi19 ? n99 : n32581;
  assign n32583 = pi21 ? n777 : n5145;
  assign n32584 = pi20 ? n27598 : n32583;
  assign n32585 = pi19 ? n32584 : n32;
  assign n32586 = pi18 ? n32582 : n32585;
  assign n32587 = pi17 ? n99 : n32586;
  assign n32588 = pi16 ? n23698 : n32587;
  assign n32589 = pi15 ? n32578 : n32588;
  assign n32590 = pi14 ? n32569 : n32589;
  assign n32591 = pi21 ? n99 : n5178;
  assign n32592 = pi20 ? n99 : n32591;
  assign n32593 = pi19 ? n32592 : n32;
  assign n32594 = pi18 ? n99 : n32593;
  assign n32595 = pi17 ? n99 : n32594;
  assign n32596 = pi16 ? n801 : n32595;
  assign n32597 = pi16 ? n201 : n32595;
  assign n32598 = pi15 ? n32596 : n32597;
  assign n32599 = pi18 ? n1508 : n30468;
  assign n32600 = pi17 ? n32 : n32599;
  assign n32601 = pi19 ? n6618 : n32;
  assign n32602 = pi18 ? n30474 : n32601;
  assign n32603 = pi17 ? n139 : n32602;
  assign n32604 = pi16 ? n32600 : n32603;
  assign n32605 = pi21 ? n14506 : n37;
  assign n32606 = pi20 ? n32 : n32605;
  assign n32607 = pi19 ? n32 : n32606;
  assign n32608 = pi21 ? n2746 : n2156;
  assign n32609 = pi19 ? n32608 : n22704;
  assign n32610 = pi18 ? n32607 : n32609;
  assign n32611 = pi17 ? n32 : n32610;
  assign n32612 = pi18 ? n139 : n32119;
  assign n32613 = pi17 ? n139 : n32612;
  assign n32614 = pi16 ? n32611 : n32613;
  assign n32615 = pi15 ? n32604 : n32614;
  assign n32616 = pi14 ? n32598 : n32615;
  assign n32617 = pi13 ? n32590 : n32616;
  assign n32618 = pi20 ? n37 : n820;
  assign n32619 = pi19 ? n37 : n32618;
  assign n32620 = pi18 ? n374 : n32619;
  assign n32621 = pi17 ? n32 : n32620;
  assign n32622 = pi18 ? n139 : n31041;
  assign n32623 = pi17 ? n139 : n32622;
  assign n32624 = pi16 ? n32621 : n32623;
  assign n32625 = pi21 ? n916 : n37;
  assign n32626 = pi20 ? n29537 : n32625;
  assign n32627 = pi19 ? n139 : n32626;
  assign n32628 = pi18 ? n8766 : n32627;
  assign n32629 = pi21 ? n4445 : n1018;
  assign n32630 = pi20 ? n139 : n32629;
  assign n32631 = pi19 ? n13093 : n32630;
  assign n32632 = pi18 ? n32631 : n31041;
  assign n32633 = pi17 ? n32628 : n32632;
  assign n32634 = pi16 ? n439 : n32633;
  assign n32635 = pi15 ? n32624 : n32634;
  assign n32636 = pi20 ? n37 : n21732;
  assign n32637 = pi19 ? n32636 : n204;
  assign n32638 = pi18 ? n32637 : n204;
  assign n32639 = pi21 ? n921 : n1056;
  assign n32640 = pi20 ? n32639 : n204;
  assign n32641 = pi21 ? n19302 : n204;
  assign n32642 = pi20 ? n204 : n32641;
  assign n32643 = pi19 ? n32640 : n32642;
  assign n32644 = pi20 ? n1060 : n7969;
  assign n32645 = pi19 ? n32644 : n32;
  assign n32646 = pi18 ? n32643 : n32645;
  assign n32647 = pi17 ? n32638 : n32646;
  assign n32648 = pi16 ? n439 : n32647;
  assign n32649 = pi18 ? n18970 : n204;
  assign n32650 = pi17 ? n32649 : n32162;
  assign n32651 = pi16 ? n439 : n32650;
  assign n32652 = pi15 ? n32648 : n32651;
  assign n32653 = pi14 ? n32635 : n32652;
  assign n32654 = pi20 ? n1003 : n3096;
  assign n32655 = pi19 ? n37 : n32654;
  assign n32656 = pi18 ? n374 : n32655;
  assign n32657 = pi17 ? n32 : n32656;
  assign n32658 = pi19 ? n6268 : n204;
  assign n32659 = pi18 ? n32658 : n204;
  assign n32660 = pi18 ? n204 : n24362;
  assign n32661 = pi17 ? n32659 : n32660;
  assign n32662 = pi16 ? n32657 : n32661;
  assign n32663 = pi20 ? n3096 : n1016;
  assign n32664 = pi19 ? n32663 : n204;
  assign n32665 = pi18 ? n32664 : n204;
  assign n32666 = pi17 ? n32665 : n32168;
  assign n32667 = pi16 ? n439 : n32666;
  assign n32668 = pi15 ? n32662 : n32667;
  assign n32669 = pi21 ? n297 : n233;
  assign n32670 = pi20 ? n32669 : n233;
  assign n32671 = pi19 ? n18082 : n32670;
  assign n32672 = pi18 ? n32671 : n233;
  assign n32673 = pi20 ? n16047 : n233;
  assign n32674 = pi20 ? n233 : n204;
  assign n32675 = pi19 ? n32673 : n32674;
  assign n32676 = pi21 ? n204 : n2578;
  assign n32677 = pi20 ? n204 : n32676;
  assign n32678 = pi19 ? n32677 : n32;
  assign n32679 = pi18 ? n32675 : n32678;
  assign n32680 = pi17 ? n32672 : n32679;
  assign n32681 = pi16 ? n439 : n32680;
  assign n32682 = pi18 ? n374 : n31371;
  assign n32683 = pi17 ? n32 : n32682;
  assign n32684 = pi20 ? n3096 : n997;
  assign n32685 = pi19 ? n32684 : n32670;
  assign n32686 = pi18 ? n32685 : n233;
  assign n32687 = pi21 ? n570 : n139;
  assign n32688 = pi20 ? n32687 : n233;
  assign n32689 = pi21 ? n19337 : n1079;
  assign n32690 = pi20 ? n233 : n32689;
  assign n32691 = pi19 ? n32688 : n32690;
  assign n32692 = pi22 ? n233 : n4079;
  assign n32693 = pi21 ? n32692 : n2637;
  assign n32694 = pi20 ? n23069 : n32693;
  assign n32695 = pi19 ? n32694 : n32;
  assign n32696 = pi18 ? n32691 : n32695;
  assign n32697 = pi17 ? n32686 : n32696;
  assign n32698 = pi16 ? n32683 : n32697;
  assign n32699 = pi15 ? n32681 : n32698;
  assign n32700 = pi14 ? n32668 : n32699;
  assign n32701 = pi13 ? n32653 : n32700;
  assign n32702 = pi12 ? n32617 : n32701;
  assign n32703 = pi20 ? n577 : n233;
  assign n32704 = pi19 ? n37 : n32703;
  assign n32705 = pi21 ? n12983 : n928;
  assign n32706 = pi20 ? n233 : n32705;
  assign n32707 = pi19 ? n32706 : n32;
  assign n32708 = pi18 ? n32704 : n32707;
  assign n32709 = pi17 ? n15129 : n32708;
  assign n32710 = pi16 ? n439 : n32709;
  assign n32711 = pi19 ? n25087 : n335;
  assign n32712 = pi18 ? n32711 : n335;
  assign n32713 = pi21 ? n12994 : n928;
  assign n32714 = pi20 ? n15465 : n32713;
  assign n32715 = pi19 ? n32714 : n32;
  assign n32716 = pi18 ? n12631 : n32715;
  assign n32717 = pi17 ? n32712 : n32716;
  assign n32718 = pi16 ? n439 : n32717;
  assign n32719 = pi15 ? n32710 : n32718;
  assign n32720 = pi19 ? n37 : n8894;
  assign n32721 = pi18 ? n374 : n32720;
  assign n32722 = pi17 ? n32 : n32721;
  assign n32723 = pi20 ? n335 : n37;
  assign n32724 = pi19 ? n32723 : n37;
  assign n32725 = pi18 ? n32724 : n37;
  assign n32726 = pi19 ? n37 : n7696;
  assign n32727 = pi22 ? n233 : n13314;
  assign n32728 = pi21 ? n32727 : n32;
  assign n32729 = pi20 ? n15465 : n32728;
  assign n32730 = pi19 ? n32729 : n32;
  assign n32731 = pi18 ? n32726 : n32730;
  assign n32732 = pi17 ? n32725 : n32731;
  assign n32733 = pi16 ? n32722 : n32732;
  assign n32734 = pi19 ? n6340 : n37;
  assign n32735 = pi18 ? n32734 : n37;
  assign n32736 = pi18 ? n2102 : n21789;
  assign n32737 = pi17 ? n32735 : n32736;
  assign n32738 = pi16 ? n25090 : n32737;
  assign n32739 = pi15 ? n32733 : n32738;
  assign n32740 = pi14 ? n32719 : n32739;
  assign n32741 = pi18 ? n335 : n37;
  assign n32742 = pi17 ? n32741 : n32736;
  assign n32743 = pi16 ? n439 : n32742;
  assign n32744 = pi20 ? n335 : n31764;
  assign n32745 = pi19 ? n32744 : n17533;
  assign n32746 = pi18 ? n32745 : n233;
  assign n32747 = pi20 ? n18174 : n233;
  assign n32748 = pi19 ? n32747 : n233;
  assign n32749 = pi18 ? n32748 : n32219;
  assign n32750 = pi17 ? n32746 : n32749;
  assign n32751 = pi16 ? n439 : n32750;
  assign n32752 = pi15 ? n32743 : n32751;
  assign n32753 = pi19 ? n25087 : n13535;
  assign n32754 = pi18 ? n32753 : n233;
  assign n32755 = pi20 ? n28701 : n7705;
  assign n32756 = pi19 ? n32755 : n233;
  assign n32757 = pi18 ? n32756 : n32219;
  assign n32758 = pi17 ? n32754 : n32757;
  assign n32759 = pi16 ? n439 : n32758;
  assign n32760 = pi20 ? n25146 : n233;
  assign n32761 = pi19 ? n643 : n32760;
  assign n32762 = pi18 ? n32761 : n233;
  assign n32763 = pi20 ? n2094 : n7705;
  assign n32764 = pi19 ? n32763 : n233;
  assign n32765 = pi18 ? n32764 : n20844;
  assign n32766 = pi17 ? n32762 : n32765;
  assign n32767 = pi16 ? n439 : n32766;
  assign n32768 = pi15 ? n32759 : n32767;
  assign n32769 = pi14 ? n32752 : n32768;
  assign n32770 = pi13 ? n32740 : n32769;
  assign n32771 = pi19 ? n26819 : n233;
  assign n32772 = pi19 ? n8927 : n233;
  assign n32773 = pi18 ? n32771 : n32772;
  assign n32774 = pi18 ? n233 : n20844;
  assign n32775 = pi17 ? n32773 : n32774;
  assign n32776 = pi16 ? n439 : n32775;
  assign n32777 = pi20 ? n685 : n22920;
  assign n32778 = pi19 ? n32777 : n32;
  assign n32779 = pi18 ? n2731 : n32778;
  assign n32780 = pi17 ? n37 : n32779;
  assign n32781 = pi16 ? n439 : n32780;
  assign n32782 = pi15 ? n32776 : n32781;
  assign n32783 = pi18 ? n2731 : n32243;
  assign n32784 = pi17 ? n37 : n32783;
  assign n32785 = pi16 ? n439 : n32784;
  assign n32786 = pi20 ? n99 : n28732;
  assign n32787 = pi21 ? n722 : n363;
  assign n32788 = pi21 ? n99 : n722;
  assign n32789 = pi20 ? n32787 : n32788;
  assign n32790 = pi19 ? n32786 : n32789;
  assign n32791 = pi19 ? n99 : n363;
  assign n32792 = pi18 ? n32790 : n32791;
  assign n32793 = pi20 ? n25167 : n30766;
  assign n32794 = pi20 ? n363 : n19084;
  assign n32795 = pi19 ? n32793 : n32794;
  assign n32796 = pi20 ? n18194 : n8295;
  assign n32797 = pi19 ? n32796 : n32;
  assign n32798 = pi18 ? n32795 : n32797;
  assign n32799 = pi17 ? n32792 : n32798;
  assign n32800 = pi16 ? n721 : n32799;
  assign n32801 = pi15 ? n32785 : n32800;
  assign n32802 = pi14 ? n32782 : n32801;
  assign n32803 = pi22 ? n715 : n139;
  assign n32804 = pi21 ? n32803 : n4237;
  assign n32805 = pi20 ? n32 : n32804;
  assign n32806 = pi19 ? n32 : n32805;
  assign n32807 = pi21 ? n4237 : n4247;
  assign n32808 = pi20 ? n32807 : n14846;
  assign n32809 = pi20 ? n99 : n32788;
  assign n32810 = pi19 ? n32808 : n32809;
  assign n32811 = pi18 ? n32806 : n32810;
  assign n32812 = pi17 ? n32 : n32811;
  assign n32813 = pi21 ? n99 : n22549;
  assign n32814 = pi20 ? n99 : n32813;
  assign n32815 = pi20 ? n32813 : n99;
  assign n32816 = pi19 ? n32814 : n32815;
  assign n32817 = pi22 ? n363 : n4543;
  assign n32818 = pi21 ? n99 : n32817;
  assign n32819 = pi20 ? n32818 : n25167;
  assign n32820 = pi19 ? n99 : n32819;
  assign n32821 = pi18 ? n32816 : n32820;
  assign n32822 = pi20 ? n32788 : n30766;
  assign n32823 = pi20 ? n32787 : n25167;
  assign n32824 = pi19 ? n32822 : n32823;
  assign n32825 = pi21 ? n685 : n31444;
  assign n32826 = pi21 ? n25537 : n32;
  assign n32827 = pi20 ? n32825 : n32826;
  assign n32828 = pi19 ? n32827 : n32;
  assign n32829 = pi18 ? n32824 : n32828;
  assign n32830 = pi17 ? n32821 : n32829;
  assign n32831 = pi16 ? n32812 : n32830;
  assign n32832 = pi19 ? n363 : n32794;
  assign n32833 = pi21 ? n363 : n31444;
  assign n32834 = pi20 ? n32833 : n10011;
  assign n32835 = pi19 ? n32834 : n32;
  assign n32836 = pi18 ? n32832 : n32835;
  assign n32837 = pi17 ? n363 : n32836;
  assign n32838 = pi16 ? n26887 : n32837;
  assign n32839 = pi15 ? n32831 : n32838;
  assign n32840 = pi22 ? n12652 : n363;
  assign n32841 = pi21 ? n32840 : n363;
  assign n32842 = pi20 ? n32 : n32841;
  assign n32843 = pi19 ? n32 : n32842;
  assign n32844 = pi18 ? n32843 : n363;
  assign n32845 = pi17 ? n32 : n32844;
  assign n32846 = pi22 ? n685 : n5061;
  assign n32847 = pi21 ? n2721 : n32846;
  assign n32848 = pi20 ? n32847 : n1822;
  assign n32849 = pi19 ? n32848 : n32;
  assign n32850 = pi18 ? n32832 : n32849;
  assign n32851 = pi17 ? n363 : n32850;
  assign n32852 = pi16 ? n32845 : n32851;
  assign n32853 = pi22 ? n685 : n1457;
  assign n32854 = pi21 ? n685 : n32853;
  assign n32855 = pi20 ? n32854 : n32;
  assign n32856 = pi19 ? n32855 : n32;
  assign n32857 = pi18 ? n32832 : n32856;
  assign n32858 = pi17 ? n363 : n32857;
  assign n32859 = pi16 ? n29768 : n32858;
  assign n32860 = pi15 ? n32852 : n32859;
  assign n32861 = pi14 ? n32839 : n32860;
  assign n32862 = pi13 ? n32802 : n32861;
  assign n32863 = pi12 ? n32770 : n32862;
  assign n32864 = pi11 ? n32702 : n32863;
  assign n32865 = pi10 ? n32546 : n32864;
  assign n32866 = pi09 ? n32312 : n32865;
  assign n32867 = pi18 ? n30137 : n32275;
  assign n32868 = pi17 ? n32 : n32867;
  assign n32869 = pi16 ? n32868 : n32283;
  assign n32870 = pi15 ? n32 : n32869;
  assign n32871 = pi20 ? n32313 : n37;
  assign n32872 = pi19 ? n20563 : n32871;
  assign n32873 = pi18 ? n30119 : n32872;
  assign n32874 = pi17 ? n32 : n32873;
  assign n32875 = pi16 ? n32874 : n32292;
  assign n32876 = pi20 ? n20563 : n31925;
  assign n32877 = pi19 ? n32876 : n37;
  assign n32878 = pi18 ? n30119 : n32877;
  assign n32879 = pi17 ? n32 : n32878;
  assign n32880 = pi16 ? n32879 : n32305;
  assign n32881 = pi15 ? n32875 : n32880;
  assign n32882 = pi14 ? n32870 : n32881;
  assign n32883 = pi13 ? n32 : n32882;
  assign n32884 = pi12 ? n32 : n32883;
  assign n32885 = pi11 ? n32 : n32884;
  assign n32886 = pi10 ? n32 : n32885;
  assign n32887 = pi16 ? n32326 : n32323;
  assign n32888 = pi15 ? n32887 : n32333;
  assign n32889 = pi20 ? n37 : n220;
  assign n32890 = pi19 ? n31221 : n32889;
  assign n32891 = pi18 ? n31265 : n32890;
  assign n32892 = pi17 ? n32 : n32891;
  assign n32893 = pi20 ? n18009 : n32;
  assign n32894 = pi19 ? n99 : n32893;
  assign n32895 = pi18 ? n18854 : n32894;
  assign n32896 = pi17 ? n32341 : n32895;
  assign n32897 = pi16 ? n32892 : n32896;
  assign n32898 = pi20 ? n20563 : n30096;
  assign n32899 = pi19 ? n32898 : n37;
  assign n32900 = pi18 ? n31315 : n32899;
  assign n32901 = pi17 ? n32 : n32900;
  assign n32902 = pi16 ? n32901 : n32360;
  assign n32903 = pi15 ? n32897 : n32902;
  assign n32904 = pi14 ? n32888 : n32903;
  assign n32905 = pi23 ? n11117 : n204;
  assign n32906 = pi22 ? n32905 : n32;
  assign n32907 = pi21 ? n32906 : n32;
  assign n32908 = pi20 ? n32907 : n32;
  assign n32909 = pi19 ? n37 : n32908;
  assign n32910 = pi18 ? n37 : n32909;
  assign n32911 = pi17 ? n37 : n32910;
  assign n32912 = pi16 ? n32351 : n32911;
  assign n32913 = pi15 ? n32368 : n32912;
  assign n32914 = pi18 ? n31938 : n32377;
  assign n32915 = pi17 ? n32 : n32914;
  assign n32916 = pi19 ? n8765 : n3972;
  assign n32917 = pi18 ? n37 : n32916;
  assign n32918 = pi17 ? n37 : n32917;
  assign n32919 = pi16 ? n32915 : n32918;
  assign n32920 = pi16 ? n31941 : n32918;
  assign n32921 = pi15 ? n32919 : n32920;
  assign n32922 = pi14 ? n32913 : n32921;
  assign n32923 = pi13 ? n32904 : n32922;
  assign n32924 = pi19 ? n30097 : n37;
  assign n32925 = pi18 ? n31315 : n32924;
  assign n32926 = pi17 ? n32 : n32925;
  assign n32927 = pi21 ? n25265 : n32;
  assign n32928 = pi20 ? n32927 : n32;
  assign n32929 = pi19 ? n8765 : n32928;
  assign n32930 = pi18 ? n37 : n32929;
  assign n32931 = pi17 ? n37 : n32930;
  assign n32932 = pi16 ? n32926 : n32931;
  assign n32933 = pi20 ? n31903 : n37;
  assign n32934 = pi19 ? n32933 : n37;
  assign n32935 = pi18 ? n31315 : n32934;
  assign n32936 = pi17 ? n32 : n32935;
  assign n32937 = pi19 ? n9769 : n32928;
  assign n32938 = pi18 ? n37 : n32937;
  assign n32939 = pi17 ? n37 : n32938;
  assign n32940 = pi16 ? n32936 : n32939;
  assign n32941 = pi15 ? n32932 : n32940;
  assign n32942 = pi21 ? n25276 : n32;
  assign n32943 = pi20 ? n32942 : n32;
  assign n32944 = pi19 ? n139 : n32943;
  assign n32945 = pi18 ? n37 : n32944;
  assign n32946 = pi17 ? n37 : n32945;
  assign n32947 = pi16 ? n32936 : n32946;
  assign n32948 = pi21 ? n31293 : n30843;
  assign n32949 = pi20 ? n32 : n32948;
  assign n32950 = pi19 ? n32 : n32949;
  assign n32951 = pi18 ? n32950 : n37;
  assign n32952 = pi17 ? n32 : n32951;
  assign n32953 = pi19 ? n32416 : n6383;
  assign n32954 = pi18 ? n37 : n32953;
  assign n32955 = pi17 ? n37 : n32954;
  assign n32956 = pi16 ? n32952 : n32955;
  assign n32957 = pi15 ? n32947 : n32956;
  assign n32958 = pi14 ? n32941 : n32957;
  assign n32959 = pi22 ? n705 : n32;
  assign n32960 = pi21 ? n32959 : n32;
  assign n32961 = pi20 ? n32960 : n32;
  assign n32962 = pi19 ? n10681 : n32961;
  assign n32963 = pi18 ? n37 : n32962;
  assign n32964 = pi17 ? n37 : n32963;
  assign n32965 = pi16 ? n32415 : n32964;
  assign n32966 = pi22 ? n30865 : n30195;
  assign n32967 = pi21 ? n32966 : n37;
  assign n32968 = pi20 ? n32 : n32967;
  assign n32969 = pi19 ? n32 : n32968;
  assign n32970 = pi18 ? n32969 : n37;
  assign n32971 = pi17 ? n32 : n32970;
  assign n32972 = pi20 ? n17591 : n32;
  assign n32973 = pi19 ? n12628 : n32972;
  assign n32974 = pi18 ? n37 : n32973;
  assign n32975 = pi17 ? n37 : n32974;
  assign n32976 = pi16 ? n32971 : n32975;
  assign n32977 = pi15 ? n32965 : n32976;
  assign n32978 = pi19 ? n37 : n5815;
  assign n32979 = pi18 ? n37 : n32978;
  assign n32980 = pi17 ? n37 : n32979;
  assign n32981 = pi16 ? n32971 : n32980;
  assign n32982 = pi19 ? n37 : n4111;
  assign n32983 = pi18 ? n37 : n32982;
  assign n32984 = pi17 ? n37 : n32983;
  assign n32985 = pi16 ? n439 : n32984;
  assign n32986 = pi15 ? n32981 : n32985;
  assign n32987 = pi14 ? n32977 : n32986;
  assign n32988 = pi13 ? n32958 : n32987;
  assign n32989 = pi12 ? n32923 : n32988;
  assign n32990 = pi23 ? n6960 : n687;
  assign n32991 = pi22 ? n32990 : n32;
  assign n32992 = pi21 ? n32991 : n32;
  assign n32993 = pi20 ? n32992 : n32;
  assign n32994 = pi19 ? n37 : n32993;
  assign n32995 = pi18 ? n37 : n32994;
  assign n32996 = pi17 ? n37 : n32995;
  assign n32997 = pi16 ? n439 : n32996;
  assign n32998 = pi19 ? n32453 : n3341;
  assign n32999 = pi18 ? n32452 : n32998;
  assign n33000 = pi17 ? n15070 : n32999;
  assign n33001 = pi16 ? n439 : n33000;
  assign n33002 = pi15 ? n32997 : n33001;
  assign n33003 = pi14 ? n33002 : n32469;
  assign n33004 = pi19 ? n6391 : n2580;
  assign n33005 = pi18 ? n37 : n33004;
  assign n33006 = pi17 ? n37 : n33005;
  assign n33007 = pi16 ? n439 : n33006;
  assign n33008 = pi15 ? n33007 : n32482;
  assign n33009 = pi14 ? n33008 : n32491;
  assign n33010 = pi13 ? n33003 : n33009;
  assign n33011 = pi19 ? n24494 : n2680;
  assign n33012 = pi18 ? n37 : n33011;
  assign n33013 = pi17 ? n37 : n33012;
  assign n33014 = pi16 ? n439 : n33013;
  assign n33015 = pi19 ? n6443 : n2680;
  assign n33016 = pi18 ? n37 : n33015;
  assign n33017 = pi17 ? n37 : n33016;
  assign n33018 = pi16 ? n439 : n33017;
  assign n33019 = pi15 ? n33014 : n33018;
  assign n33020 = pi14 ? n33019 : n32507;
  assign n33021 = pi21 ? n37 : n17764;
  assign n33022 = pi20 ? n37 : n33021;
  assign n33023 = pi19 ? n33022 : n1823;
  assign n33024 = pi18 ? n37 : n33023;
  assign n33025 = pi17 ? n37 : n33024;
  assign n33026 = pi16 ? n439 : n33025;
  assign n33027 = pi19 ? n2108 : n32;
  assign n33028 = pi18 ? n37 : n33027;
  assign n33029 = pi17 ? n37 : n33028;
  assign n33030 = pi16 ? n439 : n33029;
  assign n33031 = pi15 ? n33026 : n33030;
  assign n33032 = pi21 ? n37 : n20460;
  assign n33033 = pi20 ? n37 : n33032;
  assign n33034 = pi19 ? n33033 : n32;
  assign n33035 = pi18 ? n37 : n33034;
  assign n33036 = pi17 ? n37 : n33035;
  assign n33037 = pi16 ? n439 : n33036;
  assign n33038 = pi21 ? n272 : n20460;
  assign n33039 = pi20 ? n157 : n33038;
  assign n33040 = pi19 ? n33039 : n32;
  assign n33041 = pi18 ? n32535 : n33040;
  assign n33042 = pi17 ? n37 : n33041;
  assign n33043 = pi16 ? n439 : n33042;
  assign n33044 = pi15 ? n33037 : n33043;
  assign n33045 = pi14 ? n33031 : n33044;
  assign n33046 = pi13 ? n33020 : n33045;
  assign n33047 = pi12 ? n33010 : n33046;
  assign n33048 = pi11 ? n32989 : n33047;
  assign n33049 = pi19 ? n7839 : n32;
  assign n33050 = pi18 ? n32549 : n33049;
  assign n33051 = pi17 ? n32547 : n33050;
  assign n33052 = pi16 ? n439 : n33051;
  assign n33053 = pi19 ? n9035 : n32;
  assign n33054 = pi18 ? n32564 : n33053;
  assign n33055 = pi17 ? n32561 : n33054;
  assign n33056 = pi16 ? n32558 : n33055;
  assign n33057 = pi15 ? n33052 : n33056;
  assign n33058 = pi22 ? n157 : n2299;
  assign n33059 = pi21 ? n157 : n33058;
  assign n33060 = pi20 ? n157 : n33059;
  assign n33061 = pi19 ? n33060 : n32;
  assign n33062 = pi18 ? n32571 : n33061;
  assign n33063 = pi17 ? n99 : n33062;
  assign n33064 = pi16 ? n23698 : n33063;
  assign n33065 = pi20 ? n27598 : n6536;
  assign n33066 = pi19 ? n33065 : n32;
  assign n33067 = pi18 ? n32582 : n33066;
  assign n33068 = pi17 ? n99 : n33067;
  assign n33069 = pi16 ? n23698 : n33068;
  assign n33070 = pi15 ? n33064 : n33069;
  assign n33071 = pi14 ? n33057 : n33070;
  assign n33072 = pi21 ? n99 : n397;
  assign n33073 = pi20 ? n99 : n33072;
  assign n33074 = pi19 ? n33073 : n32;
  assign n33075 = pi18 ? n99 : n33074;
  assign n33076 = pi17 ? n99 : n33075;
  assign n33077 = pi16 ? n801 : n33076;
  assign n33078 = pi16 ? n201 : n33076;
  assign n33079 = pi15 ? n33077 : n33078;
  assign n33080 = pi18 ? n799 : n30468;
  assign n33081 = pi17 ? n32 : n33080;
  assign n33082 = pi19 ? n7914 : n32;
  assign n33083 = pi18 ? n30474 : n33082;
  assign n33084 = pi17 ? n139 : n33083;
  assign n33085 = pi16 ? n33081 : n33084;
  assign n33086 = pi19 ? n3033 : n23728;
  assign n33087 = pi18 ? n374 : n33086;
  assign n33088 = pi17 ? n32 : n33087;
  assign n33089 = pi18 ? n139 : n32601;
  assign n33090 = pi17 ? n139 : n33089;
  assign n33091 = pi16 ? n33088 : n33090;
  assign n33092 = pi15 ? n33085 : n33091;
  assign n33093 = pi14 ? n33079 : n33092;
  assign n33094 = pi13 ? n33071 : n33093;
  assign n33095 = pi22 ? n316 : n14363;
  assign n33096 = pi21 ? n316 : n33095;
  assign n33097 = pi20 ? n316 : n33096;
  assign n33098 = pi19 ? n33097 : n32;
  assign n33099 = pi18 ? n139 : n33098;
  assign n33100 = pi17 ? n139 : n33099;
  assign n33101 = pi16 ? n32621 : n33100;
  assign n33102 = pi15 ? n33101 : n32634;
  assign n33103 = pi20 ? n204 : n1050;
  assign n33104 = pi19 ? n32640 : n33103;
  assign n33105 = pi22 ? n21511 : n32;
  assign n33106 = pi21 ? n204 : n33105;
  assign n33107 = pi20 ? n1060 : n33106;
  assign n33108 = pi19 ? n33107 : n32;
  assign n33109 = pi18 ? n33104 : n33108;
  assign n33110 = pi17 ? n32638 : n33109;
  assign n33111 = pi16 ? n439 : n33110;
  assign n33112 = pi18 ? n204 : n25288;
  assign n33113 = pi17 ? n32649 : n33112;
  assign n33114 = pi16 ? n439 : n33113;
  assign n33115 = pi15 ? n33111 : n33114;
  assign n33116 = pi14 ? n33102 : n33115;
  assign n33117 = pi17 ? n32659 : n33112;
  assign n33118 = pi16 ? n32657 : n33117;
  assign n33119 = pi21 ? n204 : n3302;
  assign n33120 = pi20 ? n204 : n33119;
  assign n33121 = pi19 ? n33120 : n32;
  assign n33122 = pi18 ? n204 : n33121;
  assign n33123 = pi17 ? n32665 : n33122;
  assign n33124 = pi16 ? n439 : n33123;
  assign n33125 = pi15 ? n33118 : n33124;
  assign n33126 = pi21 ? n204 : n4109;
  assign n33127 = pi20 ? n204 : n33126;
  assign n33128 = pi19 ? n33127 : n32;
  assign n33129 = pi18 ? n32675 : n33128;
  assign n33130 = pi17 ? n32672 : n33129;
  assign n33131 = pi16 ? n439 : n33130;
  assign n33132 = pi21 ? n32692 : n6416;
  assign n33133 = pi20 ? n23069 : n33132;
  assign n33134 = pi19 ? n33133 : n32;
  assign n33135 = pi18 ? n32691 : n33134;
  assign n33136 = pi17 ? n32686 : n33135;
  assign n33137 = pi16 ? n32683 : n33136;
  assign n33138 = pi15 ? n33131 : n33137;
  assign n33139 = pi14 ? n33125 : n33138;
  assign n33140 = pi13 ? n33116 : n33139;
  assign n33141 = pi12 ? n33094 : n33140;
  assign n33142 = pi20 ? n233 : n22158;
  assign n33143 = pi19 ? n33142 : n32;
  assign n33144 = pi18 ? n32704 : n33143;
  assign n33145 = pi17 ? n15129 : n33144;
  assign n33146 = pi16 ? n439 : n33145;
  assign n33147 = pi21 ? n12659 : n882;
  assign n33148 = pi20 ? n15465 : n33147;
  assign n33149 = pi19 ? n33148 : n32;
  assign n33150 = pi18 ? n12631 : n33149;
  assign n33151 = pi17 ? n32712 : n33150;
  assign n33152 = pi16 ? n439 : n33151;
  assign n33153 = pi15 ? n33146 : n33152;
  assign n33154 = pi20 ? n15465 : n21565;
  assign n33155 = pi19 ? n33154 : n32;
  assign n33156 = pi18 ? n32726 : n33155;
  assign n33157 = pi17 ? n32725 : n33156;
  assign n33158 = pi16 ? n32722 : n33157;
  assign n33159 = pi23 ? n233 : n21112;
  assign n33160 = pi22 ? n233 : n33159;
  assign n33161 = pi21 ? n33160 : n32;
  assign n33162 = pi20 ? n233 : n33161;
  assign n33163 = pi19 ? n33162 : n32;
  assign n33164 = pi18 ? n2102 : n33163;
  assign n33165 = pi17 ? n32735 : n33164;
  assign n33166 = pi16 ? n25090 : n33165;
  assign n33167 = pi15 ? n33158 : n33166;
  assign n33168 = pi14 ? n33153 : n33167;
  assign n33169 = pi20 ? n233 : n10297;
  assign n33170 = pi19 ? n33169 : n32;
  assign n33171 = pi18 ? n2102 : n33170;
  assign n33172 = pi17 ? n32741 : n33171;
  assign n33173 = pi16 ? n439 : n33172;
  assign n33174 = pi22 ? n233 : n10784;
  assign n33175 = pi21 ? n33174 : n32;
  assign n33176 = pi20 ? n233 : n33175;
  assign n33177 = pi19 ? n33176 : n32;
  assign n33178 = pi18 ? n32748 : n33177;
  assign n33179 = pi17 ? n32746 : n33178;
  assign n33180 = pi16 ? n439 : n33179;
  assign n33181 = pi15 ? n33173 : n33180;
  assign n33182 = pi20 ? n233 : n19727;
  assign n33183 = pi19 ? n33182 : n32;
  assign n33184 = pi18 ? n32756 : n33183;
  assign n33185 = pi17 ? n32754 : n33184;
  assign n33186 = pi16 ? n439 : n33185;
  assign n33187 = pi20 ? n233 : n30006;
  assign n33188 = pi19 ? n33187 : n32;
  assign n33189 = pi18 ? n32764 : n33188;
  assign n33190 = pi17 ? n32762 : n33189;
  assign n33191 = pi16 ? n439 : n33190;
  assign n33192 = pi15 ? n33186 : n33191;
  assign n33193 = pi14 ? n33181 : n33192;
  assign n33194 = pi13 ? n33168 : n33193;
  assign n33195 = pi18 ? n233 : n33188;
  assign n33196 = pi17 ? n32773 : n33195;
  assign n33197 = pi16 ? n439 : n33196;
  assign n33198 = pi20 ? n685 : n9456;
  assign n33199 = pi19 ? n33198 : n32;
  assign n33200 = pi18 ? n2731 : n33199;
  assign n33201 = pi17 ? n37 : n33200;
  assign n33202 = pi16 ? n439 : n33201;
  assign n33203 = pi15 ? n33197 : n33202;
  assign n33204 = pi20 ? n18194 : n9963;
  assign n33205 = pi19 ? n33204 : n32;
  assign n33206 = pi18 ? n32795 : n33205;
  assign n33207 = pi17 ? n32792 : n33206;
  assign n33208 = pi16 ? n721 : n33207;
  assign n33209 = pi15 ? n33202 : n33208;
  assign n33210 = pi14 ? n33203 : n33209;
  assign n33211 = pi20 ? n32825 : n5667;
  assign n33212 = pi19 ? n33211 : n32;
  assign n33213 = pi18 ? n32824 : n33212;
  assign n33214 = pi17 ? n32821 : n33213;
  assign n33215 = pi16 ? n32812 : n33214;
  assign n33216 = pi23 ? n316 : n20004;
  assign n33217 = pi22 ? n33216 : n32;
  assign n33218 = pi21 ? n33217 : n32;
  assign n33219 = pi20 ? n32833 : n33218;
  assign n33220 = pi19 ? n33219 : n32;
  assign n33221 = pi18 ? n32832 : n33220;
  assign n33222 = pi17 ? n363 : n33221;
  assign n33223 = pi16 ? n26887 : n33222;
  assign n33224 = pi15 ? n33215 : n33223;
  assign n33225 = pi22 ? n26376 : n32;
  assign n33226 = pi21 ? n33225 : n32;
  assign n33227 = pi20 ? n32847 : n33226;
  assign n33228 = pi19 ? n33227 : n32;
  assign n33229 = pi18 ? n32832 : n33228;
  assign n33230 = pi17 ? n363 : n33229;
  assign n33231 = pi16 ? n29768 : n33230;
  assign n33232 = pi20 ? n32854 : n2701;
  assign n33233 = pi19 ? n33232 : n32;
  assign n33234 = pi18 ? n32832 : n33233;
  assign n33235 = pi17 ? n363 : n33234;
  assign n33236 = pi16 ? n29768 : n33235;
  assign n33237 = pi15 ? n33231 : n33236;
  assign n33238 = pi14 ? n33224 : n33237;
  assign n33239 = pi13 ? n33210 : n33238;
  assign n33240 = pi12 ? n33194 : n33239;
  assign n33241 = pi11 ? n33141 : n33240;
  assign n33242 = pi10 ? n33048 : n33241;
  assign n33243 = pi09 ? n32886 : n33242;
  assign n33244 = pi08 ? n32866 : n33243;
  assign n33245 = pi19 ? n20563 : n32898;
  assign n33246 = pi18 ? n30119 : n33245;
  assign n33247 = pi17 ? n32 : n33246;
  assign n33248 = pi20 ? n14844 : n219;
  assign n33249 = pi19 ? n33248 : n5121;
  assign n33250 = pi18 ? n37 : n33249;
  assign n33251 = pi19 ? n99 : n4567;
  assign n33252 = pi18 ? n99 : n33251;
  assign n33253 = pi17 ? n33250 : n33252;
  assign n33254 = pi16 ? n33247 : n33253;
  assign n33255 = pi15 ? n32 : n33254;
  assign n33256 = pi19 ? n99 : n4577;
  assign n33257 = pi18 ? n99 : n33256;
  assign n33258 = pi17 ? n32291 : n33257;
  assign n33259 = pi16 ? n33247 : n33258;
  assign n33260 = pi19 ? n20563 : n31267;
  assign n33261 = pi18 ? n30119 : n33260;
  assign n33262 = pi17 ? n32 : n33261;
  assign n33263 = pi19 ? n26407 : n3050;
  assign n33264 = pi18 ? n37 : n33263;
  assign n33265 = pi17 ? n33264 : n33257;
  assign n33266 = pi16 ? n33262 : n33265;
  assign n33267 = pi15 ? n33259 : n33266;
  assign n33268 = pi14 ? n33255 : n33267;
  assign n33269 = pi13 ? n32 : n33268;
  assign n33270 = pi12 ? n32 : n33269;
  assign n33271 = pi11 ? n32 : n33270;
  assign n33272 = pi10 ? n32 : n33271;
  assign n33273 = pi18 ? n31265 : n32872;
  assign n33274 = pi17 ? n32 : n33273;
  assign n33275 = pi20 ? n37 : n7747;
  assign n33276 = pi19 ? n33275 : n27249;
  assign n33277 = pi18 ? n37 : n33276;
  assign n33278 = pi22 ? n745 : n587;
  assign n33279 = pi21 ? n33278 : n32;
  assign n33280 = pi20 ? n33279 : n32;
  assign n33281 = pi19 ? n99 : n33280;
  assign n33282 = pi18 ? n99 : n33281;
  assign n33283 = pi17 ? n33277 : n33282;
  assign n33284 = pi16 ? n33274 : n33283;
  assign n33285 = pi19 ? n20563 : n30097;
  assign n33286 = pi18 ? n31265 : n33285;
  assign n33287 = pi17 ? n32 : n33286;
  assign n33288 = pi20 ? n37 : n221;
  assign n33289 = pi19 ? n33288 : n18853;
  assign n33290 = pi18 ? n37 : n33289;
  assign n33291 = pi22 ? n1656 : n587;
  assign n33292 = pi21 ? n33291 : n32;
  assign n33293 = pi20 ? n33292 : n32;
  assign n33294 = pi19 ? n99 : n33293;
  assign n33295 = pi18 ? n99 : n33294;
  assign n33296 = pi17 ? n33290 : n33295;
  assign n33297 = pi16 ? n33287 : n33296;
  assign n33298 = pi15 ? n33284 : n33297;
  assign n33299 = pi19 ? n20563 : n37;
  assign n33300 = pi18 ? n31265 : n33299;
  assign n33301 = pi17 ? n32 : n33300;
  assign n33302 = pi20 ? n5077 : n14887;
  assign n33303 = pi19 ? n33302 : n11415;
  assign n33304 = pi18 ? n37 : n33303;
  assign n33305 = pi19 ? n3050 : n22400;
  assign n33306 = pi21 ? n11435 : n32;
  assign n33307 = pi20 ? n33306 : n32;
  assign n33308 = pi19 ? n99 : n33307;
  assign n33309 = pi18 ? n33305 : n33308;
  assign n33310 = pi17 ? n33304 : n33309;
  assign n33311 = pi16 ? n33301 : n33310;
  assign n33312 = pi18 ? n31315 : n32295;
  assign n33313 = pi17 ? n32 : n33312;
  assign n33314 = pi21 ? n181 : n3668;
  assign n33315 = pi20 ? n33314 : n37;
  assign n33316 = pi19 ? n29138 : n33315;
  assign n33317 = pi20 ? n14524 : n11743;
  assign n33318 = pi19 ? n33317 : n32343;
  assign n33319 = pi18 ? n33316 : n33318;
  assign n33320 = pi17 ? n37 : n33319;
  assign n33321 = pi16 ? n33313 : n33320;
  assign n33322 = pi15 ? n33311 : n33321;
  assign n33323 = pi14 ? n33298 : n33322;
  assign n33324 = pi22 ? n893 : n32;
  assign n33325 = pi21 ? n33324 : n32;
  assign n33326 = pi20 ? n33325 : n32;
  assign n33327 = pi19 ? n37 : n33326;
  assign n33328 = pi18 ? n37 : n33327;
  assign n33329 = pi17 ? n37 : n33328;
  assign n33330 = pi16 ? n33313 : n33329;
  assign n33331 = pi18 ? n31938 : n32899;
  assign n33332 = pi17 ? n32 : n33331;
  assign n33333 = pi19 ? n37 : n3972;
  assign n33334 = pi18 ? n37 : n33333;
  assign n33335 = pi17 ? n37 : n33334;
  assign n33336 = pi16 ? n33332 : n33335;
  assign n33337 = pi15 ? n33330 : n33336;
  assign n33338 = pi23 ? n37 : n16890;
  assign n33339 = pi22 ? n33338 : n32;
  assign n33340 = pi21 ? n33339 : n32;
  assign n33341 = pi20 ? n33340 : n32;
  assign n33342 = pi19 ? n8765 : n33341;
  assign n33343 = pi18 ? n37 : n33342;
  assign n33344 = pi17 ? n37 : n33343;
  assign n33345 = pi16 ? n32901 : n33344;
  assign n33346 = pi14 ? n33337 : n33345;
  assign n33347 = pi13 ? n33323 : n33346;
  assign n33348 = pi19 ? n9814 : n37;
  assign n33349 = pi21 ? n25654 : n32;
  assign n33350 = pi20 ? n33349 : n32;
  assign n33351 = pi19 ? n8765 : n33350;
  assign n33352 = pi18 ? n33348 : n33351;
  assign n33353 = pi17 ? n37 : n33352;
  assign n33354 = pi16 ? n32351 : n33353;
  assign n33355 = pi23 ? n139 : n1748;
  assign n33356 = pi22 ? n33355 : n32;
  assign n33357 = pi21 ? n33356 : n32;
  assign n33358 = pi20 ? n33357 : n32;
  assign n33359 = pi19 ? n9769 : n33358;
  assign n33360 = pi18 ? n19855 : n33359;
  assign n33361 = pi17 ? n37 : n33360;
  assign n33362 = pi16 ? n32351 : n33361;
  assign n33363 = pi15 ? n33354 : n33362;
  assign n33364 = pi19 ? n37 : n3075;
  assign n33365 = pi18 ? n37 : n33364;
  assign n33366 = pi20 ? n3084 : n3083;
  assign n33367 = pi20 ? n12010 : n3086;
  assign n33368 = pi19 ? n33366 : n33367;
  assign n33369 = pi19 ? n139 : n33358;
  assign n33370 = pi18 ? n33368 : n33369;
  assign n33371 = pi17 ? n33365 : n33370;
  assign n33372 = pi16 ? n32379 : n33371;
  assign n33373 = pi18 ? n31938 : n32924;
  assign n33374 = pi17 ? n32 : n33373;
  assign n33375 = pi21 ? n37 : n9119;
  assign n33376 = pi21 ? n9143 : n335;
  assign n33377 = pi20 ? n33375 : n33376;
  assign n33378 = pi22 ? n1992 : n32;
  assign n33379 = pi21 ? n33378 : n32;
  assign n33380 = pi20 ? n33379 : n32;
  assign n33381 = pi19 ? n33377 : n33380;
  assign n33382 = pi18 ? n37 : n33381;
  assign n33383 = pi17 ? n37 : n33382;
  assign n33384 = pi16 ? n33374 : n33383;
  assign n33385 = pi15 ? n33372 : n33384;
  assign n33386 = pi14 ? n33363 : n33385;
  assign n33387 = pi18 ? n31938 : n32934;
  assign n33388 = pi17 ? n32 : n33387;
  assign n33389 = pi23 ? n335 : n10750;
  assign n33390 = pi22 ? n33389 : n32;
  assign n33391 = pi21 ? n33390 : n32;
  assign n33392 = pi20 ? n33391 : n32;
  assign n33393 = pi19 ? n10681 : n33392;
  assign n33394 = pi18 ? n37 : n33393;
  assign n33395 = pi17 ? n37 : n33394;
  assign n33396 = pi16 ? n33388 : n33395;
  assign n33397 = pi22 ? n1159 : n32;
  assign n33398 = pi21 ? n33397 : n32;
  assign n33399 = pi20 ? n33398 : n32;
  assign n33400 = pi19 ? n12628 : n33399;
  assign n33401 = pi18 ? n37 : n33400;
  assign n33402 = pi17 ? n37 : n33401;
  assign n33403 = pi16 ? n32936 : n33402;
  assign n33404 = pi15 ? n33396 : n33403;
  assign n33405 = pi21 ? n30866 : n29133;
  assign n33406 = pi20 ? n32 : n33405;
  assign n33407 = pi19 ? n32 : n33406;
  assign n33408 = pi18 ? n33407 : n37;
  assign n33409 = pi17 ? n32 : n33408;
  assign n33410 = pi21 ? n28467 : n32;
  assign n33411 = pi20 ? n33410 : n32;
  assign n33412 = pi19 ? n37 : n33411;
  assign n33413 = pi18 ? n37 : n33412;
  assign n33414 = pi17 ? n37 : n33413;
  assign n33415 = pi16 ? n33409 : n33414;
  assign n33416 = pi21 ? n11057 : n32;
  assign n33417 = pi20 ? n33416 : n32;
  assign n33418 = pi19 ? n37 : n33417;
  assign n33419 = pi18 ? n37 : n33418;
  assign n33420 = pi17 ? n37 : n33419;
  assign n33421 = pi16 ? n32432 : n33420;
  assign n33422 = pi15 ? n33415 : n33421;
  assign n33423 = pi14 ? n33404 : n33422;
  assign n33424 = pi13 ? n33386 : n33423;
  assign n33425 = pi12 ? n33347 : n33424;
  assign n33426 = pi19 ? n12478 : n4111;
  assign n33427 = pi18 ? n37 : n33426;
  assign n33428 = pi17 ? n37 : n33427;
  assign n33429 = pi16 ? n439 : n33428;
  assign n33430 = pi21 ? n2091 : n6361;
  assign n33431 = pi20 ? n571 : n33430;
  assign n33432 = pi19 ? n33431 : n4111;
  assign n33433 = pi18 ? n37 : n33432;
  assign n33434 = pi17 ? n37 : n33433;
  assign n33435 = pi16 ? n439 : n33434;
  assign n33436 = pi15 ? n33429 : n33435;
  assign n33437 = pi19 ? n32459 : n4111;
  assign n33438 = pi18 ? n37 : n33437;
  assign n33439 = pi17 ? n37 : n33438;
  assign n33440 = pi16 ? n439 : n33439;
  assign n33441 = pi20 ? n21148 : n335;
  assign n33442 = pi22 ? n21744 : n32;
  assign n33443 = pi21 ? n33442 : n32;
  assign n33444 = pi20 ? n33443 : n32;
  assign n33445 = pi19 ? n33441 : n33444;
  assign n33446 = pi18 ? n37 : n33445;
  assign n33447 = pi17 ? n37 : n33446;
  assign n33448 = pi16 ? n439 : n33447;
  assign n33449 = pi15 ? n33440 : n33448;
  assign n33450 = pi14 ? n33436 : n33449;
  assign n33451 = pi19 ? n6391 : n6418;
  assign n33452 = pi18 ? n37 : n33451;
  assign n33453 = pi17 ? n37 : n33452;
  assign n33454 = pi16 ? n439 : n33453;
  assign n33455 = pi19 ? n32478 : n4117;
  assign n33456 = pi18 ? n37 : n33455;
  assign n33457 = pi17 ? n37 : n33456;
  assign n33458 = pi16 ? n439 : n33457;
  assign n33459 = pi15 ? n33454 : n33458;
  assign n33460 = pi19 ? n6403 : n5831;
  assign n33461 = pi18 ? n37 : n33460;
  assign n33462 = pi17 ? n37 : n33461;
  assign n33463 = pi16 ? n439 : n33462;
  assign n33464 = pi14 ? n33459 : n33463;
  assign n33465 = pi13 ? n33450 : n33464;
  assign n33466 = pi21 ? n37 : n21653;
  assign n33467 = pi20 ? n37 : n33466;
  assign n33468 = pi19 ? n33467 : n2639;
  assign n33469 = pi18 ? n37 : n33468;
  assign n33470 = pi17 ? n37 : n33469;
  assign n33471 = pi16 ? n439 : n33470;
  assign n33472 = pi19 ? n5029 : n2639;
  assign n33473 = pi18 ? n37 : n33472;
  assign n33474 = pi17 ? n37 : n33473;
  assign n33475 = pi16 ? n439 : n33474;
  assign n33476 = pi15 ? n33471 : n33475;
  assign n33477 = pi19 ? n2108 : n2639;
  assign n33478 = pi18 ? n37 : n33477;
  assign n33479 = pi17 ? n37 : n33478;
  assign n33480 = pi16 ? n439 : n33479;
  assign n33481 = pi19 ? n2108 : n2654;
  assign n33482 = pi18 ? n37 : n33481;
  assign n33483 = pi17 ? n37 : n33482;
  assign n33484 = pi16 ? n439 : n33483;
  assign n33485 = pi15 ? n33480 : n33484;
  assign n33486 = pi14 ? n33476 : n33485;
  assign n33487 = pi19 ? n33022 : n2654;
  assign n33488 = pi18 ? n37 : n33487;
  assign n33489 = pi17 ? n37 : n33488;
  assign n33490 = pi16 ? n439 : n33489;
  assign n33491 = pi15 ? n33490 : n33030;
  assign n33492 = pi20 ? n37 : n2974;
  assign n33493 = pi19 ? n37 : n33492;
  assign n33494 = pi20 ? n2974 : n6500;
  assign n33495 = pi19 ? n33492 : n33494;
  assign n33496 = pi18 ? n33493 : n33495;
  assign n33497 = pi21 ? n244 : n777;
  assign n33498 = pi21 ? n2175 : n777;
  assign n33499 = pi20 ? n33497 : n33498;
  assign n33500 = pi20 ? n2176 : n273;
  assign n33501 = pi19 ? n33499 : n33500;
  assign n33502 = pi18 ? n33501 : n33049;
  assign n33503 = pi17 ? n33496 : n33502;
  assign n33504 = pi16 ? n439 : n33503;
  assign n33505 = pi15 ? n33037 : n33504;
  assign n33506 = pi14 ? n33491 : n33505;
  assign n33507 = pi13 ? n33486 : n33506;
  assign n33508 = pi12 ? n33465 : n33507;
  assign n33509 = pi11 ? n33425 : n33508;
  assign n33510 = pi20 ? n15263 : n2238;
  assign n33511 = pi19 ? n33510 : n11445;
  assign n33512 = pi18 ? n33511 : n33049;
  assign n33513 = pi17 ? n32547 : n33512;
  assign n33514 = pi16 ? n439 : n33513;
  assign n33515 = pi19 ? n99 : n6542;
  assign n33516 = pi18 ? n30851 : n33515;
  assign n33517 = pi21 ? n777 : n2981;
  assign n33518 = pi20 ? n33517 : n99;
  assign n33519 = pi19 ? n33518 : n19134;
  assign n33520 = pi18 ? n33519 : n33053;
  assign n33521 = pi17 ? n33516 : n33520;
  assign n33522 = pi16 ? n439 : n33521;
  assign n33523 = pi15 ? n33514 : n33522;
  assign n33524 = pi18 ? n99 : n33053;
  assign n33525 = pi17 ? n99 : n33524;
  assign n33526 = pi16 ? n23698 : n33525;
  assign n33527 = pi22 ? n157 : n1263;
  assign n33528 = pi21 ? n777 : n33527;
  assign n33529 = pi20 ? n20977 : n33528;
  assign n33530 = pi19 ? n33529 : n32;
  assign n33531 = pi18 ? n99 : n33530;
  assign n33532 = pi17 ? n99 : n33531;
  assign n33533 = pi16 ? n23698 : n33532;
  assign n33534 = pi15 ? n33526 : n33533;
  assign n33535 = pi14 ? n33523 : n33534;
  assign n33536 = pi21 ? n777 : n7137;
  assign n33537 = pi20 ? n2238 : n33536;
  assign n33538 = pi19 ? n33537 : n32;
  assign n33539 = pi18 ? n99 : n33538;
  assign n33540 = pi17 ? n99 : n33539;
  assign n33541 = pi16 ? n744 : n33540;
  assign n33542 = pi21 ? n99 : n10318;
  assign n33543 = pi20 ? n99 : n33542;
  assign n33544 = pi19 ? n33543 : n32;
  assign n33545 = pi18 ? n99 : n33544;
  assign n33546 = pi17 ? n99 : n33545;
  assign n33547 = pi16 ? n744 : n33546;
  assign n33548 = pi15 ? n33541 : n33547;
  assign n33549 = pi21 ? n22940 : n99;
  assign n33550 = pi20 ? n139 : n33549;
  assign n33551 = pi19 ? n139 : n33550;
  assign n33552 = pi18 ? n33551 : n33082;
  assign n33553 = pi17 ? n139 : n33552;
  assign n33554 = pi16 ? n30470 : n33553;
  assign n33555 = pi18 ? n374 : n28256;
  assign n33556 = pi17 ? n32 : n33555;
  assign n33557 = pi20 ? n139 : n4767;
  assign n33558 = pi19 ? n139 : n33557;
  assign n33559 = pi18 ? n33558 : n32601;
  assign n33560 = pi17 ? n139 : n33559;
  assign n33561 = pi16 ? n33556 : n33560;
  assign n33562 = pi15 ? n33554 : n33561;
  assign n33563 = pi14 ? n33548 : n33562;
  assign n33564 = pi13 ? n33535 : n33563;
  assign n33565 = pi21 ? n349 : n346;
  assign n33566 = pi20 ? n139 : n33565;
  assign n33567 = pi19 ? n139 : n33566;
  assign n33568 = pi18 ? n9770 : n33567;
  assign n33569 = pi19 ? n3168 : n33557;
  assign n33570 = pi18 ? n33569 : n32119;
  assign n33571 = pi17 ? n33568 : n33570;
  assign n33572 = pi16 ? n439 : n33571;
  assign n33573 = pi21 ? n916 : n4451;
  assign n33574 = pi20 ? n941 : n33573;
  assign n33575 = pi19 ? n139 : n33574;
  assign n33576 = pi18 ? n8766 : n33575;
  assign n33577 = pi21 ? n139 : n4445;
  assign n33578 = pi20 ? n33577 : n139;
  assign n33579 = pi20 ? n139 : n1056;
  assign n33580 = pi19 ? n33578 : n33579;
  assign n33581 = pi18 ? n33580 : n32119;
  assign n33582 = pi17 ? n33576 : n33581;
  assign n33583 = pi16 ? n439 : n33582;
  assign n33584 = pi15 ? n33572 : n33583;
  assign n33585 = pi20 ? n204 : n5926;
  assign n33586 = pi19 ? n13494 : n33585;
  assign n33587 = pi21 ? n204 : n4094;
  assign n33588 = pi20 ? n204 : n33587;
  assign n33589 = pi19 ? n33588 : n32;
  assign n33590 = pi18 ? n33586 : n33589;
  assign n33591 = pi17 ? n32638 : n33590;
  assign n33592 = pi16 ? n439 : n33591;
  assign n33593 = pi18 ? n18985 : n204;
  assign n33594 = pi19 ? n7970 : n32;
  assign n33595 = pi18 ? n204 : n33594;
  assign n33596 = pi17 ? n33593 : n33595;
  assign n33597 = pi16 ? n439 : n33596;
  assign n33598 = pi15 ? n33592 : n33597;
  assign n33599 = pi14 ? n33584 : n33598;
  assign n33600 = pi20 ? n31625 : n204;
  assign n33601 = pi19 ? n33600 : n204;
  assign n33602 = pi18 ? n33601 : n204;
  assign n33603 = pi17 ? n33602 : n33595;
  assign n33604 = pi16 ? n32657 : n33603;
  assign n33605 = pi23 ? n204 : n32126;
  assign n33606 = pi22 ? n33605 : n32;
  assign n33607 = pi21 ? n204 : n33606;
  assign n33608 = pi20 ? n204 : n33607;
  assign n33609 = pi19 ? n33608 : n32;
  assign n33610 = pi18 ? n204 : n33609;
  assign n33611 = pi17 ? n32665 : n33610;
  assign n33612 = pi16 ? n439 : n33611;
  assign n33613 = pi15 ? n33604 : n33612;
  assign n33614 = pi18 ? n19359 : n233;
  assign n33615 = pi20 ? n3104 : n233;
  assign n33616 = pi19 ? n33615 : n32674;
  assign n33617 = pi18 ? n33616 : n33128;
  assign n33618 = pi17 ? n33614 : n33617;
  assign n33619 = pi16 ? n439 : n33618;
  assign n33620 = pi20 ? n642 : n233;
  assign n33621 = pi19 ? n33620 : n18446;
  assign n33622 = pi22 ? n10784 : n32;
  assign n33623 = pi21 ? n233 : n33622;
  assign n33624 = pi20 ? n233 : n33623;
  assign n33625 = pi19 ? n33624 : n32;
  assign n33626 = pi18 ? n33621 : n33625;
  assign n33627 = pi17 ? n33614 : n33626;
  assign n33628 = pi16 ? n439 : n33627;
  assign n33629 = pi15 ? n33619 : n33628;
  assign n33630 = pi14 ? n33613 : n33629;
  assign n33631 = pi13 ? n33599 : n33630;
  assign n33632 = pi12 ? n33564 : n33631;
  assign n33633 = pi19 ? n37 : n27727;
  assign n33634 = pi18 ? n37 : n33633;
  assign n33635 = pi21 ? n233 : n760;
  assign n33636 = pi20 ? n233 : n33635;
  assign n33637 = pi19 ? n33636 : n32;
  assign n33638 = pi18 ? n32704 : n33637;
  assign n33639 = pi17 ? n33634 : n33638;
  assign n33640 = pi16 ? n439 : n33639;
  assign n33641 = pi21 ? n9398 : n882;
  assign n33642 = pi20 ? n233 : n33641;
  assign n33643 = pi19 ? n33642 : n32;
  assign n33644 = pi18 ? n335 : n33643;
  assign n33645 = pi17 ? n32712 : n33644;
  assign n33646 = pi16 ? n439 : n33645;
  assign n33647 = pi15 ? n33640 : n33646;
  assign n33648 = pi20 ? n649 : n647;
  assign n33649 = pi19 ? n37 : n33648;
  assign n33650 = pi18 ? n374 : n33649;
  assign n33651 = pi17 ? n32 : n33650;
  assign n33652 = pi21 ? n9405 : n928;
  assign n33653 = pi20 ? n233 : n33652;
  assign n33654 = pi19 ? n33653 : n32;
  assign n33655 = pi18 ? n17205 : n33654;
  assign n33656 = pi17 ? n32725 : n33655;
  assign n33657 = pi16 ? n33651 : n33656;
  assign n33658 = pi21 ? n12994 : n32;
  assign n33659 = pi20 ? n233 : n33658;
  assign n33660 = pi19 ? n33659 : n32;
  assign n33661 = pi18 ? n7677 : n33660;
  assign n33662 = pi17 ? n32735 : n33661;
  assign n33663 = pi16 ? n25090 : n33662;
  assign n33664 = pi15 ? n33657 : n33663;
  assign n33665 = pi14 ? n33647 : n33664;
  assign n33666 = pi20 ? n4971 : n37;
  assign n33667 = pi19 ? n37 : n33666;
  assign n33668 = pi18 ? n374 : n33667;
  assign n33669 = pi17 ? n32 : n33668;
  assign n33670 = pi16 ? n33669 : n33172;
  assign n33671 = pi20 ? n647 : n7980;
  assign n33672 = pi19 ? n10957 : n33671;
  assign n33673 = pi18 ? n33672 : n233;
  assign n33674 = pi20 ? n6358 : n4921;
  assign n33675 = pi19 ? n33674 : n233;
  assign n33676 = pi18 ? n33675 : n33170;
  assign n33677 = pi17 ? n33673 : n33676;
  assign n33678 = pi16 ? n439 : n33677;
  assign n33679 = pi15 ? n33670 : n33678;
  assign n33680 = pi19 ? n37 : n10272;
  assign n33681 = pi18 ? n374 : n33680;
  assign n33682 = pi17 ? n32 : n33681;
  assign n33683 = pi20 ? n575 : n610;
  assign n33684 = pi21 ? n335 : n4900;
  assign n33685 = pi20 ? n33684 : n233;
  assign n33686 = pi19 ? n33683 : n33685;
  assign n33687 = pi18 ? n33686 : n233;
  assign n33688 = pi21 ? n19386 : n233;
  assign n33689 = pi20 ? n7980 : n33688;
  assign n33690 = pi19 ? n33689 : n233;
  assign n33691 = pi18 ? n33690 : n33170;
  assign n33692 = pi17 ? n33687 : n33691;
  assign n33693 = pi16 ? n33682 : n33692;
  assign n33694 = pi20 ? n37 : n9912;
  assign n33695 = pi21 ? n37 : n15143;
  assign n33696 = pi20 ? n33695 : n233;
  assign n33697 = pi19 ? n33694 : n33696;
  assign n33698 = pi18 ? n33697 : n233;
  assign n33699 = pi20 ? n2092 : n4921;
  assign n33700 = pi19 ? n33699 : n233;
  assign n33701 = pi18 ? n33700 : n33170;
  assign n33702 = pi17 ? n33698 : n33701;
  assign n33703 = pi16 ? n439 : n33702;
  assign n33704 = pi15 ? n33693 : n33703;
  assign n33705 = pi14 ? n33679 : n33704;
  assign n33706 = pi13 ? n33665 : n33705;
  assign n33707 = pi18 ? n374 : n3407;
  assign n33708 = pi17 ? n32 : n33707;
  assign n33709 = pi18 ? n233 : n33177;
  assign n33710 = pi17 ? n32773 : n33709;
  assign n33711 = pi16 ? n33708 : n33710;
  assign n33712 = pi20 ? n37 : n23929;
  assign n33713 = pi19 ? n37 : n33712;
  assign n33714 = pi18 ? n37 : n33713;
  assign n33715 = pi20 ? n685 : n11695;
  assign n33716 = pi19 ? n33715 : n32;
  assign n33717 = pi18 ? n2731 : n33716;
  assign n33718 = pi17 ? n33714 : n33717;
  assign n33719 = pi16 ? n439 : n33718;
  assign n33720 = pi15 ? n33711 : n33719;
  assign n33721 = pi22 ? n685 : n2834;
  assign n33722 = pi21 ? n33721 : n32;
  assign n33723 = pi20 ? n685 : n33722;
  assign n33724 = pi19 ? n33723 : n32;
  assign n33725 = pi18 ? n2731 : n33724;
  assign n33726 = pi17 ? n37 : n33725;
  assign n33727 = pi16 ? n439 : n33726;
  assign n33728 = pi19 ? n99 : n4557;
  assign n33729 = pi18 ? n719 : n33728;
  assign n33730 = pi17 ? n32 : n33729;
  assign n33731 = pi20 ? n30778 : n722;
  assign n33732 = pi20 ? n32787 : n23162;
  assign n33733 = pi19 ? n33731 : n33732;
  assign n33734 = pi19 ? n28732 : n363;
  assign n33735 = pi18 ? n33733 : n33734;
  assign n33736 = pi21 ? n4551 : n363;
  assign n33737 = pi20 ? n33736 : n29686;
  assign n33738 = pi21 ? n363 : n14255;
  assign n33739 = pi20 ? n363 : n33738;
  assign n33740 = pi19 ? n33737 : n33739;
  assign n33741 = pi20 ? n685 : n10326;
  assign n33742 = pi19 ? n33741 : n32;
  assign n33743 = pi18 ? n33740 : n33742;
  assign n33744 = pi17 ? n33735 : n33743;
  assign n33745 = pi16 ? n33730 : n33744;
  assign n33746 = pi15 ? n33727 : n33745;
  assign n33747 = pi14 ? n33720 : n33746;
  assign n33748 = pi21 ? n823 : n29838;
  assign n33749 = pi22 ? n812 : n363;
  assign n33750 = pi21 ? n4252 : n33749;
  assign n33751 = pi20 ? n33748 : n33750;
  assign n33752 = pi19 ? n139 : n33751;
  assign n33753 = pi18 ? n23990 : n33752;
  assign n33754 = pi17 ? n32 : n33753;
  assign n33755 = pi22 ? n139 : n4543;
  assign n33756 = pi21 ? n33755 : n4234;
  assign n33757 = pi22 ? n745 : n4543;
  assign n33758 = pi22 ? n363 : n4537;
  assign n33759 = pi21 ? n33757 : n33758;
  assign n33760 = pi20 ? n33756 : n33759;
  assign n33761 = pi22 ? n812 : n4543;
  assign n33762 = pi21 ? n33761 : n33758;
  assign n33763 = pi21 ? n22557 : n33757;
  assign n33764 = pi20 ? n33762 : n33763;
  assign n33765 = pi19 ? n33760 : n33764;
  assign n33766 = pi21 ? n20228 : n823;
  assign n33767 = pi22 ? n745 : n363;
  assign n33768 = pi21 ? n20228 : n33767;
  assign n33769 = pi22 ? n363 : n745;
  assign n33770 = pi21 ? n33769 : n363;
  assign n33771 = pi20 ? n33768 : n33770;
  assign n33772 = pi19 ? n33766 : n33771;
  assign n33773 = pi18 ? n33765 : n33772;
  assign n33774 = pi21 ? n33755 : n33749;
  assign n33775 = pi21 ? n363 : n33769;
  assign n33776 = pi20 ? n33774 : n33775;
  assign n33777 = pi21 ? n33767 : n363;
  assign n33778 = pi20 ? n33777 : n33738;
  assign n33779 = pi19 ? n33776 : n33778;
  assign n33780 = pi21 ? n685 : n24222;
  assign n33781 = pi20 ? n33780 : n6935;
  assign n33782 = pi19 ? n33781 : n32;
  assign n33783 = pi18 ? n33779 : n33782;
  assign n33784 = pi17 ? n33773 : n33783;
  assign n33785 = pi16 ? n33754 : n33784;
  assign n33786 = pi20 ? n26898 : n3210;
  assign n33787 = pi19 ? n33786 : n32;
  assign n33788 = pi18 ? n32832 : n33787;
  assign n33789 = pi17 ? n363 : n33788;
  assign n33790 = pi16 ? n21219 : n33789;
  assign n33791 = pi15 ? n33785 : n33790;
  assign n33792 = pi25 ? n138 : n32;
  assign n33793 = pi24 ? n32 : n33792;
  assign n33794 = pi23 ? n33793 : n363;
  assign n33795 = pi22 ? n33794 : n363;
  assign n33796 = pi21 ? n33795 : n363;
  assign n33797 = pi20 ? n32 : n33796;
  assign n33798 = pi19 ? n32 : n33797;
  assign n33799 = pi18 ? n33798 : n363;
  assign n33800 = pi17 ? n32 : n33799;
  assign n33801 = pi23 ? n2766 : n14362;
  assign n33802 = pi22 ? n33801 : n32;
  assign n33803 = pi21 ? n33802 : n32;
  assign n33804 = pi20 ? n26890 : n33803;
  assign n33805 = pi19 ? n33804 : n32;
  assign n33806 = pi18 ? n32832 : n33805;
  assign n33807 = pi17 ? n363 : n33806;
  assign n33808 = pi16 ? n33800 : n33807;
  assign n33809 = pi20 ? n685 : n2701;
  assign n33810 = pi19 ? n33809 : n32;
  assign n33811 = pi18 ? n32832 : n33810;
  assign n33812 = pi17 ? n363 : n33811;
  assign n33813 = pi16 ? n26062 : n33812;
  assign n33814 = pi15 ? n33808 : n33813;
  assign n33815 = pi14 ? n33791 : n33814;
  assign n33816 = pi13 ? n33747 : n33815;
  assign n33817 = pi12 ? n33706 : n33816;
  assign n33818 = pi11 ? n33632 : n33817;
  assign n33819 = pi10 ? n33509 : n33818;
  assign n33820 = pi09 ? n33272 : n33819;
  assign n33821 = pi21 ? n31924 : n37;
  assign n33822 = pi20 ? n20563 : n33821;
  assign n33823 = pi19 ? n20563 : n33822;
  assign n33824 = pi18 ? n30119 : n33823;
  assign n33825 = pi17 ? n32 : n33824;
  assign n33826 = pi16 ? n33825 : n33253;
  assign n33827 = pi15 ? n32 : n33826;
  assign n33828 = pi19 ? n20563 : n31904;
  assign n33829 = pi18 ? n30119 : n33828;
  assign n33830 = pi17 ? n32 : n33829;
  assign n33831 = pi16 ? n33830 : n33265;
  assign n33832 = pi15 ? n33259 : n33831;
  assign n33833 = pi14 ? n33827 : n33832;
  assign n33834 = pi13 ? n32 : n33833;
  assign n33835 = pi12 ? n32 : n33834;
  assign n33836 = pi11 ? n32 : n33835;
  assign n33837 = pi10 ? n32 : n33836;
  assign n33838 = pi22 ? n3492 : n587;
  assign n33839 = pi21 ? n33838 : n32;
  assign n33840 = pi20 ? n33839 : n32;
  assign n33841 = pi19 ? n99 : n33840;
  assign n33842 = pi18 ? n99 : n33841;
  assign n33843 = pi17 ? n33277 : n33842;
  assign n33844 = pi16 ? n33274 : n33843;
  assign n33845 = pi21 ? n31924 : n30843;
  assign n33846 = pi20 ? n33845 : n37;
  assign n33847 = pi19 ? n20563 : n33846;
  assign n33848 = pi18 ? n31265 : n33847;
  assign n33849 = pi17 ? n32 : n33848;
  assign n33850 = pi22 ? n11963 : n587;
  assign n33851 = pi21 ? n33850 : n32;
  assign n33852 = pi20 ? n33851 : n32;
  assign n33853 = pi19 ? n99 : n33852;
  assign n33854 = pi18 ? n99 : n33853;
  assign n33855 = pi17 ? n33290 : n33854;
  assign n33856 = pi16 ? n33849 : n33855;
  assign n33857 = pi15 ? n33844 : n33856;
  assign n33858 = pi19 ? n20563 : n31299;
  assign n33859 = pi18 ? n31265 : n33858;
  assign n33860 = pi17 ? n32 : n33859;
  assign n33861 = pi19 ? n33302 : n11418;
  assign n33862 = pi18 ? n37 : n33861;
  assign n33863 = pi21 ? n11921 : n32;
  assign n33864 = pi20 ? n33863 : n32;
  assign n33865 = pi19 ? n99 : n33864;
  assign n33866 = pi18 ? n33305 : n33865;
  assign n33867 = pi17 ? n33862 : n33866;
  assign n33868 = pi16 ? n33860 : n33867;
  assign n33869 = pi19 ? n32876 : n32933;
  assign n33870 = pi18 ? n31315 : n33869;
  assign n33871 = pi17 ? n32 : n33870;
  assign n33872 = pi19 ? n37 : n33315;
  assign n33873 = pi22 ? n7024 : n32;
  assign n33874 = pi21 ? n33873 : n32;
  assign n33875 = pi20 ? n33874 : n32;
  assign n33876 = pi19 ? n33317 : n33875;
  assign n33877 = pi18 ? n33872 : n33876;
  assign n33878 = pi17 ? n37 : n33877;
  assign n33879 = pi16 ? n33871 : n33878;
  assign n33880 = pi15 ? n33868 : n33879;
  assign n33881 = pi14 ? n33857 : n33880;
  assign n33882 = pi18 ? n31315 : n32877;
  assign n33883 = pi17 ? n32 : n33882;
  assign n33884 = pi23 ? n37 : n31328;
  assign n33885 = pi22 ? n33884 : n32;
  assign n33886 = pi21 ? n33885 : n32;
  assign n33887 = pi20 ? n33886 : n32;
  assign n33888 = pi19 ? n37 : n33887;
  assign n33889 = pi18 ? n37 : n33888;
  assign n33890 = pi17 ? n37 : n33889;
  assign n33891 = pi16 ? n33883 : n33890;
  assign n33892 = pi21 ? n29133 : n31200;
  assign n33893 = pi20 ? n20563 : n33892;
  assign n33894 = pi19 ? n33893 : n37;
  assign n33895 = pi18 ? n31315 : n33894;
  assign n33896 = pi17 ? n32 : n33895;
  assign n33897 = pi22 ? n1038 : n532;
  assign n33898 = pi21 ? n33897 : n32;
  assign n33899 = pi20 ? n33898 : n32;
  assign n33900 = pi19 ? n37 : n33899;
  assign n33901 = pi18 ? n37 : n33900;
  assign n33902 = pi17 ? n37 : n33901;
  assign n33903 = pi16 ? n33896 : n33902;
  assign n33904 = pi15 ? n33891 : n33903;
  assign n33905 = pi20 ? n20563 : n33845;
  assign n33906 = pi19 ? n33905 : n37;
  assign n33907 = pi18 ? n31315 : n33906;
  assign n33908 = pi17 ? n32 : n33907;
  assign n33909 = pi22 ? n295 : n532;
  assign n33910 = pi21 ? n33909 : n32;
  assign n33911 = pi20 ? n33910 : n32;
  assign n33912 = pi19 ? n8765 : n33911;
  assign n33913 = pi18 ? n37 : n33912;
  assign n33914 = pi17 ? n37 : n33913;
  assign n33915 = pi16 ? n33908 : n33914;
  assign n33916 = pi19 ? n33822 : n37;
  assign n33917 = pi18 ? n31315 : n33916;
  assign n33918 = pi17 ? n32 : n33917;
  assign n33919 = pi16 ? n33918 : n33914;
  assign n33920 = pi15 ? n33915 : n33919;
  assign n33921 = pi14 ? n33904 : n33920;
  assign n33922 = pi13 ? n33881 : n33921;
  assign n33923 = pi20 ? n20563 : n31298;
  assign n33924 = pi19 ? n33923 : n37;
  assign n33925 = pi18 ? n31315 : n33924;
  assign n33926 = pi17 ? n32 : n33925;
  assign n33927 = pi20 ? n18906 : n32;
  assign n33928 = pi19 ? n8765 : n33927;
  assign n33929 = pi18 ? n33348 : n33928;
  assign n33930 = pi17 ? n37 : n33929;
  assign n33931 = pi16 ? n33926 : n33930;
  assign n33932 = pi18 ? n31938 : n32349;
  assign n33933 = pi17 ? n32 : n33932;
  assign n33934 = pi22 ? n25629 : n688;
  assign n33935 = pi21 ? n33934 : n32;
  assign n33936 = pi20 ? n33935 : n32;
  assign n33937 = pi19 ? n9769 : n33936;
  assign n33938 = pi18 ? n37 : n33937;
  assign n33939 = pi17 ? n37 : n33938;
  assign n33940 = pi16 ? n33933 : n33939;
  assign n33941 = pi15 ? n33931 : n33940;
  assign n33942 = pi22 ? n1038 : n688;
  assign n33943 = pi21 ? n33942 : n32;
  assign n33944 = pi20 ? n33943 : n32;
  assign n33945 = pi19 ? n139 : n33944;
  assign n33946 = pi18 ? n33368 : n33945;
  assign n33947 = pi17 ? n37 : n33946;
  assign n33948 = pi16 ? n32915 : n33947;
  assign n33949 = pi20 ? n33821 : n37;
  assign n33950 = pi19 ? n33949 : n37;
  assign n33951 = pi18 ? n31315 : n33950;
  assign n33952 = pi17 ? n32 : n33951;
  assign n33953 = pi21 ? n9119 : n335;
  assign n33954 = pi20 ? n649 : n33953;
  assign n33955 = pi22 ? n6961 : n706;
  assign n33956 = pi21 ? n33955 : n32;
  assign n33957 = pi20 ? n33956 : n32;
  assign n33958 = pi19 ? n33954 : n33957;
  assign n33959 = pi18 ? n37 : n33958;
  assign n33960 = pi17 ? n37 : n33959;
  assign n33961 = pi16 ? n33952 : n33960;
  assign n33962 = pi15 ? n33948 : n33961;
  assign n33963 = pi14 ? n33941 : n33962;
  assign n33964 = pi21 ? n30195 : n37;
  assign n33965 = pi20 ? n33964 : n37;
  assign n33966 = pi19 ? n33965 : n37;
  assign n33967 = pi18 ? n31315 : n33966;
  assign n33968 = pi17 ? n32 : n33967;
  assign n33969 = pi22 ? n2060 : n706;
  assign n33970 = pi21 ? n33969 : n32;
  assign n33971 = pi20 ? n33970 : n32;
  assign n33972 = pi19 ? n10681 : n33971;
  assign n33973 = pi18 ? n37 : n33972;
  assign n33974 = pi17 ? n37 : n33973;
  assign n33975 = pi16 ? n33968 : n33974;
  assign n33976 = pi19 ? n33846 : n37;
  assign n33977 = pi18 ? n31315 : n33976;
  assign n33978 = pi17 ? n32 : n33977;
  assign n33979 = pi19 ? n12628 : n7019;
  assign n33980 = pi18 ? n37 : n33979;
  assign n33981 = pi17 ? n37 : n33980;
  assign n33982 = pi16 ? n33978 : n33981;
  assign n33983 = pi15 ? n33975 : n33982;
  assign n33984 = pi21 ? n31293 : n31924;
  assign n33985 = pi20 ? n32 : n33984;
  assign n33986 = pi19 ? n32 : n33985;
  assign n33987 = pi18 ? n33986 : n37;
  assign n33988 = pi17 ? n32 : n33987;
  assign n33989 = pi23 ? n1342 : n233;
  assign n33990 = pi22 ? n33989 : n32;
  assign n33991 = pi21 ? n33990 : n32;
  assign n33992 = pi20 ? n33991 : n32;
  assign n33993 = pi19 ? n37 : n33992;
  assign n33994 = pi18 ? n37 : n33993;
  assign n33995 = pi17 ? n37 : n33994;
  assign n33996 = pi16 ? n33988 : n33995;
  assign n33997 = pi21 ? n30866 : n31200;
  assign n33998 = pi20 ? n32 : n33997;
  assign n33999 = pi19 ? n32 : n33998;
  assign n34000 = pi18 ? n33999 : n37;
  assign n34001 = pi17 ? n32 : n34000;
  assign n34002 = pi16 ? n34001 : n33995;
  assign n34003 = pi15 ? n33996 : n34002;
  assign n34004 = pi14 ? n33983 : n34003;
  assign n34005 = pi13 ? n33963 : n34004;
  assign n34006 = pi12 ? n33922 : n34005;
  assign n34007 = pi19 ? n12478 : n7043;
  assign n34008 = pi18 ? n37 : n34007;
  assign n34009 = pi17 ? n37 : n34008;
  assign n34010 = pi16 ? n31987 : n34009;
  assign n34011 = pi22 ? n31993 : n37;
  assign n34012 = pi21 ? n34011 : n37;
  assign n34013 = pi20 ? n32 : n34012;
  assign n34014 = pi19 ? n32 : n34013;
  assign n34015 = pi18 ? n34014 : n37;
  assign n34016 = pi17 ? n32 : n34015;
  assign n34017 = pi19 ? n33431 : n4103;
  assign n34018 = pi18 ? n37 : n34017;
  assign n34019 = pi17 ? n37 : n34018;
  assign n34020 = pi16 ? n34016 : n34019;
  assign n34021 = pi15 ? n34010 : n34020;
  assign n34022 = pi19 ? n32459 : n5815;
  assign n34023 = pi18 ? n37 : n34022;
  assign n34024 = pi17 ? n37 : n34023;
  assign n34025 = pi16 ? n439 : n34024;
  assign n34026 = pi19 ? n33441 : n6408;
  assign n34027 = pi18 ? n37 : n34026;
  assign n34028 = pi17 ? n37 : n34027;
  assign n34029 = pi16 ? n439 : n34028;
  assign n34030 = pi15 ? n34025 : n34029;
  assign n34031 = pi14 ? n34021 : n34030;
  assign n34032 = pi13 ? n34031 : n33464;
  assign n34033 = pi14 ? n33476 : n33480;
  assign n34034 = pi19 ? n33022 : n7833;
  assign n34035 = pi18 ? n37 : n34034;
  assign n34036 = pi17 ? n37 : n34035;
  assign n34037 = pi16 ? n439 : n34036;
  assign n34038 = pi15 ? n34037 : n32507;
  assign n34039 = pi19 ? n33033 : n2702;
  assign n34040 = pi18 ? n37 : n34039;
  assign n34041 = pi17 ? n37 : n34040;
  assign n34042 = pi16 ? n439 : n34041;
  assign n34043 = pi20 ? n16008 : n2968;
  assign n34044 = pi19 ? n37 : n34043;
  assign n34045 = pi20 ? n2982 : n15964;
  assign n34046 = pi20 ? n2968 : n6500;
  assign n34047 = pi19 ? n34045 : n34046;
  assign n34048 = pi18 ? n34044 : n34047;
  assign n34049 = pi21 ? n2160 : n218;
  assign n34050 = pi20 ? n34049 : n28939;
  assign n34051 = pi19 ? n33499 : n34050;
  assign n34052 = pi19 ? n7839 : n1823;
  assign n34053 = pi18 ? n34051 : n34052;
  assign n34054 = pi17 ? n34048 : n34053;
  assign n34055 = pi16 ? n439 : n34054;
  assign n34056 = pi15 ? n34042 : n34055;
  assign n34057 = pi14 ? n34038 : n34056;
  assign n34058 = pi13 ? n34033 : n34057;
  assign n34059 = pi12 ? n34032 : n34058;
  assign n34060 = pi11 ? n34006 : n34059;
  assign n34061 = pi18 ? n33511 : n34052;
  assign n34062 = pi17 ? n32547 : n34061;
  assign n34063 = pi16 ? n439 : n34062;
  assign n34064 = pi19 ? n9035 : n1823;
  assign n34065 = pi18 ? n33519 : n34064;
  assign n34066 = pi17 ? n33516 : n34065;
  assign n34067 = pi16 ? n439 : n34066;
  assign n34068 = pi15 ? n34063 : n34067;
  assign n34069 = pi21 ? n777 : n3562;
  assign n34070 = pi20 ? n20977 : n34069;
  assign n34071 = pi19 ? n34070 : n32;
  assign n34072 = pi18 ? n99 : n34071;
  assign n34073 = pi17 ? n99 : n34072;
  assign n34074 = pi16 ? n23698 : n34073;
  assign n34075 = pi15 ? n33526 : n34074;
  assign n34076 = pi14 ? n34068 : n34075;
  assign n34077 = pi21 ? n777 : n316;
  assign n34078 = pi20 ? n2238 : n34077;
  assign n34079 = pi19 ? n34078 : n32;
  assign n34080 = pi18 ? n99 : n34079;
  assign n34081 = pi17 ? n99 : n34080;
  assign n34082 = pi16 ? n744 : n34081;
  assign n34083 = pi21 ? n99 : n26256;
  assign n34084 = pi20 ? n99 : n34083;
  assign n34085 = pi19 ? n34084 : n32;
  assign n34086 = pi18 ? n99 : n34085;
  assign n34087 = pi17 ? n99 : n34086;
  assign n34088 = pi16 ? n744 : n34087;
  assign n34089 = pi15 ? n34082 : n34088;
  assign n34090 = pi19 ? n316 : n32;
  assign n34091 = pi18 ? n33551 : n34090;
  assign n34092 = pi17 ? n139 : n34091;
  assign n34093 = pi16 ? n30470 : n34092;
  assign n34094 = pi18 ? n33558 : n33082;
  assign n34095 = pi17 ? n139 : n34094;
  assign n34096 = pi16 ? n33556 : n34095;
  assign n34097 = pi15 ? n34093 : n34096;
  assign n34098 = pi14 ? n34089 : n34097;
  assign n34099 = pi13 ? n34076 : n34098;
  assign n34100 = pi20 ? n316 : n18715;
  assign n34101 = pi19 ? n34100 : n32;
  assign n34102 = pi18 ? n33569 : n34101;
  assign n34103 = pi17 ? n33568 : n34102;
  assign n34104 = pi16 ? n439 : n34103;
  assign n34105 = pi20 ? n316 : n18721;
  assign n34106 = pi19 ? n34105 : n32;
  assign n34107 = pi18 ? n33580 : n34106;
  assign n34108 = pi17 ? n33576 : n34107;
  assign n34109 = pi16 ? n439 : n34108;
  assign n34110 = pi15 ? n34104 : n34109;
  assign n34111 = pi21 ? n204 : n5746;
  assign n34112 = pi20 ? n204 : n34111;
  assign n34113 = pi19 ? n34112 : n32;
  assign n34114 = pi18 ? n33586 : n34113;
  assign n34115 = pi17 ? n32638 : n34114;
  assign n34116 = pi16 ? n439 : n34115;
  assign n34117 = pi18 ? n204 : n34113;
  assign n34118 = pi17 ? n33593 : n34117;
  assign n34119 = pi16 ? n439 : n34118;
  assign n34120 = pi15 ? n34116 : n34119;
  assign n34121 = pi14 ? n34110 : n34120;
  assign n34122 = pi18 ? n204 : n26138;
  assign n34123 = pi17 ? n33602 : n34122;
  assign n34124 = pi16 ? n32657 : n34123;
  assign n34125 = pi21 ? n204 : n14789;
  assign n34126 = pi20 ? n204 : n34125;
  assign n34127 = pi19 ? n34126 : n32;
  assign n34128 = pi18 ? n204 : n34127;
  assign n34129 = pi17 ? n32665 : n34128;
  assign n34130 = pi16 ? n439 : n34129;
  assign n34131 = pi15 ? n34124 : n34130;
  assign n34132 = pi23 ? n4882 : n685;
  assign n34133 = pi22 ? n34132 : n32;
  assign n34134 = pi21 ? n204 : n34133;
  assign n34135 = pi20 ? n204 : n34134;
  assign n34136 = pi19 ? n34135 : n32;
  assign n34137 = pi18 ? n33616 : n34136;
  assign n34138 = pi17 ? n33614 : n34137;
  assign n34139 = pi16 ? n439 : n34138;
  assign n34140 = pi20 ? n233 : n22089;
  assign n34141 = pi19 ? n34140 : n32;
  assign n34142 = pi18 ? n33621 : n34141;
  assign n34143 = pi17 ? n33614 : n34142;
  assign n34144 = pi16 ? n439 : n34143;
  assign n34145 = pi15 ? n34139 : n34144;
  assign n34146 = pi14 ? n34131 : n34145;
  assign n34147 = pi13 ? n34121 : n34146;
  assign n34148 = pi12 ? n34099 : n34147;
  assign n34149 = pi21 ? n233 : n7048;
  assign n34150 = pi20 ? n233 : n34149;
  assign n34151 = pi19 ? n34150 : n32;
  assign n34152 = pi18 ? n32704 : n34151;
  assign n34153 = pi17 ? n33634 : n34152;
  assign n34154 = pi16 ? n439 : n34153;
  assign n34155 = pi20 ? n233 : n22103;
  assign n34156 = pi19 ? n34155 : n32;
  assign n34157 = pi18 ? n335 : n34156;
  assign n34158 = pi17 ? n32712 : n34157;
  assign n34159 = pi16 ? n439 : n34158;
  assign n34160 = pi15 ? n34154 : n34159;
  assign n34161 = pi20 ? n233 : n24379;
  assign n34162 = pi19 ? n34161 : n32;
  assign n34163 = pi18 ? n17205 : n34162;
  assign n34164 = pi17 ? n32725 : n34163;
  assign n34165 = pi16 ? n33651 : n34164;
  assign n34166 = pi20 ? n233 : n18392;
  assign n34167 = pi19 ? n34166 : n32;
  assign n34168 = pi18 ? n7677 : n34167;
  assign n34169 = pi17 ? n32735 : n34168;
  assign n34170 = pi16 ? n25090 : n34169;
  assign n34171 = pi15 ? n34165 : n34170;
  assign n34172 = pi14 ? n34160 : n34171;
  assign n34173 = pi20 ? n233 : n17898;
  assign n34174 = pi19 ? n34173 : n32;
  assign n34175 = pi18 ? n2102 : n34174;
  assign n34176 = pi17 ? n32741 : n34175;
  assign n34177 = pi16 ? n33669 : n34176;
  assign n34178 = pi18 ? n33675 : n34174;
  assign n34179 = pi17 ? n33673 : n34178;
  assign n34180 = pi16 ? n439 : n34179;
  assign n34181 = pi15 ? n34177 : n34180;
  assign n34182 = pi18 ? n33690 : n33660;
  assign n34183 = pi17 ? n33687 : n34182;
  assign n34184 = pi16 ? n33682 : n34183;
  assign n34185 = pi20 ? n1921 : n233;
  assign n34186 = pi19 ? n33694 : n34185;
  assign n34187 = pi18 ? n34186 : n233;
  assign n34188 = pi20 ? n233 : n17905;
  assign n34189 = pi19 ? n34188 : n32;
  assign n34190 = pi18 ? n33700 : n34189;
  assign n34191 = pi17 ? n34187 : n34190;
  assign n34192 = pi16 ? n439 : n34191;
  assign n34193 = pi15 ? n34184 : n34192;
  assign n34194 = pi14 ? n34181 : n34193;
  assign n34195 = pi13 ? n34172 : n34194;
  assign n34196 = pi24 ? n32 : n30868;
  assign n34197 = pi23 ? n34196 : n139;
  assign n34198 = pi22 ? n34197 : n139;
  assign n34199 = pi21 ? n34198 : n139;
  assign n34200 = pi20 ? n32 : n34199;
  assign n34201 = pi19 ? n32 : n34200;
  assign n34202 = pi21 ? n139 : n20228;
  assign n34203 = pi20 ? n29839 : n34202;
  assign n34204 = pi19 ? n139 : n34203;
  assign n34205 = pi18 ? n34201 : n34204;
  assign n34206 = pi17 ? n32 : n34205;
  assign n34207 = pi22 ? n139 : n18795;
  assign n34208 = pi21 ? n34207 : n139;
  assign n34209 = pi21 ? n34207 : n22236;
  assign n34210 = pi20 ? n34208 : n34209;
  assign n34211 = pi21 ? n20600 : n34207;
  assign n34212 = pi20 ? n34209 : n34211;
  assign n34213 = pi19 ? n34210 : n34212;
  assign n34214 = pi21 ? n20228 : n139;
  assign n34215 = pi20 ? n20228 : n23182;
  assign n34216 = pi19 ? n34214 : n34215;
  assign n34217 = pi18 ? n34213 : n34216;
  assign n34218 = pi21 ? n34207 : n20228;
  assign n34219 = pi21 ? n363 : n20605;
  assign n34220 = pi20 ? n34218 : n34219;
  assign n34221 = pi21 ? n20228 : n363;
  assign n34222 = pi20 ? n34221 : n33738;
  assign n34223 = pi19 ? n34220 : n34222;
  assign n34224 = pi18 ? n34223 : n33782;
  assign n34225 = pi17 ? n34217 : n34224;
  assign n34226 = pi16 ? n34206 : n34225;
  assign n34227 = pi15 ? n34226 : n33790;
  assign n34228 = pi20 ? n26890 : n2638;
  assign n34229 = pi19 ? n34228 : n32;
  assign n34230 = pi18 ? n32832 : n34229;
  assign n34231 = pi17 ? n363 : n34230;
  assign n34232 = pi16 ? n21561 : n34231;
  assign n34233 = pi18 ? n32832 : n19946;
  assign n34234 = pi17 ? n363 : n34233;
  assign n34235 = pi16 ? n21561 : n34234;
  assign n34236 = pi15 ? n34232 : n34235;
  assign n34237 = pi14 ? n34227 : n34236;
  assign n34238 = pi13 ? n33747 : n34237;
  assign n34239 = pi12 ? n34195 : n34238;
  assign n34240 = pi11 ? n34148 : n34239;
  assign n34241 = pi10 ? n34060 : n34240;
  assign n34242 = pi09 ? n33837 : n34241;
  assign n34243 = pi08 ? n33820 : n34242;
  assign n34244 = pi07 ? n33244 : n34243;
  assign n34245 = pi06 ? n32274 : n34244;
  assign n34246 = pi20 ? n20563 : n31913;
  assign n34247 = pi19 ? n20563 : n34246;
  assign n34248 = pi18 ? n30119 : n34247;
  assign n34249 = pi17 ? n32 : n34248;
  assign n34250 = pi20 ? n3824 : n4202;
  assign n34251 = pi19 ? n34250 : n99;
  assign n34252 = pi18 ? n37 : n34251;
  assign n34253 = pi19 ? n99 : n5431;
  assign n34254 = pi18 ? n99 : n34253;
  assign n34255 = pi17 ? n34252 : n34254;
  assign n34256 = pi16 ? n34249 : n34255;
  assign n34257 = pi15 ? n32 : n34256;
  assign n34258 = pi19 ? n20563 : n32294;
  assign n34259 = pi18 ? n30119 : n34258;
  assign n34260 = pi17 ? n32 : n34259;
  assign n34261 = pi20 ? n37 : n14844;
  assign n34262 = pi19 ? n37 : n34261;
  assign n34263 = pi18 ? n34262 : n99;
  assign n34264 = pi19 ? n99 : n5439;
  assign n34265 = pi18 ? n99 : n34264;
  assign n34266 = pi17 ? n34263 : n34265;
  assign n34267 = pi16 ? n34260 : n34266;
  assign n34268 = pi16 ? n33825 : n34266;
  assign n34269 = pi15 ? n34267 : n34268;
  assign n34270 = pi14 ? n34257 : n34269;
  assign n34271 = pi13 ? n32 : n34270;
  assign n34272 = pi12 ? n32 : n34271;
  assign n34273 = pi11 ? n32 : n34272;
  assign n34274 = pi10 ? n32 : n34273;
  assign n34275 = pi18 ? n31265 : n33245;
  assign n34276 = pi17 ? n32 : n34275;
  assign n34277 = pi19 ? n34261 : n99;
  assign n34278 = pi18 ? n37 : n34277;
  assign n34279 = pi19 ? n15543 : n5446;
  assign n34280 = pi18 ? n99 : n34279;
  assign n34281 = pi17 ? n34278 : n34280;
  assign n34282 = pi16 ? n34276 : n34281;
  assign n34283 = pi18 ? n31265 : n33828;
  assign n34284 = pi17 ? n32 : n34283;
  assign n34285 = pi19 ? n6046 : n99;
  assign n34286 = pi18 ? n37 : n34285;
  assign n34287 = pi22 ? n99 : n1370;
  assign n34288 = pi21 ? n34287 : n32;
  assign n34289 = pi20 ? n34288 : n32;
  assign n34290 = pi19 ? n99 : n34289;
  assign n34291 = pi18 ? n99 : n34290;
  assign n34292 = pi17 ? n34286 : n34291;
  assign n34293 = pi16 ? n34284 : n34292;
  assign n34294 = pi15 ? n34282 : n34293;
  assign n34295 = pi19 ? n20563 : n32348;
  assign n34296 = pi18 ? n31265 : n34295;
  assign n34297 = pi17 ? n32 : n34296;
  assign n34298 = pi18 ? n30851 : n99;
  assign n34299 = pi21 ? n12267 : n32;
  assign n34300 = pi20 ? n34299 : n32;
  assign n34301 = pi19 ? n99 : n34300;
  assign n34302 = pi18 ? n99 : n34301;
  assign n34303 = pi17 ? n34298 : n34302;
  assign n34304 = pi16 ? n34297 : n34303;
  assign n34305 = pi18 ? n31315 : n33260;
  assign n34306 = pi17 ? n32 : n34305;
  assign n34307 = pi19 ? n37 : n31363;
  assign n34308 = pi20 ? n376 : n14038;
  assign n34309 = pi22 ? n295 : n5631;
  assign n34310 = pi21 ? n34309 : n32;
  assign n34311 = pi20 ? n34310 : n32;
  assign n34312 = pi19 ? n34308 : n34311;
  assign n34313 = pi18 ? n34307 : n34312;
  assign n34314 = pi17 ? n37 : n34313;
  assign n34315 = pi16 ? n34306 : n34314;
  assign n34316 = pi15 ? n34304 : n34315;
  assign n34317 = pi14 ? n34294 : n34316;
  assign n34318 = pi18 ? n31938 : n32275;
  assign n34319 = pi17 ? n32 : n34318;
  assign n34320 = pi22 ? n295 : n2468;
  assign n34321 = pi21 ? n34320 : n32;
  assign n34322 = pi20 ? n34321 : n32;
  assign n34323 = pi19 ? n37 : n34322;
  assign n34324 = pi18 ? n37 : n34323;
  assign n34325 = pi17 ? n37 : n34324;
  assign n34326 = pi16 ? n34319 : n34325;
  assign n34327 = pi18 ? n31315 : n33285;
  assign n34328 = pi17 ? n32 : n34327;
  assign n34329 = pi19 ? n9814 : n4738;
  assign n34330 = pi18 ? n37 : n34329;
  assign n34331 = pi17 ? n37 : n34330;
  assign n34332 = pi16 ? n34328 : n34331;
  assign n34333 = pi15 ? n34326 : n34332;
  assign n34334 = pi18 ? n31315 : n33299;
  assign n34335 = pi17 ? n32 : n34334;
  assign n34336 = pi20 ? n992 : n37;
  assign n34337 = pi19 ? n3083 : n34336;
  assign n34338 = pi19 ? n8765 : n4738;
  assign n34339 = pi18 ? n34337 : n34338;
  assign n34340 = pi17 ? n37 : n34339;
  assign n34341 = pi16 ? n34335 : n34340;
  assign n34342 = pi18 ? n37 : n13167;
  assign n34343 = pi19 ? n8765 : n2307;
  assign n34344 = pi19 ? n9769 : n33927;
  assign n34345 = pi18 ? n34343 : n34344;
  assign n34346 = pi17 ? n34342 : n34345;
  assign n34347 = pi16 ? n34335 : n34346;
  assign n34348 = pi15 ? n34341 : n34347;
  assign n34349 = pi14 ? n34333 : n34348;
  assign n34350 = pi13 ? n34317 : n34349;
  assign n34351 = pi18 ? n31938 : n32295;
  assign n34352 = pi17 ? n32 : n34351;
  assign n34353 = pi20 ? n13139 : n37;
  assign n34354 = pi19 ? n9814 : n34353;
  assign n34355 = pi18 ? n34354 : n33928;
  assign n34356 = pi17 ? n37 : n34355;
  assign n34357 = pi16 ? n34352 : n34356;
  assign n34358 = pi19 ? n31221 : n37;
  assign n34359 = pi18 ? n31315 : n34358;
  assign n34360 = pi17 ? n32 : n34359;
  assign n34361 = pi19 ? n37 : n18070;
  assign n34362 = pi20 ? n18917 : n32;
  assign n34363 = pi19 ? n8765 : n34362;
  assign n34364 = pi18 ? n34361 : n34363;
  assign n34365 = pi17 ? n37 : n34364;
  assign n34366 = pi16 ? n34360 : n34365;
  assign n34367 = pi15 ? n34357 : n34366;
  assign n34368 = pi21 ? n139 : n335;
  assign n34369 = pi20 ? n3087 : n34368;
  assign n34370 = pi19 ? n34369 : n34362;
  assign n34371 = pi18 ? n34361 : n34370;
  assign n34372 = pi17 ? n37 : n34371;
  assign n34373 = pi16 ? n34360 : n34372;
  assign n34374 = pi22 ? n335 : n706;
  assign n34375 = pi21 ? n34374 : n32;
  assign n34376 = pi20 ? n34375 : n32;
  assign n34377 = pi19 ? n17204 : n34376;
  assign n34378 = pi18 ? n37 : n34377;
  assign n34379 = pi17 ? n37 : n34378;
  assign n34380 = pi16 ? n32901 : n34379;
  assign n34381 = pi15 ? n34373 : n34380;
  assign n34382 = pi14 ? n34367 : n34381;
  assign n34383 = pi22 ? n363 : n706;
  assign n34384 = pi21 ? n34383 : n32;
  assign n34385 = pi20 ? n34384 : n32;
  assign n34386 = pi19 ? n12628 : n34385;
  assign n34387 = pi18 ? n37 : n34386;
  assign n34388 = pi17 ? n37 : n34387;
  assign n34389 = pi16 ? n32901 : n34388;
  assign n34390 = pi21 ? n11026 : n32;
  assign n34391 = pi20 ? n34390 : n32;
  assign n34392 = pi19 ? n25087 : n34391;
  assign n34393 = pi18 ? n37 : n34392;
  assign n34394 = pi17 ? n37 : n34393;
  assign n34395 = pi16 ? n32379 : n34394;
  assign n34396 = pi15 ? n34389 : n34395;
  assign n34397 = pi22 ? n448 : n32;
  assign n34398 = pi21 ? n34397 : n32;
  assign n34399 = pi20 ? n34398 : n32;
  assign n34400 = pi19 ? n37 : n34399;
  assign n34401 = pi18 ? n37 : n34400;
  assign n34402 = pi17 ? n37 : n34401;
  assign n34403 = pi16 ? n33374 : n34402;
  assign n34404 = pi20 ? n37 : n25125;
  assign n34405 = pi19 ? n34404 : n4853;
  assign n34406 = pi18 ? n37 : n34405;
  assign n34407 = pi17 ? n37 : n34406;
  assign n34408 = pi16 ? n32388 : n34407;
  assign n34409 = pi15 ? n34403 : n34408;
  assign n34410 = pi14 ? n34396 : n34409;
  assign n34411 = pi13 ? n34382 : n34410;
  assign n34412 = pi12 ? n34350 : n34411;
  assign n34413 = pi20 ? n577 : n16544;
  assign n34414 = pi19 ? n34413 : n7036;
  assign n34415 = pi18 ? n37 : n34414;
  assign n34416 = pi17 ? n37 : n34415;
  assign n34417 = pi16 ? n31317 : n34416;
  assign n34418 = pi19 ? n37 : n3289;
  assign n34419 = pi18 ? n37 : n34418;
  assign n34420 = pi20 ? n3292 : n639;
  assign n34421 = pi20 ? n24105 : n37;
  assign n34422 = pi19 ? n34420 : n34421;
  assign n34423 = pi20 ? n577 : n26846;
  assign n34424 = pi19 ? n34423 : n7036;
  assign n34425 = pi18 ? n34422 : n34424;
  assign n34426 = pi17 ? n34419 : n34425;
  assign n34427 = pi16 ? n32388 : n34426;
  assign n34428 = pi15 ? n34417 : n34427;
  assign n34429 = pi19 ? n603 : n5773;
  assign n34430 = pi18 ? n37 : n34429;
  assign n34431 = pi17 ? n37 : n34430;
  assign n34432 = pi16 ? n31317 : n34431;
  assign n34433 = pi20 ? n20157 : n24865;
  assign n34434 = pi19 ? n34433 : n5773;
  assign n34435 = pi18 ? n37 : n34434;
  assign n34436 = pi17 ? n37 : n34435;
  assign n34437 = pi16 ? n33409 : n34436;
  assign n34438 = pi15 ? n34432 : n34437;
  assign n34439 = pi14 ? n34428 : n34438;
  assign n34440 = pi21 ? n31293 : n37;
  assign n34441 = pi20 ? n32 : n34440;
  assign n34442 = pi19 ? n32 : n34441;
  assign n34443 = pi18 ? n34442 : n37;
  assign n34444 = pi17 ? n32 : n34443;
  assign n34445 = pi20 ? n7730 : n23175;
  assign n34446 = pi20 ? n21388 : n32;
  assign n34447 = pi19 ? n34445 : n34446;
  assign n34448 = pi18 ? n37 : n34447;
  assign n34449 = pi17 ? n37 : n34448;
  assign n34450 = pi16 ? n34444 : n34449;
  assign n34451 = pi19 ? n5029 : n7725;
  assign n34452 = pi18 ? n37 : n34451;
  assign n34453 = pi17 ? n37 : n34452;
  assign n34454 = pi16 ? n32415 : n34453;
  assign n34455 = pi15 ? n34450 : n34454;
  assign n34456 = pi19 ? n6403 : n3211;
  assign n34457 = pi18 ? n37 : n34456;
  assign n34458 = pi17 ? n37 : n34457;
  assign n34459 = pi16 ? n32014 : n34458;
  assign n34460 = pi14 ? n34455 : n34459;
  assign n34461 = pi13 ? n34439 : n34460;
  assign n34462 = pi20 ? n20902 : n32;
  assign n34463 = pi19 ? n5029 : n34462;
  assign n34464 = pi18 ? n37 : n34463;
  assign n34465 = pi17 ? n37 : n34464;
  assign n34466 = pi16 ? n32014 : n34465;
  assign n34467 = pi19 ? n6403 : n3321;
  assign n34468 = pi18 ? n37 : n34467;
  assign n34469 = pi17 ? n37 : n34468;
  assign n34470 = pi16 ? n439 : n34469;
  assign n34471 = pi15 ? n34466 : n34470;
  assign n34472 = pi19 ? n6403 : n4117;
  assign n34473 = pi18 ? n37 : n34472;
  assign n34474 = pi17 ? n37 : n34473;
  assign n34475 = pi16 ? n439 : n34474;
  assign n34476 = pi15 ? n34475 : n33463;
  assign n34477 = pi14 ? n34471 : n34476;
  assign n34478 = pi21 ? n19958 : n19933;
  assign n34479 = pi20 ? n37 : n34478;
  assign n34480 = pi19 ? n34479 : n10012;
  assign n34481 = pi18 ? n37 : n34480;
  assign n34482 = pi17 ? n37 : n34481;
  assign n34483 = pi16 ? n439 : n34482;
  assign n34484 = pi19 ? n34479 : n2680;
  assign n34485 = pi18 ? n37 : n34484;
  assign n34486 = pi17 ? n37 : n34485;
  assign n34487 = pi16 ? n439 : n34486;
  assign n34488 = pi15 ? n34483 : n34487;
  assign n34489 = pi19 ? n37 : n24494;
  assign n34490 = pi21 ? n272 : n37;
  assign n34491 = pi20 ? n279 : n34490;
  assign n34492 = pi20 ? n30414 : n278;
  assign n34493 = pi19 ? n34491 : n34492;
  assign n34494 = pi19 ? n157 : n2702;
  assign n34495 = pi18 ? n34493 : n34494;
  assign n34496 = pi17 ? n34489 : n34495;
  assign n34497 = pi16 ? n439 : n34496;
  assign n34498 = pi20 ? n2243 : n157;
  assign n34499 = pi19 ? n21611 : n34498;
  assign n34500 = pi18 ? n34499 : n157;
  assign n34501 = pi20 ? n157 : n6508;
  assign n34502 = pi19 ? n34501 : n157;
  assign n34503 = pi18 ? n34502 : n34494;
  assign n34504 = pi17 ? n34500 : n34503;
  assign n34505 = pi16 ? n439 : n34504;
  assign n34506 = pi15 ? n34497 : n34505;
  assign n34507 = pi14 ? n34488 : n34506;
  assign n34508 = pi13 ? n34477 : n34507;
  assign n34509 = pi12 ? n34461 : n34508;
  assign n34510 = pi11 ? n34412 : n34509;
  assign n34511 = pi20 ? n7745 : n2238;
  assign n34512 = pi19 ? n37 : n34511;
  assign n34513 = pi21 ? n37 : n159;
  assign n34514 = pi20 ? n15263 : n34513;
  assign n34515 = pi21 ? n157 : n5899;
  assign n34516 = pi20 ? n9997 : n34515;
  assign n34517 = pi19 ? n34514 : n34516;
  assign n34518 = pi18 ? n34512 : n34517;
  assign n34519 = pi19 ? n19137 : n157;
  assign n34520 = pi19 ? n157 : n1823;
  assign n34521 = pi18 ? n34519 : n34520;
  assign n34522 = pi17 ? n34518 : n34521;
  assign n34523 = pi16 ? n439 : n34522;
  assign n34524 = pi20 ? n7745 : n99;
  assign n34525 = pi19 ? n37 : n34524;
  assign n34526 = pi19 ? n14844 : n7845;
  assign n34527 = pi18 ? n34525 : n34526;
  assign n34528 = pi21 ? n14461 : n99;
  assign n34529 = pi20 ? n776 : n34528;
  assign n34530 = pi20 ? n802 : n2243;
  assign n34531 = pi19 ? n34529 : n34530;
  assign n34532 = pi18 ? n34531 : n34064;
  assign n34533 = pi17 ? n34527 : n34532;
  assign n34534 = pi16 ? n439 : n34533;
  assign n34535 = pi15 ? n34523 : n34534;
  assign n34536 = pi19 ? n14285 : n7845;
  assign n34537 = pi21 ? n157 : n316;
  assign n34538 = pi21 ? n316 : n3562;
  assign n34539 = pi20 ? n34537 : n34538;
  assign n34540 = pi19 ? n34539 : n32;
  assign n34541 = pi18 ? n34536 : n34540;
  assign n34542 = pi17 ? n99 : n34541;
  assign n34543 = pi16 ? n201 : n34542;
  assign n34544 = pi20 ? n34077 : n20978;
  assign n34545 = pi19 ? n34544 : n32;
  assign n34546 = pi18 ? n99 : n34545;
  assign n34547 = pi17 ? n99 : n34546;
  assign n34548 = pi16 ? n25610 : n34547;
  assign n34549 = pi15 ? n34543 : n34548;
  assign n34550 = pi14 ? n34535 : n34549;
  assign n34551 = pi21 ? n99 : n33058;
  assign n34552 = pi20 ? n99 : n34551;
  assign n34553 = pi19 ? n34552 : n32;
  assign n34554 = pi18 ? n99 : n34553;
  assign n34555 = pi17 ? n99 : n34554;
  assign n34556 = pi16 ? n1510 : n34555;
  assign n34557 = pi23 ? n3491 : n204;
  assign n34558 = pi22 ? n34557 : n316;
  assign n34559 = pi21 ? n99 : n34558;
  assign n34560 = pi20 ? n99 : n34559;
  assign n34561 = pi19 ? n34560 : n32;
  assign n34562 = pi18 ? n99 : n34561;
  assign n34563 = pi17 ? n99 : n34562;
  assign n34564 = pi16 ? n23698 : n34563;
  assign n34565 = pi15 ? n34556 : n34564;
  assign n34566 = pi20 ? n226 : n219;
  assign n34567 = pi19 ? n34566 : n17972;
  assign n34568 = pi18 ? n799 : n34567;
  assign n34569 = pi17 ? n32 : n34568;
  assign n34570 = pi21 ? n4247 : n139;
  assign n34571 = pi20 ? n34570 : n139;
  assign n34572 = pi19 ? n34571 : n139;
  assign n34573 = pi18 ? n34572 : n139;
  assign n34574 = pi21 ? n139 : n4247;
  assign n34575 = pi20 ? n139 : n34574;
  assign n34576 = pi19 ? n139 : n34575;
  assign n34577 = pi20 ? n20978 : n316;
  assign n34578 = pi19 ? n34577 : n32;
  assign n34579 = pi18 ? n34576 : n34578;
  assign n34580 = pi17 ? n34573 : n34579;
  assign n34581 = pi16 ? n34569 : n34580;
  assign n34582 = pi19 ? n37 : n14033;
  assign n34583 = pi18 ? n374 : n34582;
  assign n34584 = pi17 ? n32 : n34583;
  assign n34585 = pi19 ? n13192 : n139;
  assign n34586 = pi18 ? n34585 : n139;
  assign n34587 = pi21 ? n139 : n3693;
  assign n34588 = pi20 ? n139 : n34587;
  assign n34589 = pi19 ? n139 : n34588;
  assign n34590 = pi19 ? n5288 : n32;
  assign n34591 = pi18 ? n34589 : n34590;
  assign n34592 = pi17 ? n34586 : n34591;
  assign n34593 = pi16 ? n34584 : n34592;
  assign n34594 = pi15 ? n34581 : n34593;
  assign n34595 = pi14 ? n34565 : n34594;
  assign n34596 = pi13 ? n34550 : n34595;
  assign n34597 = pi19 ? n12370 : n139;
  assign n34598 = pi18 ? n34597 : n139;
  assign n34599 = pi20 ? n1001 : n19249;
  assign n34600 = pi19 ? n34599 : n32;
  assign n34601 = pi18 ? n31565 : n34600;
  assign n34602 = pi17 ? n34598 : n34601;
  assign n34603 = pi16 ? n439 : n34602;
  assign n34604 = pi20 ? n139 : n16493;
  assign n34605 = pi19 ? n139 : n34604;
  assign n34606 = pi18 ? n14115 : n34605;
  assign n34607 = pi20 ? n1582 : n3096;
  assign n34608 = pi19 ? n34607 : n32663;
  assign n34609 = pi21 ? n204 : n4748;
  assign n34610 = pi20 ? n204 : n34609;
  assign n34611 = pi19 ? n34610 : n32;
  assign n34612 = pi18 ? n34608 : n34611;
  assign n34613 = pi17 ? n34606 : n34612;
  assign n34614 = pi16 ? n439 : n34613;
  assign n34615 = pi15 ? n34603 : n34614;
  assign n34616 = pi20 ? n28575 : n1906;
  assign n34617 = pi19 ? n37 : n34616;
  assign n34618 = pi21 ? n139 : n499;
  assign n34619 = pi20 ? n34618 : n1016;
  assign n34620 = pi19 ? n34619 : n204;
  assign n34621 = pi18 ? n34617 : n34620;
  assign n34622 = pi20 ? n204 : n1016;
  assign n34623 = pi19 ? n34622 : n204;
  assign n34624 = pi20 ? n2316 : n34609;
  assign n34625 = pi19 ? n34624 : n32;
  assign n34626 = pi18 ? n34623 : n34625;
  assign n34627 = pi17 ? n34621 : n34626;
  assign n34628 = pi16 ? n439 : n34627;
  assign n34629 = pi20 ? n1056 : n1057;
  assign n34630 = pi19 ? n37 : n34629;
  assign n34631 = pi18 ? n34630 : n204;
  assign n34632 = pi18 ? n204 : n34611;
  assign n34633 = pi17 ? n34631 : n34632;
  assign n34634 = pi16 ? n439 : n34633;
  assign n34635 = pi15 ? n34628 : n34634;
  assign n34636 = pi14 ? n34615 : n34635;
  assign n34637 = pi20 ? n3086 : n1003;
  assign n34638 = pi19 ? n37 : n34637;
  assign n34639 = pi18 ? n374 : n34638;
  assign n34640 = pi17 ? n32 : n34639;
  assign n34641 = pi20 ? n5199 : n204;
  assign n34642 = pi19 ? n14962 : n34641;
  assign n34643 = pi18 ? n34642 : n204;
  assign n34644 = pi22 ? n4079 : n532;
  assign n34645 = pi21 ? n204 : n34644;
  assign n34646 = pi20 ? n204 : n34645;
  assign n34647 = pi19 ? n34646 : n32;
  assign n34648 = pi18 ? n204 : n34647;
  assign n34649 = pi17 ? n34643 : n34648;
  assign n34650 = pi16 ? n34640 : n34649;
  assign n34651 = pi19 ? n1017 : n204;
  assign n34652 = pi18 ? n14963 : n34651;
  assign n34653 = pi21 ? n204 : n26303;
  assign n34654 = pi20 ? n204 : n34653;
  assign n34655 = pi19 ? n34654 : n32;
  assign n34656 = pi18 ? n204 : n34655;
  assign n34657 = pi17 ? n34652 : n34656;
  assign n34658 = pi16 ? n439 : n34657;
  assign n34659 = pi15 ? n34650 : n34658;
  assign n34660 = pi22 ? n233 : n139;
  assign n34661 = pi21 ? n37 : n34660;
  assign n34662 = pi20 ? n3083 : n34661;
  assign n34663 = pi19 ? n34662 : n19358;
  assign n34664 = pi18 ? n37 : n34663;
  assign n34665 = pi21 ? n3073 : n28649;
  assign n34666 = pi20 ? n233 : n34665;
  assign n34667 = pi19 ? n34666 : n233;
  assign n34668 = pi21 ? n1039 : n19337;
  assign n34669 = pi21 ? n19337 : n7002;
  assign n34670 = pi20 ? n34668 : n34669;
  assign n34671 = pi19 ? n34670 : n32;
  assign n34672 = pi18 ? n34667 : n34671;
  assign n34673 = pi17 ? n34664 : n34672;
  assign n34674 = pi16 ? n439 : n34673;
  assign n34675 = pi19 ? n23844 : n19358;
  assign n34676 = pi18 ? n37 : n34675;
  assign n34677 = pi20 ? n233 : n8857;
  assign n34678 = pi20 ? n25957 : n233;
  assign n34679 = pi19 ? n34677 : n34678;
  assign n34680 = pi21 ? n233 : n7002;
  assign n34681 = pi20 ? n233 : n34680;
  assign n34682 = pi19 ? n34681 : n32;
  assign n34683 = pi18 ? n34679 : n34682;
  assign n34684 = pi17 ? n34676 : n34683;
  assign n34685 = pi16 ? n439 : n34684;
  assign n34686 = pi15 ? n34674 : n34685;
  assign n34687 = pi14 ? n34659 : n34686;
  assign n34688 = pi13 ? n34636 : n34687;
  assign n34689 = pi12 ? n34596 : n34688;
  assign n34690 = pi20 ? n233 : n24629;
  assign n34691 = pi19 ? n34690 : n32;
  assign n34692 = pi18 ? n17205 : n34691;
  assign n34693 = pi17 ? n6339 : n34692;
  assign n34694 = pi16 ? n439 : n34693;
  assign n34695 = pi19 ? n7685 : n10681;
  assign n34696 = pi18 ? n37 : n34695;
  assign n34697 = pi19 ? n335 : n10681;
  assign n34698 = pi20 ? n33688 : n14657;
  assign n34699 = pi19 ? n34698 : n32;
  assign n34700 = pi18 ? n34697 : n34699;
  assign n34701 = pi17 ? n34696 : n34700;
  assign n34702 = pi16 ? n439 : n34701;
  assign n34703 = pi15 ? n34694 : n34702;
  assign n34704 = pi18 ? n374 : n7686;
  assign n34705 = pi17 ? n32 : n34704;
  assign n34706 = pi18 ? n34697 : n32724;
  assign n34707 = pi19 ? n577 : n6340;
  assign n34708 = pi21 ? n4920 : n19386;
  assign n34709 = pi21 ? n233 : n882;
  assign n34710 = pi20 ? n34708 : n34709;
  assign n34711 = pi19 ? n34710 : n32;
  assign n34712 = pi18 ? n34707 : n34711;
  assign n34713 = pi17 ? n34706 : n34712;
  assign n34714 = pi16 ? n34705 : n34713;
  assign n34715 = pi19 ? n335 : n14166;
  assign n34716 = pi19 ? n17500 : n37;
  assign n34717 = pi18 ? n34715 : n34716;
  assign n34718 = pi20 ? n577 : n642;
  assign n34719 = pi20 ? n647 : n1921;
  assign n34720 = pi19 ? n34718 : n34719;
  assign n34721 = pi20 ? n233 : n18756;
  assign n34722 = pi19 ? n34721 : n32;
  assign n34723 = pi18 ? n34720 : n34722;
  assign n34724 = pi17 ? n34717 : n34723;
  assign n34725 = pi16 ? n34705 : n34724;
  assign n34726 = pi15 ? n34714 : n34725;
  assign n34727 = pi14 ? n34703 : n34726;
  assign n34728 = pi20 ? n335 : n8927;
  assign n34729 = pi19 ? n10957 : n34728;
  assign n34730 = pi18 ? n34729 : n34167;
  assign n34731 = pi17 ? n335 : n34730;
  assign n34732 = pi16 ? n3351 : n34731;
  assign n34733 = pi19 ? n8914 : n30698;
  assign n34734 = pi18 ? n335 : n34733;
  assign n34735 = pi19 ? n21154 : n30698;
  assign n34736 = pi18 ? n34735 : n34167;
  assign n34737 = pi17 ? n34734 : n34736;
  assign n34738 = pi16 ? n2035 : n34737;
  assign n34739 = pi15 ? n34732 : n34738;
  assign n34740 = pi19 ? n37 : n11632;
  assign n34741 = pi18 ? n374 : n34740;
  assign n34742 = pi17 ? n32 : n34741;
  assign n34743 = pi20 ? n27730 : n571;
  assign n34744 = pi19 ? n639 : n34743;
  assign n34745 = pi20 ? n610 : n25947;
  assign n34746 = pi19 ? n34745 : n233;
  assign n34747 = pi18 ? n34744 : n34746;
  assign n34748 = pi18 ? n21155 : n34167;
  assign n34749 = pi17 ? n34747 : n34748;
  assign n34750 = pi16 ? n34742 : n34749;
  assign n34751 = pi20 ? n27501 : n363;
  assign n34752 = pi19 ? n22883 : n34751;
  assign n34753 = pi18 ? n34752 : n22156;
  assign n34754 = pi19 ? n25188 : n233;
  assign n34755 = pi18 ? n34754 : n34167;
  assign n34756 = pi17 ? n34753 : n34755;
  assign n34757 = pi16 ? n439 : n34756;
  assign n34758 = pi15 ? n34750 : n34757;
  assign n34759 = pi14 ? n34739 : n34758;
  assign n34760 = pi13 ? n34727 : n34759;
  assign n34761 = pi18 ? n374 : n363;
  assign n34762 = pi17 ? n32 : n34761;
  assign n34763 = pi20 ? n363 : n27796;
  assign n34764 = pi20 ? n25199 : n685;
  assign n34765 = pi19 ? n34763 : n34764;
  assign n34766 = pi18 ? n363 : n34765;
  assign n34767 = pi20 ? n685 : n25199;
  assign n34768 = pi20 ? n18194 : n685;
  assign n34769 = pi19 ? n34767 : n34768;
  assign n34770 = pi20 ? n685 : n11674;
  assign n34771 = pi19 ? n34770 : n32;
  assign n34772 = pi18 ? n34769 : n34771;
  assign n34773 = pi17 ? n34766 : n34772;
  assign n34774 = pi16 ? n34762 : n34773;
  assign n34775 = pi20 ? n18194 : n11674;
  assign n34776 = pi19 ? n34775 : n32;
  assign n34777 = pi18 ? n2731 : n34776;
  assign n34778 = pi17 ? n29350 : n34777;
  assign n34779 = pi16 ? n439 : n34778;
  assign n34780 = pi15 ? n34774 : n34779;
  assign n34781 = pi19 ? n37 : n24866;
  assign n34782 = pi20 ? n24220 : n13398;
  assign n34783 = pi19 ? n34782 : n32;
  assign n34784 = pi18 ? n34781 : n34783;
  assign n34785 = pi17 ? n29350 : n34784;
  assign n34786 = pi16 ? n439 : n34785;
  assign n34787 = pi21 ? n4548 : n99;
  assign n34788 = pi20 ? n99 : n34787;
  assign n34789 = pi19 ? n99 : n34788;
  assign n34790 = pi18 ? n719 : n34789;
  assign n34791 = pi17 ? n32 : n34790;
  assign n34792 = pi20 ? n32788 : n25167;
  assign n34793 = pi21 ? n722 : n4551;
  assign n34794 = pi20 ? n34793 : n363;
  assign n34795 = pi19 ? n34792 : n34794;
  assign n34796 = pi20 ? n32787 : n363;
  assign n34797 = pi20 ? n25167 : n363;
  assign n34798 = pi19 ? n34796 : n34797;
  assign n34799 = pi18 ? n34795 : n34798;
  assign n34800 = pi20 ? n24220 : n12514;
  assign n34801 = pi19 ? n34800 : n32;
  assign n34802 = pi18 ? n363 : n34801;
  assign n34803 = pi17 ? n34799 : n34802;
  assign n34804 = pi16 ? n34791 : n34803;
  assign n34805 = pi15 ? n34786 : n34804;
  assign n34806 = pi14 ? n34780 : n34805;
  assign n34807 = pi18 ? n966 : n363;
  assign n34808 = pi17 ? n32 : n34807;
  assign n34809 = pi20 ? n24220 : n6935;
  assign n34810 = pi19 ? n34809 : n32;
  assign n34811 = pi18 ? n363 : n34810;
  assign n34812 = pi17 ? n363 : n34811;
  assign n34813 = pi16 ? n34808 : n34812;
  assign n34814 = pi20 ? n363 : n3210;
  assign n34815 = pi19 ? n34814 : n32;
  assign n34816 = pi18 ? n363 : n34815;
  assign n34817 = pi17 ? n363 : n34816;
  assign n34818 = pi16 ? n21219 : n34817;
  assign n34819 = pi15 ? n34813 : n34818;
  assign n34820 = pi20 ? n25199 : n2638;
  assign n34821 = pi19 ? n34820 : n32;
  assign n34822 = pi18 ? n363 : n34821;
  assign n34823 = pi17 ? n363 : n34822;
  assign n34824 = pi16 ? n26062 : n34823;
  assign n34825 = pi22 ? n26056 : n157;
  assign n34826 = pi21 ? n34825 : n157;
  assign n34827 = pi20 ? n32 : n34826;
  assign n34828 = pi19 ? n32 : n34827;
  assign n34829 = pi18 ? n34828 : n157;
  assign n34830 = pi17 ? n32 : n34829;
  assign n34831 = pi21 ? n5054 : n157;
  assign n34832 = pi20 ? n157 : n34831;
  assign n34833 = pi22 ? n157 : n363;
  assign n34834 = pi21 ? n157 : n34833;
  assign n34835 = pi20 ? n34831 : n34834;
  assign n34836 = pi19 ? n34832 : n34835;
  assign n34837 = pi21 ? n34833 : n157;
  assign n34838 = pi21 ? n34833 : n5054;
  assign n34839 = pi20 ? n34837 : n34838;
  assign n34840 = pi21 ? n157 : n5054;
  assign n34841 = pi21 ? n363 : n34833;
  assign n34842 = pi20 ? n34840 : n34841;
  assign n34843 = pi19 ? n34839 : n34842;
  assign n34844 = pi18 ? n34836 : n34843;
  assign n34845 = pi20 ? n34831 : n34838;
  assign n34846 = pi21 ? n157 : n363;
  assign n34847 = pi20 ? n34846 : n363;
  assign n34848 = pi19 ? n34845 : n34847;
  assign n34849 = pi18 ? n34848 : n19946;
  assign n34850 = pi17 ? n34844 : n34849;
  assign n34851 = pi16 ? n34830 : n34850;
  assign n34852 = pi15 ? n34824 : n34851;
  assign n34853 = pi14 ? n34819 : n34852;
  assign n34854 = pi13 ? n34806 : n34853;
  assign n34855 = pi12 ? n34760 : n34854;
  assign n34856 = pi11 ? n34689 : n34855;
  assign n34857 = pi10 ? n34510 : n34856;
  assign n34858 = pi09 ? n34274 : n34857;
  assign n34859 = pi18 ? n30119 : n20563;
  assign n34860 = pi17 ? n32 : n34859;
  assign n34861 = pi18 ? n33966 : n34251;
  assign n34862 = pi17 ? n34861 : n34254;
  assign n34863 = pi16 ? n34860 : n34862;
  assign n34864 = pi15 ? n32 : n34863;
  assign n34865 = pi19 ? n20563 : n32876;
  assign n34866 = pi18 ? n30119 : n34865;
  assign n34867 = pi17 ? n32 : n34866;
  assign n34868 = pi16 ? n34867 : n34266;
  assign n34869 = pi19 ? n20563 : n31221;
  assign n34870 = pi18 ? n30119 : n34869;
  assign n34871 = pi17 ? n32 : n34870;
  assign n34872 = pi16 ? n34871 : n34266;
  assign n34873 = pi15 ? n34868 : n34872;
  assign n34874 = pi14 ? n34864 : n34873;
  assign n34875 = pi13 ? n32 : n34874;
  assign n34876 = pi12 ? n32 : n34875;
  assign n34877 = pi11 ? n32 : n34876;
  assign n34878 = pi10 ? n32 : n34877;
  assign n34879 = pi18 ? n31265 : n33823;
  assign n34880 = pi17 ? n32 : n34879;
  assign n34881 = pi16 ? n34880 : n34281;
  assign n34882 = pi15 ? n34881 : n34293;
  assign n34883 = pi18 ? n31938 : n33260;
  assign n34884 = pi17 ? n32 : n34883;
  assign n34885 = pi16 ? n34884 : n34314;
  assign n34886 = pi15 ? n34304 : n34885;
  assign n34887 = pi14 ? n34882 : n34886;
  assign n34888 = pi18 ? n31315 : n32275;
  assign n34889 = pi17 ? n32 : n34888;
  assign n34890 = pi16 ? n34889 : n34325;
  assign n34891 = pi19 ? n20563 : n33949;
  assign n34892 = pi18 ? n31315 : n34891;
  assign n34893 = pi17 ? n32 : n34892;
  assign n34894 = pi19 ? n9814 : n6186;
  assign n34895 = pi18 ? n37 : n34894;
  assign n34896 = pi17 ? n37 : n34895;
  assign n34897 = pi16 ? n34893 : n34896;
  assign n34898 = pi15 ? n34890 : n34897;
  assign n34899 = pi19 ? n20563 : n33965;
  assign n34900 = pi18 ? n31315 : n34899;
  assign n34901 = pi17 ? n32 : n34900;
  assign n34902 = pi19 ? n8765 : n6186;
  assign n34903 = pi18 ? n34337 : n34902;
  assign n34904 = pi17 ? n37 : n34903;
  assign n34905 = pi16 ? n34901 : n34904;
  assign n34906 = pi21 ? n26965 : n32;
  assign n34907 = pi20 ? n34906 : n32;
  assign n34908 = pi19 ? n9769 : n34907;
  assign n34909 = pi18 ? n34343 : n34908;
  assign n34910 = pi17 ? n34342 : n34909;
  assign n34911 = pi16 ? n34335 : n34910;
  assign n34912 = pi15 ? n34905 : n34911;
  assign n34913 = pi14 ? n34898 : n34912;
  assign n34914 = pi13 ? n34887 : n34913;
  assign n34915 = pi19 ? n8765 : n34907;
  assign n34916 = pi18 ? n34354 : n34915;
  assign n34917 = pi17 ? n37 : n34916;
  assign n34918 = pi16 ? n33883 : n34917;
  assign n34919 = pi21 ? n20563 : n30195;
  assign n34920 = pi20 ? n20563 : n34919;
  assign n34921 = pi19 ? n34920 : n37;
  assign n34922 = pi18 ? n31315 : n34921;
  assign n34923 = pi17 ? n32 : n34922;
  assign n34924 = pi21 ? n26972 : n32;
  assign n34925 = pi20 ? n34924 : n32;
  assign n34926 = pi19 ? n8765 : n34925;
  assign n34927 = pi18 ? n34361 : n34926;
  assign n34928 = pi17 ? n37 : n34927;
  assign n34929 = pi16 ? n34923 : n34928;
  assign n34930 = pi15 ? n34918 : n34929;
  assign n34931 = pi20 ? n19523 : n32;
  assign n34932 = pi19 ? n34369 : n34931;
  assign n34933 = pi18 ? n34361 : n34932;
  assign n34934 = pi17 ? n37 : n34933;
  assign n34935 = pi16 ? n34360 : n34934;
  assign n34936 = pi19 ? n17204 : n6215;
  assign n34937 = pi18 ? n37 : n34936;
  assign n34938 = pi17 ? n37 : n34937;
  assign n34939 = pi16 ? n34360 : n34938;
  assign n34940 = pi15 ? n34935 : n34939;
  assign n34941 = pi14 ? n34930 : n34940;
  assign n34942 = pi22 ? n363 : n317;
  assign n34943 = pi21 ? n34942 : n32;
  assign n34944 = pi20 ? n34943 : n32;
  assign n34945 = pi19 ? n12628 : n34944;
  assign n34946 = pi18 ? n37 : n34945;
  assign n34947 = pi17 ? n37 : n34946;
  assign n34948 = pi16 ? n33332 : n34947;
  assign n34949 = pi19 ? n31914 : n37;
  assign n34950 = pi18 ? n31938 : n34949;
  assign n34951 = pi17 ? n32 : n34950;
  assign n34952 = pi21 ? n11928 : n32;
  assign n34953 = pi20 ? n34952 : n32;
  assign n34954 = pi19 ? n25087 : n34953;
  assign n34955 = pi18 ? n37 : n34954;
  assign n34956 = pi17 ? n37 : n34955;
  assign n34957 = pi16 ? n34951 : n34956;
  assign n34958 = pi15 ? n34948 : n34957;
  assign n34959 = pi22 ? n456 : n532;
  assign n34960 = pi21 ? n34959 : n32;
  assign n34961 = pi20 ? n34960 : n32;
  assign n34962 = pi19 ? n37 : n34961;
  assign n34963 = pi18 ? n37 : n34962;
  assign n34964 = pi17 ? n37 : n34963;
  assign n34965 = pi16 ? n33978 : n34964;
  assign n34966 = pi18 ? n31938 : n31300;
  assign n34967 = pi17 ? n32 : n34966;
  assign n34968 = pi16 ? n34967 : n34407;
  assign n34969 = pi15 ? n34965 : n34968;
  assign n34970 = pi14 ? n34958 : n34969;
  assign n34971 = pi13 ? n34941 : n34970;
  assign n34972 = pi12 ? n34914 : n34971;
  assign n34973 = pi19 ? n34413 : n15447;
  assign n34974 = pi18 ? n37 : n34973;
  assign n34975 = pi17 ? n37 : n34974;
  assign n34976 = pi16 ? n34967 : n34975;
  assign n34977 = pi19 ? n34423 : n5760;
  assign n34978 = pi18 ? n34422 : n34977;
  assign n34979 = pi17 ? n37 : n34978;
  assign n34980 = pi16 ? n32936 : n34979;
  assign n34981 = pi15 ? n34976 : n34980;
  assign n34982 = pi20 ? n649 : n24865;
  assign n34983 = pi19 ? n34982 : n5773;
  assign n34984 = pi18 ? n37 : n34983;
  assign n34985 = pi17 ? n37 : n34984;
  assign n34986 = pi16 ? n32404 : n34985;
  assign n34987 = pi15 ? n34432 : n34986;
  assign n34988 = pi14 ? n34981 : n34987;
  assign n34989 = pi21 ? n30866 : n30867;
  assign n34990 = pi20 ? n32 : n34989;
  assign n34991 = pi19 ? n32 : n34990;
  assign n34992 = pi18 ? n34991 : n37;
  assign n34993 = pi17 ? n32 : n34992;
  assign n34994 = pi16 ? n34993 : n34449;
  assign n34995 = pi21 ? n30866 : n30195;
  assign n34996 = pi20 ? n32 : n34995;
  assign n34997 = pi19 ? n32 : n34996;
  assign n34998 = pi18 ? n34997 : n37;
  assign n34999 = pi17 ? n32 : n34998;
  assign n35000 = pi16 ? n34999 : n34453;
  assign n35001 = pi15 ? n34994 : n35000;
  assign n35002 = pi21 ? n32966 : n30843;
  assign n35003 = pi20 ? n32 : n35002;
  assign n35004 = pi19 ? n32 : n35003;
  assign n35005 = pi18 ? n35004 : n37;
  assign n35006 = pi17 ? n32 : n35005;
  assign n35007 = pi16 ? n35006 : n34458;
  assign n35008 = pi15 ? n35007 : n34459;
  assign n35009 = pi14 ? n35001 : n35008;
  assign n35010 = pi13 ? n34988 : n35009;
  assign n35011 = pi22 ? n30865 : n37;
  assign n35012 = pi21 ? n35011 : n37;
  assign n35013 = pi20 ? n32 : n35012;
  assign n35014 = pi19 ? n32 : n35013;
  assign n35015 = pi18 ? n35014 : n37;
  assign n35016 = pi17 ? n32 : n35015;
  assign n35017 = pi21 ? n748 : n32;
  assign n35018 = pi20 ? n35017 : n32;
  assign n35019 = pi19 ? n5029 : n35018;
  assign n35020 = pi18 ? n37 : n35019;
  assign n35021 = pi17 ? n37 : n35020;
  assign n35022 = pi16 ? n35016 : n35021;
  assign n35023 = pi16 ? n34016 : n34469;
  assign n35024 = pi15 ? n35022 : n35023;
  assign n35025 = pi14 ? n35024 : n34475;
  assign n35026 = pi19 ? n34479 : n2639;
  assign n35027 = pi18 ? n37 : n35026;
  assign n35028 = pi17 ? n37 : n35027;
  assign n35029 = pi16 ? n439 : n35028;
  assign n35030 = pi15 ? n34483 : n35029;
  assign n35031 = pi19 ? n157 : n2639;
  assign n35032 = pi18 ? n34493 : n35031;
  assign n35033 = pi17 ? n34489 : n35032;
  assign n35034 = pi16 ? n439 : n35033;
  assign n35035 = pi19 ? n157 : n2654;
  assign n35036 = pi18 ? n34502 : n35035;
  assign n35037 = pi17 ? n34500 : n35036;
  assign n35038 = pi16 ? n439 : n35037;
  assign n35039 = pi15 ? n35034 : n35038;
  assign n35040 = pi14 ? n35030 : n35039;
  assign n35041 = pi13 ? n35025 : n35040;
  assign n35042 = pi12 ? n35010 : n35041;
  assign n35043 = pi11 ? n34972 : n35042;
  assign n35044 = pi18 ? n34519 : n35035;
  assign n35045 = pi17 ? n34518 : n35044;
  assign n35046 = pi16 ? n439 : n35045;
  assign n35047 = pi19 ? n9035 : n2654;
  assign n35048 = pi18 ? n34531 : n35047;
  assign n35049 = pi17 ? n34527 : n35048;
  assign n35050 = pi16 ? n439 : n35049;
  assign n35051 = pi15 ? n35046 : n35050;
  assign n35052 = pi19 ? n34539 : n2654;
  assign n35053 = pi18 ? n34536 : n35052;
  assign n35054 = pi17 ? n99 : n35053;
  assign n35055 = pi16 ? n201 : n35054;
  assign n35056 = pi19 ? n34544 : n2680;
  assign n35057 = pi18 ? n99 : n35056;
  assign n35058 = pi17 ? n99 : n35057;
  assign n35059 = pi16 ? n25610 : n35058;
  assign n35060 = pi15 ? n35055 : n35059;
  assign n35061 = pi14 ? n35051 : n35060;
  assign n35062 = pi20 ? n99 : n20468;
  assign n35063 = pi19 ? n35062 : n1823;
  assign n35064 = pi18 ? n99 : n35063;
  assign n35065 = pi17 ? n99 : n35064;
  assign n35066 = pi16 ? n801 : n35065;
  assign n35067 = pi21 ? n99 : n3207;
  assign n35068 = pi20 ? n99 : n35067;
  assign n35069 = pi19 ? n35068 : n2702;
  assign n35070 = pi18 ? n99 : n35069;
  assign n35071 = pi17 ? n99 : n35070;
  assign n35072 = pi16 ? n23698 : n35071;
  assign n35073 = pi15 ? n35066 : n35072;
  assign n35074 = pi19 ? n34577 : n1823;
  assign n35075 = pi18 ? n34576 : n35074;
  assign n35076 = pi17 ? n34573 : n35075;
  assign n35077 = pi16 ? n34569 : n35076;
  assign n35078 = pi15 ? n35077 : n34593;
  assign n35079 = pi14 ? n35073 : n35078;
  assign n35080 = pi13 ? n35061 : n35079;
  assign n35081 = pi22 ? n204 : n31630;
  assign n35082 = pi21 ? n204 : n35081;
  assign n35083 = pi20 ? n204 : n35082;
  assign n35084 = pi19 ? n35083 : n32;
  assign n35085 = pi18 ? n34608 : n35084;
  assign n35086 = pi17 ? n34606 : n35085;
  assign n35087 = pi16 ? n439 : n35086;
  assign n35088 = pi15 ? n34603 : n35087;
  assign n35089 = pi21 ? n204 : n10106;
  assign n35090 = pi20 ? n2316 : n35089;
  assign n35091 = pi19 ? n35090 : n32;
  assign n35092 = pi18 ? n34623 : n35091;
  assign n35093 = pi17 ? n34621 : n35092;
  assign n35094 = pi16 ? n439 : n35093;
  assign n35095 = pi18 ? n204 : n26998;
  assign n35096 = pi17 ? n34631 : n35095;
  assign n35097 = pi16 ? n439 : n35096;
  assign n35098 = pi15 ? n35094 : n35097;
  assign n35099 = pi14 ? n35088 : n35098;
  assign n35100 = pi21 ? n204 : n15439;
  assign n35101 = pi20 ? n204 : n35100;
  assign n35102 = pi19 ? n35101 : n32;
  assign n35103 = pi18 ? n204 : n35102;
  assign n35104 = pi17 ? n34643 : n35103;
  assign n35105 = pi16 ? n34640 : n35104;
  assign n35106 = pi15 ? n35105 : n34658;
  assign n35107 = pi21 ? n916 : n19337;
  assign n35108 = pi22 ? n233 : n1038;
  assign n35109 = pi21 ? n35108 : n7002;
  assign n35110 = pi20 ? n35107 : n35109;
  assign n35111 = pi19 ? n35110 : n32;
  assign n35112 = pi18 ? n34667 : n35111;
  assign n35113 = pi17 ? n34664 : n35112;
  assign n35114 = pi16 ? n439 : n35113;
  assign n35115 = pi15 ? n35114 : n34685;
  assign n35116 = pi14 ? n35106 : n35115;
  assign n35117 = pi13 ? n35099 : n35116;
  assign n35118 = pi12 ? n35080 : n35117;
  assign n35119 = pi20 ? n233 : n19361;
  assign n35120 = pi19 ? n35119 : n32;
  assign n35121 = pi18 ? n34720 : n35120;
  assign n35122 = pi17 ? n34717 : n35121;
  assign n35123 = pi16 ? n34705 : n35122;
  assign n35124 = pi15 ? n34714 : n35123;
  assign n35125 = pi14 ? n34703 : n35124;
  assign n35126 = pi20 ? n233 : n24432;
  assign n35127 = pi19 ? n35126 : n32;
  assign n35128 = pi18 ? n34729 : n35127;
  assign n35129 = pi17 ? n335 : n35128;
  assign n35130 = pi16 ? n3351 : n35129;
  assign n35131 = pi18 ? n34735 : n35127;
  assign n35132 = pi17 ? n34734 : n35131;
  assign n35133 = pi16 ? n2035 : n35132;
  assign n35134 = pi15 ? n35130 : n35133;
  assign n35135 = pi18 ? n21155 : n34722;
  assign n35136 = pi17 ? n34747 : n35135;
  assign n35137 = pi16 ? n34742 : n35136;
  assign n35138 = pi18 ? n34754 : n34722;
  assign n35139 = pi17 ? n34753 : n35138;
  assign n35140 = pi16 ? n439 : n35139;
  assign n35141 = pi15 ? n35137 : n35140;
  assign n35142 = pi14 ? n35134 : n35141;
  assign n35143 = pi13 ? n35125 : n35142;
  assign n35144 = pi20 ? n25199 : n4116;
  assign n35145 = pi19 ? n35144 : n32;
  assign n35146 = pi18 ? n363 : n35145;
  assign n35147 = pi17 ? n363 : n35146;
  assign n35148 = pi16 ? n26062 : n35147;
  assign n35149 = pi18 ? n34848 : n20419;
  assign n35150 = pi17 ? n34844 : n35149;
  assign n35151 = pi16 ? n34830 : n35150;
  assign n35152 = pi15 ? n35148 : n35151;
  assign n35153 = pi14 ? n34819 : n35152;
  assign n35154 = pi13 ? n34806 : n35153;
  assign n35155 = pi12 ? n35143 : n35154;
  assign n35156 = pi11 ? n35118 : n35155;
  assign n35157 = pi10 ? n35043 : n35156;
  assign n35158 = pi09 ? n34878 : n35157;
  assign n35159 = pi08 ? n34858 : n35158;
  assign n35160 = pi19 ? n31914 : n34261;
  assign n35161 = pi18 ? n35160 : n99;
  assign n35162 = pi21 ? n27251 : n32;
  assign n35163 = pi20 ? n35162 : n32;
  assign n35164 = pi19 ? n99 : n35163;
  assign n35165 = pi18 ? n99 : n35164;
  assign n35166 = pi17 ? n35161 : n35165;
  assign n35167 = pi16 ? n34860 : n35166;
  assign n35168 = pi15 ? n32 : n35167;
  assign n35169 = pi19 ? n30097 : n34261;
  assign n35170 = pi18 ? n35169 : n99;
  assign n35171 = pi20 ? n19760 : n32;
  assign n35172 = pi19 ? n99 : n35171;
  assign n35173 = pi18 ? n99 : n35172;
  assign n35174 = pi17 ? n35170 : n35173;
  assign n35175 = pi16 ? n34860 : n35174;
  assign n35176 = pi17 ? n34263 : n35173;
  assign n35177 = pi16 ? n34860 : n35176;
  assign n35178 = pi15 ? n35175 : n35177;
  assign n35179 = pi14 ? n35168 : n35178;
  assign n35180 = pi13 ? n32 : n35179;
  assign n35181 = pi12 ? n32 : n35180;
  assign n35182 = pi11 ? n32 : n35181;
  assign n35183 = pi10 ? n32 : n35182;
  assign n35184 = pi18 ? n31265 : n34258;
  assign n35185 = pi17 ? n32 : n35184;
  assign n35186 = pi23 ? n3491 : n586;
  assign n35187 = pi22 ? n99 : n35186;
  assign n35188 = pi21 ? n35187 : n32;
  assign n35189 = pi20 ? n35188 : n32;
  assign n35190 = pi19 ? n15543 : n35189;
  assign n35191 = pi18 ? n99 : n35190;
  assign n35192 = pi17 ? n34278 : n35191;
  assign n35193 = pi16 ? n35185 : n35192;
  assign n35194 = pi18 ? n31265 : n34865;
  assign n35195 = pi17 ? n32 : n35194;
  assign n35196 = pi19 ? n17013 : n37;
  assign n35197 = pi18 ? n35196 : n18854;
  assign n35198 = pi23 ? n11962 : n5630;
  assign n35199 = pi22 ? n99 : n35198;
  assign n35200 = pi21 ? n35199 : n32;
  assign n35201 = pi20 ? n35200 : n32;
  assign n35202 = pi19 ? n99 : n35201;
  assign n35203 = pi18 ? n99 : n35202;
  assign n35204 = pi17 ? n35197 : n35203;
  assign n35205 = pi16 ? n35195 : n35204;
  assign n35206 = pi15 ? n35193 : n35205;
  assign n35207 = pi18 ? n31265 : n34869;
  assign n35208 = pi17 ? n32 : n35207;
  assign n35209 = pi20 ? n37 : n226;
  assign n35210 = pi19 ? n35209 : n99;
  assign n35211 = pi18 ? n35210 : n99;
  assign n35212 = pi22 ? n99 : n24295;
  assign n35213 = pi21 ? n35212 : n32;
  assign n35214 = pi20 ? n35213 : n32;
  assign n35215 = pi19 ? n99 : n35214;
  assign n35216 = pi18 ? n99 : n35215;
  assign n35217 = pi17 ? n35211 : n35216;
  assign n35218 = pi16 ? n35208 : n35217;
  assign n35219 = pi18 ? n31315 : n33245;
  assign n35220 = pi17 ? n32 : n35219;
  assign n35221 = pi22 ? n37 : n17582;
  assign n35222 = pi21 ? n35221 : n32;
  assign n35223 = pi20 ? n35222 : n32;
  assign n35224 = pi19 ? n37 : n35223;
  assign n35225 = pi18 ? n37 : n35224;
  assign n35226 = pi17 ? n37 : n35225;
  assign n35227 = pi16 ? n35220 : n35226;
  assign n35228 = pi15 ? n35218 : n35227;
  assign n35229 = pi14 ? n35206 : n35228;
  assign n35230 = pi22 ? n37 : n30195;
  assign n35231 = pi21 ? n35230 : n37;
  assign n35232 = pi20 ? n20563 : n35231;
  assign n35233 = pi19 ? n20563 : n35232;
  assign n35234 = pi18 ? n31315 : n35233;
  assign n35235 = pi17 ? n32 : n35234;
  assign n35236 = pi22 ? n37 : n31329;
  assign n35237 = pi21 ? n35236 : n32;
  assign n35238 = pi20 ? n35237 : n32;
  assign n35239 = pi19 ? n37 : n35238;
  assign n35240 = pi18 ? n37 : n35239;
  assign n35241 = pi17 ? n37 : n35240;
  assign n35242 = pi16 ? n35235 : n35241;
  assign n35243 = pi18 ? n31315 : n34295;
  assign n35244 = pi17 ? n32 : n35243;
  assign n35245 = pi16 ? n35244 : n34896;
  assign n35246 = pi15 ? n35242 : n35245;
  assign n35247 = pi19 ? n37 : n9769;
  assign n35248 = pi18 ? n37 : n35247;
  assign n35249 = pi18 ? n139 : n34902;
  assign n35250 = pi17 ? n35248 : n35249;
  assign n35251 = pi16 ? n34306 : n35250;
  assign n35252 = pi20 ? n3086 : n939;
  assign n35253 = pi19 ? n37 : n35252;
  assign n35254 = pi18 ? n37 : n35253;
  assign n35255 = pi20 ? n19516 : n32;
  assign n35256 = pi19 ? n9769 : n35255;
  assign n35257 = pi18 ? n139 : n35256;
  assign n35258 = pi17 ? n35254 : n35257;
  assign n35259 = pi16 ? n34319 : n35258;
  assign n35260 = pi15 ? n35251 : n35259;
  assign n35261 = pi14 ? n35246 : n35260;
  assign n35262 = pi13 ? n35229 : n35261;
  assign n35263 = pi20 ? n139 : n3083;
  assign n35264 = pi19 ? n9765 : n35263;
  assign n35265 = pi19 ? n8765 : n35255;
  assign n35266 = pi18 ? n35264 : n35265;
  assign n35267 = pi17 ? n37 : n35266;
  assign n35268 = pi16 ? n34889 : n35267;
  assign n35269 = pi20 ? n139 : n9354;
  assign n35270 = pi19 ? n30265 : n35269;
  assign n35271 = pi19 ? n4733 : n34931;
  assign n35272 = pi18 ? n35270 : n35271;
  assign n35273 = pi17 ? n37 : n35272;
  assign n35274 = pi16 ? n34901 : n35273;
  assign n35275 = pi15 ? n35268 : n35274;
  assign n35276 = pi19 ? n37 : n34336;
  assign n35277 = pi20 ? n942 : n34368;
  assign n35278 = pi19 ? n35277 : n34931;
  assign n35279 = pi18 ? n35276 : n35278;
  assign n35280 = pi17 ? n37 : n35279;
  assign n35281 = pi16 ? n34889 : n35280;
  assign n35282 = pi18 ? n31938 : n33299;
  assign n35283 = pi17 ? n32 : n35282;
  assign n35284 = pi16 ? n35283 : n34938;
  assign n35285 = pi15 ? n35281 : n35284;
  assign n35286 = pi14 ? n35275 : n35285;
  assign n35287 = pi16 ? n34923 : n34947;
  assign n35288 = pi22 ? n5011 : n2468;
  assign n35289 = pi21 ? n35288 : n32;
  assign n35290 = pi20 ? n35289 : n32;
  assign n35291 = pi19 ? n3332 : n35290;
  assign n35292 = pi18 ? n37 : n35291;
  assign n35293 = pi17 ? n37 : n35292;
  assign n35294 = pi16 ? n34360 : n35293;
  assign n35295 = pi15 ? n35287 : n35294;
  assign n35296 = pi19 ? n37 : n8948;
  assign n35297 = pi18 ? n37 : n35296;
  assign n35298 = pi17 ? n37 : n35297;
  assign n35299 = pi16 ? n34360 : n35298;
  assign n35300 = pi19 ? n31904 : n37;
  assign n35301 = pi18 ? n31315 : n35300;
  assign n35302 = pi17 ? n32 : n35301;
  assign n35303 = pi19 ? n7706 : n9442;
  assign n35304 = pi18 ? n37 : n35303;
  assign n35305 = pi17 ? n37 : n35304;
  assign n35306 = pi16 ? n35302 : n35305;
  assign n35307 = pi15 ? n35299 : n35306;
  assign n35308 = pi14 ? n35295 : n35307;
  assign n35309 = pi13 ? n35286 : n35308;
  assign n35310 = pi12 ? n35262 : n35309;
  assign n35311 = pi20 ? n577 : n16530;
  assign n35312 = pi19 ? n35311 : n6985;
  assign n35313 = pi18 ? n14149 : n35312;
  assign n35314 = pi17 ? n37 : n35313;
  assign n35315 = pi16 ? n32379 : n35314;
  assign n35316 = pi21 ? n20563 : n31200;
  assign n35317 = pi20 ? n35316 : n37;
  assign n35318 = pi19 ? n35317 : n37;
  assign n35319 = pi18 ? n31315 : n35318;
  assign n35320 = pi17 ? n32 : n35319;
  assign n35321 = pi19 ? n6373 : n8802;
  assign n35322 = pi20 ? n577 : n571;
  assign n35323 = pi19 ? n35322 : n6985;
  assign n35324 = pi18 ? n35321 : n35323;
  assign n35325 = pi17 ? n37 : n35324;
  assign n35326 = pi16 ? n35320 : n35325;
  assign n35327 = pi15 ? n35315 : n35326;
  assign n35328 = pi18 ? n31938 : n33976;
  assign n35329 = pi17 ? n32 : n35328;
  assign n35330 = pi19 ? n7676 : n37;
  assign n35331 = pi19 ? n10681 : n6985;
  assign n35332 = pi18 ? n35330 : n35331;
  assign n35333 = pi17 ? n37 : n35332;
  assign n35334 = pi16 ? n35329 : n35333;
  assign n35335 = pi22 ? n673 : n688;
  assign n35336 = pi21 ? n35335 : n32;
  assign n35337 = pi20 ? n35336 : n32;
  assign n35338 = pi19 ? n24866 : n35337;
  assign n35339 = pi18 ? n37 : n35338;
  assign n35340 = pi17 ? n37 : n35339;
  assign n35341 = pi16 ? n35329 : n35340;
  assign n35342 = pi15 ? n35334 : n35341;
  assign n35343 = pi14 ? n35327 : n35342;
  assign n35344 = pi19 ? n22883 : n9473;
  assign n35345 = pi18 ? n37 : n35344;
  assign n35346 = pi17 ? n37 : n35345;
  assign n35347 = pi16 ? n32926 : n35346;
  assign n35348 = pi19 ? n6403 : n8959;
  assign n35349 = pi18 ? n37 : n35348;
  assign n35350 = pi17 ? n37 : n35349;
  assign n35351 = pi16 ? n33374 : n35350;
  assign n35352 = pi15 ? n35347 : n35351;
  assign n35353 = pi19 ? n37 : n8959;
  assign n35354 = pi18 ? n37 : n35353;
  assign n35355 = pi17 ? n37 : n35354;
  assign n35356 = pi16 ? n32926 : n35355;
  assign n35357 = pi19 ? n6403 : n34446;
  assign n35358 = pi18 ? n37 : n35357;
  assign n35359 = pi17 ? n37 : n35358;
  assign n35360 = pi16 ? n32936 : n35359;
  assign n35361 = pi15 ? n35356 : n35360;
  assign n35362 = pi14 ? n35352 : n35361;
  assign n35363 = pi13 ? n35343 : n35362;
  assign n35364 = pi19 ? n5029 : n34446;
  assign n35365 = pi18 ? n37 : n35364;
  assign n35366 = pi17 ? n37 : n35365;
  assign n35367 = pi16 ? n31317 : n35366;
  assign n35368 = pi19 ? n6403 : n7725;
  assign n35369 = pi18 ? n37 : n35368;
  assign n35370 = pi17 ? n37 : n35369;
  assign n35371 = pi16 ? n33409 : n35370;
  assign n35372 = pi15 ? n35367 : n35371;
  assign n35373 = pi19 ? n8743 : n7725;
  assign n35374 = pi18 ? n37 : n35373;
  assign n35375 = pi17 ? n37 : n35374;
  assign n35376 = pi16 ? n33409 : n35375;
  assign n35377 = pi19 ? n37 : n19091;
  assign n35378 = pi18 ? n37 : n35377;
  assign n35379 = pi21 ? n6401 : n37;
  assign n35380 = pi20 ? n35379 : n37;
  assign n35381 = pi19 ? n15174 : n35380;
  assign n35382 = pi19 ? n8802 : n3211;
  assign n35383 = pi18 ? n35381 : n35382;
  assign n35384 = pi17 ? n35378 : n35383;
  assign n35385 = pi16 ? n33409 : n35384;
  assign n35386 = pi15 ? n35376 : n35385;
  assign n35387 = pi14 ? n35372 : n35386;
  assign n35388 = pi21 ? n32427 : n30843;
  assign n35389 = pi20 ? n32 : n35388;
  assign n35390 = pi19 ? n32 : n35389;
  assign n35391 = pi18 ? n35390 : n37;
  assign n35392 = pi17 ? n32 : n35391;
  assign n35393 = pi19 ? n34479 : n3211;
  assign n35394 = pi18 ? n37 : n35393;
  assign n35395 = pi17 ? n37 : n35394;
  assign n35396 = pi16 ? n35392 : n35395;
  assign n35397 = pi20 ? n37 : n19934;
  assign n35398 = pi19 ? n35397 : n2639;
  assign n35399 = pi18 ? n37 : n35398;
  assign n35400 = pi17 ? n37 : n35399;
  assign n35401 = pi16 ? n34444 : n35400;
  assign n35402 = pi15 ? n35396 : n35401;
  assign n35403 = pi18 ? n32413 : n18519;
  assign n35404 = pi17 ? n32 : n35403;
  assign n35405 = pi20 ? n23939 : n24502;
  assign n35406 = pi19 ? n18522 : n35405;
  assign n35407 = pi22 ? n889 : n112;
  assign n35408 = pi21 ? n22379 : n35407;
  assign n35409 = pi21 ? n8654 : n23932;
  assign n35410 = pi20 ? n35408 : n35409;
  assign n35411 = pi21 ? n5877 : n23932;
  assign n35412 = pi19 ? n35410 : n35411;
  assign n35413 = pi18 ? n35406 : n35412;
  assign n35414 = pi21 ? n22379 : n157;
  assign n35415 = pi21 ? n157 : n24501;
  assign n35416 = pi20 ? n35414 : n35415;
  assign n35417 = pi21 ? n23932 : n157;
  assign n35418 = pi20 ? n28939 : n35417;
  assign n35419 = pi19 ? n35416 : n35418;
  assign n35420 = pi18 ? n35419 : n35035;
  assign n35421 = pi17 ? n35413 : n35420;
  assign n35422 = pi16 ? n35404 : n35421;
  assign n35423 = pi18 ? n157 : n35035;
  assign n35424 = pi17 ? n34500 : n35423;
  assign n35425 = pi16 ? n32014 : n35424;
  assign n35426 = pi15 ? n35422 : n35425;
  assign n35427 = pi14 ? n35402 : n35426;
  assign n35428 = pi13 ? n35387 : n35427;
  assign n35429 = pi12 ? n35363 : n35428;
  assign n35430 = pi11 ? n35310 : n35429;
  assign n35431 = pi20 ? n15263 : n3039;
  assign n35432 = pi21 ? n157 : n218;
  assign n35433 = pi20 ? n35432 : n6508;
  assign n35434 = pi19 ? n35431 : n35433;
  assign n35435 = pi18 ? n34512 : n35434;
  assign n35436 = pi20 ? n18265 : n157;
  assign n35437 = pi19 ? n19137 : n35436;
  assign n35438 = pi18 ? n35437 : n35031;
  assign n35439 = pi17 ? n35435 : n35438;
  assign n35440 = pi16 ? n30201 : n35439;
  assign n35441 = pi18 ? n34262 : n34277;
  assign n35442 = pi21 ? n157 : n181;
  assign n35443 = pi20 ? n99 : n35442;
  assign n35444 = pi19 ? n35443 : n7845;
  assign n35445 = pi18 ? n35444 : n35047;
  assign n35446 = pi17 ? n35441 : n35445;
  assign n35447 = pi16 ? n439 : n35446;
  assign n35448 = pi15 ? n35440 : n35447;
  assign n35449 = pi20 ? n99 : n19171;
  assign n35450 = pi19 ? n14285 : n35449;
  assign n35451 = pi20 ? n9752 : n34538;
  assign n35452 = pi19 ? n35451 : n2654;
  assign n35453 = pi18 ? n35450 : n35452;
  assign n35454 = pi17 ? n99 : n35453;
  assign n35455 = pi16 ? n29201 : n35454;
  assign n35456 = pi20 ? n19208 : n9747;
  assign n35457 = pi19 ? n35456 : n2654;
  assign n35458 = pi18 ? n99 : n35457;
  assign n35459 = pi17 ? n99 : n35458;
  assign n35460 = pi16 ? n23698 : n35459;
  assign n35461 = pi15 ? n35455 : n35460;
  assign n35462 = pi14 ? n35448 : n35461;
  assign n35463 = pi20 ? n22965 : n20930;
  assign n35464 = pi19 ? n35463 : n2654;
  assign n35465 = pi18 ? n99 : n35464;
  assign n35466 = pi17 ? n99 : n35465;
  assign n35467 = pi16 ? n186 : n35466;
  assign n35468 = pi20 ? n99 : n24957;
  assign n35469 = pi19 ? n99 : n35468;
  assign n35470 = pi19 ? n316 : n2654;
  assign n35471 = pi18 ? n35469 : n35470;
  assign n35472 = pi17 ? n99 : n35471;
  assign n35473 = pi16 ? n23698 : n35472;
  assign n35474 = pi15 ? n35467 : n35473;
  assign n35475 = pi18 ? n1821 : n35470;
  assign n35476 = pi17 ? n22747 : n35475;
  assign n35477 = pi16 ? n439 : n35476;
  assign n35478 = pi20 ? n976 : n34587;
  assign n35479 = pi19 ? n1022 : n35478;
  assign n35480 = pi21 ? n10084 : n316;
  assign n35481 = pi20 ? n35480 : n316;
  assign n35482 = pi20 ? n20953 : n32;
  assign n35483 = pi19 ? n35481 : n35482;
  assign n35484 = pi18 ? n35479 : n35483;
  assign n35485 = pi17 ? n9797 : n35484;
  assign n35486 = pi16 ? n439 : n35485;
  assign n35487 = pi15 ? n35477 : n35486;
  assign n35488 = pi14 ? n35474 : n35487;
  assign n35489 = pi13 ? n35462 : n35488;
  assign n35490 = pi19 ? n37 : n998;
  assign n35491 = pi18 ? n35490 : n139;
  assign n35492 = pi21 ? n3990 : n397;
  assign n35493 = pi20 ? n9082 : n35492;
  assign n35494 = pi19 ? n35493 : n32;
  assign n35495 = pi18 ? n139 : n35494;
  assign n35496 = pi17 ? n35491 : n35495;
  assign n35497 = pi16 ? n439 : n35496;
  assign n35498 = pi20 ? n139 : n1912;
  assign n35499 = pi19 ? n139 : n35498;
  assign n35500 = pi18 ? n14115 : n35499;
  assign n35501 = pi20 ? n1582 : n18978;
  assign n35502 = pi20 ? n18978 : n1016;
  assign n35503 = pi19 ? n35501 : n35502;
  assign n35504 = pi21 ? n204 : n6194;
  assign n35505 = pi20 ? n204 : n35504;
  assign n35506 = pi19 ? n35505 : n32;
  assign n35507 = pi18 ? n35503 : n35506;
  assign n35508 = pi17 ? n35500 : n35507;
  assign n35509 = pi16 ? n439 : n35508;
  assign n35510 = pi15 ? n35497 : n35509;
  assign n35511 = pi20 ? n941 : n1016;
  assign n35512 = pi19 ? n35511 : n204;
  assign n35513 = pi18 ? n12371 : n35512;
  assign n35514 = pi20 ? n204 : n17130;
  assign n35515 = pi20 ? n204 : n31588;
  assign n35516 = pi19 ? n35514 : n35515;
  assign n35517 = pi18 ? n35516 : n35506;
  assign n35518 = pi17 ? n35513 : n35517;
  assign n35519 = pi16 ? n439 : n35518;
  assign n35520 = pi18 ? n37 : n18109;
  assign n35521 = pi21 ? n204 : n6270;
  assign n35522 = pi20 ? n204 : n35521;
  assign n35523 = pi19 ? n35522 : n32;
  assign n35524 = pi18 ? n204 : n35523;
  assign n35525 = pi17 ? n35520 : n35524;
  assign n35526 = pi16 ? n439 : n35525;
  assign n35527 = pi15 ? n35519 : n35526;
  assign n35528 = pi14 ? n35510 : n35527;
  assign n35529 = pi18 ? n374 : n13110;
  assign n35530 = pi17 ? n32 : n35529;
  assign n35531 = pi20 ? n6568 : n8710;
  assign n35532 = pi19 ? n8765 : n35531;
  assign n35533 = pi21 ? n1056 : n4709;
  assign n35534 = pi21 ? n2876 : n204;
  assign n35535 = pi20 ? n35533 : n35534;
  assign n35536 = pi19 ? n35535 : n204;
  assign n35537 = pi18 ? n35532 : n35536;
  assign n35538 = pi17 ? n35537 : n35524;
  assign n35539 = pi16 ? n35530 : n35538;
  assign n35540 = pi18 ? n15029 : n34651;
  assign n35541 = pi21 ? n204 : n15874;
  assign n35542 = pi20 ? n204 : n35541;
  assign n35543 = pi19 ? n35542 : n32;
  assign n35544 = pi18 ? n204 : n35543;
  assign n35545 = pi17 ? n35540 : n35544;
  assign n35546 = pi16 ? n439 : n35545;
  assign n35547 = pi15 ? n35539 : n35546;
  assign n35548 = pi21 ? n37 : n3411;
  assign n35549 = pi20 ? n37 : n35548;
  assign n35550 = pi19 ? n35549 : n19358;
  assign n35551 = pi18 ? n37 : n35550;
  assign n35552 = pi20 ? n233 : n2094;
  assign n35553 = pi19 ? n35552 : n233;
  assign n35554 = pi20 ? n16544 : n24117;
  assign n35555 = pi19 ? n35554 : n32;
  assign n35556 = pi18 ? n35553 : n35555;
  assign n35557 = pi17 ? n35551 : n35556;
  assign n35558 = pi16 ? n439 : n35557;
  assign n35559 = pi19 ? n6373 : n19358;
  assign n35560 = pi18 ? n37 : n35559;
  assign n35561 = pi20 ? n233 : n649;
  assign n35562 = pi19 ? n35561 : n34678;
  assign n35563 = pi21 ? n233 : n15889;
  assign n35564 = pi20 ? n233 : n35563;
  assign n35565 = pi19 ? n35564 : n32;
  assign n35566 = pi18 ? n35562 : n35565;
  assign n35567 = pi17 ? n35560 : n35566;
  assign n35568 = pi16 ? n439 : n35567;
  assign n35569 = pi15 ? n35558 : n35568;
  assign n35570 = pi14 ? n35547 : n35569;
  assign n35571 = pi13 ? n35528 : n35570;
  assign n35572 = pi12 ? n35489 : n35571;
  assign n35573 = pi20 ? n233 : n24135;
  assign n35574 = pi19 ? n35573 : n32;
  assign n35575 = pi18 ? n17205 : n35574;
  assign n35576 = pi17 ? n6375 : n35575;
  assign n35577 = pi16 ? n439 : n35576;
  assign n35578 = pi20 ? n16544 : n14657;
  assign n35579 = pi19 ? n35578 : n32;
  assign n35580 = pi18 ? n34697 : n35579;
  assign n35581 = pi17 ? n34696 : n35580;
  assign n35582 = pi16 ? n439 : n35581;
  assign n35583 = pi15 ? n35577 : n35582;
  assign n35584 = pi21 ? n6376 : n316;
  assign n35585 = pi21 ? n25977 : n882;
  assign n35586 = pi20 ? n35584 : n35585;
  assign n35587 = pi19 ? n35586 : n32;
  assign n35588 = pi18 ? n34707 : n35587;
  assign n35589 = pi17 ? n34706 : n35588;
  assign n35590 = pi16 ? n34705 : n35589;
  assign n35591 = pi19 ? n612 : n22046;
  assign n35592 = pi18 ? n335 : n35591;
  assign n35593 = pi20 ? n610 : n37;
  assign n35594 = pi19 ? n30712 : n35593;
  assign n35595 = pi18 ? n35594 : n35120;
  assign n35596 = pi17 ? n35592 : n35595;
  assign n35597 = pi16 ? n34705 : n35596;
  assign n35598 = pi15 ? n35590 : n35597;
  assign n35599 = pi14 ? n35583 : n35598;
  assign n35600 = pi18 ? n34729 : n35120;
  assign n35601 = pi17 ? n335 : n35600;
  assign n35602 = pi16 ? n3351 : n35601;
  assign n35603 = pi19 ? n31719 : n18432;
  assign n35604 = pi18 ? n335 : n35603;
  assign n35605 = pi20 ? n6362 : n2075;
  assign n35606 = pi19 ? n35605 : n19405;
  assign n35607 = pi18 ? n35606 : n35120;
  assign n35608 = pi17 ? n35604 : n35607;
  assign n35609 = pi16 ? n2035 : n35608;
  assign n35610 = pi15 ? n35602 : n35609;
  assign n35611 = pi22 ? n335 : n7326;
  assign n35612 = pi21 ? n37 : n35611;
  assign n35613 = pi20 ? n35612 : n13289;
  assign n35614 = pi22 ? n18461 : n37;
  assign n35615 = pi21 ? n35614 : n1943;
  assign n35616 = pi21 ? n5015 : n18462;
  assign n35617 = pi20 ? n35615 : n35616;
  assign n35618 = pi19 ? n35613 : n35617;
  assign n35619 = pi22 ? n583 : n363;
  assign n35620 = pi21 ? n17548 : n35619;
  assign n35621 = pi22 ? n10400 : n583;
  assign n35622 = pi21 ? n35621 : n22142;
  assign n35623 = pi20 ? n35620 : n35622;
  assign n35624 = pi19 ? n35623 : n233;
  assign n35625 = pi18 ? n35618 : n35624;
  assign n35626 = pi21 ? n2048 : n4998;
  assign n35627 = pi20 ? n233 : n35626;
  assign n35628 = pi19 ? n35627 : n233;
  assign n35629 = pi18 ? n35628 : n35120;
  assign n35630 = pi17 ? n35625 : n35629;
  assign n35631 = pi16 ? n439 : n35630;
  assign n35632 = pi21 ? n935 : n37;
  assign n35633 = pi20 ? n32 : n35632;
  assign n35634 = pi19 ? n32 : n35633;
  assign n35635 = pi18 ? n35634 : n37;
  assign n35636 = pi17 ? n32 : n35635;
  assign n35637 = pi19 ? n22883 : n363;
  assign n35638 = pi20 ? n363 : n23155;
  assign n35639 = pi19 ? n35638 : n233;
  assign n35640 = pi18 ? n35637 : n35639;
  assign n35641 = pi21 ? n363 : n1920;
  assign n35642 = pi20 ? n233 : n35641;
  assign n35643 = pi19 ? n35642 : n233;
  assign n35644 = pi18 ? n35643 : n35127;
  assign n35645 = pi17 ? n35640 : n35644;
  assign n35646 = pi16 ? n35636 : n35645;
  assign n35647 = pi15 ? n35631 : n35646;
  assign n35648 = pi14 ? n35610 : n35647;
  assign n35649 = pi13 ? n35599 : n35648;
  assign n35650 = pi21 ? n12608 : n37;
  assign n35651 = pi20 ? n32 : n35650;
  assign n35652 = pi19 ? n32 : n35651;
  assign n35653 = pi18 ? n35652 : n363;
  assign n35654 = pi17 ? n32 : n35653;
  assign n35655 = pi20 ? n19084 : n685;
  assign n35656 = pi19 ? n363 : n35655;
  assign n35657 = pi18 ? n363 : n35656;
  assign n35658 = pi21 ? n363 : n19933;
  assign n35659 = pi20 ? n25199 : n35658;
  assign n35660 = pi20 ? n26891 : n685;
  assign n35661 = pi19 ? n35659 : n35660;
  assign n35662 = pi20 ? n685 : n7407;
  assign n35663 = pi19 ? n35662 : n32;
  assign n35664 = pi18 ? n35661 : n35663;
  assign n35665 = pi17 ? n35657 : n35664;
  assign n35666 = pi16 ? n35654 : n35665;
  assign n35667 = pi20 ? n37 : n3392;
  assign n35668 = pi19 ? n37 : n35667;
  assign n35669 = pi18 ? n37 : n35668;
  assign n35670 = pi20 ? n19091 : n37;
  assign n35671 = pi19 ? n35670 : n2730;
  assign n35672 = pi20 ? n18194 : n13793;
  assign n35673 = pi19 ? n35672 : n32;
  assign n35674 = pi18 ? n35671 : n35673;
  assign n35675 = pi17 ? n35669 : n35674;
  assign n35676 = pi16 ? n439 : n35675;
  assign n35677 = pi15 ? n35666 : n35676;
  assign n35678 = pi18 ? n20569 : n99;
  assign n35679 = pi17 ? n32 : n35678;
  assign n35680 = pi20 ? n32788 : n30773;
  assign n35681 = pi19 ? n99 : n35680;
  assign n35682 = pi20 ? n25167 : n99;
  assign n35683 = pi20 ? n30766 : n363;
  assign n35684 = pi19 ? n35682 : n35683;
  assign n35685 = pi18 ? n35681 : n35684;
  assign n35686 = pi21 ? n22549 : n722;
  assign n35687 = pi20 ? n32787 : n35686;
  assign n35688 = pi19 ? n35687 : n29738;
  assign n35689 = pi20 ? n24220 : n1010;
  assign n35690 = pi19 ? n35689 : n32;
  assign n35691 = pi18 ? n35688 : n35690;
  assign n35692 = pi17 ? n35685 : n35691;
  assign n35693 = pi16 ? n35679 : n35692;
  assign n35694 = pi21 ? n29690 : n363;
  assign n35695 = pi20 ? n99 : n35694;
  assign n35696 = pi20 ? n30778 : n363;
  assign n35697 = pi19 ? n35695 : n35696;
  assign n35698 = pi21 ? n22557 : n363;
  assign n35699 = pi20 ? n35698 : n23162;
  assign n35700 = pi19 ? n35699 : n34797;
  assign n35701 = pi18 ? n35697 : n35700;
  assign n35702 = pi17 ? n35701 : n34802;
  assign n35703 = pi16 ? n721 : n35702;
  assign n35704 = pi15 ? n35693 : n35703;
  assign n35705 = pi14 ? n35677 : n35704;
  assign n35706 = pi20 ? n363 : n7049;
  assign n35707 = pi19 ? n35706 : n32;
  assign n35708 = pi18 ? n363 : n35707;
  assign n35709 = pi17 ? n363 : n35708;
  assign n35710 = pi16 ? n21561 : n35709;
  assign n35711 = pi15 ? n34813 : n35710;
  assign n35712 = pi23 ? n1590 : n157;
  assign n35713 = pi22 ? n35712 : n363;
  assign n35714 = pi22 ? n10400 : n363;
  assign n35715 = pi21 ? n35713 : n35714;
  assign n35716 = pi20 ? n32 : n35715;
  assign n35717 = pi19 ? n32 : n35716;
  assign n35718 = pi18 ? n35717 : n363;
  assign n35719 = pi17 ? n32 : n35718;
  assign n35720 = pi20 ? n19084 : n20902;
  assign n35721 = pi19 ? n35720 : n32;
  assign n35722 = pi18 ? n363 : n35721;
  assign n35723 = pi17 ? n363 : n35722;
  assign n35724 = pi16 ? n35719 : n35723;
  assign n35725 = pi21 ? n7781 : n157;
  assign n35726 = pi20 ? n35725 : n26641;
  assign n35727 = pi19 ? n35726 : n157;
  assign n35728 = pi18 ? n157 : n35727;
  assign n35729 = pi20 ? n685 : n3320;
  assign n35730 = pi19 ? n35729 : n32;
  assign n35731 = pi18 ? n157 : n35730;
  assign n35732 = pi17 ? n35728 : n35731;
  assign n35733 = pi16 ? n7793 : n35732;
  assign n35734 = pi15 ? n35724 : n35733;
  assign n35735 = pi14 ? n35711 : n35734;
  assign n35736 = pi13 ? n35705 : n35735;
  assign n35737 = pi12 ? n35649 : n35736;
  assign n35738 = pi11 ? n35572 : n35737;
  assign n35739 = pi10 ? n35430 : n35738;
  assign n35740 = pi09 ? n35183 : n35739;
  assign n35741 = pi19 ? n31904 : n34261;
  assign n35742 = pi18 ? n35741 : n99;
  assign n35743 = pi17 ? n35742 : n35165;
  assign n35744 = pi16 ? n34860 : n35743;
  assign n35745 = pi15 ? n32 : n35744;
  assign n35746 = pi19 ? n31299 : n34261;
  assign n35747 = pi18 ? n35746 : n99;
  assign n35748 = pi17 ? n35747 : n35173;
  assign n35749 = pi16 ? n34860 : n35748;
  assign n35750 = pi15 ? n35175 : n35749;
  assign n35751 = pi14 ? n35745 : n35750;
  assign n35752 = pi13 ? n32 : n35751;
  assign n35753 = pi12 ? n32 : n35752;
  assign n35754 = pi11 ? n32 : n35753;
  assign n35755 = pi10 ? n32 : n35754;
  assign n35756 = pi18 ? n33966 : n34277;
  assign n35757 = pi22 ? n99 : n2026;
  assign n35758 = pi21 ? n35757 : n32;
  assign n35759 = pi20 ? n35758 : n32;
  assign n35760 = pi19 ? n15543 : n35759;
  assign n35761 = pi18 ? n99 : n35760;
  assign n35762 = pi17 ? n35756 : n35761;
  assign n35763 = pi16 ? n35195 : n35762;
  assign n35764 = pi18 ? n31265 : n20563;
  assign n35765 = pi17 ? n32 : n35764;
  assign n35766 = pi22 ? n99 : n8198;
  assign n35767 = pi21 ? n35766 : n32;
  assign n35768 = pi20 ? n35767 : n32;
  assign n35769 = pi19 ? n99 : n35768;
  assign n35770 = pi18 ? n99 : n35769;
  assign n35771 = pi17 ? n35197 : n35770;
  assign n35772 = pi16 ? n35765 : n35771;
  assign n35773 = pi15 ? n35763 : n35772;
  assign n35774 = pi17 ? n35211 : n34291;
  assign n35775 = pi16 ? n35208 : n35774;
  assign n35776 = pi20 ? n20563 : n32286;
  assign n35777 = pi19 ? n20563 : n35776;
  assign n35778 = pi18 ? n31315 : n35777;
  assign n35779 = pi17 ? n32 : n35778;
  assign n35780 = pi20 ? n19794 : n32;
  assign n35781 = pi19 ? n37 : n35780;
  assign n35782 = pi18 ? n37 : n35781;
  assign n35783 = pi17 ? n37 : n35782;
  assign n35784 = pi16 ? n35779 : n35783;
  assign n35785 = pi15 ? n35775 : n35784;
  assign n35786 = pi14 ? n35773 : n35785;
  assign n35787 = pi20 ? n20563 : n31948;
  assign n35788 = pi19 ? n20563 : n35787;
  assign n35789 = pi18 ? n31315 : n35788;
  assign n35790 = pi17 ? n32 : n35789;
  assign n35791 = pi22 ? n37 : n1378;
  assign n35792 = pi21 ? n35791 : n32;
  assign n35793 = pi20 ? n35792 : n32;
  assign n35794 = pi19 ? n37 : n35793;
  assign n35795 = pi18 ? n37 : n35794;
  assign n35796 = pi17 ? n37 : n35795;
  assign n35797 = pi16 ? n35790 : n35796;
  assign n35798 = pi20 ? n20563 : n33964;
  assign n35799 = pi19 ? n20563 : n35798;
  assign n35800 = pi18 ? n31315 : n35799;
  assign n35801 = pi17 ? n32 : n35800;
  assign n35802 = pi20 ? n21726 : n32;
  assign n35803 = pi19 ? n9814 : n35802;
  assign n35804 = pi18 ? n37 : n35803;
  assign n35805 = pi17 ? n37 : n35804;
  assign n35806 = pi16 ? n35801 : n35805;
  assign n35807 = pi15 ? n35797 : n35806;
  assign n35808 = pi19 ? n8765 : n7503;
  assign n35809 = pi18 ? n139 : n35808;
  assign n35810 = pi17 ? n35248 : n35809;
  assign n35811 = pi16 ? n34884 : n35810;
  assign n35812 = pi19 ? n20563 : n35317;
  assign n35813 = pi18 ? n31315 : n35812;
  assign n35814 = pi17 ? n32 : n35813;
  assign n35815 = pi20 ? n20301 : n32;
  assign n35816 = pi19 ? n9769 : n35815;
  assign n35817 = pi18 ? n139 : n35816;
  assign n35818 = pi17 ? n35254 : n35817;
  assign n35819 = pi16 ? n35814 : n35818;
  assign n35820 = pi15 ? n35811 : n35819;
  assign n35821 = pi14 ? n35807 : n35820;
  assign n35822 = pi13 ? n35786 : n35821;
  assign n35823 = pi19 ? n8765 : n35815;
  assign n35824 = pi18 ? n35264 : n35823;
  assign n35825 = pi17 ? n37 : n35824;
  assign n35826 = pi16 ? n34889 : n35825;
  assign n35827 = pi20 ? n20309 : n32;
  assign n35828 = pi19 ? n4733 : n35827;
  assign n35829 = pi18 ? n35270 : n35828;
  assign n35830 = pi17 ? n37 : n35829;
  assign n35831 = pi16 ? n34889 : n35830;
  assign n35832 = pi15 ? n35826 : n35831;
  assign n35833 = pi21 ? n27868 : n32;
  assign n35834 = pi20 ? n35833 : n32;
  assign n35835 = pi19 ? n35277 : n35834;
  assign n35836 = pi18 ? n35276 : n35835;
  assign n35837 = pi17 ? n37 : n35836;
  assign n35838 = pi16 ? n34889 : n35837;
  assign n35839 = pi22 ? n335 : n396;
  assign n35840 = pi21 ? n35839 : n32;
  assign n35841 = pi20 ? n35840 : n32;
  assign n35842 = pi19 ? n17204 : n35841;
  assign n35843 = pi18 ? n37 : n35842;
  assign n35844 = pi17 ? n37 : n35843;
  assign n35845 = pi16 ? n34335 : n35844;
  assign n35846 = pi15 ? n35838 : n35845;
  assign n35847 = pi14 ? n35832 : n35846;
  assign n35848 = pi21 ? n30390 : n32;
  assign n35849 = pi20 ? n35848 : n32;
  assign n35850 = pi19 ? n12628 : n35849;
  assign n35851 = pi18 ? n37 : n35850;
  assign n35852 = pi17 ? n37 : n35851;
  assign n35853 = pi16 ? n33883 : n35852;
  assign n35854 = pi20 ? n20563 : n35316;
  assign n35855 = pi19 ? n35854 : n37;
  assign n35856 = pi18 ? n31315 : n35855;
  assign n35857 = pi17 ? n32 : n35856;
  assign n35858 = pi22 ? n5011 : n1378;
  assign n35859 = pi21 ? n35858 : n32;
  assign n35860 = pi20 ? n35859 : n32;
  assign n35861 = pi19 ? n3332 : n35860;
  assign n35862 = pi18 ? n37 : n35861;
  assign n35863 = pi17 ? n37 : n35862;
  assign n35864 = pi16 ? n35857 : n35863;
  assign n35865 = pi15 ? n35853 : n35864;
  assign n35866 = pi21 ? n14155 : n32;
  assign n35867 = pi20 ? n35866 : n32;
  assign n35868 = pi19 ? n37 : n35867;
  assign n35869 = pi18 ? n37 : n35868;
  assign n35870 = pi17 ? n37 : n35869;
  assign n35871 = pi16 ? n34360 : n35870;
  assign n35872 = pi16 ? n33332 : n35305;
  assign n35873 = pi15 ? n35871 : n35872;
  assign n35874 = pi14 ? n35865 : n35873;
  assign n35875 = pi13 ? n35847 : n35874;
  assign n35876 = pi12 ? n35822 : n35875;
  assign n35877 = pi19 ? n35311 : n8262;
  assign n35878 = pi18 ? n14149 : n35877;
  assign n35879 = pi17 ? n37 : n35878;
  assign n35880 = pi16 ? n32915 : n35879;
  assign n35881 = pi18 ? n31938 : n32369;
  assign n35882 = pi17 ? n32 : n35881;
  assign n35883 = pi19 ? n35322 : n7680;
  assign n35884 = pi18 ? n35321 : n35883;
  assign n35885 = pi17 ? n37 : n35884;
  assign n35886 = pi16 ? n35882 : n35885;
  assign n35887 = pi15 ? n35880 : n35886;
  assign n35888 = pi22 ? n19715 : n625;
  assign n35889 = pi21 ? n35888 : n32;
  assign n35890 = pi20 ? n35889 : n32;
  assign n35891 = pi19 ? n10681 : n35890;
  assign n35892 = pi18 ? n35330 : n35891;
  assign n35893 = pi17 ? n37 : n35892;
  assign n35894 = pi16 ? n32371 : n35893;
  assign n35895 = pi20 ? n22333 : n32;
  assign n35896 = pi19 ? n24866 : n35895;
  assign n35897 = pi18 ? n37 : n35896;
  assign n35898 = pi17 ? n37 : n35897;
  assign n35899 = pi16 ? n32371 : n35898;
  assign n35900 = pi15 ? n35894 : n35899;
  assign n35901 = pi14 ? n35887 : n35900;
  assign n35902 = pi23 ? n363 : n8310;
  assign n35903 = pi22 ? n35902 : n688;
  assign n35904 = pi21 ? n35903 : n32;
  assign n35905 = pi20 ? n35904 : n32;
  assign n35906 = pi19 ? n22883 : n35905;
  assign n35907 = pi18 ? n37 : n35906;
  assign n35908 = pi17 ? n37 : n35907;
  assign n35909 = pi16 ? n33374 : n35908;
  assign n35910 = pi18 ? n31938 : n33950;
  assign n35911 = pi17 ? n32 : n35910;
  assign n35912 = pi23 ? n363 : n7420;
  assign n35913 = pi22 ? n35912 : n706;
  assign n35914 = pi21 ? n35913 : n32;
  assign n35915 = pi20 ? n35914 : n32;
  assign n35916 = pi19 ? n6403 : n35915;
  assign n35917 = pi18 ? n37 : n35916;
  assign n35918 = pi17 ? n37 : n35917;
  assign n35919 = pi16 ? n35911 : n35918;
  assign n35920 = pi15 ? n35909 : n35919;
  assign n35921 = pi22 ? n10341 : n706;
  assign n35922 = pi21 ? n35921 : n32;
  assign n35923 = pi20 ? n35922 : n32;
  assign n35924 = pi19 ? n37 : n35923;
  assign n35925 = pi18 ? n37 : n35924;
  assign n35926 = pi17 ? n37 : n35925;
  assign n35927 = pi16 ? n35911 : n35926;
  assign n35928 = pi22 ? n35912 : n32;
  assign n35929 = pi21 ? n35928 : n32;
  assign n35930 = pi20 ? n35929 : n32;
  assign n35931 = pi19 ? n6403 : n35930;
  assign n35932 = pi18 ? n37 : n35931;
  assign n35933 = pi17 ? n37 : n35932;
  assign n35934 = pi16 ? n32926 : n35933;
  assign n35935 = pi15 ? n35927 : n35934;
  assign n35936 = pi14 ? n35920 : n35935;
  assign n35937 = pi13 ? n35901 : n35936;
  assign n35938 = pi24 ? n157 : n233;
  assign n35939 = pi23 ? n363 : n35938;
  assign n35940 = pi22 ? n35939 : n32;
  assign n35941 = pi21 ? n35940 : n32;
  assign n35942 = pi20 ? n35941 : n32;
  assign n35943 = pi19 ? n5029 : n35942;
  assign n35944 = pi18 ? n37 : n35943;
  assign n35945 = pi17 ? n37 : n35944;
  assign n35946 = pi16 ? n31317 : n35945;
  assign n35947 = pi21 ? n31293 : n29133;
  assign n35948 = pi20 ? n32 : n35947;
  assign n35949 = pi19 ? n32 : n35948;
  assign n35950 = pi18 ? n35949 : n32934;
  assign n35951 = pi17 ? n32 : n35950;
  assign n35952 = pi19 ? n6403 : n8296;
  assign n35953 = pi18 ? n37 : n35952;
  assign n35954 = pi17 ? n37 : n35953;
  assign n35955 = pi16 ? n35951 : n35954;
  assign n35956 = pi15 ? n35946 : n35955;
  assign n35957 = pi21 ? n30866 : n31924;
  assign n35958 = pi20 ? n32 : n35957;
  assign n35959 = pi19 ? n32 : n35958;
  assign n35960 = pi18 ? n35959 : n32934;
  assign n35961 = pi17 ? n32 : n35960;
  assign n35962 = pi19 ? n8743 : n8296;
  assign n35963 = pi18 ? n37 : n35962;
  assign n35964 = pi17 ? n37 : n35963;
  assign n35965 = pi16 ? n35961 : n35964;
  assign n35966 = pi19 ? n8802 : n4009;
  assign n35967 = pi18 ? n35381 : n35966;
  assign n35968 = pi17 ? n35378 : n35967;
  assign n35969 = pi16 ? n35961 : n35968;
  assign n35970 = pi15 ? n35965 : n35969;
  assign n35971 = pi14 ? n35956 : n35970;
  assign n35972 = pi19 ? n34479 : n4009;
  assign n35973 = pi18 ? n37 : n35972;
  assign n35974 = pi17 ? n37 : n35973;
  assign n35975 = pi16 ? n33409 : n35974;
  assign n35976 = pi19 ? n35397 : n4117;
  assign n35977 = pi18 ? n37 : n35976;
  assign n35978 = pi17 ? n37 : n35977;
  assign n35979 = pi16 ? n32415 : n35978;
  assign n35980 = pi15 ? n35975 : n35979;
  assign n35981 = pi18 ? n34997 : n17982;
  assign n35982 = pi17 ? n32 : n35981;
  assign n35983 = pi21 ? n8654 : n3002;
  assign n35984 = pi22 ? n893 : n2160;
  assign n35985 = pi21 ? n35984 : n3002;
  assign n35986 = pi20 ? n35983 : n35985;
  assign n35987 = pi19 ? n5502 : n35986;
  assign n35988 = pi22 ? n164 : n112;
  assign n35989 = pi21 ? n22379 : n35988;
  assign n35990 = pi22 ? n2160 : n889;
  assign n35991 = pi21 ? n35990 : n3002;
  assign n35992 = pi20 ? n35989 : n35991;
  assign n35993 = pi21 ? n5877 : n3002;
  assign n35994 = pi19 ? n35992 : n35993;
  assign n35995 = pi18 ? n35987 : n35994;
  assign n35996 = pi21 ? n157 : n35984;
  assign n35997 = pi20 ? n6523 : n35996;
  assign n35998 = pi20 ? n28939 : n9015;
  assign n35999 = pi19 ? n35997 : n35998;
  assign n36000 = pi19 ? n157 : n10012;
  assign n36001 = pi18 ? n35999 : n36000;
  assign n36002 = pi17 ? n35995 : n36001;
  assign n36003 = pi16 ? n35982 : n36002;
  assign n36004 = pi18 ? n157 : n36000;
  assign n36005 = pi17 ? n34500 : n36004;
  assign n36006 = pi16 ? n35006 : n36005;
  assign n36007 = pi15 ? n36003 : n36006;
  assign n36008 = pi14 ? n35980 : n36007;
  assign n36009 = pi13 ? n35971 : n36008;
  assign n36010 = pi12 ? n35937 : n36009;
  assign n36011 = pi11 ? n35876 : n36010;
  assign n36012 = pi19 ? n157 : n5831;
  assign n36013 = pi18 ? n35437 : n36012;
  assign n36014 = pi17 ? n35435 : n36013;
  assign n36015 = pi16 ? n32415 : n36014;
  assign n36016 = pi19 ? n9035 : n10012;
  assign n36017 = pi18 ? n35444 : n36016;
  assign n36018 = pi17 ? n35441 : n36017;
  assign n36019 = pi16 ? n32014 : n36018;
  assign n36020 = pi15 ? n36015 : n36019;
  assign n36021 = pi18 ? n32012 : n18854;
  assign n36022 = pi17 ? n32 : n36021;
  assign n36023 = pi16 ? n36022 : n35454;
  assign n36024 = pi18 ? n34014 : n21612;
  assign n36025 = pi17 ? n32 : n36024;
  assign n36026 = pi16 ? n36025 : n35459;
  assign n36027 = pi15 ? n36023 : n36026;
  assign n36028 = pi14 ? n36020 : n36027;
  assign n36029 = pi23 ? n38 : n30868;
  assign n36030 = pi22 ? n36029 : n37;
  assign n36031 = pi21 ? n36030 : n37;
  assign n36032 = pi20 ? n32 : n36031;
  assign n36033 = pi19 ? n32 : n36032;
  assign n36034 = pi18 ? n36033 : n37;
  assign n36035 = pi17 ? n32 : n36034;
  assign n36036 = pi16 ? n36035 : n35485;
  assign n36037 = pi15 ? n35477 : n36036;
  assign n36038 = pi14 ? n35474 : n36037;
  assign n36039 = pi13 ? n36028 : n36038;
  assign n36040 = pi21 ? n1785 : n4780;
  assign n36041 = pi22 ? n316 : n3301;
  assign n36042 = pi21 ? n3188 : n36041;
  assign n36043 = pi20 ? n36040 : n36042;
  assign n36044 = pi19 ? n36043 : n32;
  assign n36045 = pi18 ? n139 : n36044;
  assign n36046 = pi17 ? n35491 : n36045;
  assign n36047 = pi16 ? n439 : n36046;
  assign n36048 = pi21 ? n204 : n16933;
  assign n36049 = pi20 ? n204 : n36048;
  assign n36050 = pi19 ? n36049 : n32;
  assign n36051 = pi18 ? n35503 : n36050;
  assign n36052 = pi17 ? n35500 : n36051;
  assign n36053 = pi16 ? n439 : n36052;
  assign n36054 = pi15 ? n36047 : n36053;
  assign n36055 = pi18 ? n35516 : n36050;
  assign n36056 = pi17 ? n35513 : n36055;
  assign n36057 = pi16 ? n439 : n36056;
  assign n36058 = pi22 ? n204 : n3338;
  assign n36059 = pi21 ? n204 : n36058;
  assign n36060 = pi20 ? n204 : n36059;
  assign n36061 = pi19 ? n36060 : n32;
  assign n36062 = pi18 ? n204 : n36061;
  assign n36063 = pi17 ? n35520 : n36062;
  assign n36064 = pi16 ? n439 : n36063;
  assign n36065 = pi15 ? n36057 : n36064;
  assign n36066 = pi14 ? n36054 : n36065;
  assign n36067 = pi17 ? n35537 : n36062;
  assign n36068 = pi16 ? n35530 : n36067;
  assign n36069 = pi15 ? n36068 : n35546;
  assign n36070 = pi14 ? n36069 : n35569;
  assign n36071 = pi13 ? n36066 : n36070;
  assign n36072 = pi12 ? n36039 : n36071;
  assign n36073 = pi18 ? n17205 : n35565;
  assign n36074 = pi17 ? n6375 : n36073;
  assign n36075 = pi16 ? n439 : n36074;
  assign n36076 = pi21 ? n233 : n9202;
  assign n36077 = pi20 ? n16544 : n36076;
  assign n36078 = pi19 ? n36077 : n32;
  assign n36079 = pi18 ? n34697 : n36078;
  assign n36080 = pi17 ? n34696 : n36079;
  assign n36081 = pi16 ? n439 : n36080;
  assign n36082 = pi15 ? n36075 : n36081;
  assign n36083 = pi20 ? n233 : n24817;
  assign n36084 = pi19 ? n36083 : n32;
  assign n36085 = pi18 ? n35594 : n36084;
  assign n36086 = pi17 ? n35592 : n36085;
  assign n36087 = pi16 ? n34705 : n36086;
  assign n36088 = pi15 ? n35590 : n36087;
  assign n36089 = pi14 ? n36082 : n36088;
  assign n36090 = pi18 ? n34729 : n36084;
  assign n36091 = pi17 ? n335 : n36090;
  assign n36092 = pi16 ? n3351 : n36091;
  assign n36093 = pi21 ? n233 : n3397;
  assign n36094 = pi20 ? n233 : n36093;
  assign n36095 = pi19 ? n36094 : n32;
  assign n36096 = pi18 ? n35606 : n36095;
  assign n36097 = pi17 ? n35604 : n36096;
  assign n36098 = pi16 ? n2035 : n36097;
  assign n36099 = pi15 ? n36092 : n36098;
  assign n36100 = pi20 ? n35612 : n639;
  assign n36101 = pi21 ? n7334 : n1943;
  assign n36102 = pi20 ? n36101 : n35616;
  assign n36103 = pi19 ? n36100 : n36102;
  assign n36104 = pi22 ? n7326 : n233;
  assign n36105 = pi21 ? n35621 : n36104;
  assign n36106 = pi20 ? n35620 : n36105;
  assign n36107 = pi19 ? n36106 : n233;
  assign n36108 = pi18 ? n36103 : n36107;
  assign n36109 = pi20 ? n233 : n31811;
  assign n36110 = pi19 ? n36109 : n233;
  assign n36111 = pi20 ? n233 : n19352;
  assign n36112 = pi19 ? n36111 : n32;
  assign n36113 = pi18 ? n36110 : n36112;
  assign n36114 = pi17 ? n36108 : n36113;
  assign n36115 = pi16 ? n439 : n36114;
  assign n36116 = pi15 ? n36115 : n35646;
  assign n36117 = pi14 ? n36099 : n36116;
  assign n36118 = pi13 ? n36089 : n36117;
  assign n36119 = pi16 ? n721 : n35692;
  assign n36120 = pi22 ? n685 : n11681;
  assign n36121 = pi21 ? n36120 : n32;
  assign n36122 = pi20 ? n24220 : n36121;
  assign n36123 = pi19 ? n36122 : n32;
  assign n36124 = pi18 ? n363 : n36123;
  assign n36125 = pi17 ? n35701 : n36124;
  assign n36126 = pi16 ? n721 : n36125;
  assign n36127 = pi15 ? n36119 : n36126;
  assign n36128 = pi14 ? n35677 : n36127;
  assign n36129 = pi16 ? n21219 : n35709;
  assign n36130 = pi15 ? n34813 : n36129;
  assign n36131 = pi22 ? n3935 : n363;
  assign n36132 = pi21 ? n35713 : n36131;
  assign n36133 = pi20 ? n32 : n36132;
  assign n36134 = pi19 ? n32 : n36133;
  assign n36135 = pi18 ? n36134 : n363;
  assign n36136 = pi17 ? n32 : n36135;
  assign n36137 = pi20 ? n19084 : n8967;
  assign n36138 = pi19 ? n36137 : n32;
  assign n36139 = pi18 ? n363 : n36138;
  assign n36140 = pi17 ? n363 : n36139;
  assign n36141 = pi16 ? n36136 : n36140;
  assign n36142 = pi22 ? n35712 : n157;
  assign n36143 = pi21 ? n36142 : n157;
  assign n36144 = pi20 ? n32 : n36143;
  assign n36145 = pi19 ? n32 : n36144;
  assign n36146 = pi18 ? n36145 : n157;
  assign n36147 = pi17 ? n32 : n36146;
  assign n36148 = pi20 ? n685 : n3977;
  assign n36149 = pi19 ? n36148 : n32;
  assign n36150 = pi18 ? n157 : n36149;
  assign n36151 = pi17 ? n35728 : n36150;
  assign n36152 = pi16 ? n36147 : n36151;
  assign n36153 = pi15 ? n36141 : n36152;
  assign n36154 = pi14 ? n36130 : n36153;
  assign n36155 = pi13 ? n36128 : n36154;
  assign n36156 = pi12 ? n36118 : n36155;
  assign n36157 = pi11 ? n36072 : n36156;
  assign n36158 = pi10 ? n36011 : n36157;
  assign n36159 = pi09 ? n35755 : n36158;
  assign n36160 = pi08 ? n35740 : n36159;
  assign n36161 = pi07 ? n35159 : n36160;
  assign n36162 = pi18 ? n28159 : n20563;
  assign n36163 = pi17 ? n32 : n36162;
  assign n36164 = pi19 ? n31221 : n34261;
  assign n36165 = pi18 ? n36164 : n99;
  assign n36166 = pi19 ? n99 : n7301;
  assign n36167 = pi18 ? n99 : n36166;
  assign n36168 = pi17 ? n36165 : n36167;
  assign n36169 = pi16 ? n36163 : n36168;
  assign n36170 = pi15 ? n32 : n36169;
  assign n36171 = pi20 ? n37 : n23686;
  assign n36172 = pi19 ? n32348 : n36171;
  assign n36173 = pi18 ? n36172 : n99;
  assign n36174 = pi21 ? n746 : n32;
  assign n36175 = pi20 ? n36174 : n32;
  assign n36176 = pi19 ? n99 : n36175;
  assign n36177 = pi18 ? n99 : n36176;
  assign n36178 = pi17 ? n36173 : n36177;
  assign n36179 = pi16 ? n34860 : n36178;
  assign n36180 = pi19 ? n32348 : n34261;
  assign n36181 = pi18 ? n36180 : n99;
  assign n36182 = pi21 ? n4237 : n32;
  assign n36183 = pi20 ? n36182 : n32;
  assign n36184 = pi19 ? n99 : n36183;
  assign n36185 = pi18 ? n99 : n36184;
  assign n36186 = pi17 ? n36181 : n36185;
  assign n36187 = pi16 ? n34860 : n36186;
  assign n36188 = pi15 ? n36179 : n36187;
  assign n36189 = pi14 ? n36170 : n36188;
  assign n36190 = pi13 ? n32 : n36189;
  assign n36191 = pi12 ? n32 : n36190;
  assign n36192 = pi11 ? n32 : n36191;
  assign n36193 = pi10 ? n32 : n36192;
  assign n36194 = pi19 ? n31267 : n34261;
  assign n36195 = pi18 ? n36194 : n99;
  assign n36196 = pi20 ? n21276 : n32;
  assign n36197 = pi19 ? n99 : n36196;
  assign n36198 = pi18 ? n99 : n36197;
  assign n36199 = pi17 ? n36195 : n36198;
  assign n36200 = pi16 ? n35765 : n36199;
  assign n36201 = pi19 ? n30097 : n23648;
  assign n36202 = pi18 ? n36201 : n18854;
  assign n36203 = pi21 ? n4548 : n32;
  assign n36204 = pi20 ? n36203 : n32;
  assign n36205 = pi19 ? n99 : n36204;
  assign n36206 = pi18 ? n99 : n36205;
  assign n36207 = pi17 ? n36202 : n36206;
  assign n36208 = pi16 ? n35765 : n36207;
  assign n36209 = pi15 ? n36200 : n36208;
  assign n36210 = pi18 ? n32924 : n37;
  assign n36211 = pi19 ? n37 : n6030;
  assign n36212 = pi18 ? n37 : n36211;
  assign n36213 = pi17 ? n36210 : n36212;
  assign n36214 = pi16 ? n35765 : n36213;
  assign n36215 = pi18 ? n31315 : n20563;
  assign n36216 = pi17 ? n32 : n36215;
  assign n36217 = pi16 ? n36216 : n36213;
  assign n36218 = pi15 ? n36214 : n36217;
  assign n36219 = pi14 ? n36209 : n36218;
  assign n36220 = pi21 ? n28267 : n32;
  assign n36221 = pi20 ? n36220 : n32;
  assign n36222 = pi19 ? n9824 : n36221;
  assign n36223 = pi18 ? n37 : n36222;
  assign n36224 = pi17 ? n37 : n36223;
  assign n36225 = pi16 ? n36216 : n36224;
  assign n36226 = pi18 ? n31315 : n34258;
  assign n36227 = pi17 ? n32 : n36226;
  assign n36228 = pi18 ? n37 : n139;
  assign n36229 = pi19 ? n139 : n7503;
  assign n36230 = pi18 ? n139 : n36229;
  assign n36231 = pi17 ? n36228 : n36230;
  assign n36232 = pi16 ? n36227 : n36231;
  assign n36233 = pi15 ? n36225 : n36232;
  assign n36234 = pi18 ? n31315 : n34869;
  assign n36235 = pi17 ? n32 : n36234;
  assign n36236 = pi19 ? n16023 : n7503;
  assign n36237 = pi18 ? n139 : n36236;
  assign n36238 = pi17 ? n9816 : n36237;
  assign n36239 = pi16 ? n36235 : n36238;
  assign n36240 = pi19 ? n37 : n30225;
  assign n36241 = pi18 ? n36240 : n139;
  assign n36242 = pi19 ? n139 : n35815;
  assign n36243 = pi18 ? n139 : n36242;
  assign n36244 = pi17 ? n36241 : n36243;
  assign n36245 = pi16 ? n36227 : n36244;
  assign n36246 = pi15 ? n36239 : n36245;
  assign n36247 = pi14 ? n36233 : n36246;
  assign n36248 = pi13 ? n36219 : n36247;
  assign n36249 = pi22 ? n37 : n20563;
  assign n36250 = pi21 ? n36249 : n37;
  assign n36251 = pi20 ? n20563 : n36250;
  assign n36252 = pi19 ? n20563 : n36251;
  assign n36253 = pi18 ? n31315 : n36252;
  assign n36254 = pi17 ? n32 : n36253;
  assign n36255 = pi19 ? n9814 : n35252;
  assign n36256 = pi18 ? n37 : n36255;
  assign n36257 = pi17 ? n36256 : n35817;
  assign n36258 = pi16 ? n36254 : n36257;
  assign n36259 = pi19 ? n13125 : n3096;
  assign n36260 = pi18 ? n37 : n36259;
  assign n36261 = pi19 ? n9769 : n35827;
  assign n36262 = pi18 ? n139 : n36261;
  assign n36263 = pi17 ? n36260 : n36262;
  assign n36264 = pi16 ? n35220 : n36263;
  assign n36265 = pi15 ? n36258 : n36264;
  assign n36266 = pi18 ? n31938 : n34295;
  assign n36267 = pi17 ? n32 : n36266;
  assign n36268 = pi22 ? n37 : n20317;
  assign n36269 = pi21 ? n36268 : n32;
  assign n36270 = pi20 ? n36269 : n32;
  assign n36271 = pi19 ? n11827 : n36270;
  assign n36272 = pi18 ? n22047 : n36271;
  assign n36273 = pi17 ? n37 : n36272;
  assign n36274 = pi16 ? n36267 : n36273;
  assign n36275 = pi22 ? n37 : n1333;
  assign n36276 = pi21 ? n36275 : n32;
  assign n36277 = pi20 ? n36276 : n32;
  assign n36278 = pi19 ? n17204 : n36277;
  assign n36279 = pi18 ? n37 : n36278;
  assign n36280 = pi17 ? n37 : n36279;
  assign n36281 = pi16 ? n35244 : n36280;
  assign n36282 = pi15 ? n36274 : n36281;
  assign n36283 = pi14 ? n36265 : n36282;
  assign n36284 = pi22 ? n99 : n3124;
  assign n36285 = pi21 ? n36284 : n32;
  assign n36286 = pi20 ? n36285 : n32;
  assign n36287 = pi19 ? n17204 : n36286;
  assign n36288 = pi18 ? n37 : n36287;
  assign n36289 = pi17 ? n37 : n36288;
  assign n36290 = pi16 ? n34889 : n36289;
  assign n36291 = pi22 ? n112 : n1378;
  assign n36292 = pi21 ? n36291 : n32;
  assign n36293 = pi20 ? n36292 : n32;
  assign n36294 = pi19 ? n37 : n36293;
  assign n36295 = pi18 ? n37 : n36294;
  assign n36296 = pi17 ? n37 : n36295;
  assign n36297 = pi16 ? n34889 : n36296;
  assign n36298 = pi15 ? n36290 : n36297;
  assign n36299 = pi19 ? n2095 : n9442;
  assign n36300 = pi18 ? n37 : n36299;
  assign n36301 = pi17 ? n37 : n36300;
  assign n36302 = pi16 ? n34319 : n36301;
  assign n36303 = pi21 ? n30168 : n20563;
  assign n36304 = pi20 ? n32 : n36303;
  assign n36305 = pi19 ? n32 : n36304;
  assign n36306 = pi18 ? n36305 : n32295;
  assign n36307 = pi17 ? n32 : n36306;
  assign n36308 = pi20 ? n21760 : n32;
  assign n36309 = pi19 ? n17204 : n36308;
  assign n36310 = pi18 ? n37 : n36309;
  assign n36311 = pi17 ? n37 : n36310;
  assign n36312 = pi16 ? n36307 : n36311;
  assign n36313 = pi15 ? n36302 : n36312;
  assign n36314 = pi14 ? n36298 : n36313;
  assign n36315 = pi13 ? n36283 : n36314;
  assign n36316 = pi12 ? n36248 : n36315;
  assign n36317 = pi19 ? n37 : n639;
  assign n36318 = pi18 ? n37 : n36317;
  assign n36319 = pi20 ? n639 : n25064;
  assign n36320 = pi20 ? n610 : n22076;
  assign n36321 = pi19 ? n36319 : n36320;
  assign n36322 = pi19 ? n335 : n7660;
  assign n36323 = pi18 ? n36321 : n36322;
  assign n36324 = pi17 ? n36318 : n36323;
  assign n36325 = pi16 ? n35283 : n36324;
  assign n36326 = pi19 ? n22812 : n335;
  assign n36327 = pi18 ? n37 : n36326;
  assign n36328 = pi20 ? n20801 : n32;
  assign n36329 = pi19 ? n335 : n36328;
  assign n36330 = pi18 ? n335 : n36329;
  assign n36331 = pi17 ? n36327 : n36330;
  assign n36332 = pi16 ? n35857 : n36331;
  assign n36333 = pi15 ? n36325 : n36332;
  assign n36334 = pi21 ? n7986 : n1943;
  assign n36335 = pi20 ? n7646 : n36334;
  assign n36336 = pi19 ? n36335 : n9944;
  assign n36337 = pi18 ? n32452 : n36336;
  assign n36338 = pi17 ? n37 : n36337;
  assign n36339 = pi16 ? n34360 : n36338;
  assign n36340 = pi19 ? n23917 : n9950;
  assign n36341 = pi18 ? n37 : n36340;
  assign n36342 = pi17 ? n37 : n36341;
  assign n36343 = pi16 ? n32901 : n36342;
  assign n36344 = pi15 ? n36339 : n36343;
  assign n36345 = pi14 ? n36333 : n36344;
  assign n36346 = pi21 ? n7327 : n37;
  assign n36347 = pi20 ? n37 : n36346;
  assign n36348 = pi19 ? n36347 : n8042;
  assign n36349 = pi19 ? n22897 : n9950;
  assign n36350 = pi18 ? n36348 : n36349;
  assign n36351 = pi17 ? n37 : n36350;
  assign n36352 = pi16 ? n32901 : n36351;
  assign n36353 = pi19 ? n37 : n9950;
  assign n36354 = pi18 ? n37 : n36353;
  assign n36355 = pi17 ? n37 : n36354;
  assign n36356 = pi16 ? n32901 : n36355;
  assign n36357 = pi15 ? n36352 : n36356;
  assign n36358 = pi19 ? n37 : n34944;
  assign n36359 = pi18 ? n37 : n36358;
  assign n36360 = pi17 ? n37 : n36359;
  assign n36361 = pi16 ? n32901 : n36360;
  assign n36362 = pi20 ? n34919 : n37;
  assign n36363 = pi19 ? n36362 : n37;
  assign n36364 = pi18 ? n31938 : n36363;
  assign n36365 = pi17 ? n32 : n36364;
  assign n36366 = pi19 ? n17275 : n34944;
  assign n36367 = pi18 ? n37 : n36366;
  assign n36368 = pi17 ? n37 : n36367;
  assign n36369 = pi16 ? n36365 : n36368;
  assign n36370 = pi15 ? n36361 : n36369;
  assign n36371 = pi14 ? n36357 : n36370;
  assign n36372 = pi13 ? n36345 : n36371;
  assign n36373 = pi18 ? n31938 : n35318;
  assign n36374 = pi17 ? n32 : n36373;
  assign n36375 = pi19 ? n37 : n8296;
  assign n36376 = pi18 ? n37 : n36375;
  assign n36377 = pi17 ? n37 : n36376;
  assign n36378 = pi16 ? n36374 : n36377;
  assign n36379 = pi16 ? n35320 : n36377;
  assign n36380 = pi15 ? n36378 : n36379;
  assign n36381 = pi16 ? n31941 : n36377;
  assign n36382 = pi21 ? n685 : n19933;
  assign n36383 = pi20 ? n19934 : n36382;
  assign n36384 = pi19 ? n36383 : n9483;
  assign n36385 = pi18 ? n37 : n36384;
  assign n36386 = pi17 ? n37 : n36385;
  assign n36387 = pi16 ? n35911 : n36386;
  assign n36388 = pi15 ? n36381 : n36387;
  assign n36389 = pi14 ? n36380 : n36388;
  assign n36390 = pi20 ? n2107 : n36382;
  assign n36391 = pi20 ? n32826 : n32;
  assign n36392 = pi19 ? n36390 : n36391;
  assign n36393 = pi18 ? n37 : n36392;
  assign n36394 = pi17 ? n37 : n36393;
  assign n36395 = pi16 ? n33952 : n36394;
  assign n36396 = pi21 ? n2106 : n428;
  assign n36397 = pi20 ? n19106 : n36396;
  assign n36398 = pi19 ? n36397 : n34462;
  assign n36399 = pi18 ? n37 : n36398;
  assign n36400 = pi17 ? n37 : n36399;
  assign n36401 = pi16 ? n32926 : n36400;
  assign n36402 = pi15 ? n36395 : n36401;
  assign n36403 = pi19 ? n31280 : n21611;
  assign n36404 = pi18 ? n31315 : n36403;
  assign n36405 = pi17 ? n32 : n36404;
  assign n36406 = pi20 ? n1665 : n14464;
  assign n36407 = pi19 ? n13069 : n36406;
  assign n36408 = pi20 ? n23980 : n32;
  assign n36409 = pi19 ? n157 : n36408;
  assign n36410 = pi18 ? n36407 : n36409;
  assign n36411 = pi17 ? n99 : n36410;
  assign n36412 = pi16 ? n36405 : n36411;
  assign n36413 = pi20 ? n14478 : n787;
  assign n36414 = pi19 ? n31280 : n36413;
  assign n36415 = pi18 ? n31315 : n36414;
  assign n36416 = pi17 ? n32 : n36415;
  assign n36417 = pi20 ? n6523 : n6508;
  assign n36418 = pi20 ? n802 : n6500;
  assign n36419 = pi19 ? n36417 : n36418;
  assign n36420 = pi20 ? n787 : n802;
  assign n36421 = pi19 ? n36420 : n1492;
  assign n36422 = pi18 ? n36419 : n36421;
  assign n36423 = pi20 ? n160 : n6523;
  assign n36424 = pi20 ? n2243 : n2238;
  assign n36425 = pi19 ? n36423 : n36424;
  assign n36426 = pi20 ? n24033 : n32;
  assign n36427 = pi19 ? n157 : n36426;
  assign n36428 = pi18 ? n36425 : n36427;
  assign n36429 = pi17 ? n36422 : n36428;
  assign n36430 = pi16 ? n36416 : n36429;
  assign n36431 = pi15 ? n36412 : n36430;
  assign n36432 = pi14 ? n36402 : n36431;
  assign n36433 = pi13 ? n36389 : n36432;
  assign n36434 = pi12 ? n36372 : n36433;
  assign n36435 = pi11 ? n36316 : n36434;
  assign n36436 = pi19 ? n33965 : n3050;
  assign n36437 = pi18 ? n31315 : n36436;
  assign n36438 = pi17 ? n32 : n36437;
  assign n36439 = pi20 ? n2238 : n10526;
  assign n36440 = pi21 ? n3013 : n168;
  assign n36441 = pi20 ? n36440 : n10534;
  assign n36442 = pi19 ? n36439 : n36441;
  assign n36443 = pi20 ? n9015 : n36440;
  assign n36444 = pi19 ? n36443 : n5881;
  assign n36445 = pi18 ? n36442 : n36444;
  assign n36446 = pi20 ? n7824 : n10532;
  assign n36447 = pi21 ? n159 : n3002;
  assign n36448 = pi21 ? n168 : n2998;
  assign n36449 = pi20 ? n36447 : n36448;
  assign n36450 = pi19 ? n36446 : n36449;
  assign n36451 = pi19 ? n6529 : n36426;
  assign n36452 = pi18 ? n36450 : n36451;
  assign n36453 = pi17 ? n36445 : n36452;
  assign n36454 = pi16 ? n36438 : n36453;
  assign n36455 = pi20 ? n5077 : n3046;
  assign n36456 = pi19 ? n17013 : n36455;
  assign n36457 = pi20 ? n6500 : n226;
  assign n36458 = pi19 ? n36457 : n1492;
  assign n36459 = pi18 ? n36456 : n36458;
  assign n36460 = pi21 ? n165 : n99;
  assign n36461 = pi20 ? n36460 : n157;
  assign n36462 = pi22 ? n112 : n158;
  assign n36463 = pi21 ? n36462 : n777;
  assign n36464 = pi20 ? n36463 : n2238;
  assign n36465 = pi19 ? n36461 : n36464;
  assign n36466 = pi19 ? n15271 : n10012;
  assign n36467 = pi18 ? n36465 : n36466;
  assign n36468 = pi17 ? n36459 : n36467;
  assign n36469 = pi16 ? n33968 : n36468;
  assign n36470 = pi15 ? n36454 : n36469;
  assign n36471 = pi18 ? n31315 : n14842;
  assign n36472 = pi17 ? n32 : n36471;
  assign n36473 = pi20 ? n7779 : n99;
  assign n36474 = pi19 ? n36473 : n2242;
  assign n36475 = pi21 ? n777 : n8640;
  assign n36476 = pi20 ? n36475 : n316;
  assign n36477 = pi19 ? n36476 : n10012;
  assign n36478 = pi18 ? n36474 : n36477;
  assign n36479 = pi17 ? n99 : n36478;
  assign n36480 = pi16 ? n36472 : n36479;
  assign n36481 = pi19 ? n20973 : n99;
  assign n36482 = pi20 ? n19171 : n316;
  assign n36483 = pi19 ? n36482 : n10012;
  assign n36484 = pi18 ? n36481 : n36483;
  assign n36485 = pi17 ? n99 : n36484;
  assign n36486 = pi16 ? n36472 : n36485;
  assign n36487 = pi15 ? n36480 : n36486;
  assign n36488 = pi14 ? n36470 : n36487;
  assign n36489 = pi22 ? n20563 : n30868;
  assign n36490 = pi21 ? n30866 : n36489;
  assign n36491 = pi20 ? n32 : n36490;
  assign n36492 = pi19 ? n32 : n36491;
  assign n36493 = pi20 ? n2974 : n99;
  assign n36494 = pi19 ? n36493 : n99;
  assign n36495 = pi18 ? n36492 : n36494;
  assign n36496 = pi17 ? n32 : n36495;
  assign n36497 = pi20 ? n24957 : n316;
  assign n36498 = pi19 ? n36497 : n10012;
  assign n36499 = pi18 ? n99 : n36498;
  assign n36500 = pi17 ? n99 : n36499;
  assign n36501 = pi16 ? n36496 : n36500;
  assign n36502 = pi18 ? n35959 : n37;
  assign n36503 = pi17 ? n32 : n36502;
  assign n36504 = pi18 ? n30851 : n22703;
  assign n36505 = pi21 ? n17375 : n316;
  assign n36506 = pi20 ? n36505 : n316;
  assign n36507 = pi19 ? n36506 : n10012;
  assign n36508 = pi18 ? n139 : n36507;
  assign n36509 = pi17 ? n36504 : n36508;
  assign n36510 = pi16 ? n36503 : n36509;
  assign n36511 = pi15 ? n36501 : n36510;
  assign n36512 = pi19 ? n5305 : n2654;
  assign n36513 = pi18 ? n139 : n36512;
  assign n36514 = pi17 ? n8767 : n36513;
  assign n36515 = pi16 ? n36503 : n36514;
  assign n36516 = pi22 ? n30868 : n37;
  assign n36517 = pi21 ? n31293 : n36516;
  assign n36518 = pi20 ? n32 : n36517;
  assign n36519 = pi19 ? n32 : n36518;
  assign n36520 = pi18 ? n36519 : n15003;
  assign n36521 = pi17 ? n32 : n36520;
  assign n36522 = pi18 ? n9770 : n139;
  assign n36523 = pi19 ? n4003 : n1823;
  assign n36524 = pi18 ? n139 : n36523;
  assign n36525 = pi17 ? n36522 : n36524;
  assign n36526 = pi16 ? n36521 : n36525;
  assign n36527 = pi15 ? n36515 : n36526;
  assign n36528 = pi14 ? n36511 : n36527;
  assign n36529 = pi13 ? n36488 : n36528;
  assign n36530 = pi18 ? n14115 : n139;
  assign n36531 = pi21 ? n204 : n7621;
  assign n36532 = pi20 ? n1016 : n36531;
  assign n36533 = pi19 ? n36532 : n32;
  assign n36534 = pi18 ? n139 : n36533;
  assign n36535 = pi17 ? n36530 : n36534;
  assign n36536 = pi16 ? n33409 : n36535;
  assign n36537 = pi19 ? n37 : n20722;
  assign n36538 = pi19 ? n139 : n21060;
  assign n36539 = pi18 ? n36537 : n36538;
  assign n36540 = pi20 ? n204 : n5204;
  assign n36541 = pi20 ? n139 : n6568;
  assign n36542 = pi19 ? n36540 : n36541;
  assign n36543 = pi20 ? n5926 : n36531;
  assign n36544 = pi19 ? n36543 : n32;
  assign n36545 = pi18 ? n36542 : n36544;
  assign n36546 = pi17 ? n36539 : n36545;
  assign n36547 = pi16 ? n33409 : n36546;
  assign n36548 = pi15 ? n36536 : n36547;
  assign n36549 = pi18 ? n9815 : n30556;
  assign n36550 = pi20 ? n2318 : n922;
  assign n36551 = pi19 ? n15405 : n36550;
  assign n36552 = pi21 ? n204 : n21337;
  assign n36553 = pi20 ? n204 : n36552;
  assign n36554 = pi19 ? n36553 : n32;
  assign n36555 = pi18 ? n36551 : n36554;
  assign n36556 = pi17 ? n36549 : n36555;
  assign n36557 = pi16 ? n33409 : n36556;
  assign n36558 = pi20 ? n3075 : n139;
  assign n36559 = pi19 ? n29273 : n36558;
  assign n36560 = pi18 ? n36559 : n30556;
  assign n36561 = pi19 ? n15405 : n13462;
  assign n36562 = pi21 ? n204 : n7637;
  assign n36563 = pi20 ? n204 : n36562;
  assign n36564 = pi19 ? n36563 : n32;
  assign n36565 = pi18 ? n36561 : n36564;
  assign n36566 = pi17 ? n36560 : n36565;
  assign n36567 = pi16 ? n32952 : n36566;
  assign n36568 = pi15 ? n36557 : n36567;
  assign n36569 = pi14 ? n36548 : n36568;
  assign n36570 = pi19 ? n139 : n204;
  assign n36571 = pi18 ? n17061 : n36570;
  assign n36572 = pi21 ? n204 : n21980;
  assign n36573 = pi20 ? n204 : n36572;
  assign n36574 = pi19 ? n36573 : n32;
  assign n36575 = pi18 ? n204 : n36574;
  assign n36576 = pi17 ? n36571 : n36575;
  assign n36577 = pi16 ? n32952 : n36576;
  assign n36578 = pi21 ? n9122 : n139;
  assign n36579 = pi20 ? n36578 : n139;
  assign n36580 = pi19 ? n16516 : n36579;
  assign n36581 = pi18 ? n37 : n36580;
  assign n36582 = pi22 ? n1038 : n233;
  assign n36583 = pi21 ? n139 : n36582;
  assign n36584 = pi22 ? n233 : n918;
  assign n36585 = pi21 ? n36584 : n19726;
  assign n36586 = pi20 ? n36583 : n36585;
  assign n36587 = pi19 ? n36586 : n32;
  assign n36588 = pi18 ? n139 : n36587;
  assign n36589 = pi17 ? n36581 : n36588;
  assign n36590 = pi16 ? n32952 : n36589;
  assign n36591 = pi15 ? n36577 : n36590;
  assign n36592 = pi18 ? n37 : n7707;
  assign n36593 = pi20 ? n233 : n37;
  assign n36594 = pi21 ? n4938 : n233;
  assign n36595 = pi20 ? n36594 : n233;
  assign n36596 = pi19 ? n36593 : n36595;
  assign n36597 = pi20 ? n233 : n26021;
  assign n36598 = pi19 ? n36597 : n32;
  assign n36599 = pi18 ? n36596 : n36598;
  assign n36600 = pi17 ? n36592 : n36599;
  assign n36601 = pi16 ? n32432 : n36600;
  assign n36602 = pi21 ? n4938 : n570;
  assign n36603 = pi20 ? n36602 : n8927;
  assign n36604 = pi19 ? n7695 : n36603;
  assign n36605 = pi21 ? n685 : n25174;
  assign n36606 = pi20 ? n233 : n36605;
  assign n36607 = pi19 ? n36606 : n32;
  assign n36608 = pi18 ? n36604 : n36607;
  assign n36609 = pi17 ? n37 : n36608;
  assign n36610 = pi16 ? n32415 : n36609;
  assign n36611 = pi15 ? n36601 : n36610;
  assign n36612 = pi14 ? n36591 : n36611;
  assign n36613 = pi13 ? n36569 : n36612;
  assign n36614 = pi12 ? n36529 : n36613;
  assign n36615 = pi23 ? n33792 : n20563;
  assign n36616 = pi22 ? n30865 : n36615;
  assign n36617 = pi23 ? n37 : n33792;
  assign n36618 = pi22 ? n36617 : n37;
  assign n36619 = pi21 ? n36616 : n36618;
  assign n36620 = pi20 ? n32 : n36619;
  assign n36621 = pi19 ? n32 : n36620;
  assign n36622 = pi18 ? n36621 : n37;
  assign n36623 = pi17 ? n32 : n36622;
  assign n36624 = pi19 ? n7695 : n37;
  assign n36625 = pi20 ? n13527 : n24135;
  assign n36626 = pi19 ? n36625 : n32;
  assign n36627 = pi18 ? n36624 : n36626;
  assign n36628 = pi17 ? n37 : n36627;
  assign n36629 = pi16 ? n36623 : n36628;
  assign n36630 = pi19 ? n6340 : n335;
  assign n36631 = pi21 ? n316 : n9202;
  assign n36632 = pi20 ? n6377 : n36631;
  assign n36633 = pi19 ? n36632 : n32;
  assign n36634 = pi18 ? n36630 : n36633;
  assign n36635 = pi17 ? n14165 : n36634;
  assign n36636 = pi16 ? n32014 : n36635;
  assign n36637 = pi15 ? n36629 : n36636;
  assign n36638 = pi18 ? n374 : n9856;
  assign n36639 = pi17 ? n32 : n36638;
  assign n36640 = pi20 ? n13527 : n20548;
  assign n36641 = pi19 ? n36640 : n32;
  assign n36642 = pi18 ? n335 : n36641;
  assign n36643 = pi17 ? n335 : n36642;
  assign n36644 = pi16 ? n36639 : n36643;
  assign n36645 = pi19 ? n17224 : n335;
  assign n36646 = pi18 ? n374 : n36645;
  assign n36647 = pi17 ? n32 : n36646;
  assign n36648 = pi20 ? n13527 : n13339;
  assign n36649 = pi19 ? n36648 : n32;
  assign n36650 = pi18 ? n335 : n36649;
  assign n36651 = pi17 ? n335 : n36650;
  assign n36652 = pi16 ? n36647 : n36651;
  assign n36653 = pi15 ? n36644 : n36652;
  assign n36654 = pi14 ? n36637 : n36653;
  assign n36655 = pi19 ? n6341 : n335;
  assign n36656 = pi18 ? n32012 : n36655;
  assign n36657 = pi17 ? n32 : n36656;
  assign n36658 = pi16 ? n36657 : n36651;
  assign n36659 = pi25 ? n334 : n32;
  assign n36660 = pi23 ? n36659 : n37;
  assign n36661 = pi22 ? n31292 : n36660;
  assign n36662 = pi21 ? n36661 : n37;
  assign n36663 = pi20 ? n32 : n36662;
  assign n36664 = pi19 ? n32 : n36663;
  assign n36665 = pi19 ? n27685 : n335;
  assign n36666 = pi18 ? n36664 : n36665;
  assign n36667 = pi17 ? n32 : n36666;
  assign n36668 = pi20 ? n233 : n13339;
  assign n36669 = pi19 ? n36668 : n32;
  assign n36670 = pi18 ? n335 : n36669;
  assign n36671 = pi17 ? n335 : n36670;
  assign n36672 = pi16 ? n36667 : n36671;
  assign n36673 = pi15 ? n36658 : n36672;
  assign n36674 = pi19 ? n37 : n24865;
  assign n36675 = pi20 ? n21220 : n233;
  assign n36676 = pi19 ? n363 : n36675;
  assign n36677 = pi18 ? n36674 : n36676;
  assign n36678 = pi20 ? n23179 : n21222;
  assign n36679 = pi19 ? n36678 : n19434;
  assign n36680 = pi20 ? n30361 : n27076;
  assign n36681 = pi19 ? n36680 : n32;
  assign n36682 = pi18 ? n36679 : n36681;
  assign n36683 = pi17 ? n36677 : n36682;
  assign n36684 = pi16 ? n30201 : n36683;
  assign n36685 = pi23 ? n38 : n33792;
  assign n36686 = pi22 ? n36685 : n30195;
  assign n36687 = pi21 ? n36686 : n375;
  assign n36688 = pi20 ? n32 : n36687;
  assign n36689 = pi19 ? n32 : n36688;
  assign n36690 = pi18 ? n36689 : n37;
  assign n36691 = pi17 ? n32 : n36690;
  assign n36692 = pi20 ? n7730 : n22881;
  assign n36693 = pi19 ? n36692 : n363;
  assign n36694 = pi20 ? n363 : n26890;
  assign n36695 = pi19 ? n363 : n36694;
  assign n36696 = pi18 ? n36693 : n36695;
  assign n36697 = pi20 ? n26891 : n363;
  assign n36698 = pi20 ? n24220 : n25199;
  assign n36699 = pi19 ? n36697 : n36698;
  assign n36700 = pi20 ? n685 : n27076;
  assign n36701 = pi19 ? n36700 : n32;
  assign n36702 = pi18 ? n36699 : n36701;
  assign n36703 = pi17 ? n36696 : n36702;
  assign n36704 = pi16 ? n36691 : n36703;
  assign n36705 = pi15 ? n36684 : n36704;
  assign n36706 = pi14 ? n36673 : n36705;
  assign n36707 = pi13 ? n36654 : n36706;
  assign n36708 = pi23 ? n38 : n36659;
  assign n36709 = pi22 ? n36708 : n30195;
  assign n36710 = pi23 ? n36659 : n335;
  assign n36711 = pi22 ? n36710 : n37;
  assign n36712 = pi21 ? n36709 : n36711;
  assign n36713 = pi20 ? n32 : n36712;
  assign n36714 = pi19 ? n32 : n36713;
  assign n36715 = pi19 ? n19092 : n363;
  assign n36716 = pi18 ? n36714 : n36715;
  assign n36717 = pi17 ? n32 : n36716;
  assign n36718 = pi20 ? n26905 : n363;
  assign n36719 = pi20 ? n20866 : n25199;
  assign n36720 = pi19 ? n36718 : n36719;
  assign n36721 = pi20 ? n685 : n14723;
  assign n36722 = pi19 ? n36721 : n32;
  assign n36723 = pi18 ? n36720 : n36722;
  assign n36724 = pi17 ? n363 : n36723;
  assign n36725 = pi16 ? n36717 : n36724;
  assign n36726 = pi18 ? n37 : n36722;
  assign n36727 = pi17 ? n37 : n36726;
  assign n36728 = pi16 ? n32014 : n36727;
  assign n36729 = pi15 ? n36725 : n36728;
  assign n36730 = pi23 ? n714 : n30868;
  assign n36731 = pi22 ? n36730 : n99;
  assign n36732 = pi21 ? n36731 : n99;
  assign n36733 = pi20 ? n32 : n36732;
  assign n36734 = pi19 ? n32 : n36733;
  assign n36735 = pi18 ? n36734 : n99;
  assign n36736 = pi17 ? n32 : n36735;
  assign n36737 = pi21 ? n363 : n4551;
  assign n36738 = pi20 ? n36737 : n25167;
  assign n36739 = pi19 ? n36738 : n29738;
  assign n36740 = pi18 ? n99 : n36739;
  assign n36741 = pi20 ? n363 : n25181;
  assign n36742 = pi20 ? n29686 : n25167;
  assign n36743 = pi19 ? n36741 : n36742;
  assign n36744 = pi20 ? n685 : n12925;
  assign n36745 = pi19 ? n36744 : n32;
  assign n36746 = pi18 ? n36743 : n36745;
  assign n36747 = pi17 ? n36740 : n36746;
  assign n36748 = pi16 ? n36736 : n36747;
  assign n36749 = pi20 ? n29686 : n363;
  assign n36750 = pi19 ? n25167 : n36749;
  assign n36751 = pi18 ? n99 : n36750;
  assign n36752 = pi20 ? n363 : n25167;
  assign n36753 = pi20 ? n685 : n13398;
  assign n36754 = pi19 ? n36753 : n32;
  assign n36755 = pi18 ? n36752 : n36754;
  assign n36756 = pi17 ? n36751 : n36755;
  assign n36757 = pi16 ? n36736 : n36756;
  assign n36758 = pi15 ? n36748 : n36757;
  assign n36759 = pi14 ? n36729 : n36758;
  assign n36760 = pi23 ? n961 : n33792;
  assign n36761 = pi22 ? n36760 : n33792;
  assign n36762 = pi23 ? n33792 : n139;
  assign n36763 = pi22 ? n36762 : n139;
  assign n36764 = pi21 ? n36761 : n36763;
  assign n36765 = pi20 ? n32 : n36764;
  assign n36766 = pi19 ? n32 : n36765;
  assign n36767 = pi18 ? n36766 : n139;
  assign n36768 = pi17 ? n32 : n36767;
  assign n36769 = pi20 ? n139 : n20605;
  assign n36770 = pi19 ? n36769 : n36697;
  assign n36771 = pi20 ? n363 : n26891;
  assign n36772 = pi20 ? n29741 : n25199;
  assign n36773 = pi19 ? n36771 : n36772;
  assign n36774 = pi18 ? n36770 : n36773;
  assign n36775 = pi21 ? n685 : n27813;
  assign n36776 = pi20 ? n2721 : n36775;
  assign n36777 = pi19 ? n25200 : n36776;
  assign n36778 = pi18 ? n36777 : n33742;
  assign n36779 = pi17 ? n36774 : n36778;
  assign n36780 = pi16 ? n36768 : n36779;
  assign n36781 = pi25 ? n362 : n32;
  assign n36782 = pi24 ? n32 : n36781;
  assign n36783 = pi23 ? n36782 : n36781;
  assign n36784 = pi22 ? n36783 : n36781;
  assign n36785 = pi23 ? n36781 : n139;
  assign n36786 = pi22 ? n36781 : n36785;
  assign n36787 = pi21 ? n36784 : n36786;
  assign n36788 = pi20 ? n32 : n36787;
  assign n36789 = pi19 ? n32 : n36788;
  assign n36790 = pi18 ? n36789 : n363;
  assign n36791 = pi17 ? n32 : n36790;
  assign n36792 = pi20 ? n25199 : n7724;
  assign n36793 = pi19 ? n36792 : n32;
  assign n36794 = pi18 ? n363 : n36793;
  assign n36795 = pi17 ? n363 : n36794;
  assign n36796 = pi16 ? n36791 : n36795;
  assign n36797 = pi15 ? n36780 : n36796;
  assign n36798 = pi25 ? n156 : n32;
  assign n36799 = pi23 ? n1590 : n36798;
  assign n36800 = pi22 ? n36799 : n36781;
  assign n36801 = pi23 ? n36781 : n335;
  assign n36802 = pi22 ? n36710 : n36801;
  assign n36803 = pi21 ? n36800 : n36802;
  assign n36804 = pi20 ? n32 : n36803;
  assign n36805 = pi19 ? n32 : n36804;
  assign n36806 = pi21 ? n7986 : n363;
  assign n36807 = pi20 ? n36806 : n363;
  assign n36808 = pi21 ? n5054 : n363;
  assign n36809 = pi20 ? n36808 : n34841;
  assign n36810 = pi19 ? n36807 : n36809;
  assign n36811 = pi18 ? n36805 : n36810;
  assign n36812 = pi17 ? n32 : n36811;
  assign n36813 = pi21 ? n363 : n5054;
  assign n36814 = pi20 ? n36813 : n363;
  assign n36815 = pi21 ? n5054 : n34833;
  assign n36816 = pi20 ? n5054 : n36815;
  assign n36817 = pi19 ? n36814 : n36816;
  assign n36818 = pi20 ? n36808 : n20866;
  assign n36819 = pi21 ? n14277 : n363;
  assign n36820 = pi20 ? n36819 : n25199;
  assign n36821 = pi19 ? n36818 : n36820;
  assign n36822 = pi18 ? n36817 : n36821;
  assign n36823 = pi21 ? n363 : n14277;
  assign n36824 = pi20 ? n36823 : n25199;
  assign n36825 = pi20 ? n20866 : n36808;
  assign n36826 = pi19 ? n36824 : n36825;
  assign n36827 = pi18 ? n36826 : n36793;
  assign n36828 = pi17 ? n36822 : n36827;
  assign n36829 = pi16 ? n36812 : n36828;
  assign n36830 = pi24 ? n32 : n36798;
  assign n36831 = pi23 ? n36830 : n36798;
  assign n36832 = pi22 ? n36831 : n36781;
  assign n36833 = pi22 ? n36798 : n36801;
  assign n36834 = pi21 ? n36832 : n36833;
  assign n36835 = pi20 ? n32 : n36834;
  assign n36836 = pi19 ? n32 : n36835;
  assign n36837 = pi22 ? n335 : n157;
  assign n36838 = pi21 ? n36837 : n157;
  assign n36839 = pi20 ? n335 : n36838;
  assign n36840 = pi19 ? n36839 : n157;
  assign n36841 = pi18 ? n36836 : n36840;
  assign n36842 = pi17 ? n32 : n36841;
  assign n36843 = pi21 ? n6461 : n157;
  assign n36844 = pi20 ? n157 : n36843;
  assign n36845 = pi19 ? n157 : n36844;
  assign n36846 = pi20 ? n35725 : n15272;
  assign n36847 = pi21 ? n685 : n6461;
  assign n36848 = pi20 ? n685 : n36847;
  assign n36849 = pi19 ? n36846 : n36848;
  assign n36850 = pi18 ? n36845 : n36849;
  assign n36851 = pi21 ? n14277 : n685;
  assign n36852 = pi20 ? n15272 : n36851;
  assign n36853 = pi19 ? n685 : n36852;
  assign n36854 = pi21 ? n20460 : n685;
  assign n36855 = pi20 ? n36854 : n7724;
  assign n36856 = pi19 ? n36855 : n32;
  assign n36857 = pi18 ? n36853 : n36856;
  assign n36858 = pi17 ? n36850 : n36857;
  assign n36859 = pi16 ? n36842 : n36858;
  assign n36860 = pi15 ? n36829 : n36859;
  assign n36861 = pi14 ? n36797 : n36860;
  assign n36862 = pi13 ? n36759 : n36861;
  assign n36863 = pi12 ? n36707 : n36862;
  assign n36864 = pi11 ? n36614 : n36863;
  assign n36865 = pi10 ? n36435 : n36864;
  assign n36866 = pi09 ? n36193 : n36865;
  assign n36867 = pi21 ? n32 : n30116;
  assign n36868 = pi20 ? n32 : n36867;
  assign n36869 = pi19 ? n32 : n36868;
  assign n36870 = pi18 ? n36869 : n20563;
  assign n36871 = pi17 ? n32 : n36870;
  assign n36872 = pi21 ? n20563 : n35230;
  assign n36873 = pi20 ? n20563 : n36872;
  assign n36874 = pi19 ? n36873 : n34261;
  assign n36875 = pi18 ? n36874 : n99;
  assign n36876 = pi17 ? n36875 : n36167;
  assign n36877 = pi16 ? n36871 : n36876;
  assign n36878 = pi15 ? n32 : n36877;
  assign n36879 = pi21 ? n31890 : n37;
  assign n36880 = pi20 ? n20563 : n36879;
  assign n36881 = pi19 ? n36880 : n36171;
  assign n36882 = pi18 ? n36881 : n99;
  assign n36883 = pi17 ? n36882 : n36177;
  assign n36884 = pi16 ? n34860 : n36883;
  assign n36885 = pi21 ? n30867 : n37;
  assign n36886 = pi20 ? n20563 : n36885;
  assign n36887 = pi19 ? n36886 : n34261;
  assign n36888 = pi18 ? n36887 : n99;
  assign n36889 = pi17 ? n36888 : n36185;
  assign n36890 = pi16 ? n34860 : n36889;
  assign n36891 = pi15 ? n36884 : n36890;
  assign n36892 = pi14 ? n36878 : n36891;
  assign n36893 = pi13 ? n32 : n36892;
  assign n36894 = pi12 ? n32 : n36893;
  assign n36895 = pi11 ? n32 : n36894;
  assign n36896 = pi10 ? n32 : n36895;
  assign n36897 = pi20 ? n31925 : n31903;
  assign n36898 = pi19 ? n36897 : n34261;
  assign n36899 = pi18 ? n36898 : n99;
  assign n36900 = pi17 ? n36899 : n36198;
  assign n36901 = pi16 ? n35765 : n36900;
  assign n36902 = pi19 ? n32287 : n23648;
  assign n36903 = pi18 ? n36902 : n18854;
  assign n36904 = pi17 ? n36903 : n36206;
  assign n36905 = pi16 ? n35765 : n36904;
  assign n36906 = pi15 ? n36901 : n36905;
  assign n36907 = pi18 ? n33976 : n37;
  assign n36908 = pi17 ? n36907 : n36212;
  assign n36909 = pi16 ? n35765 : n36908;
  assign n36910 = pi22 ? n37 : n13969;
  assign n36911 = pi21 ? n36910 : n32;
  assign n36912 = pi20 ? n36911 : n32;
  assign n36913 = pi19 ? n37 : n36912;
  assign n36914 = pi18 ? n37 : n36913;
  assign n36915 = pi17 ? n36210 : n36914;
  assign n36916 = pi16 ? n36216 : n36915;
  assign n36917 = pi15 ? n36909 : n36916;
  assign n36918 = pi14 ? n36906 : n36917;
  assign n36919 = pi18 ? n31300 : n37;
  assign n36920 = pi17 ? n36919 : n36223;
  assign n36921 = pi16 ? n36216 : n36920;
  assign n36922 = pi18 ? n31315 : n34865;
  assign n36923 = pi17 ? n32 : n36922;
  assign n36924 = pi19 ? n139 : n8749;
  assign n36925 = pi18 ? n139 : n36924;
  assign n36926 = pi17 ? n36228 : n36925;
  assign n36927 = pi16 ? n36923 : n36926;
  assign n36928 = pi15 ? n36921 : n36927;
  assign n36929 = pi21 ? n20563 : n30867;
  assign n36930 = pi20 ? n20563 : n36929;
  assign n36931 = pi19 ? n20563 : n36930;
  assign n36932 = pi18 ? n31315 : n36931;
  assign n36933 = pi17 ? n32 : n36932;
  assign n36934 = pi19 ? n16023 : n8749;
  assign n36935 = pi18 ? n139 : n36934;
  assign n36936 = pi17 ? n9816 : n36935;
  assign n36937 = pi16 ? n36933 : n36936;
  assign n36938 = pi20 ? n21305 : n32;
  assign n36939 = pi19 ? n139 : n36938;
  assign n36940 = pi18 ? n139 : n36939;
  assign n36941 = pi17 ? n36241 : n36940;
  assign n36942 = pi16 ? n36227 : n36941;
  assign n36943 = pi15 ? n36937 : n36942;
  assign n36944 = pi14 ? n36928 : n36943;
  assign n36945 = pi13 ? n36918 : n36944;
  assign n36946 = pi21 ? n31885 : n30843;
  assign n36947 = pi20 ? n20563 : n36946;
  assign n36948 = pi19 ? n20563 : n36947;
  assign n36949 = pi18 ? n31315 : n36948;
  assign n36950 = pi17 ? n32 : n36949;
  assign n36951 = pi19 ? n9769 : n36938;
  assign n36952 = pi18 ? n139 : n36951;
  assign n36953 = pi17 ? n36256 : n36952;
  assign n36954 = pi16 ? n36950 : n36953;
  assign n36955 = pi18 ? n31938 : n33245;
  assign n36956 = pi17 ? n32 : n36955;
  assign n36957 = pi20 ? n21320 : n32;
  assign n36958 = pi19 ? n9769 : n36957;
  assign n36959 = pi18 ? n139 : n36958;
  assign n36960 = pi17 ? n36260 : n36959;
  assign n36961 = pi16 ? n36956 : n36960;
  assign n36962 = pi15 ? n36954 : n36961;
  assign n36963 = pi21 ? n17755 : n32;
  assign n36964 = pi20 ? n36963 : n32;
  assign n36965 = pi19 ? n11827 : n36964;
  assign n36966 = pi18 ? n22047 : n36965;
  assign n36967 = pi17 ? n37 : n36966;
  assign n36968 = pi16 ? n35244 : n36967;
  assign n36969 = pi21 ? n17741 : n32;
  assign n36970 = pi20 ? n36969 : n32;
  assign n36971 = pi19 ? n17204 : n36970;
  assign n36972 = pi18 ? n37 : n36971;
  assign n36973 = pi17 ? n37 : n36972;
  assign n36974 = pi16 ? n35244 : n36973;
  assign n36975 = pi15 ? n36968 : n36974;
  assign n36976 = pi14 ? n36962 : n36975;
  assign n36977 = pi21 ? n20563 : n31890;
  assign n36978 = pi20 ? n36977 : n37;
  assign n36979 = pi19 ? n20563 : n36978;
  assign n36980 = pi18 ? n31315 : n36979;
  assign n36981 = pi17 ? n32 : n36980;
  assign n36982 = pi22 ? n99 : n705;
  assign n36983 = pi21 ? n36982 : n32;
  assign n36984 = pi20 ? n36983 : n32;
  assign n36985 = pi19 ? n17204 : n36984;
  assign n36986 = pi18 ? n37 : n36985;
  assign n36987 = pi17 ? n37 : n36986;
  assign n36988 = pi16 ? n36981 : n36987;
  assign n36989 = pi22 ? n112 : n6114;
  assign n36990 = pi21 ? n36989 : n32;
  assign n36991 = pi20 ? n36990 : n32;
  assign n36992 = pi19 ? n37 : n36991;
  assign n36993 = pi18 ? n37 : n36992;
  assign n36994 = pi17 ? n37 : n36993;
  assign n36995 = pi16 ? n34889 : n36994;
  assign n36996 = pi15 ? n36988 : n36995;
  assign n36997 = pi19 ? n2095 : n10298;
  assign n36998 = pi18 ? n37 : n36997;
  assign n36999 = pi17 ? n37 : n36998;
  assign n37000 = pi16 ? n34319 : n36999;
  assign n37001 = pi22 ? n31993 : n20563;
  assign n37002 = pi21 ? n37001 : n20563;
  assign n37003 = pi20 ? n32 : n37002;
  assign n37004 = pi19 ? n32 : n37003;
  assign n37005 = pi18 ? n37004 : n32295;
  assign n37006 = pi17 ? n32 : n37005;
  assign n37007 = pi16 ? n37006 : n36311;
  assign n37008 = pi15 ? n37000 : n37007;
  assign n37009 = pi14 ? n36996 : n37008;
  assign n37010 = pi13 ? n36976 : n37009;
  assign n37011 = pi12 ? n36945 : n37010;
  assign n37012 = pi16 ? n34335 : n36324;
  assign n37013 = pi21 ? n28879 : n32;
  assign n37014 = pi20 ? n37013 : n32;
  assign n37015 = pi19 ? n335 : n37014;
  assign n37016 = pi18 ? n335 : n37015;
  assign n37017 = pi17 ? n36327 : n37016;
  assign n37018 = pi16 ? n33883 : n37017;
  assign n37019 = pi15 ? n37012 : n37018;
  assign n37020 = pi21 ? n35619 : n2007;
  assign n37021 = pi20 ? n7646 : n37020;
  assign n37022 = pi19 ? n37021 : n9944;
  assign n37023 = pi18 ? n32452 : n37022;
  assign n37024 = pi17 ? n37 : n37023;
  assign n37025 = pi16 ? n34360 : n37024;
  assign n37026 = pi16 ? n33332 : n36342;
  assign n37027 = pi15 ? n37025 : n37026;
  assign n37028 = pi14 ? n37019 : n37027;
  assign n37029 = pi19 ? n35776 : n37;
  assign n37030 = pi18 ? n31315 : n37029;
  assign n37031 = pi17 ? n32 : n37030;
  assign n37032 = pi16 ? n37031 : n36351;
  assign n37033 = pi16 ? n33918 : n36355;
  assign n37034 = pi15 ? n37032 : n37033;
  assign n37035 = pi16 ? n32351 : n36368;
  assign n37036 = pi15 ? n36361 : n37035;
  assign n37037 = pi14 ? n37034 : n37036;
  assign n37038 = pi13 ? n37028 : n37037;
  assign n37039 = pi19 ? n37 : n9457;
  assign n37040 = pi18 ? n37 : n37039;
  assign n37041 = pi17 ? n37 : n37040;
  assign n37042 = pi16 ? n32351 : n37041;
  assign n37043 = pi16 ? n31941 : n37041;
  assign n37044 = pi19 ? n36383 : n9964;
  assign n37045 = pi18 ? n37 : n37044;
  assign n37046 = pi17 ? n37 : n37045;
  assign n37047 = pi16 ? n31941 : n37046;
  assign n37048 = pi15 ? n37043 : n37047;
  assign n37049 = pi14 ? n37042 : n37048;
  assign n37050 = pi19 ? n36390 : n9964;
  assign n37051 = pi18 ? n37 : n37050;
  assign n37052 = pi17 ? n37 : n37051;
  assign n37053 = pi16 ? n31941 : n37052;
  assign n37054 = pi19 ? n32287 : n37;
  assign n37055 = pi18 ? n31315 : n37054;
  assign n37056 = pi17 ? n32 : n37055;
  assign n37057 = pi20 ? n37 : n36396;
  assign n37058 = pi19 ? n37057 : n7734;
  assign n37059 = pi18 ? n37 : n37058;
  assign n37060 = pi17 ? n37 : n37059;
  assign n37061 = pi16 ? n37056 : n37060;
  assign n37062 = pi15 ? n37053 : n37061;
  assign n37063 = pi19 ? n157 : n7734;
  assign n37064 = pi18 ? n36407 : n37063;
  assign n37065 = pi17 ? n99 : n37064;
  assign n37066 = pi16 ? n36405 : n37065;
  assign n37067 = pi20 ? n4625 : n787;
  assign n37068 = pi19 ? n31280 : n37067;
  assign n37069 = pi18 ? n31315 : n37068;
  assign n37070 = pi17 ? n32 : n37069;
  assign n37071 = pi19 ? n157 : n3978;
  assign n37072 = pi18 ? n36425 : n37071;
  assign n37073 = pi17 ? n36422 : n37072;
  assign n37074 = pi16 ? n37070 : n37073;
  assign n37075 = pi15 ? n37066 : n37074;
  assign n37076 = pi14 ? n37062 : n37075;
  assign n37077 = pi13 ? n37049 : n37076;
  assign n37078 = pi12 ? n37038 : n37077;
  assign n37079 = pi11 ? n37011 : n37078;
  assign n37080 = pi19 ? n31280 : n3050;
  assign n37081 = pi18 ? n31938 : n37080;
  assign n37082 = pi17 ? n32 : n37081;
  assign n37083 = pi21 ? n35988 : n168;
  assign n37084 = pi19 ? n36443 : n37083;
  assign n37085 = pi18 ? n36442 : n37084;
  assign n37086 = pi20 ? n7104 : n10532;
  assign n37087 = pi21 ? n99 : n3002;
  assign n37088 = pi20 ? n37087 : n36448;
  assign n37089 = pi19 ? n37086 : n37088;
  assign n37090 = pi19 ? n6529 : n3978;
  assign n37091 = pi18 ? n37089 : n37090;
  assign n37092 = pi17 ? n37085 : n37091;
  assign n37093 = pi16 ? n37082 : n37092;
  assign n37094 = pi19 ? n19134 : n36464;
  assign n37095 = pi19 ? n15271 : n3211;
  assign n37096 = pi18 ? n37094 : n37095;
  assign n37097 = pi17 ? n36459 : n37096;
  assign n37098 = pi16 ? n33952 : n37097;
  assign n37099 = pi15 ? n37093 : n37098;
  assign n37100 = pi19 ? n31299 : n99;
  assign n37101 = pi18 ? n31315 : n37100;
  assign n37102 = pi17 ? n32 : n37101;
  assign n37103 = pi19 ? n36476 : n12193;
  assign n37104 = pi18 ? n36474 : n37103;
  assign n37105 = pi17 ? n99 : n37104;
  assign n37106 = pi16 ? n37102 : n37105;
  assign n37107 = pi19 ? n32933 : n99;
  assign n37108 = pi18 ? n31938 : n37107;
  assign n37109 = pi17 ? n32 : n37108;
  assign n37110 = pi19 ? n36482 : n12193;
  assign n37111 = pi18 ? n36481 : n37110;
  assign n37112 = pi17 ? n99 : n37111;
  assign n37113 = pi16 ? n37109 : n37112;
  assign n37114 = pi15 ? n37106 : n37113;
  assign n37115 = pi14 ? n37099 : n37114;
  assign n37116 = pi20 ? n31903 : n99;
  assign n37117 = pi19 ? n37116 : n99;
  assign n37118 = pi18 ? n36492 : n37117;
  assign n37119 = pi17 ? n32 : n37118;
  assign n37120 = pi16 ? n37119 : n36500;
  assign n37121 = pi16 ? n32936 : n36509;
  assign n37122 = pi15 ? n37120 : n37121;
  assign n37123 = pi16 ? n32936 : n36514;
  assign n37124 = pi22 ? n30868 : n30867;
  assign n37125 = pi21 ? n30866 : n37124;
  assign n37126 = pi20 ? n32 : n37125;
  assign n37127 = pi19 ? n32 : n37126;
  assign n37128 = pi18 ? n37127 : n15003;
  assign n37129 = pi17 ? n32 : n37128;
  assign n37130 = pi16 ? n37129 : n36525;
  assign n37131 = pi15 ? n37123 : n37130;
  assign n37132 = pi14 ? n37122 : n37131;
  assign n37133 = pi13 ? n37115 : n37132;
  assign n37134 = pi20 ? n1016 : n25056;
  assign n37135 = pi19 ? n37134 : n32;
  assign n37136 = pi18 ? n139 : n37135;
  assign n37137 = pi17 ? n36530 : n37136;
  assign n37138 = pi16 ? n31317 : n37137;
  assign n37139 = pi20 ? n5926 : n25056;
  assign n37140 = pi19 ? n37139 : n32;
  assign n37141 = pi18 ? n36542 : n37140;
  assign n37142 = pi17 ? n36539 : n37141;
  assign n37143 = pi16 ? n31317 : n37142;
  assign n37144 = pi15 ? n37138 : n37143;
  assign n37145 = pi20 ? n204 : n24067;
  assign n37146 = pi19 ? n37145 : n32;
  assign n37147 = pi18 ? n36551 : n37146;
  assign n37148 = pi17 ? n36549 : n37147;
  assign n37149 = pi16 ? n36503 : n37148;
  assign n37150 = pi21 ? n204 : n1071;
  assign n37151 = pi20 ? n204 : n37150;
  assign n37152 = pi19 ? n37151 : n32;
  assign n37153 = pi18 ? n36561 : n37152;
  assign n37154 = pi17 ? n36560 : n37153;
  assign n37155 = pi16 ? n34999 : n37154;
  assign n37156 = pi15 ? n37149 : n37155;
  assign n37157 = pi14 ? n37144 : n37156;
  assign n37158 = pi16 ? n36503 : n36576;
  assign n37159 = pi21 ? n139 : n28649;
  assign n37160 = pi21 ? n34660 : n19726;
  assign n37161 = pi20 ? n37159 : n37160;
  assign n37162 = pi19 ? n37161 : n32;
  assign n37163 = pi18 ? n139 : n37162;
  assign n37164 = pi17 ? n36581 : n37163;
  assign n37165 = pi16 ? n36503 : n37164;
  assign n37166 = pi15 ? n37158 : n37165;
  assign n37167 = pi16 ? n34001 : n36600;
  assign n37168 = pi16 ? n33409 : n36609;
  assign n37169 = pi15 ? n37167 : n37168;
  assign n37170 = pi14 ? n37166 : n37169;
  assign n37171 = pi13 ? n37157 : n37170;
  assign n37172 = pi12 ? n37133 : n37171;
  assign n37173 = pi23 ? n20563 : n33792;
  assign n37174 = pi22 ? n37173 : n37;
  assign n37175 = pi21 ? n30866 : n37174;
  assign n37176 = pi20 ? n32 : n37175;
  assign n37177 = pi19 ? n32 : n37176;
  assign n37178 = pi18 ? n37177 : n37;
  assign n37179 = pi17 ? n32 : n37178;
  assign n37180 = pi16 ? n37179 : n36628;
  assign n37181 = pi16 ? n35006 : n36635;
  assign n37182 = pi15 ? n37180 : n37181;
  assign n37183 = pi18 ? n30199 : n9856;
  assign n37184 = pi17 ? n32 : n37183;
  assign n37185 = pi20 ? n13527 : n21182;
  assign n37186 = pi19 ? n37185 : n32;
  assign n37187 = pi18 ? n335 : n37186;
  assign n37188 = pi17 ? n335 : n37187;
  assign n37189 = pi16 ? n37184 : n37188;
  assign n37190 = pi18 ? n32430 : n36645;
  assign n37191 = pi17 ? n32 : n37190;
  assign n37192 = pi16 ? n37191 : n37188;
  assign n37193 = pi15 ? n37189 : n37192;
  assign n37194 = pi14 ? n37182 : n37193;
  assign n37195 = pi18 ? n35004 : n36655;
  assign n37196 = pi17 ? n32 : n37195;
  assign n37197 = pi16 ? n37196 : n36643;
  assign n37198 = pi22 ? n30865 : n36660;
  assign n37199 = pi21 ? n37198 : n30843;
  assign n37200 = pi20 ? n32 : n37199;
  assign n37201 = pi19 ? n32 : n37200;
  assign n37202 = pi18 ? n37201 : n36665;
  assign n37203 = pi17 ? n32 : n37202;
  assign n37204 = pi20 ? n233 : n20548;
  assign n37205 = pi19 ? n37204 : n32;
  assign n37206 = pi18 ? n335 : n37205;
  assign n37207 = pi17 ? n335 : n37206;
  assign n37208 = pi16 ? n37203 : n37207;
  assign n37209 = pi15 ? n37197 : n37208;
  assign n37210 = pi21 ? n37001 : n30843;
  assign n37211 = pi20 ? n32 : n37210;
  assign n37212 = pi19 ? n32 : n37211;
  assign n37213 = pi18 ? n37212 : n37;
  assign n37214 = pi17 ? n32 : n37213;
  assign n37215 = pi16 ? n37214 : n36683;
  assign n37216 = pi23 ? n20564 : n33792;
  assign n37217 = pi22 ? n37216 : n20563;
  assign n37218 = pi23 ? n20563 : n139;
  assign n37219 = pi22 ? n37218 : n37;
  assign n37220 = pi21 ? n37217 : n37219;
  assign n37221 = pi20 ? n32 : n37220;
  assign n37222 = pi19 ? n32 : n37221;
  assign n37223 = pi18 ? n37222 : n37;
  assign n37224 = pi17 ? n32 : n37223;
  assign n37225 = pi16 ? n37224 : n36703;
  assign n37226 = pi15 ? n37215 : n37225;
  assign n37227 = pi14 ? n37209 : n37226;
  assign n37228 = pi13 ? n37194 : n37227;
  assign n37229 = pi23 ? n20564 : n36659;
  assign n37230 = pi22 ? n37229 : n20563;
  assign n37231 = pi22 ? n36659 : n37;
  assign n37232 = pi21 ? n37230 : n37231;
  assign n37233 = pi20 ? n32 : n37232;
  assign n37234 = pi19 ? n32 : n37233;
  assign n37235 = pi18 ? n37234 : n36715;
  assign n37236 = pi17 ? n32 : n37235;
  assign n37237 = pi16 ? n37236 : n36724;
  assign n37238 = pi16 ? n31987 : n36727;
  assign n37239 = pi15 ? n37237 : n37238;
  assign n37240 = pi23 ? n99 : n30868;
  assign n37241 = pi22 ? n36730 : n37240;
  assign n37242 = pi21 ? n37241 : n99;
  assign n37243 = pi20 ? n32 : n37242;
  assign n37244 = pi19 ? n32 : n37243;
  assign n37245 = pi18 ? n37244 : n99;
  assign n37246 = pi17 ? n32 : n37245;
  assign n37247 = pi16 ? n37246 : n36747;
  assign n37248 = pi16 ? n37246 : n36756;
  assign n37249 = pi15 ? n37247 : n37248;
  assign n37250 = pi14 ? n37239 : n37249;
  assign n37251 = pi23 ? n33793 : n33792;
  assign n37252 = pi22 ? n37251 : n33792;
  assign n37253 = pi22 ? n33792 : n36762;
  assign n37254 = pi21 ? n37252 : n37253;
  assign n37255 = pi20 ? n32 : n37254;
  assign n37256 = pi19 ? n32 : n37255;
  assign n37257 = pi18 ? n37256 : n139;
  assign n37258 = pi17 ? n32 : n37257;
  assign n37259 = pi16 ? n37258 : n36779;
  assign n37260 = pi23 ? n33793 : n36781;
  assign n37261 = pi22 ? n37260 : n36781;
  assign n37262 = pi21 ? n37261 : n36781;
  assign n37263 = pi20 ? n32 : n37262;
  assign n37264 = pi19 ? n32 : n37263;
  assign n37265 = pi18 ? n37264 : n363;
  assign n37266 = pi17 ? n32 : n37265;
  assign n37267 = pi20 ? n25199 : n8295;
  assign n37268 = pi19 ? n37267 : n32;
  assign n37269 = pi18 ? n363 : n37268;
  assign n37270 = pi17 ? n363 : n37269;
  assign n37271 = pi16 ? n37266 : n37270;
  assign n37272 = pi15 ? n37259 : n37271;
  assign n37273 = pi24 ? n32 : n36659;
  assign n37274 = pi23 ? n37273 : n36798;
  assign n37275 = pi22 ? n37274 : n36781;
  assign n37276 = pi23 ? n36659 : n36798;
  assign n37277 = pi22 ? n37276 : n36781;
  assign n37278 = pi21 ? n37275 : n37277;
  assign n37279 = pi20 ? n32 : n37278;
  assign n37280 = pi19 ? n32 : n37279;
  assign n37281 = pi18 ? n37280 : n36810;
  assign n37282 = pi17 ? n32 : n37281;
  assign n37283 = pi20 ? n25199 : n9482;
  assign n37284 = pi19 ? n37283 : n32;
  assign n37285 = pi18 ? n36826 : n37284;
  assign n37286 = pi17 ? n36822 : n37285;
  assign n37287 = pi16 ? n37282 : n37286;
  assign n37288 = pi23 ? n36781 : n36659;
  assign n37289 = pi22 ? n36798 : n37288;
  assign n37290 = pi21 ? n37275 : n37289;
  assign n37291 = pi20 ? n32 : n37290;
  assign n37292 = pi19 ? n32 : n37291;
  assign n37293 = pi18 ? n37292 : n36840;
  assign n37294 = pi17 ? n32 : n37293;
  assign n37295 = pi20 ? n36854 : n9482;
  assign n37296 = pi19 ? n37295 : n32;
  assign n37297 = pi18 ? n36853 : n37296;
  assign n37298 = pi17 ? n36850 : n37297;
  assign n37299 = pi16 ? n37294 : n37298;
  assign n37300 = pi15 ? n37287 : n37299;
  assign n37301 = pi14 ? n37272 : n37300;
  assign n37302 = pi13 ? n37250 : n37301;
  assign n37303 = pi12 ? n37228 : n37302;
  assign n37304 = pi11 ? n37172 : n37303;
  assign n37305 = pi10 ? n37079 : n37304;
  assign n37306 = pi09 ? n36896 : n37305;
  assign n37307 = pi08 ? n36866 : n37306;
  assign n37308 = pi21 ? n20563 : n36249;
  assign n37309 = pi20 ? n20563 : n37308;
  assign n37310 = pi20 ? n30096 : n14844;
  assign n37311 = pi19 ? n37309 : n37310;
  assign n37312 = pi18 ? n37311 : n99;
  assign n37313 = pi21 ? n99 : n8008;
  assign n37314 = pi20 ? n37313 : n32;
  assign n37315 = pi19 ? n99 : n37314;
  assign n37316 = pi18 ? n99 : n37315;
  assign n37317 = pi17 ? n37312 : n37316;
  assign n37318 = pi16 ? n36871 : n37317;
  assign n37319 = pi15 ? n32 : n37318;
  assign n37320 = pi21 ? n32 : n20563;
  assign n37321 = pi20 ? n32 : n37320;
  assign n37322 = pi19 ? n32 : n37321;
  assign n37323 = pi18 ? n37322 : n20563;
  assign n37324 = pi17 ? n32 : n37323;
  assign n37325 = pi20 ? n30096 : n226;
  assign n37326 = pi19 ? n20563 : n37325;
  assign n37327 = pi18 ? n37326 : n99;
  assign n37328 = pi19 ? n99 : n8017;
  assign n37329 = pi18 ? n99 : n37328;
  assign n37330 = pi17 ? n37327 : n37329;
  assign n37331 = pi16 ? n37324 : n37330;
  assign n37332 = pi22 ? n32 : n30115;
  assign n37333 = pi21 ? n37332 : n20563;
  assign n37334 = pi20 ? n32 : n37333;
  assign n37335 = pi19 ? n32 : n37334;
  assign n37336 = pi18 ? n37335 : n20563;
  assign n37337 = pi17 ? n32 : n37336;
  assign n37338 = pi20 ? n37 : n3879;
  assign n37339 = pi19 ? n20563 : n37338;
  assign n37340 = pi18 ? n37339 : n99;
  assign n37341 = pi21 ? n746 : n8015;
  assign n37342 = pi20 ? n37341 : n32;
  assign n37343 = pi19 ? n99 : n37342;
  assign n37344 = pi18 ? n99 : n37343;
  assign n37345 = pi17 ? n37340 : n37344;
  assign n37346 = pi16 ? n37337 : n37345;
  assign n37347 = pi15 ? n37331 : n37346;
  assign n37348 = pi14 ? n37319 : n37347;
  assign n37349 = pi13 ? n32 : n37348;
  assign n37350 = pi12 ? n32 : n37349;
  assign n37351 = pi11 ? n32 : n37350;
  assign n37352 = pi10 ? n32 : n37351;
  assign n37353 = pi19 ? n20563 : n34261;
  assign n37354 = pi18 ? n37353 : n99;
  assign n37355 = pi21 ? n1657 : n8557;
  assign n37356 = pi20 ? n37355 : n32;
  assign n37357 = pi19 ? n99 : n37356;
  assign n37358 = pi18 ? n99 : n37357;
  assign n37359 = pi17 ? n37354 : n37358;
  assign n37360 = pi16 ? n34860 : n37359;
  assign n37361 = pi20 ? n31266 : n31220;
  assign n37362 = pi19 ? n37361 : n35209;
  assign n37363 = pi18 ? n37362 : n99;
  assign n37364 = pi22 ? n99 : n583;
  assign n37365 = pi21 ? n37364 : n8044;
  assign n37366 = pi20 ? n37365 : n32;
  assign n37367 = pi19 ? n99 : n37366;
  assign n37368 = pi18 ? n99 : n37367;
  assign n37369 = pi17 ? n37363 : n37368;
  assign n37370 = pi16 ? n35765 : n37369;
  assign n37371 = pi15 ? n37360 : n37370;
  assign n37372 = pi18 ? n34358 : n37;
  assign n37373 = pi19 ? n37 : n6808;
  assign n37374 = pi18 ? n37 : n37373;
  assign n37375 = pi17 ? n37372 : n37374;
  assign n37376 = pi16 ? n35765 : n37375;
  assign n37377 = pi18 ? n32349 : n37;
  assign n37378 = pi21 ? n6433 : n32;
  assign n37379 = pi20 ? n37378 : n32;
  assign n37380 = pi19 ? n37 : n37379;
  assign n37381 = pi18 ? n37 : n37380;
  assign n37382 = pi17 ? n37377 : n37381;
  assign n37383 = pi16 ? n36216 : n37382;
  assign n37384 = pi15 ? n37376 : n37383;
  assign n37385 = pi14 ? n37371 : n37384;
  assign n37386 = pi18 ? n31939 : n37;
  assign n37387 = pi23 ? n139 : n3145;
  assign n37388 = pi22 ? n139 : n37387;
  assign n37389 = pi21 ? n37388 : n32;
  assign n37390 = pi20 ? n37389 : n32;
  assign n37391 = pi19 ? n9814 : n37390;
  assign n37392 = pi18 ? n37 : n37391;
  assign n37393 = pi17 ? n37386 : n37392;
  assign n37394 = pi16 ? n36216 : n37393;
  assign n37395 = pi20 ? n37 : n1697;
  assign n37396 = pi19 ? n31267 : n37395;
  assign n37397 = pi18 ? n37396 : n139;
  assign n37398 = pi22 ? n139 : n25629;
  assign n37399 = pi21 ? n37398 : n32;
  assign n37400 = pi20 ? n37399 : n32;
  assign n37401 = pi19 ? n139 : n37400;
  assign n37402 = pi18 ? n139 : n37401;
  assign n37403 = pi17 ? n37397 : n37402;
  assign n37404 = pi16 ? n36216 : n37403;
  assign n37405 = pi15 ? n37394 : n37404;
  assign n37406 = pi19 ? n18912 : n139;
  assign n37407 = pi18 ? n32924 : n37406;
  assign n37408 = pi17 ? n37407 : n37402;
  assign n37409 = pi16 ? n36216 : n37408;
  assign n37410 = pi19 ? n29248 : n139;
  assign n37411 = pi18 ? n31300 : n37410;
  assign n37412 = pi22 ? n139 : n25653;
  assign n37413 = pi21 ? n37412 : n32;
  assign n37414 = pi20 ? n37413 : n32;
  assign n37415 = pi19 ? n139 : n37414;
  assign n37416 = pi18 ? n139 : n37415;
  assign n37417 = pi17 ? n37411 : n37416;
  assign n37418 = pi16 ? n36216 : n37417;
  assign n37419 = pi15 ? n37409 : n37418;
  assign n37420 = pi14 ? n37405 : n37419;
  assign n37421 = pi13 ? n37385 : n37420;
  assign n37422 = pi19 ? n9769 : n37414;
  assign n37423 = pi18 ? n139 : n37422;
  assign n37424 = pi17 ? n35254 : n37423;
  assign n37425 = pi16 ? n36216 : n37424;
  assign n37426 = pi18 ? n37 : n11551;
  assign n37427 = pi22 ? n139 : n33355;
  assign n37428 = pi21 ? n37427 : n32;
  assign n37429 = pi20 ? n37428 : n32;
  assign n37430 = pi19 ? n9769 : n37429;
  assign n37431 = pi18 ? n139 : n37430;
  assign n37432 = pi17 ? n37426 : n37431;
  assign n37433 = pi16 ? n36216 : n37432;
  assign n37434 = pi15 ? n37425 : n37433;
  assign n37435 = pi19 ? n28367 : n36964;
  assign n37436 = pi18 ? n22047 : n37435;
  assign n37437 = pi17 ? n37 : n37436;
  assign n37438 = pi16 ? n36235 : n37437;
  assign n37439 = pi21 ? n36249 : n29133;
  assign n37440 = pi20 ? n20563 : n37439;
  assign n37441 = pi19 ? n20563 : n37440;
  assign n37442 = pi18 ? n31315 : n37441;
  assign n37443 = pi17 ? n32 : n37442;
  assign n37444 = pi16 ? n37443 : n36973;
  assign n37445 = pi15 ? n37438 : n37444;
  assign n37446 = pi14 ? n37434 : n37445;
  assign n37447 = pi20 ? n638 : n4971;
  assign n37448 = pi19 ? n37 : n37447;
  assign n37449 = pi19 ? n17204 : n35768;
  assign n37450 = pi18 ? n37448 : n37449;
  assign n37451 = pi17 ? n37 : n37450;
  assign n37452 = pi16 ? n35220 : n37451;
  assign n37453 = pi19 ? n8928 : n18393;
  assign n37454 = pi18 ? n37 : n37453;
  assign n37455 = pi17 ? n37 : n37454;
  assign n37456 = pi16 ? n34884 : n37455;
  assign n37457 = pi15 ? n37452 : n37456;
  assign n37458 = pi21 ? n37 : n19386;
  assign n37459 = pi20 ? n37 : n37458;
  assign n37460 = pi19 ? n37459 : n18393;
  assign n37461 = pi18 ? n37 : n37460;
  assign n37462 = pi17 ? n37 : n37461;
  assign n37463 = pi16 ? n34889 : n37462;
  assign n37464 = pi19 ? n17204 : n8850;
  assign n37465 = pi18 ? n37 : n37464;
  assign n37466 = pi17 ? n37 : n37465;
  assign n37467 = pi16 ? n34335 : n37466;
  assign n37468 = pi15 ? n37463 : n37467;
  assign n37469 = pi14 ? n37457 : n37468;
  assign n37470 = pi13 ? n37446 : n37469;
  assign n37471 = pi12 ? n37421 : n37470;
  assign n37472 = pi19 ? n17224 : n577;
  assign n37473 = pi18 ? n37 : n37472;
  assign n37474 = pi19 ? n16516 : n31719;
  assign n37475 = pi20 ? n22836 : n32;
  assign n37476 = pi19 ? n335 : n37475;
  assign n37477 = pi18 ? n37474 : n37476;
  assign n37478 = pi17 ? n37473 : n37477;
  assign n37479 = pi16 ? n34889 : n37478;
  assign n37480 = pi18 ? n37 : n4985;
  assign n37481 = pi21 ? n3693 : n32;
  assign n37482 = pi20 ? n37481 : n32;
  assign n37483 = pi19 ? n335 : n37482;
  assign n37484 = pi18 ? n335 : n37483;
  assign n37485 = pi17 ? n37480 : n37484;
  assign n37486 = pi16 ? n34335 : n37485;
  assign n37487 = pi15 ? n37479 : n37486;
  assign n37488 = pi18 ? n31938 : n33285;
  assign n37489 = pi17 ? n32 : n37488;
  assign n37490 = pi22 ? n363 : n6405;
  assign n37491 = pi21 ? n37490 : n32;
  assign n37492 = pi20 ? n37491 : n32;
  assign n37493 = pi19 ? n29357 : n37492;
  assign n37494 = pi18 ? n37 : n37493;
  assign n37495 = pi17 ? n37 : n37494;
  assign n37496 = pi16 ? n37489 : n37495;
  assign n37497 = pi20 ? n24466 : n32;
  assign n37498 = pi19 ? n23917 : n37497;
  assign n37499 = pi18 ? n37 : n37498;
  assign n37500 = pi17 ? n37 : n37499;
  assign n37501 = pi16 ? n34889 : n37500;
  assign n37502 = pi15 ? n37496 : n37501;
  assign n37503 = pi14 ? n37487 : n37502;
  assign n37504 = pi19 ? n27443 : n5013;
  assign n37505 = pi18 ? n37 : n37504;
  assign n37506 = pi21 ? n3392 : n5012;
  assign n37507 = pi20 ? n37506 : n15173;
  assign n37508 = pi20 ? n9654 : n19091;
  assign n37509 = pi19 ? n37507 : n37508;
  assign n37510 = pi20 ? n3392 : n363;
  assign n37511 = pi19 ? n37510 : n37497;
  assign n37512 = pi18 ? n37509 : n37511;
  assign n37513 = pi17 ? n37505 : n37512;
  assign n37514 = pi16 ? n34335 : n37513;
  assign n37515 = pi22 ? n363 : n3318;
  assign n37516 = pi21 ? n37515 : n32;
  assign n37517 = pi20 ? n37516 : n32;
  assign n37518 = pi19 ? n37 : n37517;
  assign n37519 = pi18 ? n37 : n37518;
  assign n37520 = pi17 ? n37 : n37519;
  assign n37521 = pi16 ? n33313 : n37520;
  assign n37522 = pi15 ? n37514 : n37521;
  assign n37523 = pi22 ? n363 : n430;
  assign n37524 = pi21 ? n37523 : n32;
  assign n37525 = pi20 ? n37524 : n32;
  assign n37526 = pi19 ? n37 : n37525;
  assign n37527 = pi18 ? n37 : n37526;
  assign n37528 = pi17 ? n37 : n37527;
  assign n37529 = pi16 ? n34335 : n37528;
  assign n37530 = pi19 ? n27535 : n9944;
  assign n37531 = pi18 ? n37 : n37530;
  assign n37532 = pi17 ? n37 : n37531;
  assign n37533 = pi16 ? n34923 : n37532;
  assign n37534 = pi15 ? n37529 : n37533;
  assign n37535 = pi14 ? n37522 : n37534;
  assign n37536 = pi13 ? n37503 : n37535;
  assign n37537 = pi16 ? n34360 : n37041;
  assign n37538 = pi16 ? n33918 : n37041;
  assign n37539 = pi21 ? n685 : n37;
  assign n37540 = pi20 ? n37 : n37539;
  assign n37541 = pi19 ? n37540 : n9964;
  assign n37542 = pi18 ? n37 : n37541;
  assign n37543 = pi17 ? n37 : n37542;
  assign n37544 = pi16 ? n33918 : n37543;
  assign n37545 = pi15 ? n37538 : n37544;
  assign n37546 = pi14 ? n37537 : n37545;
  assign n37547 = pi22 ? n685 : n14363;
  assign n37548 = pi21 ? n37547 : n32;
  assign n37549 = pi20 ? n37548 : n32;
  assign n37550 = pi19 ? n37540 : n37549;
  assign n37551 = pi18 ? n37 : n37550;
  assign n37552 = pi17 ? n37 : n37551;
  assign n37553 = pi16 ? n32901 : n37552;
  assign n37554 = pi19 ? n37 : n3211;
  assign n37555 = pi18 ? n37 : n37554;
  assign n37556 = pi17 ? n37 : n37555;
  assign n37557 = pi16 ? n34951 : n37556;
  assign n37558 = pi15 ? n37553 : n37557;
  assign n37559 = pi19 ? n32898 : n21611;
  assign n37560 = pi18 ? n31938 : n37559;
  assign n37561 = pi17 ? n32 : n37560;
  assign n37562 = pi20 ? n2238 : n2243;
  assign n37563 = pi19 ? n37562 : n99;
  assign n37564 = pi18 ? n37563 : n37063;
  assign n37565 = pi17 ? n99 : n37564;
  assign n37566 = pi16 ? n37561 : n37565;
  assign n37567 = pi19 ? n33923 : n18853;
  assign n37568 = pi18 ? n31315 : n37567;
  assign n37569 = pi17 ? n32 : n37568;
  assign n37570 = pi18 ? n99 : n9716;
  assign n37571 = pi19 ? n6532 : n3211;
  assign n37572 = pi18 ? n19145 : n37571;
  assign n37573 = pi17 ? n37570 : n37572;
  assign n37574 = pi16 ? n37569 : n37573;
  assign n37575 = pi15 ? n37566 : n37574;
  assign n37576 = pi14 ? n37558 : n37575;
  assign n37577 = pi13 ? n37546 : n37576;
  assign n37578 = pi12 ? n37536 : n37577;
  assign n37579 = pi11 ? n37471 : n37578;
  assign n37580 = pi19 ? n31267 : n21611;
  assign n37581 = pi18 ? n31315 : n37580;
  assign n37582 = pi17 ? n32 : n37581;
  assign n37583 = pi19 ? n2242 : n99;
  assign n37584 = pi19 ? n13069 : n3978;
  assign n37585 = pi18 ? n37583 : n37584;
  assign n37586 = pi17 ? n37570 : n37585;
  assign n37587 = pi16 ? n37582 : n37586;
  assign n37588 = pi19 ? n31267 : n18853;
  assign n37589 = pi18 ? n31938 : n37588;
  assign n37590 = pi17 ? n32 : n37589;
  assign n37591 = pi21 ? n8640 : n157;
  assign n37592 = pi20 ? n2243 : n37591;
  assign n37593 = pi19 ? n37592 : n3211;
  assign n37594 = pi18 ? n37583 : n37593;
  assign n37595 = pi17 ? n99 : n37594;
  assign n37596 = pi16 ? n37590 : n37595;
  assign n37597 = pi15 ? n37587 : n37596;
  assign n37598 = pi19 ? n31267 : n99;
  assign n37599 = pi18 ? n31938 : n37598;
  assign n37600 = pi17 ? n32 : n37599;
  assign n37601 = pi22 ? n19177 : n99;
  assign n37602 = pi23 ? n316 : n99;
  assign n37603 = pi22 ? n37602 : n157;
  assign n37604 = pi21 ? n37601 : n37603;
  assign n37605 = pi20 ? n37604 : n316;
  assign n37606 = pi19 ? n37605 : n3211;
  assign n37607 = pi18 ? n99 : n37606;
  assign n37608 = pi17 ? n99 : n37607;
  assign n37609 = pi16 ? n37600 : n37608;
  assign n37610 = pi18 ? n31315 : n37598;
  assign n37611 = pi17 ? n32 : n37610;
  assign n37612 = pi19 ? n36497 : n3211;
  assign n37613 = pi18 ? n99 : n37612;
  assign n37614 = pi17 ? n99 : n37613;
  assign n37615 = pi16 ? n37611 : n37614;
  assign n37616 = pi15 ? n37609 : n37615;
  assign n37617 = pi14 ? n37597 : n37616;
  assign n37618 = pi20 ? n31266 : n14844;
  assign n37619 = pi19 ? n37618 : n99;
  assign n37620 = pi18 ? n31315 : n37619;
  assign n37621 = pi17 ? n32 : n37620;
  assign n37622 = pi16 ? n37621 : n37614;
  assign n37623 = pi21 ? n218 : n139;
  assign n37624 = pi20 ? n37623 : n139;
  assign n37625 = pi19 ? n37 : n37624;
  assign n37626 = pi21 ? n4237 : n139;
  assign n37627 = pi20 ? n139 : n37626;
  assign n37628 = pi19 ? n37627 : n139;
  assign n37629 = pi18 ? n37625 : n37628;
  assign n37630 = pi19 ? n5305 : n10012;
  assign n37631 = pi18 ? n139 : n37630;
  assign n37632 = pi17 ? n37629 : n37631;
  assign n37633 = pi16 ? n32379 : n37632;
  assign n37634 = pi15 ? n37622 : n37633;
  assign n37635 = pi16 ? n36365 : n36514;
  assign n37636 = pi19 ? n36362 : n8765;
  assign n37637 = pi18 ? n31315 : n37636;
  assign n37638 = pi17 ? n32 : n37637;
  assign n37639 = pi22 ? n21502 : n32;
  assign n37640 = pi21 ? n37639 : n32;
  assign n37641 = pi20 ? n37640 : n32;
  assign n37642 = pi19 ? n30527 : n37641;
  assign n37643 = pi18 ? n139 : n37642;
  assign n37644 = pi17 ? n139 : n37643;
  assign n37645 = pi16 ? n37638 : n37644;
  assign n37646 = pi15 ? n37635 : n37645;
  assign n37647 = pi14 ? n37634 : n37646;
  assign n37648 = pi13 ? n37617 : n37647;
  assign n37649 = pi19 ? n32871 : n37;
  assign n37650 = pi18 ? n31315 : n37649;
  assign n37651 = pi17 ? n32 : n37650;
  assign n37652 = pi19 ? n26742 : n32;
  assign n37653 = pi18 ? n6652 : n37652;
  assign n37654 = pi17 ? n36530 : n37653;
  assign n37655 = pi16 ? n37651 : n37654;
  assign n37656 = pi18 ? n14115 : n36538;
  assign n37657 = pi19 ? n36540 : n139;
  assign n37658 = pi19 ? n34641 : n32;
  assign n37659 = pi18 ? n37657 : n37658;
  assign n37660 = pi17 ? n37656 : n37659;
  assign n37661 = pi16 ? n32379 : n37660;
  assign n37662 = pi15 ? n37655 : n37661;
  assign n37663 = pi20 ? n6158 : n922;
  assign n37664 = pi19 ? n7454 : n37663;
  assign n37665 = pi19 ? n11810 : n32;
  assign n37666 = pi18 ? n37664 : n37665;
  assign n37667 = pi17 ? n36549 : n37666;
  assign n37668 = pi16 ? n35320 : n37667;
  assign n37669 = pi18 ? n14115 : n30556;
  assign n37670 = pi18 ? n36561 : n37665;
  assign n37671 = pi17 ? n37669 : n37670;
  assign n37672 = pi16 ? n32382 : n37671;
  assign n37673 = pi15 ? n37668 : n37672;
  assign n37674 = pi14 ? n37662 : n37673;
  assign n37675 = pi19 ? n13124 : n3086;
  assign n37676 = pi18 ? n37675 : n36570;
  assign n37677 = pi21 ? n204 : n29992;
  assign n37678 = pi20 ? n204 : n37677;
  assign n37679 = pi19 ? n37678 : n32;
  assign n37680 = pi18 ? n204 : n37679;
  assign n37681 = pi17 ? n37676 : n37680;
  assign n37682 = pi16 ? n37651 : n37681;
  assign n37683 = pi19 ? n16516 : n13535;
  assign n37684 = pi18 ? n37 : n37683;
  assign n37685 = pi20 ? n233 : n25965;
  assign n37686 = pi19 ? n37685 : n32;
  assign n37687 = pi18 ? n233 : n37686;
  assign n37688 = pi17 ? n37684 : n37687;
  assign n37689 = pi16 ? n33978 : n37688;
  assign n37690 = pi15 ? n37682 : n37689;
  assign n37691 = pi19 ? n36593 : n19358;
  assign n37692 = pi20 ? n233 : n25978;
  assign n37693 = pi19 ? n37692 : n32;
  assign n37694 = pi18 ? n37691 : n37693;
  assign n37695 = pi17 ? n36592 : n37694;
  assign n37696 = pi16 ? n33952 : n37695;
  assign n37697 = pi20 ? n639 : n8927;
  assign n37698 = pi19 ? n6340 : n37697;
  assign n37699 = pi21 ? n28746 : n19438;
  assign n37700 = pi20 ? n233 : n37699;
  assign n37701 = pi19 ? n37700 : n32;
  assign n37702 = pi18 ? n37698 : n37701;
  assign n37703 = pi17 ? n37 : n37702;
  assign n37704 = pi16 ? n33952 : n37703;
  assign n37705 = pi15 ? n37696 : n37704;
  assign n37706 = pi14 ? n37690 : n37705;
  assign n37707 = pi13 ? n37674 : n37706;
  assign n37708 = pi12 ? n37648 : n37707;
  assign n37709 = pi21 ? n233 : n10325;
  assign n37710 = pi20 ? n13527 : n37709;
  assign n37711 = pi19 ? n37710 : n32;
  assign n37712 = pi18 ? n37 : n37711;
  assign n37713 = pi17 ? n37 : n37712;
  assign n37714 = pi16 ? n32382 : n37713;
  assign n37715 = pi22 ? n316 : n233;
  assign n37716 = pi21 ? n37715 : n5178;
  assign n37717 = pi20 ? n6377 : n37716;
  assign n37718 = pi19 ? n37717 : n32;
  assign n37719 = pi18 ? n36630 : n37718;
  assign n37720 = pi17 ? n14165 : n37719;
  assign n37721 = pi16 ? n31317 : n37720;
  assign n37722 = pi15 ? n37714 : n37721;
  assign n37723 = pi18 ? n31315 : n9856;
  assign n37724 = pi17 ? n32 : n37723;
  assign n37725 = pi20 ? n6377 : n13743;
  assign n37726 = pi19 ? n37725 : n32;
  assign n37727 = pi18 ? n335 : n37726;
  assign n37728 = pi17 ? n335 : n37727;
  assign n37729 = pi16 ? n37724 : n37728;
  assign n37730 = pi19 ? n30097 : n335;
  assign n37731 = pi18 ? n31315 : n37730;
  assign n37732 = pi17 ? n32 : n37731;
  assign n37733 = pi20 ? n13527 : n13743;
  assign n37734 = pi19 ? n37733 : n32;
  assign n37735 = pi18 ? n335 : n37734;
  assign n37736 = pi17 ? n335 : n37735;
  assign n37737 = pi16 ? n37732 : n37736;
  assign n37738 = pi15 ? n37729 : n37737;
  assign n37739 = pi14 ? n37722 : n37738;
  assign n37740 = pi20 ? n30096 : n3299;
  assign n37741 = pi19 ? n37740 : n335;
  assign n37742 = pi18 ? n31315 : n37741;
  assign n37743 = pi17 ? n32 : n37742;
  assign n37744 = pi16 ? n37743 : n37728;
  assign n37745 = pi20 ? n30096 : n25064;
  assign n37746 = pi19 ? n37745 : n335;
  assign n37747 = pi18 ? n31315 : n37746;
  assign n37748 = pi17 ? n32 : n37747;
  assign n37749 = pi18 ? n335 : n25696;
  assign n37750 = pi17 ? n335 : n37749;
  assign n37751 = pi16 ? n37748 : n37750;
  assign n37752 = pi15 ? n37744 : n37751;
  assign n37753 = pi20 ? n363 : n24865;
  assign n37754 = pi19 ? n37 : n37753;
  assign n37755 = pi19 ? n363 : n27521;
  assign n37756 = pi18 ? n37754 : n37755;
  assign n37757 = pi20 ? n27520 : n20860;
  assign n37758 = pi21 ? n5015 : n560;
  assign n37759 = pi21 ? n5014 : n3392;
  assign n37760 = pi20 ? n37758 : n37759;
  assign n37761 = pi19 ? n37757 : n37760;
  assign n37762 = pi21 ? n685 : n6416;
  assign n37763 = pi20 ? n685 : n37762;
  assign n37764 = pi19 ? n37763 : n32;
  assign n37765 = pi18 ? n37761 : n37764;
  assign n37766 = pi17 ? n37756 : n37765;
  assign n37767 = pi16 ? n32382 : n37766;
  assign n37768 = pi22 ? n37173 : n20563;
  assign n37769 = pi21 ? n30866 : n37768;
  assign n37770 = pi20 ? n32 : n37769;
  assign n37771 = pi19 ? n32 : n37770;
  assign n37772 = pi18 ? n37771 : n31939;
  assign n37773 = pi17 ? n32 : n37772;
  assign n37774 = pi18 ? n36693 : n363;
  assign n37775 = pi20 ? n685 : n28002;
  assign n37776 = pi19 ? n37775 : n32;
  assign n37777 = pi18 ? n32832 : n37776;
  assign n37778 = pi17 ? n37774 : n37777;
  assign n37779 = pi16 ? n37773 : n37778;
  assign n37780 = pi15 ? n37767 : n37779;
  assign n37781 = pi14 ? n37752 : n37780;
  assign n37782 = pi13 ? n37739 : n37781;
  assign n37783 = pi23 ? n20563 : n36659;
  assign n37784 = pi22 ? n37783 : n20563;
  assign n37785 = pi21 ? n30866 : n37784;
  assign n37786 = pi20 ? n32 : n37785;
  assign n37787 = pi19 ? n32 : n37786;
  assign n37788 = pi19 ? n31280 : n29403;
  assign n37789 = pi18 ? n37787 : n37788;
  assign n37790 = pi17 ? n32 : n37789;
  assign n37791 = pi19 ? n363 : n27797;
  assign n37792 = pi20 ? n29741 : n14262;
  assign n37793 = pi19 ? n37792 : n32;
  assign n37794 = pi18 ? n37791 : n37793;
  assign n37795 = pi17 ? n363 : n37794;
  assign n37796 = pi16 ? n37790 : n37795;
  assign n37797 = pi21 ? n685 : n882;
  assign n37798 = pi20 ? n685 : n37797;
  assign n37799 = pi19 ? n37798 : n32;
  assign n37800 = pi18 ? n37 : n37799;
  assign n37801 = pi17 ? n37 : n37800;
  assign n37802 = pi16 ? n33952 : n37801;
  assign n37803 = pi15 ? n37796 : n37802;
  assign n37804 = pi23 ? n34196 : n30868;
  assign n37805 = pi22 ? n37804 : n30868;
  assign n37806 = pi21 ? n37805 : n30868;
  assign n37807 = pi20 ? n32 : n37806;
  assign n37808 = pi19 ? n32 : n37807;
  assign n37809 = pi23 ? n30868 : n99;
  assign n37810 = pi22 ? n30868 : n37809;
  assign n37811 = pi21 ? n37810 : n99;
  assign n37812 = pi20 ? n37811 : n99;
  assign n37813 = pi19 ? n37812 : n99;
  assign n37814 = pi18 ? n37808 : n37813;
  assign n37815 = pi17 ? n32 : n37814;
  assign n37816 = pi19 ? n25182 : n29738;
  assign n37817 = pi18 ? n99 : n37816;
  assign n37818 = pi20 ? n25199 : n25167;
  assign n37819 = pi19 ? n36741 : n37818;
  assign n37820 = pi21 ? n3445 : n928;
  assign n37821 = pi20 ? n685 : n37820;
  assign n37822 = pi19 ? n37821 : n32;
  assign n37823 = pi18 ? n37819 : n37822;
  assign n37824 = pi17 ? n37817 : n37823;
  assign n37825 = pi16 ? n37815 : n37824;
  assign n37826 = pi20 ? n30778 : n32813;
  assign n37827 = pi19 ? n99 : n37826;
  assign n37828 = pi20 ? n25167 : n33736;
  assign n37829 = pi19 ? n37828 : n36749;
  assign n37830 = pi18 ? n37827 : n37829;
  assign n37831 = pi19 ? n23151 : n36752;
  assign n37832 = pi20 ? n685 : n1010;
  assign n37833 = pi19 ? n37832 : n32;
  assign n37834 = pi18 ? n37831 : n37833;
  assign n37835 = pi17 ? n37830 : n37834;
  assign n37836 = pi16 ? n37815 : n37835;
  assign n37837 = pi15 ? n37825 : n37836;
  assign n37838 = pi14 ? n37803 : n37837;
  assign n37839 = pi21 ? n37252 : n33792;
  assign n37840 = pi20 ? n32 : n37839;
  assign n37841 = pi19 ? n32 : n37840;
  assign n37842 = pi21 ? n33792 : n36763;
  assign n37843 = pi20 ? n37842 : n139;
  assign n37844 = pi19 ? n37843 : n139;
  assign n37845 = pi18 ? n37841 : n37844;
  assign n37846 = pi17 ? n32 : n37845;
  assign n37847 = pi20 ? n18194 : n363;
  assign n37848 = pi19 ? n139 : n37847;
  assign n37849 = pi20 ? n26905 : n18194;
  assign n37850 = pi19 ? n37849 : n29741;
  assign n37851 = pi18 ? n37848 : n37850;
  assign n37852 = pi20 ? n24220 : n26890;
  assign n37853 = pi20 ? n24220 : n18194;
  assign n37854 = pi19 ? n37852 : n37853;
  assign n37855 = pi20 ? n685 : n12514;
  assign n37856 = pi19 ? n37855 : n32;
  assign n37857 = pi18 ? n37854 : n37856;
  assign n37858 = pi17 ? n37851 : n37857;
  assign n37859 = pi16 ? n37846 : n37858;
  assign n37860 = pi22 ? n37251 : n36781;
  assign n37861 = pi22 ? n36781 : n33792;
  assign n37862 = pi21 ? n37860 : n37861;
  assign n37863 = pi20 ? n32 : n37862;
  assign n37864 = pi19 ? n32 : n37863;
  assign n37865 = pi22 ? n36762 : n36785;
  assign n37866 = pi21 ? n36781 : n37865;
  assign n37867 = pi20 ? n37866 : n34221;
  assign n37868 = pi19 ? n37867 : n363;
  assign n37869 = pi18 ? n37864 : n37868;
  assign n37870 = pi17 ? n32 : n37869;
  assign n37871 = pi16 ? n37870 : n37270;
  assign n37872 = pi15 ? n37859 : n37871;
  assign n37873 = pi23 ? n37273 : n36659;
  assign n37874 = pi22 ? n37873 : n36781;
  assign n37875 = pi21 ? n37874 : n36659;
  assign n37876 = pi20 ? n32 : n37875;
  assign n37877 = pi19 ? n32 : n37876;
  assign n37878 = pi22 ? n36659 : n36781;
  assign n37879 = pi21 ? n37878 : n36802;
  assign n37880 = pi20 ? n37879 : n34837;
  assign n37881 = pi20 ? n34840 : n34834;
  assign n37882 = pi19 ? n37880 : n37881;
  assign n37883 = pi18 ? n37877 : n37882;
  assign n37884 = pi17 ? n32 : n37883;
  assign n37885 = pi20 ? n16279 : n9021;
  assign n37886 = pi19 ? n34832 : n37885;
  assign n37887 = pi21 ? n14277 : n6461;
  assign n37888 = pi20 ? n37887 : n685;
  assign n37889 = pi20 ? n36851 : n685;
  assign n37890 = pi19 ? n37888 : n37889;
  assign n37891 = pi18 ? n37886 : n37890;
  assign n37892 = pi21 ? n685 : n14277;
  assign n37893 = pi20 ? n37892 : n685;
  assign n37894 = pi20 ? n685 : n37887;
  assign n37895 = pi19 ? n37893 : n37894;
  assign n37896 = pi18 ? n37895 : n32243;
  assign n37897 = pi17 ? n37891 : n37896;
  assign n37898 = pi16 ? n37884 : n37897;
  assign n37899 = pi22 ? n36798 : n36659;
  assign n37900 = pi21 ? n37874 : n37899;
  assign n37901 = pi20 ? n32 : n37900;
  assign n37902 = pi19 ? n32 : n37901;
  assign n37903 = pi21 ? n36659 : n36710;
  assign n37904 = pi20 ? n37903 : n36838;
  assign n37905 = pi19 ? n37904 : n157;
  assign n37906 = pi18 ? n37902 : n37905;
  assign n37907 = pi17 ? n32 : n37906;
  assign n37908 = pi21 ? n685 : n27554;
  assign n37909 = pi20 ? n157 : n37908;
  assign n37910 = pi20 ? n36851 : n15272;
  assign n37911 = pi19 ? n37909 : n37910;
  assign n37912 = pi18 ? n157 : n37911;
  assign n37913 = pi19 ? n37892 : n36852;
  assign n37914 = pi20 ? n27551 : n8295;
  assign n37915 = pi19 ? n37914 : n32;
  assign n37916 = pi18 ? n37913 : n37915;
  assign n37917 = pi17 ? n37912 : n37916;
  assign n37918 = pi16 ? n37907 : n37917;
  assign n37919 = pi15 ? n37898 : n37918;
  assign n37920 = pi14 ? n37872 : n37919;
  assign n37921 = pi13 ? n37838 : n37920;
  assign n37922 = pi12 ? n37782 : n37921;
  assign n37923 = pi11 ? n37708 : n37922;
  assign n37924 = pi10 ? n37579 : n37923;
  assign n37925 = pi09 ? n37352 : n37924;
  assign n37926 = pi21 ? n32 : n37332;
  assign n37927 = pi20 ? n32 : n37926;
  assign n37928 = pi19 ? n32 : n37927;
  assign n37929 = pi18 ? n37928 : n20563;
  assign n37930 = pi17 ? n32 : n37929;
  assign n37931 = pi16 ? n37930 : n37317;
  assign n37932 = pi15 ? n32 : n37931;
  assign n37933 = pi21 ? n32 : n28156;
  assign n37934 = pi20 ? n32 : n37933;
  assign n37935 = pi19 ? n32 : n37934;
  assign n37936 = pi18 ? n37935 : n20563;
  assign n37937 = pi17 ? n32 : n37936;
  assign n37938 = pi20 ? n32286 : n226;
  assign n37939 = pi19 ? n20563 : n37938;
  assign n37940 = pi18 ? n37939 : n99;
  assign n37941 = pi17 ? n37940 : n37329;
  assign n37942 = pi16 ? n37937 : n37941;
  assign n37943 = pi21 ? n3493 : n8015;
  assign n37944 = pi20 ? n37943 : n32;
  assign n37945 = pi19 ? n99 : n37944;
  assign n37946 = pi18 ? n99 : n37945;
  assign n37947 = pi17 ? n37340 : n37946;
  assign n37948 = pi16 ? n36871 : n37947;
  assign n37949 = pi15 ? n37942 : n37948;
  assign n37950 = pi14 ? n37932 : n37949;
  assign n37951 = pi13 ? n32 : n37950;
  assign n37952 = pi12 ? n32 : n37951;
  assign n37953 = pi11 ? n32 : n37952;
  assign n37954 = pi10 ? n32 : n37953;
  assign n37955 = pi21 ? n32 : n30155;
  assign n37956 = pi20 ? n32 : n37955;
  assign n37957 = pi19 ? n32 : n37956;
  assign n37958 = pi18 ? n37957 : n20563;
  assign n37959 = pi17 ? n32 : n37958;
  assign n37960 = pi22 ? n99 : n11963;
  assign n37961 = pi21 ? n37960 : n8557;
  assign n37962 = pi20 ? n37961 : n32;
  assign n37963 = pi19 ? n99 : n37962;
  assign n37964 = pi18 ? n99 : n37963;
  assign n37965 = pi17 ? n37354 : n37964;
  assign n37966 = pi16 ? n37959 : n37965;
  assign n37967 = pi22 ? n99 : n7024;
  assign n37968 = pi21 ? n37967 : n8044;
  assign n37969 = pi20 ? n37968 : n32;
  assign n37970 = pi19 ? n99 : n37969;
  assign n37971 = pi18 ? n99 : n37970;
  assign n37972 = pi17 ? n37363 : n37971;
  assign n37973 = pi16 ? n35765 : n37972;
  assign n37974 = pi15 ? n37966 : n37973;
  assign n37975 = pi21 ? n7025 : n32;
  assign n37976 = pi20 ? n37975 : n32;
  assign n37977 = pi19 ? n37 : n37976;
  assign n37978 = pi18 ? n37 : n37977;
  assign n37979 = pi17 ? n37372 : n37978;
  assign n37980 = pi16 ? n35765 : n37979;
  assign n37981 = pi19 ? n36886 : n37;
  assign n37982 = pi18 ? n37981 : n37;
  assign n37983 = pi22 ? n37 : n33884;
  assign n37984 = pi21 ? n37983 : n32;
  assign n37985 = pi20 ? n37984 : n32;
  assign n37986 = pi19 ? n37 : n37985;
  assign n37987 = pi18 ? n37 : n37986;
  assign n37988 = pi17 ? n37982 : n37987;
  assign n37989 = pi16 ? n36216 : n37988;
  assign n37990 = pi15 ? n37980 : n37989;
  assign n37991 = pi14 ? n37974 : n37990;
  assign n37992 = pi20 ? n31220 : n31903;
  assign n37993 = pi19 ? n37992 : n37;
  assign n37994 = pi18 ? n37993 : n37;
  assign n37995 = pi19 ? n9814 : n7309;
  assign n37996 = pi18 ? n37 : n37995;
  assign n37997 = pi17 ? n37994 : n37996;
  assign n37998 = pi16 ? n36216 : n37997;
  assign n37999 = pi19 ? n31926 : n37395;
  assign n38000 = pi18 ? n37999 : n139;
  assign n38001 = pi19 ? n139 : n9799;
  assign n38002 = pi18 ? n139 : n38001;
  assign n38003 = pi17 ? n38000 : n38002;
  assign n38004 = pi16 ? n36216 : n38003;
  assign n38005 = pi15 ? n37998 : n38004;
  assign n38006 = pi17 ? n37407 : n38002;
  assign n38007 = pi16 ? n36216 : n38006;
  assign n38008 = pi18 ? n32924 : n37410;
  assign n38009 = pi17 ? n38008 : n38002;
  assign n38010 = pi16 ? n36216 : n38009;
  assign n38011 = pi15 ? n38007 : n38010;
  assign n38012 = pi14 ? n38005 : n38011;
  assign n38013 = pi13 ? n37991 : n38012;
  assign n38014 = pi20 ? n22214 : n32;
  assign n38015 = pi19 ? n9769 : n38014;
  assign n38016 = pi18 ? n139 : n38015;
  assign n38017 = pi17 ? n35254 : n38016;
  assign n38018 = pi16 ? n36216 : n38017;
  assign n38019 = pi17 ? n37426 : n38016;
  assign n38020 = pi16 ? n36216 : n38019;
  assign n38021 = pi15 ? n38018 : n38020;
  assign n38022 = pi21 ? n17755 : n2700;
  assign n38023 = pi20 ? n38022 : n32;
  assign n38024 = pi19 ? n28367 : n38023;
  assign n38025 = pi18 ? n22047 : n38024;
  assign n38026 = pi17 ? n37 : n38025;
  assign n38027 = pi16 ? n36235 : n38026;
  assign n38028 = pi21 ? n31885 : n29133;
  assign n38029 = pi20 ? n20563 : n38028;
  assign n38030 = pi19 ? n20563 : n38029;
  assign n38031 = pi18 ? n31315 : n38030;
  assign n38032 = pi17 ? n32 : n38031;
  assign n38033 = pi21 ? n17741 : n2700;
  assign n38034 = pi20 ? n38033 : n32;
  assign n38035 = pi19 ? n17204 : n38034;
  assign n38036 = pi18 ? n37 : n38035;
  assign n38037 = pi17 ? n37 : n38036;
  assign n38038 = pi16 ? n38032 : n38037;
  assign n38039 = pi15 ? n38027 : n38038;
  assign n38040 = pi14 ? n38021 : n38039;
  assign n38041 = pi22 ? n99 : n10400;
  assign n38042 = pi21 ? n38041 : n1009;
  assign n38043 = pi20 ? n38042 : n32;
  assign n38044 = pi19 ? n17204 : n38043;
  assign n38045 = pi18 ? n37448 : n38044;
  assign n38046 = pi17 ? n37 : n38045;
  assign n38047 = pi16 ? n36956 : n38046;
  assign n38048 = pi16 ? n34306 : n37455;
  assign n38049 = pi15 ? n38047 : n38048;
  assign n38050 = pi16 ? n35283 : n37466;
  assign n38051 = pi15 ? n37463 : n38050;
  assign n38052 = pi14 ? n38049 : n38051;
  assign n38053 = pi13 ? n38040 : n38052;
  assign n38054 = pi12 ? n38013 : n38053;
  assign n38055 = pi16 ? n34328 : n37495;
  assign n38056 = pi15 ? n38055 : n37501;
  assign n38057 = pi14 ? n37487 : n38056;
  assign n38058 = pi16 ? n34352 : n37520;
  assign n38059 = pi15 ? n37514 : n38058;
  assign n38060 = pi16 ? n34335 : n37520;
  assign n38061 = pi21 ? n30820 : n32;
  assign n38062 = pi20 ? n38061 : n32;
  assign n38063 = pi19 ? n27535 : n38062;
  assign n38064 = pi18 ? n37 : n38063;
  assign n38065 = pi17 ? n37 : n38064;
  assign n38066 = pi16 ? n34335 : n38065;
  assign n38067 = pi15 ? n38060 : n38066;
  assign n38068 = pi14 ? n38059 : n38067;
  assign n38069 = pi13 ? n38057 : n38068;
  assign n38070 = pi18 ? n31938 : n34358;
  assign n38071 = pi17 ? n32 : n38070;
  assign n38072 = pi19 ? n37 : n11696;
  assign n38073 = pi18 ? n37 : n38072;
  assign n38074 = pi17 ? n37 : n38073;
  assign n38075 = pi16 ? n38071 : n38074;
  assign n38076 = pi19 ? n37 : n11244;
  assign n38077 = pi18 ? n37 : n38076;
  assign n38078 = pi17 ? n37 : n38077;
  assign n38079 = pi16 ? n33908 : n38078;
  assign n38080 = pi16 ? n33908 : n37543;
  assign n38081 = pi15 ? n38079 : n38080;
  assign n38082 = pi14 ? n38075 : n38081;
  assign n38083 = pi21 ? n26377 : n32;
  assign n38084 = pi20 ? n38083 : n32;
  assign n38085 = pi19 ? n37540 : n38084;
  assign n38086 = pi18 ? n37 : n38085;
  assign n38087 = pi17 ? n37 : n38086;
  assign n38088 = pi16 ? n32901 : n38087;
  assign n38089 = pi19 ? n37 : n4009;
  assign n38090 = pi18 ? n37 : n38089;
  assign n38091 = pi17 ? n37 : n38090;
  assign n38092 = pi16 ? n32901 : n38091;
  assign n38093 = pi15 ? n38088 : n38092;
  assign n38094 = pi19 ? n33822 : n21611;
  assign n38095 = pi18 ? n31315 : n38094;
  assign n38096 = pi17 ? n32 : n38095;
  assign n38097 = pi20 ? n24937 : n32;
  assign n38098 = pi19 ? n157 : n38097;
  assign n38099 = pi18 ? n37563 : n38098;
  assign n38100 = pi17 ? n99 : n38099;
  assign n38101 = pi16 ? n38096 : n38100;
  assign n38102 = pi19 ? n33822 : n18853;
  assign n38103 = pi18 ? n31315 : n38102;
  assign n38104 = pi17 ? n32 : n38103;
  assign n38105 = pi19 ? n6532 : n4009;
  assign n38106 = pi18 ? n19145 : n38105;
  assign n38107 = pi17 ? n37570 : n38106;
  assign n38108 = pi16 ? n38104 : n38107;
  assign n38109 = pi15 ? n38101 : n38108;
  assign n38110 = pi14 ? n38093 : n38109;
  assign n38111 = pi13 ? n38082 : n38110;
  assign n38112 = pi12 ? n38069 : n38111;
  assign n38113 = pi11 ? n38054 : n38112;
  assign n38114 = pi19 ? n13069 : n13467;
  assign n38115 = pi18 ? n37583 : n38114;
  assign n38116 = pi17 ? n37570 : n38115;
  assign n38117 = pi16 ? n37582 : n38116;
  assign n38118 = pi19 ? n31914 : n18853;
  assign n38119 = pi18 ? n31315 : n38118;
  assign n38120 = pi17 ? n32 : n38119;
  assign n38121 = pi16 ? n38120 : n37595;
  assign n38122 = pi15 ? n38117 : n38121;
  assign n38123 = pi19 ? n31914 : n99;
  assign n38124 = pi18 ? n31315 : n38123;
  assign n38125 = pi17 ? n32 : n38124;
  assign n38126 = pi16 ? n38125 : n37608;
  assign n38127 = pi18 ? n31315 : n31927;
  assign n38128 = pi17 ? n32 : n38127;
  assign n38129 = pi16 ? n38128 : n37614;
  assign n38130 = pi15 ? n38126 : n38129;
  assign n38131 = pi14 ? n38122 : n38130;
  assign n38132 = pi20 ? n31925 : n14844;
  assign n38133 = pi19 ? n38132 : n99;
  assign n38134 = pi18 ? n31315 : n38133;
  assign n38135 = pi17 ? n32 : n38134;
  assign n38136 = pi16 ? n38135 : n37614;
  assign n38137 = pi16 ? n32371 : n37632;
  assign n38138 = pi15 ? n38136 : n38137;
  assign n38139 = pi16 ? n32371 : n36514;
  assign n38140 = pi19 ? n32348 : n8765;
  assign n38141 = pi18 ? n31315 : n38140;
  assign n38142 = pi17 ? n32 : n38141;
  assign n38143 = pi19 ? n30527 : n2680;
  assign n38144 = pi18 ? n139 : n38143;
  assign n38145 = pi17 ? n139 : n38144;
  assign n38146 = pi16 ? n38142 : n38145;
  assign n38147 = pi15 ? n38139 : n38146;
  assign n38148 = pi14 ? n38138 : n38147;
  assign n38149 = pi13 ? n38131 : n38148;
  assign n38150 = pi18 ? n31315 : n34949;
  assign n38151 = pi17 ? n32 : n38150;
  assign n38152 = pi20 ? n2512 : n139;
  assign n38153 = pi19 ? n38152 : n139;
  assign n38154 = pi19 ? n26742 : n2702;
  assign n38155 = pi18 ? n38153 : n38154;
  assign n38156 = pi17 ? n36530 : n38155;
  assign n38157 = pi16 ? n38151 : n38156;
  assign n38158 = pi19 ? n34641 : n2702;
  assign n38159 = pi18 ? n37657 : n38158;
  assign n38160 = pi17 ? n37656 : n38159;
  assign n38161 = pi16 ? n32915 : n38160;
  assign n38162 = pi15 ? n38157 : n38161;
  assign n38163 = pi19 ? n11810 : n1823;
  assign n38164 = pi18 ? n37664 : n38163;
  assign n38165 = pi17 ? n36549 : n38164;
  assign n38166 = pi16 ? n32371 : n38165;
  assign n38167 = pi18 ? n31315 : n36363;
  assign n38168 = pi17 ? n32 : n38167;
  assign n38169 = pi16 ? n38168 : n37671;
  assign n38170 = pi15 ? n38166 : n38169;
  assign n38171 = pi14 ? n38162 : n38170;
  assign n38172 = pi16 ? n38168 : n37681;
  assign n38173 = pi16 ? n37651 : n37688;
  assign n38174 = pi15 ? n38172 : n38173;
  assign n38175 = pi16 ? n35320 : n37695;
  assign n38176 = pi21 ? n28746 : n10981;
  assign n38177 = pi20 ? n233 : n38176;
  assign n38178 = pi19 ? n38177 : n32;
  assign n38179 = pi18 ? n37698 : n38178;
  assign n38180 = pi17 ? n37 : n38179;
  assign n38181 = pi16 ? n35320 : n38180;
  assign n38182 = pi15 ? n38175 : n38181;
  assign n38183 = pi14 ? n38174 : n38182;
  assign n38184 = pi13 ? n38171 : n38183;
  assign n38185 = pi12 ? n38149 : n38184;
  assign n38186 = pi18 ? n37 : n36626;
  assign n38187 = pi17 ? n37 : n38186;
  assign n38188 = pi16 ? n32382 : n38187;
  assign n38189 = pi21 ? n37715 : n3523;
  assign n38190 = pi20 ? n6377 : n38189;
  assign n38191 = pi19 ? n38190 : n32;
  assign n38192 = pi18 ? n36630 : n38191;
  assign n38193 = pi17 ? n14165 : n38192;
  assign n38194 = pi16 ? n32936 : n38193;
  assign n38195 = pi15 ? n38188 : n38194;
  assign n38196 = pi19 ? n33965 : n335;
  assign n38197 = pi18 ? n31315 : n38196;
  assign n38198 = pi17 ? n32 : n38197;
  assign n38199 = pi20 ? n6377 : n26514;
  assign n38200 = pi19 ? n38199 : n32;
  assign n38201 = pi18 ? n335 : n38200;
  assign n38202 = pi17 ? n335 : n38201;
  assign n38203 = pi16 ? n38198 : n38202;
  assign n38204 = pi19 ? n33949 : n335;
  assign n38205 = pi18 ? n31315 : n38204;
  assign n38206 = pi17 ? n32 : n38205;
  assign n38207 = pi20 ? n13527 : n26514;
  assign n38208 = pi19 ? n38207 : n32;
  assign n38209 = pi18 ? n335 : n38208;
  assign n38210 = pi17 ? n335 : n38209;
  assign n38211 = pi16 ? n38206 : n38210;
  assign n38212 = pi15 ? n38203 : n38211;
  assign n38213 = pi14 ? n38195 : n38212;
  assign n38214 = pi21 ? n233 : n4101;
  assign n38215 = pi20 ? n6377 : n38214;
  assign n38216 = pi19 ? n38215 : n32;
  assign n38217 = pi18 ? n335 : n38216;
  assign n38218 = pi17 ? n335 : n38217;
  assign n38219 = pi16 ? n38206 : n38218;
  assign n38220 = pi22 ? n36660 : n37;
  assign n38221 = pi21 ? n31924 : n38220;
  assign n38222 = pi20 ? n38221 : n604;
  assign n38223 = pi19 ? n38222 : n335;
  assign n38224 = pi18 ? n31315 : n38223;
  assign n38225 = pi17 ? n32 : n38224;
  assign n38226 = pi16 ? n38225 : n37750;
  assign n38227 = pi15 ? n38219 : n38226;
  assign n38228 = pi20 ? n32313 : n13147;
  assign n38229 = pi19 ? n38228 : n37;
  assign n38230 = pi18 ? n31315 : n38229;
  assign n38231 = pi17 ? n32 : n38230;
  assign n38232 = pi16 ? n38231 : n37766;
  assign n38233 = pi18 ? n37771 : n38229;
  assign n38234 = pi17 ? n32 : n38233;
  assign n38235 = pi16 ? n38234 : n37778;
  assign n38236 = pi15 ? n38232 : n38235;
  assign n38237 = pi14 ? n38227 : n38236;
  assign n38238 = pi13 ? n38213 : n38237;
  assign n38239 = pi20 ? n32313 : n24105;
  assign n38240 = pi19 ? n38239 : n29403;
  assign n38241 = pi18 ? n37787 : n38240;
  assign n38242 = pi17 ? n32 : n38241;
  assign n38243 = pi16 ? n38242 : n37795;
  assign n38244 = pi16 ? n32382 : n36727;
  assign n38245 = pi15 ? n38243 : n38244;
  assign n38246 = pi22 ? n36730 : n30868;
  assign n38247 = pi21 ? n38246 : n30868;
  assign n38248 = pi20 ? n32 : n38247;
  assign n38249 = pi19 ? n32 : n38248;
  assign n38250 = pi21 ? n30868 : n99;
  assign n38251 = pi20 ? n38250 : n99;
  assign n38252 = pi19 ? n38251 : n99;
  assign n38253 = pi18 ? n38249 : n38252;
  assign n38254 = pi17 ? n32 : n38253;
  assign n38255 = pi18 ? n37819 : n36745;
  assign n38256 = pi17 ? n37817 : n38255;
  assign n38257 = pi16 ? n38254 : n38256;
  assign n38258 = pi18 ? n37831 : n36754;
  assign n38259 = pi17 ? n37830 : n38258;
  assign n38260 = pi16 ? n38254 : n38259;
  assign n38261 = pi15 ? n38257 : n38260;
  assign n38262 = pi14 ? n38245 : n38261;
  assign n38263 = pi21 ? n33792 : n36762;
  assign n38264 = pi20 ? n38263 : n139;
  assign n38265 = pi19 ? n38264 : n139;
  assign n38266 = pi18 ? n37841 : n38265;
  assign n38267 = pi17 ? n32 : n38266;
  assign n38268 = pi18 ? n37854 : n33742;
  assign n38269 = pi17 ? n37851 : n38268;
  assign n38270 = pi16 ? n38267 : n38269;
  assign n38271 = pi23 ? n36781 : n33792;
  assign n38272 = pi22 ? n33792 : n38271;
  assign n38273 = pi21 ? n36781 : n38272;
  assign n38274 = pi20 ? n38273 : n34221;
  assign n38275 = pi19 ? n38274 : n363;
  assign n38276 = pi18 ? n37864 : n38275;
  assign n38277 = pi17 ? n32 : n38276;
  assign n38278 = pi20 ? n25199 : n9963;
  assign n38279 = pi19 ? n38278 : n32;
  assign n38280 = pi18 ? n363 : n38279;
  assign n38281 = pi17 ? n363 : n38280;
  assign n38282 = pi16 ? n38277 : n38281;
  assign n38283 = pi15 ? n38270 : n38282;
  assign n38284 = pi23 ? n36659 : n36781;
  assign n38285 = pi22 ? n38284 : n36781;
  assign n38286 = pi21 ? n37878 : n38285;
  assign n38287 = pi20 ? n38286 : n34837;
  assign n38288 = pi19 ? n38287 : n37881;
  assign n38289 = pi18 ? n37877 : n38288;
  assign n38290 = pi17 ? n32 : n38289;
  assign n38291 = pi18 ? n37895 : n32778;
  assign n38292 = pi17 ? n37891 : n38291;
  assign n38293 = pi16 ? n38290 : n38292;
  assign n38294 = pi20 ? n36659 : n36838;
  assign n38295 = pi19 ? n38294 : n157;
  assign n38296 = pi18 ? n37902 : n38295;
  assign n38297 = pi17 ? n32 : n38296;
  assign n38298 = pi20 ? n27551 : n22920;
  assign n38299 = pi19 ? n38298 : n32;
  assign n38300 = pi18 ? n37913 : n38299;
  assign n38301 = pi17 ? n37912 : n38300;
  assign n38302 = pi16 ? n38297 : n38301;
  assign n38303 = pi15 ? n38293 : n38302;
  assign n38304 = pi14 ? n38283 : n38303;
  assign n38305 = pi13 ? n38262 : n38304;
  assign n38306 = pi12 ? n38238 : n38305;
  assign n38307 = pi11 ? n38185 : n38306;
  assign n38308 = pi10 ? n38113 : n38307;
  assign n38309 = pi09 ? n37954 : n38308;
  assign n38310 = pi08 ? n37925 : n38309;
  assign n38311 = pi07 ? n37307 : n38310;
  assign n38312 = pi06 ? n36161 : n38311;
  assign n38313 = pi05 ? n34245 : n38312;
  assign n38314 = pi04 ? n30095 : n38313;
  assign n38315 = pi20 ? n31313 : n20563;
  assign n38316 = pi19 ? n38315 : n20563;
  assign n38317 = pi18 ? n32 : n38316;
  assign n38318 = pi17 ? n32 : n38317;
  assign n38319 = pi20 ? n37 : n7346;
  assign n38320 = pi19 ? n37 : n38319;
  assign n38321 = pi18 ? n34869 : n38320;
  assign n38322 = pi19 ? n22685 : n99;
  assign n38323 = pi21 ? n99 : n2989;
  assign n38324 = pi20 ? n38323 : n32;
  assign n38325 = pi19 ? n8074 : n38324;
  assign n38326 = pi18 ? n38322 : n38325;
  assign n38327 = pi17 ? n38321 : n38326;
  assign n38328 = pi16 ? n38318 : n38327;
  assign n38329 = pi15 ? n32 : n38328;
  assign n38330 = pi18 ? n32 : n20563;
  assign n38331 = pi17 ? n32 : n38330;
  assign n38332 = pi21 ? n36489 : n37;
  assign n38333 = pi20 ? n20563 : n38332;
  assign n38334 = pi19 ? n20563 : n38333;
  assign n38335 = pi18 ? n38334 : n34262;
  assign n38336 = pi19 ? n99 : n38324;
  assign n38337 = pi18 ? n99 : n38336;
  assign n38338 = pi17 ? n38335 : n38337;
  assign n38339 = pi16 ? n38331 : n38338;
  assign n38340 = pi21 ? n29133 : n31877;
  assign n38341 = pi20 ? n38340 : n37;
  assign n38342 = pi19 ? n34246 : n38341;
  assign n38343 = pi21 ? n2175 : n1143;
  assign n38344 = pi20 ? n38343 : n226;
  assign n38345 = pi19 ? n38344 : n99;
  assign n38346 = pi18 ? n38342 : n38345;
  assign n38347 = pi19 ? n99 : n8537;
  assign n38348 = pi18 ? n99 : n38347;
  assign n38349 = pi17 ? n38346 : n38348;
  assign n38350 = pi16 ? n36871 : n38349;
  assign n38351 = pi15 ? n38339 : n38350;
  assign n38352 = pi14 ? n38329 : n38351;
  assign n38353 = pi13 ? n32 : n38352;
  assign n38354 = pi12 ? n32 : n38353;
  assign n38355 = pi11 ? n32 : n38354;
  assign n38356 = pi10 ? n32 : n38355;
  assign n38357 = pi20 ? n7346 : n22644;
  assign n38358 = pi20 ? n3814 : n3884;
  assign n38359 = pi19 ? n38357 : n38358;
  assign n38360 = pi18 ? n34295 : n38359;
  assign n38361 = pi20 ? n221 : n2961;
  assign n38362 = pi19 ? n38361 : n6046;
  assign n38363 = pi21 ? n1143 : n3066;
  assign n38364 = pi20 ? n38363 : n32;
  assign n38365 = pi19 ? n17972 : n38364;
  assign n38366 = pi18 ? n38362 : n38365;
  assign n38367 = pi17 ? n38360 : n38366;
  assign n38368 = pi16 ? n37959 : n38367;
  assign n38369 = pi18 ? n32872 : n37;
  assign n38370 = pi19 ? n3105 : n9240;
  assign n38371 = pi18 ? n37 : n38370;
  assign n38372 = pi17 ? n38369 : n38371;
  assign n38373 = pi16 ? n37337 : n38372;
  assign n38374 = pi15 ? n38368 : n38373;
  assign n38375 = pi22 ? n32 : n30154;
  assign n38376 = pi21 ? n38375 : n20563;
  assign n38377 = pi20 ? n32 : n38376;
  assign n38378 = pi19 ? n32 : n38377;
  assign n38379 = pi18 ? n38378 : n20563;
  assign n38380 = pi17 ? n32 : n38379;
  assign n38381 = pi21 ? n20563 : n36516;
  assign n38382 = pi20 ? n38381 : n37;
  assign n38383 = pi19 ? n20563 : n38382;
  assign n38384 = pi18 ? n38383 : n37;
  assign n38385 = pi19 ? n37 : n8572;
  assign n38386 = pi18 ? n37 : n38385;
  assign n38387 = pi17 ? n38384 : n38386;
  assign n38388 = pi16 ? n38380 : n38387;
  assign n38389 = pi18 ? n33299 : n37;
  assign n38390 = pi17 ? n38389 : n38386;
  assign n38391 = pi16 ? n35765 : n38390;
  assign n38392 = pi15 ? n38388 : n38391;
  assign n38393 = pi14 ? n38374 : n38392;
  assign n38394 = pi19 ? n31221 : n30097;
  assign n38395 = pi18 ? n38394 : n37;
  assign n38396 = pi20 ? n13143 : n3922;
  assign n38397 = pi20 ? n947 : n1003;
  assign n38398 = pi19 ? n38396 : n38397;
  assign n38399 = pi19 ? n9795 : n9799;
  assign n38400 = pi18 ? n38398 : n38399;
  assign n38401 = pi17 ? n38395 : n38400;
  assign n38402 = pi16 ? n36216 : n38401;
  assign n38403 = pi20 ? n1705 : n1694;
  assign n38404 = pi20 ? n1697 : n12014;
  assign n38405 = pi19 ? n38403 : n38404;
  assign n38406 = pi18 ? n33299 : n38405;
  assign n38407 = pi20 ? n3572 : n11579;
  assign n38408 = pi20 ? n14039 : n1757;
  assign n38409 = pi19 ? n38407 : n38408;
  assign n38410 = pi20 ? n8707 : n139;
  assign n38411 = pi19 ? n38410 : n9799;
  assign n38412 = pi18 ? n38409 : n38411;
  assign n38413 = pi17 ? n38406 : n38412;
  assign n38414 = pi16 ? n36216 : n38413;
  assign n38415 = pi15 ? n38402 : n38414;
  assign n38416 = pi20 ? n37 : n14038;
  assign n38417 = pi19 ? n37 : n38416;
  assign n38418 = pi18 ? n32295 : n38417;
  assign n38419 = pi20 ? n30255 : n139;
  assign n38420 = pi20 ? n139 : n14068;
  assign n38421 = pi19 ? n38419 : n38420;
  assign n38422 = pi18 ? n38421 : n38411;
  assign n38423 = pi17 ? n38418 : n38422;
  assign n38424 = pi16 ? n36216 : n38423;
  assign n38425 = pi18 ? n32295 : n37;
  assign n38426 = pi19 ? n9814 : n9799;
  assign n38427 = pi18 ? n34307 : n38426;
  assign n38428 = pi17 ? n38425 : n38427;
  assign n38429 = pi16 ? n36216 : n38428;
  assign n38430 = pi15 ? n38424 : n38429;
  assign n38431 = pi14 ? n38415 : n38430;
  assign n38432 = pi13 ? n38393 : n38431;
  assign n38433 = pi18 ? n34358 : n16056;
  assign n38434 = pi20 ? n942 : n3083;
  assign n38435 = pi19 ? n38434 : n13156;
  assign n38436 = pi20 ? n376 : n139;
  assign n38437 = pi21 ? n335 : n2678;
  assign n38438 = pi20 ? n38437 : n32;
  assign n38439 = pi19 ? n38436 : n38438;
  assign n38440 = pi18 ? n38435 : n38439;
  assign n38441 = pi17 ? n38433 : n38440;
  assign n38442 = pi16 ? n36216 : n38441;
  assign n38443 = pi18 ? n35300 : n37;
  assign n38444 = pi19 ? n7676 : n38438;
  assign n38445 = pi18 ? n37 : n38444;
  assign n38446 = pi17 ? n38443 : n38445;
  assign n38447 = pi16 ? n36216 : n38446;
  assign n38448 = pi15 ? n38442 : n38447;
  assign n38449 = pi18 ? n32377 : n37;
  assign n38450 = pi20 ? n22230 : n32;
  assign n38451 = pi19 ? n3332 : n38450;
  assign n38452 = pi18 ? n37 : n38451;
  assign n38453 = pi17 ? n38449 : n38452;
  assign n38454 = pi16 ? n36216 : n38453;
  assign n38455 = pi18 ? n37649 : n37;
  assign n38456 = pi21 ? n335 : n1009;
  assign n38457 = pi20 ? n38456 : n32;
  assign n38458 = pi19 ? n37 : n38457;
  assign n38459 = pi18 ? n37 : n38458;
  assign n38460 = pi17 ? n38455 : n38459;
  assign n38461 = pi16 ? n36216 : n38460;
  assign n38462 = pi15 ? n38454 : n38461;
  assign n38463 = pi14 ? n38448 : n38462;
  assign n38464 = pi20 ? n25766 : n32;
  assign n38465 = pi19 ? n37 : n38464;
  assign n38466 = pi18 ? n37 : n38465;
  assign n38467 = pi17 ? n36210 : n38466;
  assign n38468 = pi16 ? n36216 : n38467;
  assign n38469 = pi21 ? n37 : n4920;
  assign n38470 = pi20 ? n37 : n38469;
  assign n38471 = pi19 ? n38470 : n19362;
  assign n38472 = pi18 ? n37 : n38471;
  assign n38473 = pi17 ? n37 : n38472;
  assign n38474 = pi16 ? n36235 : n38473;
  assign n38475 = pi15 ? n38468 : n38474;
  assign n38476 = pi16 ? n36956 : n38473;
  assign n38477 = pi21 ? n29133 : n20563;
  assign n38478 = pi20 ? n20563 : n38477;
  assign n38479 = pi19 ? n20563 : n38478;
  assign n38480 = pi18 ? n31315 : n38479;
  assign n38481 = pi17 ? n32 : n38480;
  assign n38482 = pi19 ? n7685 : n19362;
  assign n38483 = pi18 ? n37 : n38482;
  assign n38484 = pi17 ? n37 : n38483;
  assign n38485 = pi16 ? n38481 : n38484;
  assign n38486 = pi15 ? n38476 : n38485;
  assign n38487 = pi14 ? n38475 : n38486;
  assign n38488 = pi13 ? n38463 : n38487;
  assign n38489 = pi12 ? n38432 : n38488;
  assign n38490 = pi19 ? n37 : n3299;
  assign n38491 = pi18 ? n37 : n38490;
  assign n38492 = pi20 ? n638 : n7646;
  assign n38493 = pi19 ? n37 : n38492;
  assign n38494 = pi20 ? n37 : n604;
  assign n38495 = pi21 ? n6376 : n2700;
  assign n38496 = pi20 ? n38495 : n32;
  assign n38497 = pi19 ? n38494 : n38496;
  assign n38498 = pi18 ? n38493 : n38497;
  assign n38499 = pi17 ? n38491 : n38498;
  assign n38500 = pi16 ? n36235 : n38499;
  assign n38501 = pi19 ? n37 : n34421;
  assign n38502 = pi20 ? n37 : n27730;
  assign n38503 = pi19 ? n38502 : n11186;
  assign n38504 = pi18 ? n38501 : n38503;
  assign n38505 = pi17 ? n37 : n38504;
  assign n38506 = pi16 ? n37443 : n38505;
  assign n38507 = pi15 ? n38500 : n38506;
  assign n38508 = pi19 ? n22878 : n11216;
  assign n38509 = pi18 ? n37 : n38508;
  assign n38510 = pi17 ? n37 : n38509;
  assign n38511 = pi16 ? n36235 : n38510;
  assign n38512 = pi19 ? n7731 : n11216;
  assign n38513 = pi18 ? n37 : n38512;
  assign n38514 = pi17 ? n37 : n38513;
  assign n38515 = pi16 ? n36227 : n38514;
  assign n38516 = pi15 ? n38511 : n38515;
  assign n38517 = pi14 ? n38507 : n38516;
  assign n38518 = pi19 ? n24866 : n11216;
  assign n38519 = pi18 ? n37 : n38518;
  assign n38520 = pi17 ? n37 : n38519;
  assign n38521 = pi16 ? n36254 : n38520;
  assign n38522 = pi20 ? n31266 : n30096;
  assign n38523 = pi19 ? n20563 : n38522;
  assign n38524 = pi18 ? n31315 : n38523;
  assign n38525 = pi17 ? n32 : n38524;
  assign n38526 = pi20 ? n20729 : n32;
  assign n38527 = pi19 ? n37 : n38526;
  assign n38528 = pi18 ? n37 : n38527;
  assign n38529 = pi17 ? n37 : n38528;
  assign n38530 = pi16 ? n38525 : n38529;
  assign n38531 = pi15 ? n38521 : n38530;
  assign n38532 = pi21 ? n20977 : n32;
  assign n38533 = pi20 ? n38532 : n32;
  assign n38534 = pi19 ? n27443 : n38533;
  assign n38535 = pi18 ? n37 : n38534;
  assign n38536 = pi17 ? n37 : n38535;
  assign n38537 = pi16 ? n35220 : n38536;
  assign n38538 = pi19 ? n27443 : n37492;
  assign n38539 = pi18 ? n37 : n38538;
  assign n38540 = pi17 ? n37 : n38539;
  assign n38541 = pi16 ? n34306 : n38540;
  assign n38542 = pi15 ? n38537 : n38541;
  assign n38543 = pi14 ? n38531 : n38542;
  assign n38544 = pi13 ? n38517 : n38543;
  assign n38545 = pi16 ? n34306 : n38074;
  assign n38546 = pi16 ? n38525 : n38078;
  assign n38547 = pi15 ? n38545 : n38546;
  assign n38548 = pi16 ? n34889 : n38078;
  assign n38549 = pi19 ? n20563 : n32933;
  assign n38550 = pi18 ? n31315 : n38549;
  assign n38551 = pi17 ? n32 : n38550;
  assign n38552 = pi19 ? n27535 : n9457;
  assign n38553 = pi18 ? n37 : n38552;
  assign n38554 = pi17 ? n37 : n38553;
  assign n38555 = pi16 ? n38551 : n38554;
  assign n38556 = pi15 ? n38548 : n38555;
  assign n38557 = pi14 ? n38547 : n38556;
  assign n38558 = pi22 ? n316 : n21078;
  assign n38559 = pi21 ? n38558 : n32;
  assign n38560 = pi20 ? n38559 : n32;
  assign n38561 = pi19 ? n37 : n38560;
  assign n38562 = pi18 ? n37 : n38561;
  assign n38563 = pi17 ? n37 : n38562;
  assign n38564 = pi16 ? n34328 : n38563;
  assign n38565 = pi20 ? n36250 : n14844;
  assign n38566 = pi19 ? n20563 : n38565;
  assign n38567 = pi18 ? n31315 : n38566;
  assign n38568 = pi17 ? n32 : n38567;
  assign n38569 = pi19 ? n20972 : n4009;
  assign n38570 = pi18 ? n19124 : n38569;
  assign n38571 = pi17 ? n99 : n38570;
  assign n38572 = pi16 ? n38568 : n38571;
  assign n38573 = pi15 ? n38564 : n38572;
  assign n38574 = pi20 ? n30096 : n30859;
  assign n38575 = pi19 ? n20563 : n38574;
  assign n38576 = pi18 ? n31315 : n38575;
  assign n38577 = pi17 ? n32 : n38576;
  assign n38578 = pi19 ? n29428 : n99;
  assign n38579 = pi19 ? n99 : n776;
  assign n38580 = pi18 ? n38578 : n38579;
  assign n38581 = pi20 ? n10539 : n15263;
  assign n38582 = pi19 ? n38581 : n2243;
  assign n38583 = pi18 ? n38582 : n38098;
  assign n38584 = pi17 ? n38580 : n38583;
  assign n38585 = pi16 ? n38577 : n38584;
  assign n38586 = pi20 ? n31220 : n226;
  assign n38587 = pi19 ? n20563 : n38586;
  assign n38588 = pi18 ? n31315 : n38587;
  assign n38589 = pi17 ? n32 : n38588;
  assign n38590 = pi20 ? n775 : n2243;
  assign n38591 = pi19 ? n26685 : n38590;
  assign n38592 = pi19 ? n157 : n14353;
  assign n38593 = pi18 ? n38591 : n38592;
  assign n38594 = pi17 ? n99 : n38593;
  assign n38595 = pi16 ? n38589 : n38594;
  assign n38596 = pi15 ? n38585 : n38595;
  assign n38597 = pi14 ? n38573 : n38596;
  assign n38598 = pi13 ? n38557 : n38597;
  assign n38599 = pi12 ? n38544 : n38598;
  assign n38600 = pi11 ? n38489 : n38599;
  assign n38601 = pi20 ? n37 : n5405;
  assign n38602 = pi19 ? n32314 : n38601;
  assign n38603 = pi18 ? n31315 : n38602;
  assign n38604 = pi17 ? n32 : n38603;
  assign n38605 = pi20 ? n99 : n5881;
  assign n38606 = pi20 ? n3003 : n9686;
  assign n38607 = pi19 ? n38605 : n38606;
  assign n38608 = pi18 ? n38607 : n38098;
  assign n38609 = pi17 ? n99 : n38608;
  assign n38610 = pi16 ? n38604 : n38609;
  assign n38611 = pi19 ? n34920 : n26407;
  assign n38612 = pi18 ? n31315 : n38611;
  assign n38613 = pi17 ? n32 : n38612;
  assign n38614 = pi19 ? n157 : n4009;
  assign n38615 = pi18 ? n22958 : n38614;
  assign n38616 = pi17 ? n99 : n38615;
  assign n38617 = pi16 ? n38613 : n38616;
  assign n38618 = pi15 ? n38610 : n38617;
  assign n38619 = pi19 ? n32876 : n21611;
  assign n38620 = pi18 ? n31315 : n38619;
  assign n38621 = pi17 ? n32 : n38620;
  assign n38622 = pi21 ? n3759 : n5899;
  assign n38623 = pi20 ? n38622 : n316;
  assign n38624 = pi19 ? n38623 : n4009;
  assign n38625 = pi18 ? n99 : n38624;
  assign n38626 = pi17 ? n99 : n38625;
  assign n38627 = pi16 ? n38621 : n38626;
  assign n38628 = pi20 ? n14844 : n14887;
  assign n38629 = pi19 ? n38628 : n99;
  assign n38630 = pi18 ? n34262 : n38629;
  assign n38631 = pi20 ? n99 : n316;
  assign n38632 = pi19 ? n38631 : n4009;
  assign n38633 = pi18 ? n99 : n38632;
  assign n38634 = pi17 ? n38630 : n38633;
  assign n38635 = pi16 ? n38071 : n38634;
  assign n38636 = pi15 ? n38627 : n38635;
  assign n38637 = pi14 ? n38618 : n38636;
  assign n38638 = pi20 ? n3039 : n99;
  assign n38639 = pi19 ? n35776 : n38638;
  assign n38640 = pi18 ? n31938 : n38639;
  assign n38641 = pi17 ? n32 : n38640;
  assign n38642 = pi17 ? n99 : n38633;
  assign n38643 = pi16 ? n38641 : n38642;
  assign n38644 = pi19 ? n32314 : n34261;
  assign n38645 = pi18 ? n31938 : n38644;
  assign n38646 = pi17 ? n32 : n38645;
  assign n38647 = pi18 ? n15029 : n139;
  assign n38648 = pi19 ? n18327 : n3211;
  assign n38649 = pi18 ? n139 : n38648;
  assign n38650 = pi17 ? n38647 : n38649;
  assign n38651 = pi16 ? n38646 : n38650;
  assign n38652 = pi15 ? n38643 : n38651;
  assign n38653 = pi19 ? n32314 : n9795;
  assign n38654 = pi18 ? n31315 : n38653;
  assign n38655 = pi17 ? n32 : n38654;
  assign n38656 = pi20 ? n139 : n1027;
  assign n38657 = pi19 ? n38656 : n10012;
  assign n38658 = pi18 ? n139 : n38657;
  assign n38659 = pi17 ? n139 : n38658;
  assign n38660 = pi16 ? n38655 : n38659;
  assign n38661 = pi19 ? n32898 : n27331;
  assign n38662 = pi18 ? n31315 : n38661;
  assign n38663 = pi17 ? n32 : n38662;
  assign n38664 = pi20 ? n992 : n3086;
  assign n38665 = pi19 ? n139 : n38664;
  assign n38666 = pi20 ? n947 : n992;
  assign n38667 = pi19 ? n38666 : n139;
  assign n38668 = pi18 ? n38665 : n38667;
  assign n38669 = pi19 ? n16473 : n2555;
  assign n38670 = pi18 ? n139 : n38669;
  assign n38671 = pi17 ? n38668 : n38670;
  assign n38672 = pi16 ? n38663 : n38671;
  assign n38673 = pi15 ? n38660 : n38672;
  assign n38674 = pi14 ? n38652 : n38673;
  assign n38675 = pi13 ? n38637 : n38674;
  assign n38676 = pi17 ? n11568 : n38670;
  assign n38677 = pi16 ? n34360 : n38676;
  assign n38678 = pi18 ? n31315 : n32315;
  assign n38679 = pi17 ? n32 : n38678;
  assign n38680 = pi18 ? n14115 : n9770;
  assign n38681 = pi20 ? n1026 : n204;
  assign n38682 = pi19 ? n38681 : n2555;
  assign n38683 = pi18 ? n139 : n38682;
  assign n38684 = pi17 ? n38680 : n38683;
  assign n38685 = pi16 ? n38679 : n38684;
  assign n38686 = pi15 ? n38677 : n38685;
  assign n38687 = pi19 ? n32314 : n20722;
  assign n38688 = pi18 ? n31315 : n38687;
  assign n38689 = pi17 ? n32 : n38688;
  assign n38690 = pi19 ? n30225 : n139;
  assign n38691 = pi18 ? n38690 : n139;
  assign n38692 = pi19 ? n26742 : n2680;
  assign n38693 = pi18 ? n139 : n38692;
  assign n38694 = pi17 ? n38691 : n38693;
  assign n38695 = pi16 ? n38689 : n38694;
  assign n38696 = pi19 ? n37 : n38434;
  assign n38697 = pi19 ? n20782 : n12589;
  assign n38698 = pi18 ? n38696 : n38697;
  assign n38699 = pi20 ? n5199 : n1016;
  assign n38700 = pi19 ? n38699 : n23039;
  assign n38701 = pi20 ? n2316 : n11809;
  assign n38702 = pi19 ? n38701 : n2680;
  assign n38703 = pi18 ? n38700 : n38702;
  assign n38704 = pi17 ? n38698 : n38703;
  assign n38705 = pi16 ? n33313 : n38704;
  assign n38706 = pi15 ? n38695 : n38705;
  assign n38707 = pi14 ? n38686 : n38706;
  assign n38708 = pi21 ? n569 : n297;
  assign n38709 = pi21 ? n139 : n6376;
  assign n38710 = pi20 ? n38708 : n38709;
  assign n38711 = pi19 ? n15020 : n38710;
  assign n38712 = pi18 ? n24735 : n38711;
  assign n38713 = pi20 ? n6362 : n32669;
  assign n38714 = pi21 ? n233 : n28649;
  assign n38715 = pi20 ? n38714 : n7980;
  assign n38716 = pi19 ? n38713 : n38715;
  assign n38717 = pi19 ? n21107 : n2702;
  assign n38718 = pi18 ? n38716 : n38717;
  assign n38719 = pi17 ? n38712 : n38718;
  assign n38720 = pi16 ? n34360 : n38719;
  assign n38721 = pi18 ? n37 : n22060;
  assign n38722 = pi21 ? n3411 : n233;
  assign n38723 = pi20 ? n38722 : n25125;
  assign n38724 = pi21 ? n2091 : n4920;
  assign n38725 = pi21 ? n6376 : n3411;
  assign n38726 = pi20 ? n38724 : n38725;
  assign n38727 = pi19 ? n38723 : n38726;
  assign n38728 = pi20 ? n16544 : n25965;
  assign n38729 = pi19 ? n38728 : n2702;
  assign n38730 = pi18 ? n38727 : n38729;
  assign n38731 = pi17 ? n38721 : n38730;
  assign n38732 = pi16 ? n34360 : n38731;
  assign n38733 = pi15 ? n38720 : n38732;
  assign n38734 = pi20 ? n233 : n2048;
  assign n38735 = pi19 ? n38734 : n34185;
  assign n38736 = pi20 ? n233 : n26369;
  assign n38737 = pi19 ? n38736 : n1823;
  assign n38738 = pi18 ? n38735 : n38737;
  assign n38739 = pi17 ? n37 : n38738;
  assign n38740 = pi16 ? n34360 : n38739;
  assign n38741 = pi19 ? n27754 : n34185;
  assign n38742 = pi18 ? n38741 : n37693;
  assign n38743 = pi17 ? n37 : n38742;
  assign n38744 = pi16 ? n34360 : n38743;
  assign n38745 = pi15 ? n38740 : n38744;
  assign n38746 = pi14 ? n38733 : n38745;
  assign n38747 = pi13 ? n38707 : n38746;
  assign n38748 = pi12 ? n38675 : n38747;
  assign n38749 = pi20 ? n233 : n23544;
  assign n38750 = pi19 ? n38749 : n32;
  assign n38751 = pi18 ? n37 : n38750;
  assign n38752 = pi17 ? n37 : n38751;
  assign n38753 = pi16 ? n33918 : n38752;
  assign n38754 = pi21 ? n20563 : n36489;
  assign n38755 = pi20 ? n38754 : n37;
  assign n38756 = pi19 ? n38755 : n23838;
  assign n38757 = pi18 ? n31938 : n38756;
  assign n38758 = pi17 ? n32 : n38757;
  assign n38759 = pi20 ? n610 : n570;
  assign n38760 = pi19 ? n606 : n38759;
  assign n38761 = pi19 ? n335 : n611;
  assign n38762 = pi18 ? n38760 : n38761;
  assign n38763 = pi22 ? n233 : n21078;
  assign n38764 = pi21 ? n6376 : n38763;
  assign n38765 = pi20 ? n335 : n38764;
  assign n38766 = pi19 ? n38765 : n32;
  assign n38767 = pi18 ? n335 : n38766;
  assign n38768 = pi17 ? n38762 : n38767;
  assign n38769 = pi16 ? n38758 : n38768;
  assign n38770 = pi15 ? n38753 : n38769;
  assign n38771 = pi19 ? n32898 : n23838;
  assign n38772 = pi18 ? n31938 : n38771;
  assign n38773 = pi17 ? n32 : n38772;
  assign n38774 = pi19 ? n606 : n3384;
  assign n38775 = pi18 ? n38774 : n335;
  assign n38776 = pi20 ? n233 : n14674;
  assign n38777 = pi19 ? n38776 : n32;
  assign n38778 = pi18 ? n335 : n38777;
  assign n38779 = pi17 ? n38775 : n38778;
  assign n38780 = pi16 ? n38773 : n38779;
  assign n38781 = pi19 ? n32898 : n17522;
  assign n38782 = pi18 ? n31938 : n38781;
  assign n38783 = pi17 ? n32 : n38782;
  assign n38784 = pi20 ? n13527 : n14674;
  assign n38785 = pi19 ? n38784 : n32;
  assign n38786 = pi18 ? n335 : n38785;
  assign n38787 = pi17 ? n335 : n38786;
  assign n38788 = pi16 ? n38783 : n38787;
  assign n38789 = pi15 ? n38780 : n38788;
  assign n38790 = pi14 ? n38770 : n38789;
  assign n38791 = pi19 ? n32898 : n22031;
  assign n38792 = pi18 ? n31315 : n38791;
  assign n38793 = pi17 ? n32 : n38792;
  assign n38794 = pi20 ? n6377 : n14674;
  assign n38795 = pi19 ? n38794 : n32;
  assign n38796 = pi18 ? n335 : n38795;
  assign n38797 = pi17 ? n335 : n38796;
  assign n38798 = pi16 ? n38793 : n38797;
  assign n38799 = pi20 ? n5013 : n363;
  assign n38800 = pi19 ? n32898 : n38799;
  assign n38801 = pi18 ? n31315 : n38800;
  assign n38802 = pi17 ? n32 : n38801;
  assign n38803 = pi19 ? n363 : n37753;
  assign n38804 = pi18 ? n38803 : n363;
  assign n38805 = pi21 ? n18411 : n7723;
  assign n38806 = pi20 ? n25965 : n38805;
  assign n38807 = pi19 ? n38806 : n32;
  assign n38808 = pi18 ? n363 : n38807;
  assign n38809 = pi17 ? n38804 : n38808;
  assign n38810 = pi16 ? n38802 : n38809;
  assign n38811 = pi15 ? n38798 : n38810;
  assign n38812 = pi19 ? n23903 : n7731;
  assign n38813 = pi18 ? n38812 : n29441;
  assign n38814 = pi17 ? n37 : n38813;
  assign n38815 = pi16 ? n32901 : n38814;
  assign n38816 = pi20 ? n7747 : n99;
  assign n38817 = pi19 ? n32898 : n38816;
  assign n38818 = pi18 ? n31315 : n38817;
  assign n38819 = pi17 ? n32 : n38818;
  assign n38820 = pi20 ? n27520 : n363;
  assign n38821 = pi19 ? n38820 : n363;
  assign n38822 = pi18 ? n27444 : n38821;
  assign n38823 = pi21 ? n685 : n2320;
  assign n38824 = pi20 ? n24220 : n38823;
  assign n38825 = pi19 ? n38824 : n32;
  assign n38826 = pi18 ? n363 : n38825;
  assign n38827 = pi17 ? n38822 : n38826;
  assign n38828 = pi16 ? n38819 : n38827;
  assign n38829 = pi15 ? n38815 : n38828;
  assign n38830 = pi14 ? n38811 : n38829;
  assign n38831 = pi13 ? n38790 : n38830;
  assign n38832 = pi20 ? n7730 : n3393;
  assign n38833 = pi20 ? n27501 : n3393;
  assign n38834 = pi19 ? n38832 : n38833;
  assign n38835 = pi18 ? n37 : n38834;
  assign n38836 = pi20 ? n15173 : n27506;
  assign n38837 = pi19 ? n27503 : n38836;
  assign n38838 = pi18 ? n38837 : n38825;
  assign n38839 = pi17 ? n38835 : n38838;
  assign n38840 = pi16 ? n32901 : n38839;
  assign n38841 = pi21 ? n2106 : n685;
  assign n38842 = pi20 ? n38841 : n37797;
  assign n38843 = pi19 ? n38842 : n32;
  assign n38844 = pi18 ? n37 : n38843;
  assign n38845 = pi17 ? n37 : n38844;
  assign n38846 = pi16 ? n33918 : n38845;
  assign n38847 = pi15 ? n38840 : n38846;
  assign n38848 = pi20 ? n30868 : n37811;
  assign n38849 = pi19 ? n38848 : n99;
  assign n38850 = pi18 ? n37808 : n38849;
  assign n38851 = pi17 ? n32 : n38850;
  assign n38852 = pi22 ? n685 : n6365;
  assign n38853 = pi21 ? n38852 : n928;
  assign n38854 = pi20 ? n685 : n38853;
  assign n38855 = pi19 ? n38854 : n32;
  assign n38856 = pi18 ? n99 : n38855;
  assign n38857 = pi17 ? n99 : n38856;
  assign n38858 = pi16 ? n38851 : n38857;
  assign n38859 = pi21 ? n2768 : n1009;
  assign n38860 = pi20 ? n7754 : n38859;
  assign n38861 = pi19 ? n38860 : n32;
  assign n38862 = pi18 ? n99 : n38861;
  assign n38863 = pi17 ? n99 : n38862;
  assign n38864 = pi16 ? n38851 : n38863;
  assign n38865 = pi15 ? n38858 : n38864;
  assign n38866 = pi14 ? n38847 : n38865;
  assign n38867 = pi22 ? n33792 : n139;
  assign n38868 = pi21 ? n33792 : n38867;
  assign n38869 = pi20 ? n36659 : n38868;
  assign n38870 = pi19 ? n38869 : n139;
  assign n38871 = pi18 ? n37841 : n38870;
  assign n38872 = pi17 ? n32 : n38871;
  assign n38873 = pi21 ? n139 : n685;
  assign n38874 = pi20 ? n139 : n38873;
  assign n38875 = pi19 ? n139 : n38874;
  assign n38876 = pi18 ? n38875 : n685;
  assign n38877 = pi23 ? n685 : n20004;
  assign n38878 = pi22 ? n685 : n38877;
  assign n38879 = pi21 ? n38878 : n32;
  assign n38880 = pi20 ? n685 : n38879;
  assign n38881 = pi19 ? n38880 : n32;
  assign n38882 = pi18 ? n685 : n38881;
  assign n38883 = pi17 ? n38876 : n38882;
  assign n38884 = pi16 ? n38872 : n38883;
  assign n38885 = pi20 ? n36659 : n36781;
  assign n38886 = pi20 ? n34202 : n363;
  assign n38887 = pi19 ? n38885 : n38886;
  assign n38888 = pi18 ? n37841 : n38887;
  assign n38889 = pi17 ? n32 : n38888;
  assign n38890 = pi20 ? n29741 : n9456;
  assign n38891 = pi19 ? n38890 : n32;
  assign n38892 = pi18 ? n363 : n38891;
  assign n38893 = pi17 ? n363 : n38892;
  assign n38894 = pi16 ? n38889 : n38893;
  assign n38895 = pi15 ? n38884 : n38894;
  assign n38896 = pi22 ? n37873 : n36798;
  assign n38897 = pi21 ? n38896 : n36798;
  assign n38898 = pi20 ? n32 : n38897;
  assign n38899 = pi19 ? n32 : n38898;
  assign n38900 = pi21 ? n36798 : n37899;
  assign n38901 = pi22 ? n36798 : n36781;
  assign n38902 = pi21 ? n38901 : n36781;
  assign n38903 = pi20 ? n38900 : n38902;
  assign n38904 = pi21 ? n335 : n157;
  assign n38905 = pi22 ? n157 : n335;
  assign n38906 = pi21 ? n38905 : n157;
  assign n38907 = pi20 ? n38904 : n38906;
  assign n38908 = pi19 ? n38903 : n38907;
  assign n38909 = pi18 ? n38899 : n38908;
  assign n38910 = pi17 ? n32 : n38909;
  assign n38911 = pi20 ? n685 : n27551;
  assign n38912 = pi19 ? n7829 : n38911;
  assign n38913 = pi18 ? n36845 : n38912;
  assign n38914 = pi20 ? n36847 : n685;
  assign n38915 = pi20 ? n27551 : n9456;
  assign n38916 = pi19 ? n38915 : n32;
  assign n38917 = pi18 ? n38914 : n38916;
  assign n38918 = pi17 ? n38913 : n38917;
  assign n38919 = pi16 ? n38910 : n38918;
  assign n38920 = pi21 ? n37874 : n36798;
  assign n38921 = pi20 ? n32 : n38920;
  assign n38922 = pi19 ? n32 : n38921;
  assign n38923 = pi21 ? n36798 : n36781;
  assign n38924 = pi21 ? n37878 : n36781;
  assign n38925 = pi20 ? n38923 : n38924;
  assign n38926 = pi23 ? n335 : n36659;
  assign n38927 = pi22 ? n38926 : n10400;
  assign n38928 = pi21 ? n38927 : n157;
  assign n38929 = pi20 ? n38928 : n157;
  assign n38930 = pi19 ? n38925 : n38929;
  assign n38931 = pi18 ? n38922 : n38930;
  assign n38932 = pi17 ? n32 : n38931;
  assign n38933 = pi22 ? n316 : n1407;
  assign n38934 = pi21 ? n38933 : n32;
  assign n38935 = pi20 ? n34537 : n38934;
  assign n38936 = pi19 ? n38935 : n32;
  assign n38937 = pi18 ? n157 : n38936;
  assign n38938 = pi17 ? n157 : n38937;
  assign n38939 = pi16 ? n38932 : n38938;
  assign n38940 = pi15 ? n38919 : n38939;
  assign n38941 = pi14 ? n38895 : n38940;
  assign n38942 = pi13 ? n38866 : n38941;
  assign n38943 = pi12 ? n38831 : n38942;
  assign n38944 = pi11 ? n38748 : n38943;
  assign n38945 = pi10 ? n38600 : n38944;
  assign n38946 = pi09 ? n38356 : n38945;
  assign n38947 = pi20 ? n37320 : n20563;
  assign n38948 = pi19 ? n38947 : n20563;
  assign n38949 = pi18 ? n32 : n38948;
  assign n38950 = pi17 ? n32 : n38949;
  assign n38951 = pi19 ? n20563 : n32314;
  assign n38952 = pi18 ? n38951 : n38320;
  assign n38953 = pi17 ? n38952 : n38326;
  assign n38954 = pi16 ? n38950 : n38953;
  assign n38955 = pi15 ? n32 : n38954;
  assign n38956 = pi20 ? n37333 : n20563;
  assign n38957 = pi19 ? n38956 : n20563;
  assign n38958 = pi18 ? n32 : n38957;
  assign n38959 = pi17 ? n32 : n38958;
  assign n38960 = pi16 ? n38959 : n38338;
  assign n38961 = pi21 ? n20563 : n31877;
  assign n38962 = pi20 ? n20563 : n38961;
  assign n38963 = pi19 ? n20563 : n38962;
  assign n38964 = pi18 ? n32 : n38963;
  assign n38965 = pi17 ? n32 : n38964;
  assign n38966 = pi21 ? n31924 : n20563;
  assign n38967 = pi20 ? n38966 : n36946;
  assign n38968 = pi19 ? n38967 : n38341;
  assign n38969 = pi21 ? n37 : n1143;
  assign n38970 = pi20 ? n38969 : n226;
  assign n38971 = pi19 ? n38970 : n99;
  assign n38972 = pi18 ? n38968 : n38971;
  assign n38973 = pi17 ? n38972 : n38348;
  assign n38974 = pi16 ? n38965 : n38973;
  assign n38975 = pi15 ? n38960 : n38974;
  assign n38976 = pi14 ? n38955 : n38975;
  assign n38977 = pi13 ? n32 : n38976;
  assign n38978 = pi12 ? n32 : n38977;
  assign n38979 = pi11 ? n32 : n38978;
  assign n38980 = pi10 ? n32 : n38979;
  assign n38981 = pi21 ? n32 : n38375;
  assign n38982 = pi20 ? n32 : n38981;
  assign n38983 = pi19 ? n32 : n38982;
  assign n38984 = pi18 ? n38983 : n20563;
  assign n38985 = pi17 ? n32 : n38984;
  assign n38986 = pi21 ? n112 : n3066;
  assign n38987 = pi20 ? n38986 : n32;
  assign n38988 = pi19 ? n17972 : n38987;
  assign n38989 = pi18 ? n38362 : n38988;
  assign n38990 = pi17 ? n38360 : n38989;
  assign n38991 = pi16 ? n38985 : n38990;
  assign n38992 = pi18 ? n33260 : n37;
  assign n38993 = pi17 ? n38992 : n38371;
  assign n38994 = pi16 ? n36871 : n38993;
  assign n38995 = pi15 ? n38991 : n38994;
  assign n38996 = pi16 ? n37959 : n38387;
  assign n38997 = pi21 ? n32 : n30866;
  assign n38998 = pi20 ? n32 : n38997;
  assign n38999 = pi19 ? n32 : n38998;
  assign n39000 = pi18 ? n38999 : n20563;
  assign n39001 = pi17 ? n32 : n39000;
  assign n39002 = pi20 ? n36879 : n37;
  assign n39003 = pi19 ? n20563 : n39002;
  assign n39004 = pi18 ? n39003 : n37;
  assign n39005 = pi17 ? n39004 : n38386;
  assign n39006 = pi16 ? n39001 : n39005;
  assign n39007 = pi15 ? n38996 : n39006;
  assign n39008 = pi14 ? n38995 : n39007;
  assign n39009 = pi19 ? n9795 : n10645;
  assign n39010 = pi18 ? n38398 : n39009;
  assign n39011 = pi17 ? n38395 : n39010;
  assign n39012 = pi16 ? n36216 : n39011;
  assign n39013 = pi19 ? n38410 : n10645;
  assign n39014 = pi18 ? n38409 : n39013;
  assign n39015 = pi17 ? n38406 : n39014;
  assign n39016 = pi16 ? n36216 : n39015;
  assign n39017 = pi15 ? n39012 : n39016;
  assign n39018 = pi18 ? n38421 : n39013;
  assign n39019 = pi17 ? n38418 : n39018;
  assign n39020 = pi16 ? n36216 : n39019;
  assign n39021 = pi19 ? n9814 : n10645;
  assign n39022 = pi18 ? n34307 : n39021;
  assign n39023 = pi17 ? n38425 : n39022;
  assign n39024 = pi16 ? n36216 : n39023;
  assign n39025 = pi15 ? n39020 : n39024;
  assign n39026 = pi14 ? n39017 : n39025;
  assign n39027 = pi13 ? n39008 : n39026;
  assign n39028 = pi20 ? n24781 : n32;
  assign n39029 = pi19 ? n38436 : n39028;
  assign n39030 = pi18 ? n38435 : n39029;
  assign n39031 = pi17 ? n38433 : n39030;
  assign n39032 = pi16 ? n36216 : n39031;
  assign n39033 = pi19 ? n7676 : n39028;
  assign n39034 = pi18 ? n37 : n39033;
  assign n39035 = pi17 ? n38443 : n39034;
  assign n39036 = pi16 ? n36216 : n39035;
  assign n39037 = pi15 ? n39032 : n39036;
  assign n39038 = pi19 ? n36897 : n37;
  assign n39039 = pi18 ? n39038 : n37;
  assign n39040 = pi21 ? n335 : n2637;
  assign n39041 = pi20 ? n39040 : n32;
  assign n39042 = pi19 ? n3332 : n39041;
  assign n39043 = pi18 ? n37 : n39042;
  assign n39044 = pi17 ? n39039 : n39043;
  assign n39045 = pi16 ? n36216 : n39044;
  assign n39046 = pi21 ? n335 : n928;
  assign n39047 = pi20 ? n39046 : n32;
  assign n39048 = pi19 ? n37 : n39047;
  assign n39049 = pi18 ? n37 : n39048;
  assign n39050 = pi17 ? n38455 : n39049;
  assign n39051 = pi16 ? n36216 : n39050;
  assign n39052 = pi15 ? n39045 : n39051;
  assign n39053 = pi14 ? n39037 : n39052;
  assign n39054 = pi20 ? n25760 : n32;
  assign n39055 = pi19 ? n37 : n39054;
  assign n39056 = pi18 ? n37 : n39055;
  assign n39057 = pi17 ? n36210 : n39056;
  assign n39058 = pi16 ? n36216 : n39057;
  assign n39059 = pi15 ? n39058 : n38474;
  assign n39060 = pi16 ? n35220 : n38473;
  assign n39061 = pi18 ? n31938 : n38479;
  assign n39062 = pi17 ? n32 : n39061;
  assign n39063 = pi16 ? n39062 : n38484;
  assign n39064 = pi15 ? n39060 : n39063;
  assign n39065 = pi14 ? n39059 : n39064;
  assign n39066 = pi13 ? n39053 : n39065;
  assign n39067 = pi12 ? n39027 : n39066;
  assign n39068 = pi19 ? n644 : n11186;
  assign n39069 = pi18 ? n37 : n39068;
  assign n39070 = pi17 ? n37 : n39069;
  assign n39071 = pi16 ? n38032 : n39070;
  assign n39072 = pi15 ? n38500 : n39071;
  assign n39073 = pi19 ? n20563 : n35854;
  assign n39074 = pi18 ? n31315 : n39073;
  assign n39075 = pi17 ? n32 : n39074;
  assign n39076 = pi16 ? n39075 : n38510;
  assign n39077 = pi15 ? n39076 : n38515;
  assign n39078 = pi14 ? n39072 : n39077;
  assign n39079 = pi20 ? n31925 : n33821;
  assign n39080 = pi19 ? n20563 : n39079;
  assign n39081 = pi18 ? n31315 : n39080;
  assign n39082 = pi17 ? n32 : n39081;
  assign n39083 = pi16 ? n39082 : n38529;
  assign n39084 = pi15 ? n38521 : n39083;
  assign n39085 = pi18 ? n31315 : n38951;
  assign n39086 = pi17 ? n32 : n39085;
  assign n39087 = pi16 ? n39086 : n38536;
  assign n39088 = pi20 ? n25336 : n32;
  assign n39089 = pi19 ? n27443 : n39088;
  assign n39090 = pi18 ? n37 : n39089;
  assign n39091 = pi17 ? n37 : n39090;
  assign n39092 = pi16 ? n34306 : n39091;
  assign n39093 = pi15 ? n39087 : n39092;
  assign n39094 = pi14 ? n39084 : n39093;
  assign n39095 = pi13 ? n39078 : n39094;
  assign n39096 = pi19 ? n37 : n11675;
  assign n39097 = pi18 ? n37 : n39096;
  assign n39098 = pi17 ? n37 : n39097;
  assign n39099 = pi16 ? n34306 : n39098;
  assign n39100 = pi19 ? n37 : n12129;
  assign n39101 = pi18 ? n37 : n39100;
  assign n39102 = pi17 ? n37 : n39101;
  assign n39103 = pi16 ? n38525 : n39102;
  assign n39104 = pi15 ? n39099 : n39103;
  assign n39105 = pi18 ? n31315 : n32872;
  assign n39106 = pi17 ? n32 : n39105;
  assign n39107 = pi16 ? n39106 : n39102;
  assign n39108 = pi19 ? n27535 : n11696;
  assign n39109 = pi18 ? n37 : n39108;
  assign n39110 = pi17 ? n37 : n39109;
  assign n39111 = pi16 ? n34328 : n39110;
  assign n39112 = pi15 ? n39107 : n39111;
  assign n39113 = pi14 ? n39104 : n39112;
  assign n39114 = pi19 ? n37 : n5668;
  assign n39115 = pi18 ? n37 : n39114;
  assign n39116 = pi17 ? n37 : n39115;
  assign n39117 = pi16 ? n34328 : n39116;
  assign n39118 = pi21 ? n31877 : n37;
  assign n39119 = pi20 ? n39118 : n14844;
  assign n39120 = pi19 ? n20563 : n39119;
  assign n39121 = pi18 ? n31315 : n39120;
  assign n39122 = pi17 ? n32 : n39121;
  assign n39123 = pi19 ? n20972 : n5668;
  assign n39124 = pi18 ? n19124 : n39123;
  assign n39125 = pi17 ? n99 : n39124;
  assign n39126 = pi16 ? n39122 : n39125;
  assign n39127 = pi15 ? n39117 : n39126;
  assign n39128 = pi20 ? n31220 : n5077;
  assign n39129 = pi19 ? n20563 : n39128;
  assign n39130 = pi18 ? n31315 : n39129;
  assign n39131 = pi17 ? n32 : n39130;
  assign n39132 = pi21 ? n16841 : n32;
  assign n39133 = pi20 ? n39132 : n32;
  assign n39134 = pi19 ? n157 : n39133;
  assign n39135 = pi18 ? n38582 : n39134;
  assign n39136 = pi17 ? n38580 : n39135;
  assign n39137 = pi16 ? n39131 : n39136;
  assign n39138 = pi19 ? n157 : n13430;
  assign n39139 = pi18 ? n38591 : n39138;
  assign n39140 = pi17 ? n99 : n39139;
  assign n39141 = pi16 ? n38589 : n39140;
  assign n39142 = pi15 ? n39137 : n39141;
  assign n39143 = pi14 ? n39127 : n39142;
  assign n39144 = pi13 ? n39113 : n39143;
  assign n39145 = pi12 ? n39095 : n39144;
  assign n39146 = pi11 ? n39067 : n39145;
  assign n39147 = pi19 ? n32876 : n35209;
  assign n39148 = pi18 ? n31315 : n39147;
  assign n39149 = pi17 ? n32 : n39148;
  assign n39150 = pi20 ? n7824 : n9686;
  assign n39151 = pi19 ? n38605 : n39150;
  assign n39152 = pi18 ? n39151 : n39134;
  assign n39153 = pi17 ? n99 : n39152;
  assign n39154 = pi16 ? n39149 : n39153;
  assign n39155 = pi19 ? n20563 : n26407;
  assign n39156 = pi18 ? n31315 : n39155;
  assign n39157 = pi17 ? n32 : n39156;
  assign n39158 = pi20 ? n26293 : n32;
  assign n39159 = pi19 ? n157 : n39158;
  assign n39160 = pi18 ? n22958 : n39159;
  assign n39161 = pi17 ? n99 : n39160;
  assign n39162 = pi16 ? n39157 : n39161;
  assign n39163 = pi15 ? n39154 : n39162;
  assign n39164 = pi22 ? n30869 : n37;
  assign n39165 = pi21 ? n39164 : n99;
  assign n39166 = pi20 ? n39165 : n99;
  assign n39167 = pi19 ? n20563 : n39166;
  assign n39168 = pi18 ? n31315 : n39167;
  assign n39169 = pi17 ? n32 : n39168;
  assign n39170 = pi16 ? n39169 : n38626;
  assign n39171 = pi16 ? n38679 : n38634;
  assign n39172 = pi15 ? n39170 : n39171;
  assign n39173 = pi14 ? n39163 : n39172;
  assign n39174 = pi23 ? n30868 : n37;
  assign n39175 = pi22 ? n30195 : n39174;
  assign n39176 = pi21 ? n20563 : n39175;
  assign n39177 = pi20 ? n20563 : n39176;
  assign n39178 = pi19 ? n39177 : n38638;
  assign n39179 = pi18 ? n31315 : n39178;
  assign n39180 = pi17 ? n32 : n39179;
  assign n39181 = pi16 ? n39180 : n38642;
  assign n39182 = pi22 ? n39174 : n37;
  assign n39183 = pi21 ? n39182 : n37;
  assign n39184 = pi20 ? n39183 : n14844;
  assign n39185 = pi19 ? n34920 : n39184;
  assign n39186 = pi18 ? n31315 : n39185;
  assign n39187 = pi17 ? n32 : n39186;
  assign n39188 = pi16 ? n39187 : n38650;
  assign n39189 = pi15 ? n39181 : n39188;
  assign n39190 = pi23 ? n20563 : n30868;
  assign n39191 = pi22 ? n20563 : n39190;
  assign n39192 = pi21 ? n20563 : n39191;
  assign n39193 = pi20 ? n20563 : n39192;
  assign n39194 = pi20 ? n31903 : n139;
  assign n39195 = pi19 ? n39193 : n39194;
  assign n39196 = pi18 ? n31315 : n39195;
  assign n39197 = pi17 ? n32 : n39196;
  assign n39198 = pi21 ? n1027 : n16438;
  assign n39199 = pi20 ? n139 : n39198;
  assign n39200 = pi19 ? n39199 : n10012;
  assign n39201 = pi18 ? n139 : n39200;
  assign n39202 = pi17 ? n139 : n39201;
  assign n39203 = pi16 ? n39197 : n39202;
  assign n39204 = pi19 ? n32898 : n9765;
  assign n39205 = pi18 ? n31938 : n39204;
  assign n39206 = pi17 ? n32 : n39205;
  assign n39207 = pi19 ? n16473 : n2580;
  assign n39208 = pi18 ? n139 : n39207;
  assign n39209 = pi17 ? n38668 : n39208;
  assign n39210 = pi16 ? n39206 : n39209;
  assign n39211 = pi15 ? n39203 : n39210;
  assign n39212 = pi14 ? n39189 : n39211;
  assign n39213 = pi13 ? n39173 : n39212;
  assign n39214 = pi18 ? n31938 : n35855;
  assign n39215 = pi17 ? n32 : n39214;
  assign n39216 = pi19 ? n16473 : n2639;
  assign n39217 = pi18 ? n139 : n39216;
  assign n39218 = pi17 ? n11568 : n39217;
  assign n39219 = pi16 ? n39215 : n39218;
  assign n39220 = pi21 ? n23795 : n32;
  assign n39221 = pi20 ? n39220 : n32;
  assign n39222 = pi19 ? n38681 : n39221;
  assign n39223 = pi18 ? n139 : n39222;
  assign n39224 = pi17 ? n38680 : n39223;
  assign n39225 = pi16 ? n33313 : n39224;
  assign n39226 = pi15 ? n39219 : n39225;
  assign n39227 = pi19 ? n32294 : n20722;
  assign n39228 = pi18 ? n31315 : n39227;
  assign n39229 = pi17 ? n32 : n39228;
  assign n39230 = pi19 ? n26742 : n2654;
  assign n39231 = pi18 ? n139 : n39230;
  assign n39232 = pi17 ? n38691 : n39231;
  assign n39233 = pi16 ? n39229 : n39232;
  assign n39234 = pi15 ? n39233 : n38705;
  assign n39235 = pi14 ? n39226 : n39234;
  assign n39236 = pi16 ? n34923 : n38719;
  assign n39237 = pi18 ? n37 : n22538;
  assign n39238 = pi21 ? n6376 : n26360;
  assign n39239 = pi20 ? n38724 : n39238;
  assign n39240 = pi19 ? n25125 : n39239;
  assign n39241 = pi19 ? n38728 : n1823;
  assign n39242 = pi18 ? n39240 : n39241;
  assign n39243 = pi17 ? n39237 : n39242;
  assign n39244 = pi16 ? n34923 : n39243;
  assign n39245 = pi15 ? n39236 : n39244;
  assign n39246 = pi16 ? n35857 : n38739;
  assign n39247 = pi16 ? n35857 : n38743;
  assign n39248 = pi15 ? n39246 : n39247;
  assign n39249 = pi14 ? n39245 : n39248;
  assign n39250 = pi13 ? n39235 : n39249;
  assign n39251 = pi12 ? n39213 : n39250;
  assign n39252 = pi16 ? n35857 : n38752;
  assign n39253 = pi20 ? n38754 : n33964;
  assign n39254 = pi19 ? n39253 : n23838;
  assign n39255 = pi18 ? n31315 : n39254;
  assign n39256 = pi17 ? n32 : n39255;
  assign n39257 = pi21 ? n6376 : n8916;
  assign n39258 = pi20 ? n335 : n39257;
  assign n39259 = pi19 ? n39258 : n32;
  assign n39260 = pi18 ? n335 : n39259;
  assign n39261 = pi17 ? n38762 : n39260;
  assign n39262 = pi16 ? n39256 : n39261;
  assign n39263 = pi15 ? n39252 : n39262;
  assign n39264 = pi19 ? n33822 : n23838;
  assign n39265 = pi18 ? n31315 : n39264;
  assign n39266 = pi17 ? n32 : n39265;
  assign n39267 = pi20 ? n233 : n15162;
  assign n39268 = pi19 ? n39267 : n32;
  assign n39269 = pi18 ? n335 : n39268;
  assign n39270 = pi17 ? n38775 : n39269;
  assign n39271 = pi16 ? n39266 : n39270;
  assign n39272 = pi19 ? n33822 : n17204;
  assign n39273 = pi18 ? n31315 : n39272;
  assign n39274 = pi17 ? n32 : n39273;
  assign n39275 = pi20 ? n13527 : n15162;
  assign n39276 = pi19 ? n39275 : n32;
  assign n39277 = pi18 ? n335 : n39276;
  assign n39278 = pi17 ? n335 : n39277;
  assign n39279 = pi16 ? n39274 : n39278;
  assign n39280 = pi15 ? n39271 : n39279;
  assign n39281 = pi14 ? n39263 : n39280;
  assign n39282 = pi19 ? n33905 : n22031;
  assign n39283 = pi18 ? n31315 : n39282;
  assign n39284 = pi17 ? n32 : n39283;
  assign n39285 = pi16 ? n39284 : n38797;
  assign n39286 = pi19 ? n33905 : n23917;
  assign n39287 = pi18 ? n31315 : n39286;
  assign n39288 = pi17 ? n32 : n39287;
  assign n39289 = pi16 ? n39288 : n38809;
  assign n39290 = pi15 ? n39285 : n39289;
  assign n39291 = pi23 ? n33792 : n37;
  assign n39292 = pi22 ? n20563 : n39291;
  assign n39293 = pi21 ? n39292 : n30843;
  assign n39294 = pi20 ? n20563 : n39293;
  assign n39295 = pi19 ? n39294 : n37;
  assign n39296 = pi18 ? n31315 : n39295;
  assign n39297 = pi17 ? n32 : n39296;
  assign n39298 = pi16 ? n39297 : n38814;
  assign n39299 = pi19 ? n39294 : n38816;
  assign n39300 = pi18 ? n31315 : n39299;
  assign n39301 = pi17 ? n32 : n39300;
  assign n39302 = pi16 ? n39301 : n38827;
  assign n39303 = pi15 ? n39298 : n39302;
  assign n39304 = pi14 ? n39290 : n39303;
  assign n39305 = pi13 ? n39281 : n39304;
  assign n39306 = pi22 ? n20563 : n36660;
  assign n39307 = pi21 ? n39306 : n30843;
  assign n39308 = pi20 ? n20563 : n39307;
  assign n39309 = pi19 ? n39308 : n37;
  assign n39310 = pi18 ? n31315 : n39309;
  assign n39311 = pi17 ? n32 : n39310;
  assign n39312 = pi16 ? n39311 : n38839;
  assign n39313 = pi16 ? n38679 : n38845;
  assign n39314 = pi15 ? n39312 : n39313;
  assign n39315 = pi22 ? n37809 : n99;
  assign n39316 = pi21 ? n30868 : n39315;
  assign n39317 = pi20 ? n30868 : n39316;
  assign n39318 = pi19 ? n39317 : n99;
  assign n39319 = pi18 ? n37808 : n39318;
  assign n39320 = pi17 ? n32 : n39319;
  assign n39321 = pi22 ? n685 : n1070;
  assign n39322 = pi21 ? n39321 : n928;
  assign n39323 = pi20 ? n685 : n39322;
  assign n39324 = pi19 ? n39323 : n32;
  assign n39325 = pi18 ? n99 : n39324;
  assign n39326 = pi17 ? n99 : n39325;
  assign n39327 = pi16 ? n39320 : n39326;
  assign n39328 = pi21 ? n5113 : n1009;
  assign n39329 = pi20 ? n7754 : n39328;
  assign n39330 = pi19 ? n39329 : n32;
  assign n39331 = pi18 ? n99 : n39330;
  assign n39332 = pi17 ? n99 : n39331;
  assign n39333 = pi16 ? n39320 : n39332;
  assign n39334 = pi15 ? n39327 : n39333;
  assign n39335 = pi14 ? n39314 : n39334;
  assign n39336 = pi21 ? n33792 : n37253;
  assign n39337 = pi20 ? n36659 : n39336;
  assign n39338 = pi19 ? n39337 : n139;
  assign n39339 = pi18 ? n37841 : n39338;
  assign n39340 = pi17 ? n32 : n39339;
  assign n39341 = pi16 ? n39340 : n38883;
  assign n39342 = pi22 ? n36785 : n139;
  assign n39343 = pi21 ? n39342 : n20228;
  assign n39344 = pi20 ? n39343 : n363;
  assign n39345 = pi19 ? n38885 : n39344;
  assign n39346 = pi18 ? n37841 : n39345;
  assign n39347 = pi17 ? n32 : n39346;
  assign n39348 = pi16 ? n39347 : n38893;
  assign n39349 = pi15 ? n39341 : n39348;
  assign n39350 = pi22 ? n36801 : n335;
  assign n39351 = pi21 ? n39350 : n157;
  assign n39352 = pi20 ? n39351 : n38906;
  assign n39353 = pi19 ? n38903 : n39352;
  assign n39354 = pi18 ? n38899 : n39353;
  assign n39355 = pi17 ? n32 : n39354;
  assign n39356 = pi16 ? n39355 : n38918;
  assign n39357 = pi22 ? n37288 : n363;
  assign n39358 = pi21 ? n39357 : n157;
  assign n39359 = pi20 ? n39358 : n157;
  assign n39360 = pi19 ? n38925 : n39359;
  assign n39361 = pi18 ? n38922 : n39360;
  assign n39362 = pi17 ? n32 : n39361;
  assign n39363 = pi16 ? n39362 : n38938;
  assign n39364 = pi15 ? n39356 : n39363;
  assign n39365 = pi14 ? n39349 : n39364;
  assign n39366 = pi13 ? n39335 : n39365;
  assign n39367 = pi12 ? n39305 : n39366;
  assign n39368 = pi11 ? n39251 : n39367;
  assign n39369 = pi10 ? n39146 : n39368;
  assign n39370 = pi09 ? n38980 : n39369;
  assign n39371 = pi08 ? n38946 : n39370;
  assign n39372 = pi20 ? n37933 : n20563;
  assign n39373 = pi19 ? n39372 : n20563;
  assign n39374 = pi18 ? n32 : n39373;
  assign n39375 = pi17 ? n32 : n39374;
  assign n39376 = pi20 ? n37 : n15964;
  assign n39377 = pi19 ? n37 : n39376;
  assign n39378 = pi18 ? n20563 : n39377;
  assign n39379 = pi20 ? n3884 : n99;
  assign n39380 = pi19 ? n39379 : n99;
  assign n39381 = pi20 ? n25235 : n32;
  assign n39382 = pi19 ? n29428 : n39381;
  assign n39383 = pi18 ? n39380 : n39382;
  assign n39384 = pi17 ? n39378 : n39383;
  assign n39385 = pi16 ? n39375 : n39384;
  assign n39386 = pi15 ? n32 : n39385;
  assign n39387 = pi20 ? n37 : n3042;
  assign n39388 = pi19 ? n37 : n39387;
  assign n39389 = pi18 ? n20563 : n39388;
  assign n39390 = pi19 ? n99 : n39381;
  assign n39391 = pi18 ? n99 : n39390;
  assign n39392 = pi17 ? n39389 : n39391;
  assign n39393 = pi16 ? n38959 : n39392;
  assign n39394 = pi22 ? n32 : n30865;
  assign n39395 = pi21 ? n39394 : n20563;
  assign n39396 = pi20 ? n39395 : n20563;
  assign n39397 = pi19 ? n39396 : n20563;
  assign n39398 = pi18 ? n32 : n39397;
  assign n39399 = pi17 ? n32 : n39398;
  assign n39400 = pi20 ? n5077 : n226;
  assign n39401 = pi19 ? n39400 : n99;
  assign n39402 = pi18 ? n34865 : n39401;
  assign n39403 = pi21 ? n99 : n18039;
  assign n39404 = pi20 ? n39403 : n32;
  assign n39405 = pi19 ? n99 : n39404;
  assign n39406 = pi18 ? n99 : n39405;
  assign n39407 = pi17 ? n39402 : n39406;
  assign n39408 = pi16 ? n39399 : n39407;
  assign n39409 = pi15 ? n39393 : n39408;
  assign n39410 = pi14 ? n39386 : n39409;
  assign n39411 = pi13 ? n32 : n39410;
  assign n39412 = pi12 ? n32 : n39411;
  assign n39413 = pi11 ? n32 : n39412;
  assign n39414 = pi10 ? n32 : n39413;
  assign n39415 = pi18 ? n34258 : n37;
  assign n39416 = pi20 ? n181 : n219;
  assign n39417 = pi19 ? n37 : n39416;
  assign n39418 = pi20 ? n2973 : n7745;
  assign n39419 = pi21 ? n37 : n18051;
  assign n39420 = pi20 ? n39419 : n32;
  assign n39421 = pi19 ? n39418 : n39420;
  assign n39422 = pi18 ? n39417 : n39421;
  assign n39423 = pi17 ? n39415 : n39422;
  assign n39424 = pi16 ? n38331 : n39423;
  assign n39425 = pi21 ? n37 : n12003;
  assign n39426 = pi20 ? n39425 : n32;
  assign n39427 = pi19 ? n37 : n39426;
  assign n39428 = pi18 ? n37 : n39427;
  assign n39429 = pi17 ? n39415 : n39428;
  assign n39430 = pi16 ? n37930 : n39429;
  assign n39431 = pi15 ? n39424 : n39430;
  assign n39432 = pi19 ? n20563 : n33905;
  assign n39433 = pi18 ? n39432 : n37;
  assign n39434 = pi21 ? n37 : n33397;
  assign n39435 = pi20 ? n39434 : n32;
  assign n39436 = pi19 ? n37 : n39435;
  assign n39437 = pi18 ? n37 : n39436;
  assign n39438 = pi17 ? n39433 : n39437;
  assign n39439 = pi16 ? n37959 : n39438;
  assign n39440 = pi18 ? n33245 : n37;
  assign n39441 = pi19 ? n37 : n9240;
  assign n39442 = pi18 ? n37 : n39441;
  assign n39443 = pi17 ? n39440 : n39442;
  assign n39444 = pi16 ? n37324 : n39443;
  assign n39445 = pi15 ? n39439 : n39444;
  assign n39446 = pi14 ? n39431 : n39445;
  assign n39447 = pi19 ? n20563 : n31926;
  assign n39448 = pi18 ? n39447 : n37;
  assign n39449 = pi20 ? n14057 : n1003;
  assign n39450 = pi19 ? n9824 : n39449;
  assign n39451 = pi18 ? n39450 : n39009;
  assign n39452 = pi17 ? n39448 : n39451;
  assign n39453 = pi16 ? n38380 : n39452;
  assign n39454 = pi20 ? n32 : n39395;
  assign n39455 = pi19 ? n32 : n39454;
  assign n39456 = pi18 ? n39455 : n20563;
  assign n39457 = pi17 ? n32 : n39456;
  assign n39458 = pi19 ? n29248 : n10645;
  assign n39459 = pi18 ? n37 : n39458;
  assign n39460 = pi17 ? n39448 : n39459;
  assign n39461 = pi16 ? n39457 : n39460;
  assign n39462 = pi15 ? n39453 : n39461;
  assign n39463 = pi18 ? n35812 : n37;
  assign n39464 = pi19 ? n20722 : n10645;
  assign n39465 = pi18 ? n37 : n39464;
  assign n39466 = pi17 ? n39463 : n39465;
  assign n39467 = pi16 ? n35765 : n39466;
  assign n39468 = pi18 ? n32275 : n37;
  assign n39469 = pi19 ? n3110 : n10645;
  assign n39470 = pi18 ? n37 : n39469;
  assign n39471 = pi17 ? n39468 : n39470;
  assign n39472 = pi16 ? n36216 : n39471;
  assign n39473 = pi15 ? n39467 : n39472;
  assign n39474 = pi14 ? n39462 : n39473;
  assign n39475 = pi13 ? n39446 : n39474;
  assign n39476 = pi18 ? n38549 : n37;
  assign n39477 = pi19 ? n13192 : n39028;
  assign n39478 = pi18 ? n37 : n39477;
  assign n39479 = pi17 ? n39476 : n39478;
  assign n39480 = pi16 ? n36216 : n39479;
  assign n39481 = pi18 ? n33285 : n37;
  assign n39482 = pi17 ? n39481 : n39034;
  assign n39483 = pi16 ? n36216 : n39482;
  assign n39484 = pi15 ? n39480 : n39483;
  assign n39485 = pi19 ? n37 : n39041;
  assign n39486 = pi18 ? n37 : n39485;
  assign n39487 = pi17 ? n39481 : n39486;
  assign n39488 = pi16 ? n36216 : n39487;
  assign n39489 = pi18 ? n32877 : n37;
  assign n39490 = pi17 ? n39489 : n39049;
  assign n39491 = pi16 ? n36216 : n39490;
  assign n39492 = pi15 ? n39488 : n39491;
  assign n39493 = pi14 ? n39484 : n39492;
  assign n39494 = pi18 ? n35855 : n37;
  assign n39495 = pi17 ? n39494 : n39056;
  assign n39496 = pi16 ? n36216 : n39495;
  assign n39497 = pi18 ? n37029 : n37;
  assign n39498 = pi19 ? n38470 : n13340;
  assign n39499 = pi18 ? n37 : n39498;
  assign n39500 = pi17 ? n39497 : n39499;
  assign n39501 = pi16 ? n36216 : n39500;
  assign n39502 = pi15 ? n39496 : n39501;
  assign n39503 = pi19 ? n2095 : n13340;
  assign n39504 = pi18 ? n37 : n39503;
  assign n39505 = pi17 ? n37377 : n39504;
  assign n39506 = pi16 ? n36216 : n39505;
  assign n39507 = pi19 ? n7685 : n13340;
  assign n39508 = pi18 ? n37 : n39507;
  assign n39509 = pi17 ? n38449 : n39508;
  assign n39510 = pi16 ? n36216 : n39509;
  assign n39511 = pi15 ? n39506 : n39510;
  assign n39512 = pi14 ? n39502 : n39511;
  assign n39513 = pi13 ? n39493 : n39512;
  assign n39514 = pi12 ? n39475 : n39513;
  assign n39515 = pi20 ? n19368 : n37;
  assign n39516 = pi19 ? n37 : n39515;
  assign n39517 = pi21 ? n6376 : n2637;
  assign n39518 = pi20 ? n39517 : n32;
  assign n39519 = pi19 ? n7685 : n39518;
  assign n39520 = pi18 ? n39516 : n39519;
  assign n39521 = pi17 ? n38449 : n39520;
  assign n39522 = pi16 ? n36216 : n39521;
  assign n39523 = pi20 ? n22759 : n32;
  assign n39524 = pi19 ? n37 : n39523;
  assign n39525 = pi18 ? n37 : n39524;
  assign n39526 = pi17 ? n38449 : n39525;
  assign n39527 = pi16 ? n36216 : n39526;
  assign n39528 = pi15 ? n39522 : n39527;
  assign n39529 = pi18 ? n33950 : n37;
  assign n39530 = pi19 ? n37 : n12102;
  assign n39531 = pi18 ? n37 : n39530;
  assign n39532 = pi17 ? n39529 : n39531;
  assign n39533 = pi16 ? n36216 : n39532;
  assign n39534 = pi18 ? n32934 : n37;
  assign n39535 = pi20 ? n26207 : n32;
  assign n39536 = pi19 ? n7731 : n39535;
  assign n39537 = pi18 ? n37 : n39536;
  assign n39538 = pi17 ? n39534 : n39537;
  assign n39539 = pi16 ? n36216 : n39538;
  assign n39540 = pi15 ? n39533 : n39539;
  assign n39541 = pi14 ? n39528 : n39540;
  assign n39542 = pi22 ? n37 : n10341;
  assign n39543 = pi21 ? n39542 : n2700;
  assign n39544 = pi20 ? n39543 : n32;
  assign n39545 = pi19 ? n7731 : n39544;
  assign n39546 = pi18 ? n37 : n39545;
  assign n39547 = pi17 ? n36919 : n39546;
  assign n39548 = pi16 ? n36216 : n39547;
  assign n39549 = pi22 ? n363 : n10341;
  assign n39550 = pi21 ? n39549 : n1009;
  assign n39551 = pi20 ? n39550 : n32;
  assign n39552 = pi19 ? n37 : n39551;
  assign n39553 = pi18 ? n37 : n39552;
  assign n39554 = pi17 ? n36210 : n39553;
  assign n39555 = pi16 ? n36216 : n39554;
  assign n39556 = pi15 ? n39548 : n39555;
  assign n39557 = pi23 ? n363 : n24414;
  assign n39558 = pi22 ? n99 : n39557;
  assign n39559 = pi21 ? n39558 : n1009;
  assign n39560 = pi20 ? n39559 : n32;
  assign n39561 = pi19 ? n37 : n39560;
  assign n39562 = pi18 ? n37 : n39561;
  assign n39563 = pi17 ? n39534 : n39562;
  assign n39564 = pi16 ? n36923 : n39563;
  assign n39565 = pi19 ? n37 : n11216;
  assign n39566 = pi18 ? n37 : n39565;
  assign n39567 = pi17 ? n37 : n39566;
  assign n39568 = pi16 ? n38032 : n39567;
  assign n39569 = pi15 ? n39564 : n39568;
  assign n39570 = pi14 ? n39556 : n39569;
  assign n39571 = pi13 ? n39541 : n39570;
  assign n39572 = pi16 ? n36227 : n39098;
  assign n39573 = pi16 ? n36216 : n39102;
  assign n39574 = pi15 ? n39572 : n39573;
  assign n39575 = pi21 ? n30867 : n30843;
  assign n39576 = pi20 ? n20563 : n39575;
  assign n39577 = pi19 ? n20563 : n39576;
  assign n39578 = pi18 ? n31315 : n39577;
  assign n39579 = pi17 ? n32 : n39578;
  assign n39580 = pi19 ? n37 : n12515;
  assign n39581 = pi18 ? n37 : n39580;
  assign n39582 = pi17 ? n37 : n39581;
  assign n39583 = pi16 ? n39579 : n39582;
  assign n39584 = pi20 ? n31925 : n30096;
  assign n39585 = pi19 ? n20563 : n39584;
  assign n39586 = pi18 ? n31315 : n39585;
  assign n39587 = pi17 ? n32 : n39586;
  assign n39588 = pi22 ? n316 : n759;
  assign n39589 = pi21 ? n39588 : n32;
  assign n39590 = pi20 ? n39589 : n32;
  assign n39591 = pi19 ? n37 : n39590;
  assign n39592 = pi18 ? n37 : n39591;
  assign n39593 = pi17 ? n37 : n39592;
  assign n39594 = pi16 ? n39587 : n39593;
  assign n39595 = pi15 ? n39583 : n39594;
  assign n39596 = pi14 ? n39574 : n39595;
  assign n39597 = pi16 ? n35220 : n39116;
  assign n39598 = pi18 ? n15541 : n99;
  assign n39599 = pi19 ? n13371 : n5668;
  assign n39600 = pi18 ? n99 : n39599;
  assign n39601 = pi17 ? n39598 : n39600;
  assign n39602 = pi16 ? n36235 : n39601;
  assign n39603 = pi15 ? n39597 : n39602;
  assign n39604 = pi20 ? n31913 : n36250;
  assign n39605 = pi19 ? n20563 : n39604;
  assign n39606 = pi18 ? n31315 : n39605;
  assign n39607 = pi17 ? n32 : n39606;
  assign n39608 = pi20 ? n2243 : n15263;
  assign n39609 = pi19 ? n39608 : n2243;
  assign n39610 = pi20 ? n25399 : n32;
  assign n39611 = pi19 ? n157 : n39610;
  assign n39612 = pi18 ? n39609 : n39611;
  assign n39613 = pi17 ? n34298 : n39612;
  assign n39614 = pi16 ? n39607 : n39613;
  assign n39615 = pi19 ? n23645 : n15543;
  assign n39616 = pi18 ? n39615 : n99;
  assign n39617 = pi19 ? n19134 : n16307;
  assign n39618 = pi18 ? n39617 : n39138;
  assign n39619 = pi17 ? n39616 : n39618;
  assign n39620 = pi16 ? n34306 : n39619;
  assign n39621 = pi15 ? n39614 : n39620;
  assign n39622 = pi14 ? n39603 : n39621;
  assign n39623 = pi13 ? n39596 : n39622;
  assign n39624 = pi12 ? n39571 : n39623;
  assign n39625 = pi11 ? n39514 : n39624;
  assign n39626 = pi19 ? n20563 : n31914;
  assign n39627 = pi18 ? n31315 : n39626;
  assign n39628 = pi17 ? n32 : n39627;
  assign n39629 = pi20 ? n99 : n2973;
  assign n39630 = pi19 ? n21611 : n39629;
  assign n39631 = pi19 ? n29428 : n29191;
  assign n39632 = pi18 ? n39630 : n39631;
  assign n39633 = pi20 ? n2976 : n157;
  assign n39634 = pi21 ? n218 : n157;
  assign n39635 = pi20 ? n157 : n39634;
  assign n39636 = pi19 ? n39633 : n39635;
  assign n39637 = pi18 ? n39636 : n39138;
  assign n39638 = pi17 ? n39632 : n39637;
  assign n39639 = pi16 ? n39628 : n39638;
  assign n39640 = pi21 ? n36516 : n181;
  assign n39641 = pi20 ? n20563 : n39640;
  assign n39642 = pi19 ? n20563 : n39641;
  assign n39643 = pi18 ? n31315 : n39642;
  assign n39644 = pi17 ? n32 : n39643;
  assign n39645 = pi19 ? n25381 : n99;
  assign n39646 = pi18 ? n39645 : n99;
  assign n39647 = pi19 ? n17367 : n5668;
  assign n39648 = pi18 ? n14286 : n39647;
  assign n39649 = pi17 ? n39646 : n39648;
  assign n39650 = pi16 ? n39644 : n39649;
  assign n39651 = pi15 ? n39639 : n39650;
  assign n39652 = pi19 ? n26431 : n39400;
  assign n39653 = pi18 ? n39652 : n99;
  assign n39654 = pi21 ? n1027 : n99;
  assign n39655 = pi20 ? n39654 : n99;
  assign n39656 = pi19 ? n27596 : n39655;
  assign n39657 = pi20 ? n9181 : n2383;
  assign n39658 = pi19 ? n39657 : n5668;
  assign n39659 = pi18 ? n39656 : n39658;
  assign n39660 = pi17 ? n39653 : n39659;
  assign n39661 = pi16 ? n34319 : n39660;
  assign n39662 = pi18 ? n37 : n14842;
  assign n39663 = pi20 ? n19208 : n316;
  assign n39664 = pi19 ? n39663 : n5668;
  assign n39665 = pi18 ? n99 : n39664;
  assign n39666 = pi17 ? n39662 : n39665;
  assign n39667 = pi16 ? n34889 : n39666;
  assign n39668 = pi15 ? n39661 : n39667;
  assign n39669 = pi14 ? n39651 : n39668;
  assign n39670 = pi20 ? n35316 : n14844;
  assign n39671 = pi19 ? n20563 : n39670;
  assign n39672 = pi18 ? n31315 : n39671;
  assign n39673 = pi17 ? n32 : n39672;
  assign n39674 = pi20 ? n99 : n3871;
  assign n39675 = pi19 ? n99 : n39674;
  assign n39676 = pi21 ? n181 : n112;
  assign n39677 = pi20 ? n39676 : n2181;
  assign n39678 = pi19 ? n39677 : n2191;
  assign n39679 = pi18 ? n39675 : n39678;
  assign n39680 = pi22 ? n99 : n22428;
  assign n39681 = pi21 ? n39680 : n99;
  assign n39682 = pi20 ? n99 : n39681;
  assign n39683 = pi20 ? n4619 : n3888;
  assign n39684 = pi19 ? n39682 : n39683;
  assign n39685 = pi21 ? n3759 : n20977;
  assign n39686 = pi20 ? n39685 : n316;
  assign n39687 = pi19 ? n39686 : n5668;
  assign n39688 = pi18 ? n39684 : n39687;
  assign n39689 = pi17 ? n39679 : n39688;
  assign n39690 = pi16 ? n39673 : n39689;
  assign n39691 = pi21 ? n36516 : n99;
  assign n39692 = pi20 ? n38754 : n39691;
  assign n39693 = pi19 ? n20563 : n39692;
  assign n39694 = pi18 ? n31315 : n39693;
  assign n39695 = pi17 ? n32 : n39694;
  assign n39696 = pi18 ? n37 : n28257;
  assign n39697 = pi20 ? n20093 : n316;
  assign n39698 = pi19 ? n39697 : n4009;
  assign n39699 = pi18 ? n139 : n39698;
  assign n39700 = pi17 ? n39696 : n39699;
  assign n39701 = pi16 ? n39695 : n39700;
  assign n39702 = pi15 ? n39690 : n39701;
  assign n39703 = pi21 ? n31924 : n39182;
  assign n39704 = pi20 ? n39703 : n37;
  assign n39705 = pi19 ? n20563 : n39704;
  assign n39706 = pi18 ? n31315 : n39705;
  assign n39707 = pi17 ? n32 : n39706;
  assign n39708 = pi19 ? n15002 : n28290;
  assign n39709 = pi18 ? n39708 : n28257;
  assign n39710 = pi21 ? n1793 : n916;
  assign n39711 = pi20 ? n39710 : n5199;
  assign n39712 = pi23 ? n204 : n20004;
  assign n39713 = pi22 ? n39712 : n32;
  assign n39714 = pi21 ? n39713 : n32;
  assign n39715 = pi20 ? n39714 : n32;
  assign n39716 = pi19 ? n39711 : n39715;
  assign n39717 = pi18 ? n139 : n39716;
  assign n39718 = pi17 ? n39709 : n39717;
  assign n39719 = pi16 ? n39707 : n39718;
  assign n39720 = pi18 ? n31315 : n33847;
  assign n39721 = pi17 ? n32 : n39720;
  assign n39722 = pi19 ? n3097 : n139;
  assign n39723 = pi18 ? n37 : n39722;
  assign n39724 = pi20 ? n39710 : n204;
  assign n39725 = pi19 ? n39724 : n2567;
  assign n39726 = pi18 ? n139 : n39725;
  assign n39727 = pi17 ? n39723 : n39726;
  assign n39728 = pi16 ? n39721 : n39727;
  assign n39729 = pi15 ? n39719 : n39728;
  assign n39730 = pi14 ? n39702 : n39729;
  assign n39731 = pi13 ? n39669 : n39730;
  assign n39732 = pi17 ? n11568 : n39726;
  assign n39733 = pi16 ? n39106 : n39732;
  assign n39734 = pi20 ? n997 : n942;
  assign n39735 = pi19 ? n39734 : n139;
  assign n39736 = pi18 ? n37 : n39735;
  assign n39737 = pi19 ? n139 : n7486;
  assign n39738 = pi19 ? n26742 : n2567;
  assign n39739 = pi18 ? n39737 : n39738;
  assign n39740 = pi17 ? n39736 : n39739;
  assign n39741 = pi16 ? n39106 : n39740;
  assign n39742 = pi15 ? n39733 : n39741;
  assign n39743 = pi18 ? n31938 : n32288;
  assign n39744 = pi17 ? n32 : n39743;
  assign n39745 = pi20 ? n1003 : n3083;
  assign n39746 = pi19 ? n39745 : n13168;
  assign n39747 = pi18 ? n39746 : n39735;
  assign n39748 = pi19 ? n26742 : n2580;
  assign n39749 = pi18 ? n139 : n39748;
  assign n39750 = pi17 ? n39747 : n39749;
  assign n39751 = pi16 ? n39744 : n39750;
  assign n39752 = pi20 ? n942 : n820;
  assign n39753 = pi19 ? n31370 : n39752;
  assign n39754 = pi18 ? n37 : n39753;
  assign n39755 = pi20 ? n1003 : n941;
  assign n39756 = pi20 ? n992 : n2318;
  assign n39757 = pi19 ? n39755 : n39756;
  assign n39758 = pi20 ? n1016 : n11809;
  assign n39759 = pi19 ? n39758 : n2639;
  assign n39760 = pi18 ? n39757 : n39759;
  assign n39761 = pi17 ? n39754 : n39760;
  assign n39762 = pi16 ? n34319 : n39761;
  assign n39763 = pi15 ? n39751 : n39762;
  assign n39764 = pi14 ? n39742 : n39763;
  assign n39765 = pi18 ? n37 : n641;
  assign n39766 = pi20 ? n6358 : n7980;
  assign n39767 = pi19 ? n22046 : n39766;
  assign n39768 = pi19 ? n13535 : n2639;
  assign n39769 = pi18 ? n39767 : n39768;
  assign n39770 = pi17 ? n39765 : n39769;
  assign n39771 = pi16 ? n34889 : n39770;
  assign n39772 = pi20 ? n37 : n26846;
  assign n39773 = pi19 ? n37 : n39772;
  assign n39774 = pi20 ? n13527 : n25965;
  assign n39775 = pi19 ? n39774 : n2654;
  assign n39776 = pi18 ? n39773 : n39775;
  assign n39777 = pi17 ? n37 : n39776;
  assign n39778 = pi16 ? n34306 : n39777;
  assign n39779 = pi15 ? n39771 : n39778;
  assign n39780 = pi19 ? n31814 : n7706;
  assign n39781 = pi19 ? n37692 : n2654;
  assign n39782 = pi18 ? n39780 : n39781;
  assign n39783 = pi17 ? n37 : n39782;
  assign n39784 = pi16 ? n34889 : n39783;
  assign n39785 = pi19 ? n37692 : n35482;
  assign n39786 = pi18 ? n7707 : n39785;
  assign n39787 = pi17 ? n37 : n39786;
  assign n39788 = pi16 ? n34328 : n39787;
  assign n39789 = pi15 ? n39784 : n39788;
  assign n39790 = pi14 ? n39779 : n39789;
  assign n39791 = pi13 ? n39764 : n39790;
  assign n39792 = pi12 ? n39731 : n39791;
  assign n39793 = pi22 ? n233 : n38877;
  assign n39794 = pi21 ? n233 : n39793;
  assign n39795 = pi20 ? n233 : n39794;
  assign n39796 = pi19 ? n39795 : n32;
  assign n39797 = pi18 ? n37 : n39796;
  assign n39798 = pi17 ? n37 : n39797;
  assign n39799 = pi16 ? n34889 : n39798;
  assign n39800 = pi22 ? n36029 : n30868;
  assign n39801 = pi22 ? n30868 : n20563;
  assign n39802 = pi21 ? n39800 : n39801;
  assign n39803 = pi20 ? n32 : n39802;
  assign n39804 = pi19 ? n32 : n39803;
  assign n39805 = pi21 ? n30868 : n36489;
  assign n39806 = pi20 ? n39805 : n39801;
  assign n39807 = pi19 ? n39806 : n37;
  assign n39808 = pi18 ? n39804 : n39807;
  assign n39809 = pi17 ? n32 : n39808;
  assign n39810 = pi20 ? n638 : n13273;
  assign n39811 = pi19 ? n644 : n39810;
  assign n39812 = pi20 ? n1944 : n335;
  assign n39813 = pi19 ? n335 : n39812;
  assign n39814 = pi18 ? n39811 : n39813;
  assign n39815 = pi22 ? n233 : n19696;
  assign n39816 = pi21 ? n6376 : n39815;
  assign n39817 = pi20 ? n335 : n39816;
  assign n39818 = pi19 ? n39817 : n32;
  assign n39819 = pi18 ? n335 : n39818;
  assign n39820 = pi17 ? n39814 : n39819;
  assign n39821 = pi16 ? n39809 : n39820;
  assign n39822 = pi15 ? n39799 : n39821;
  assign n39823 = pi19 ? n20563 : n7676;
  assign n39824 = pi18 ? n31938 : n39823;
  assign n39825 = pi17 ? n32 : n39824;
  assign n39826 = pi19 ? n644 : n22046;
  assign n39827 = pi18 ? n39826 : n38761;
  assign n39828 = pi20 ? n233 : n23093;
  assign n39829 = pi19 ? n39828 : n32;
  assign n39830 = pi18 ? n335 : n39829;
  assign n39831 = pi17 ? n39827 : n39830;
  assign n39832 = pi16 ? n39825 : n39831;
  assign n39833 = pi20 ? n30096 : n5778;
  assign n39834 = pi19 ? n20563 : n39833;
  assign n39835 = pi18 ? n31315 : n39834;
  assign n39836 = pi17 ? n32 : n39835;
  assign n39837 = pi20 ? n13527 : n23093;
  assign n39838 = pi19 ? n39837 : n32;
  assign n39839 = pi18 ? n335 : n39838;
  assign n39840 = pi17 ? n335 : n39839;
  assign n39841 = pi16 ? n39836 : n39840;
  assign n39842 = pi15 ? n39832 : n39841;
  assign n39843 = pi14 ? n39822 : n39842;
  assign n39844 = pi20 ? n30096 : n605;
  assign n39845 = pi19 ? n20563 : n39844;
  assign n39846 = pi18 ? n31315 : n39845;
  assign n39847 = pi17 ? n32 : n39846;
  assign n39848 = pi20 ? n335 : n23093;
  assign n39849 = pi19 ? n39848 : n32;
  assign n39850 = pi18 ? n335 : n39849;
  assign n39851 = pi17 ? n335 : n39850;
  assign n39852 = pi16 ? n39847 : n39851;
  assign n39853 = pi20 ? n37 : n7331;
  assign n39854 = pi19 ? n20563 : n39853;
  assign n39855 = pi18 ? n31315 : n39854;
  assign n39856 = pi17 ? n32 : n39855;
  assign n39857 = pi21 ? n9657 : n5012;
  assign n39858 = pi20 ? n39857 : n10480;
  assign n39859 = pi20 ? n10481 : n10486;
  assign n39860 = pi19 ? n39858 : n39859;
  assign n39861 = pi20 ? n24865 : n27520;
  assign n39862 = pi21 ? n5015 : n9666;
  assign n39863 = pi20 ? n39862 : n7730;
  assign n39864 = pi19 ? n39861 : n39863;
  assign n39865 = pi18 ? n39860 : n39864;
  assign n39866 = pi20 ? n27482 : n10496;
  assign n39867 = pi20 ? n22881 : n363;
  assign n39868 = pi19 ? n39866 : n39867;
  assign n39869 = pi20 ? n2107 : n15729;
  assign n39870 = pi19 ? n39869 : n32;
  assign n39871 = pi18 ? n39868 : n39870;
  assign n39872 = pi17 ? n39865 : n39871;
  assign n39873 = pi16 ? n39856 : n39872;
  assign n39874 = pi15 ? n39852 : n39873;
  assign n39875 = pi21 ? n685 : n8486;
  assign n39876 = pi20 ? n685 : n39875;
  assign n39877 = pi19 ? n39876 : n32;
  assign n39878 = pi18 ? n38812 : n39877;
  assign n39879 = pi17 ? n37 : n39878;
  assign n39880 = pi16 ? n34889 : n39879;
  assign n39881 = pi22 ? n39174 : n2160;
  assign n39882 = pi21 ? n36489 : n39881;
  assign n39883 = pi20 ? n39882 : n99;
  assign n39884 = pi19 ? n20563 : n39883;
  assign n39885 = pi18 ? n31315 : n39884;
  assign n39886 = pi17 ? n32 : n39885;
  assign n39887 = pi19 ? n22883 : n37753;
  assign n39888 = pi18 ? n37 : n39887;
  assign n39889 = pi21 ? n685 : n3523;
  assign n39890 = pi20 ? n24220 : n39889;
  assign n39891 = pi19 ? n39890 : n32;
  assign n39892 = pi18 ? n363 : n39891;
  assign n39893 = pi17 ? n39888 : n39892;
  assign n39894 = pi16 ? n39886 : n39893;
  assign n39895 = pi15 ? n39880 : n39894;
  assign n39896 = pi14 ? n39874 : n39895;
  assign n39897 = pi13 ? n39843 : n39896;
  assign n39898 = pi21 ? n37 : n9666;
  assign n39899 = pi20 ? n27501 : n39898;
  assign n39900 = pi19 ? n38832 : n39899;
  assign n39901 = pi18 ? n37 : n39900;
  assign n39902 = pi21 ? n363 : n6401;
  assign n39903 = pi20 ? n39902 : n15173;
  assign n39904 = pi21 ? n9666 : n37;
  assign n39905 = pi20 ? n39904 : n10494;
  assign n39906 = pi19 ? n39903 : n39905;
  assign n39907 = pi18 ? n39906 : n38825;
  assign n39908 = pi17 ? n39901 : n39907;
  assign n39909 = pi16 ? n34889 : n39908;
  assign n39910 = pi21 ? n685 : n33217;
  assign n39911 = pi20 ? n2107 : n39910;
  assign n39912 = pi19 ? n39911 : n32;
  assign n39913 = pi18 ? n37 : n39912;
  assign n39914 = pi17 ? n37 : n39913;
  assign n39915 = pi16 ? n34889 : n39914;
  assign n39916 = pi15 ? n39909 : n39915;
  assign n39917 = pi19 ? n30868 : n38251;
  assign n39918 = pi18 ? n38249 : n39917;
  assign n39919 = pi17 ? n32 : n39918;
  assign n39920 = pi21 ? n3445 : n19697;
  assign n39921 = pi20 ? n685 : n39920;
  assign n39922 = pi19 ? n39921 : n32;
  assign n39923 = pi18 ? n99 : n39922;
  assign n39924 = pi17 ? n99 : n39923;
  assign n39925 = pi16 ? n39919 : n39924;
  assign n39926 = pi22 ? n30868 : n99;
  assign n39927 = pi21 ? n30868 : n39926;
  assign n39928 = pi20 ? n39927 : n99;
  assign n39929 = pi19 ? n30868 : n39928;
  assign n39930 = pi18 ? n37808 : n39929;
  assign n39931 = pi17 ? n32 : n39930;
  assign n39932 = pi22 ? n21078 : n32;
  assign n39933 = pi21 ? n3445 : n39932;
  assign n39934 = pi20 ? n7754 : n39933;
  assign n39935 = pi19 ? n39934 : n32;
  assign n39936 = pi18 ? n99 : n39935;
  assign n39937 = pi17 ? n99 : n39936;
  assign n39938 = pi16 ? n39931 : n39937;
  assign n39939 = pi15 ? n39925 : n39938;
  assign n39940 = pi14 ? n39916 : n39939;
  assign n39941 = pi20 ? n36659 : n33792;
  assign n39942 = pi20 ? n39336 : n139;
  assign n39943 = pi19 ? n39941 : n39942;
  assign n39944 = pi18 ? n37841 : n39943;
  assign n39945 = pi17 ? n32 : n39944;
  assign n39946 = pi21 ? n38878 : n20952;
  assign n39947 = pi20 ? n685 : n39946;
  assign n39948 = pi19 ? n39947 : n32;
  assign n39949 = pi18 ? n685 : n39948;
  assign n39950 = pi17 ? n38876 : n39949;
  assign n39951 = pi16 ? n39945 : n39950;
  assign n39952 = pi22 ? n33792 : n36781;
  assign n39953 = pi21 ? n33792 : n39952;
  assign n39954 = pi23 ? n139 : n36781;
  assign n39955 = pi22 ? n39954 : n363;
  assign n39956 = pi21 ? n39955 : n363;
  assign n39957 = pi20 ? n39953 : n39956;
  assign n39958 = pi19 ? n38885 : n39957;
  assign n39959 = pi18 ? n37841 : n39958;
  assign n39960 = pi17 ? n32 : n39959;
  assign n39961 = pi20 ? n26890 : n29741;
  assign n39962 = pi19 ? n39961 : n685;
  assign n39963 = pi18 ? n363 : n39962;
  assign n39964 = pi18 ? n685 : n33199;
  assign n39965 = pi17 ? n39963 : n39964;
  assign n39966 = pi16 ? n39960 : n39965;
  assign n39967 = pi15 ? n39951 : n39966;
  assign n39968 = pi22 ? n37274 : n36798;
  assign n39969 = pi21 ? n39968 : n36798;
  assign n39970 = pi20 ? n32 : n39969;
  assign n39971 = pi19 ? n32 : n39970;
  assign n39972 = pi22 ? n36781 : n36798;
  assign n39973 = pi21 ? n36798 : n39972;
  assign n39974 = pi20 ? n38900 : n39973;
  assign n39975 = pi21 ? n36659 : n36781;
  assign n39976 = pi23 ? n335 : n36781;
  assign n39977 = pi22 ? n39976 : n335;
  assign n39978 = pi22 ? n157 : n3935;
  assign n39979 = pi21 ? n39977 : n39978;
  assign n39980 = pi20 ? n39975 : n39979;
  assign n39981 = pi19 ? n39974 : n39980;
  assign n39982 = pi18 ? n39971 : n39981;
  assign n39983 = pi17 ? n32 : n39982;
  assign n39984 = pi20 ? n6461 : n27551;
  assign n39985 = pi19 ? n37885 : n39984;
  assign n39986 = pi18 ? n157 : n39985;
  assign n39987 = pi20 ? n36843 : n685;
  assign n39988 = pi19 ? n37888 : n39987;
  assign n39989 = pi22 ? n7780 : n685;
  assign n39990 = pi21 ? n39989 : n685;
  assign n39991 = pi20 ? n39990 : n9456;
  assign n39992 = pi19 ? n39991 : n32;
  assign n39993 = pi18 ? n39988 : n39992;
  assign n39994 = pi17 ? n39986 : n39993;
  assign n39995 = pi16 ? n39983 : n39994;
  assign n39996 = pi23 ? n37273 : n36781;
  assign n39997 = pi22 ? n39996 : n36781;
  assign n39998 = pi21 ? n39997 : n36798;
  assign n39999 = pi20 ? n32 : n39998;
  assign n40000 = pi19 ? n32 : n39999;
  assign n40001 = pi20 ? n38923 : n36781;
  assign n40002 = pi22 ? n36781 : n38284;
  assign n40003 = pi21 ? n40002 : n36781;
  assign n40004 = pi23 ? n363 : n36781;
  assign n40005 = pi22 ? n40004 : n157;
  assign n40006 = pi21 ? n40005 : n157;
  assign n40007 = pi20 ? n40003 : n40006;
  assign n40008 = pi19 ? n40001 : n40007;
  assign n40009 = pi18 ? n40000 : n40008;
  assign n40010 = pi17 ? n32 : n40009;
  assign n40011 = pi20 ? n34537 : n5667;
  assign n40012 = pi19 ? n40011 : n32;
  assign n40013 = pi18 ? n157 : n40012;
  assign n40014 = pi17 ? n157 : n40013;
  assign n40015 = pi16 ? n40010 : n40014;
  assign n40016 = pi15 ? n39995 : n40015;
  assign n40017 = pi14 ? n39967 : n40016;
  assign n40018 = pi13 ? n39940 : n40017;
  assign n40019 = pi12 ? n39897 : n40018;
  assign n40020 = pi11 ? n39792 : n40019;
  assign n40021 = pi10 ? n39625 : n40020;
  assign n40022 = pi09 ? n39414 : n40021;
  assign n40023 = pi19 ? n28158 : n20563;
  assign n40024 = pi18 ? n32 : n40023;
  assign n40025 = pi17 ? n32 : n40024;
  assign n40026 = pi16 ? n40025 : n39384;
  assign n40027 = pi15 ? n32 : n40026;
  assign n40028 = pi19 ? n32933 : n39387;
  assign n40029 = pi18 ? n20563 : n40028;
  assign n40030 = pi17 ? n40029 : n39391;
  assign n40031 = pi16 ? n39375 : n40030;
  assign n40032 = pi18 ? n20563 : n39401;
  assign n40033 = pi17 ? n40032 : n39406;
  assign n40034 = pi16 ? n38950 : n40033;
  assign n40035 = pi15 ? n40031 : n40034;
  assign n40036 = pi14 ? n40027 : n40035;
  assign n40037 = pi13 ? n32 : n40036;
  assign n40038 = pi12 ? n32 : n40037;
  assign n40039 = pi11 ? n32 : n40038;
  assign n40040 = pi10 ? n32 : n40039;
  assign n40041 = pi18 ? n34247 : n37;
  assign n40042 = pi17 ? n40041 : n39422;
  assign n40043 = pi16 ? n38959 : n40042;
  assign n40044 = pi20 ? n38376 : n20563;
  assign n40045 = pi19 ? n40044 : n20563;
  assign n40046 = pi18 ? n32 : n40045;
  assign n40047 = pi17 ? n32 : n40046;
  assign n40048 = pi18 ? n34865 : n37;
  assign n40049 = pi17 ? n40048 : n39428;
  assign n40050 = pi16 ? n40047 : n40049;
  assign n40051 = pi15 ? n40043 : n40050;
  assign n40052 = pi17 ? n39415 : n39437;
  assign n40053 = pi16 ? n37930 : n40052;
  assign n40054 = pi21 ? n32 : n39394;
  assign n40055 = pi20 ? n32 : n40054;
  assign n40056 = pi19 ? n32 : n40055;
  assign n40057 = pi18 ? n40056 : n20563;
  assign n40058 = pi17 ? n32 : n40057;
  assign n40059 = pi16 ? n40058 : n39443;
  assign n40060 = pi15 ? n40053 : n40059;
  assign n40061 = pi14 ? n40051 : n40060;
  assign n40062 = pi18 ? n33828 : n37;
  assign n40063 = pi19 ? n9795 : n11560;
  assign n40064 = pi18 ? n39450 : n40063;
  assign n40065 = pi17 ? n40062 : n40064;
  assign n40066 = pi16 ? n37959 : n40065;
  assign n40067 = pi19 ? n20563 : n33923;
  assign n40068 = pi18 ? n40067 : n37;
  assign n40069 = pi19 ? n29248 : n11560;
  assign n40070 = pi18 ? n37 : n40069;
  assign n40071 = pi17 ? n40068 : n40070;
  assign n40072 = pi16 ? n39001 : n40071;
  assign n40073 = pi15 ? n40066 : n40072;
  assign n40074 = pi19 ? n20722 : n11560;
  assign n40075 = pi18 ? n37 : n40074;
  assign n40076 = pi17 ? n39448 : n40075;
  assign n40077 = pi16 ? n39001 : n40076;
  assign n40078 = pi19 ? n3110 : n11560;
  assign n40079 = pi18 ? n37 : n40078;
  assign n40080 = pi17 ? n38369 : n40079;
  assign n40081 = pi16 ? n36216 : n40080;
  assign n40082 = pi15 ? n40077 : n40081;
  assign n40083 = pi14 ? n40073 : n40082;
  assign n40084 = pi13 ? n40061 : n40083;
  assign n40085 = pi21 ? n335 : n17618;
  assign n40086 = pi20 ? n40085 : n32;
  assign n40087 = pi19 ? n13192 : n40086;
  assign n40088 = pi18 ? n37 : n40087;
  assign n40089 = pi17 ? n39481 : n40088;
  assign n40090 = pi16 ? n36216 : n40089;
  assign n40091 = pi22 ? n20317 : n32;
  assign n40092 = pi21 ? n335 : n40091;
  assign n40093 = pi20 ? n40092 : n32;
  assign n40094 = pi19 ? n7676 : n40093;
  assign n40095 = pi18 ? n37 : n40094;
  assign n40096 = pi17 ? n39481 : n40095;
  assign n40097 = pi16 ? n36216 : n40096;
  assign n40098 = pi15 ? n40090 : n40097;
  assign n40099 = pi18 ? n34891 : n37;
  assign n40100 = pi19 ? n37 : n40093;
  assign n40101 = pi18 ? n37 : n40100;
  assign n40102 = pi17 ? n40099 : n40101;
  assign n40103 = pi16 ? n36216 : n40102;
  assign n40104 = pi21 ? n335 : n5003;
  assign n40105 = pi20 ? n40104 : n32;
  assign n40106 = pi19 ? n37 : n40105;
  assign n40107 = pi18 ? n37 : n40106;
  assign n40108 = pi17 ? n39489 : n40107;
  assign n40109 = pi16 ? n36216 : n40108;
  assign n40110 = pi15 ? n40103 : n40109;
  assign n40111 = pi14 ? n40098 : n40110;
  assign n40112 = pi20 ? n27493 : n32;
  assign n40113 = pi19 ? n37 : n40112;
  assign n40114 = pi18 ? n37 : n40113;
  assign n40115 = pi17 ? n39494 : n40114;
  assign n40116 = pi16 ? n36216 : n40115;
  assign n40117 = pi17 ? n37372 : n39499;
  assign n40118 = pi16 ? n36216 : n40117;
  assign n40119 = pi15 ? n40116 : n40118;
  assign n40120 = pi18 ? n33924 : n37;
  assign n40121 = pi17 ? n40120 : n39504;
  assign n40122 = pi16 ? n36216 : n40121;
  assign n40123 = pi20 ? n31913 : n30096;
  assign n40124 = pi19 ? n40123 : n37;
  assign n40125 = pi18 ? n40124 : n37;
  assign n40126 = pi17 ? n40125 : n39508;
  assign n40127 = pi16 ? n36216 : n40126;
  assign n40128 = pi15 ? n40122 : n40127;
  assign n40129 = pi14 ? n40119 : n40128;
  assign n40130 = pi13 ? n40111 : n40129;
  assign n40131 = pi12 ? n40084 : n40130;
  assign n40132 = pi17 ? n39039 : n39520;
  assign n40133 = pi16 ? n36216 : n40132;
  assign n40134 = pi21 ? n363 : n2553;
  assign n40135 = pi20 ? n40134 : n32;
  assign n40136 = pi19 ? n37 : n40135;
  assign n40137 = pi18 ? n37 : n40136;
  assign n40138 = pi17 ? n39039 : n40137;
  assign n40139 = pi16 ? n36216 : n40138;
  assign n40140 = pi15 ? n40133 : n40139;
  assign n40141 = pi18 ? n35318 : n37;
  assign n40142 = pi21 ? n2721 : n2678;
  assign n40143 = pi20 ? n40142 : n32;
  assign n40144 = pi19 ? n37 : n40143;
  assign n40145 = pi18 ? n37 : n40144;
  assign n40146 = pi17 ? n40141 : n40145;
  assign n40147 = pi16 ? n36216 : n40146;
  assign n40148 = pi21 ? n31294 : n31200;
  assign n40149 = pi20 ? n40148 : n37;
  assign n40150 = pi19 ? n40149 : n37;
  assign n40151 = pi18 ? n40150 : n37;
  assign n40152 = pi17 ? n40151 : n39537;
  assign n40153 = pi16 ? n36216 : n40152;
  assign n40154 = pi15 ? n40147 : n40153;
  assign n40155 = pi14 ? n40140 : n40154;
  assign n40156 = pi21 ? n5070 : n2700;
  assign n40157 = pi20 ? n40156 : n32;
  assign n40158 = pi19 ? n7731 : n40157;
  assign n40159 = pi18 ? n37 : n40158;
  assign n40160 = pi17 ? n36907 : n40159;
  assign n40161 = pi16 ? n36216 : n40160;
  assign n40162 = pi21 ? n5062 : n2700;
  assign n40163 = pi20 ? n40162 : n32;
  assign n40164 = pi19 ? n37 : n40163;
  assign n40165 = pi18 ? n37 : n40164;
  assign n40166 = pi17 ? n39529 : n40165;
  assign n40167 = pi16 ? n36216 : n40166;
  assign n40168 = pi15 ? n40161 : n40167;
  assign n40169 = pi21 ? n11178 : n2700;
  assign n40170 = pi20 ? n40169 : n32;
  assign n40171 = pi19 ? n37 : n40170;
  assign n40172 = pi18 ? n37 : n40171;
  assign n40173 = pi17 ? n36210 : n40172;
  assign n40174 = pi16 ? n36216 : n40173;
  assign n40175 = pi18 ? n31315 : n34247;
  assign n40176 = pi17 ? n32 : n40175;
  assign n40177 = pi17 ? n36919 : n39531;
  assign n40178 = pi16 ? n40176 : n40177;
  assign n40179 = pi15 ? n40174 : n40178;
  assign n40180 = pi14 ? n40168 : n40179;
  assign n40181 = pi13 ? n40155 : n40180;
  assign n40182 = pi19 ? n37 : n7408;
  assign n40183 = pi18 ? n37 : n40182;
  assign n40184 = pi17 ? n39534 : n40183;
  assign n40185 = pi16 ? n36216 : n40184;
  assign n40186 = pi19 ? n37 : n13794;
  assign n40187 = pi18 ? n37 : n40186;
  assign n40188 = pi17 ? n37 : n40187;
  assign n40189 = pi16 ? n36216 : n40188;
  assign n40190 = pi15 ? n40185 : n40189;
  assign n40191 = pi19 ? n20563 : n34920;
  assign n40192 = pi18 ? n31315 : n40191;
  assign n40193 = pi17 ? n32 : n40192;
  assign n40194 = pi19 ? n37 : n12926;
  assign n40195 = pi18 ? n37 : n40194;
  assign n40196 = pi17 ? n37 : n40195;
  assign n40197 = pi16 ? n40193 : n40196;
  assign n40198 = pi20 ? n20563 : n40148;
  assign n40199 = pi19 ? n20563 : n40198;
  assign n40200 = pi18 ? n31315 : n40199;
  assign n40201 = pi17 ? n32 : n40200;
  assign n40202 = pi22 ? n316 : n1475;
  assign n40203 = pi21 ? n40202 : n32;
  assign n40204 = pi20 ? n40203 : n32;
  assign n40205 = pi19 ? n37 : n40204;
  assign n40206 = pi18 ? n37 : n40205;
  assign n40207 = pi17 ? n37 : n40206;
  assign n40208 = pi16 ? n40201 : n40207;
  assign n40209 = pi15 ? n40197 : n40208;
  assign n40210 = pi14 ? n40190 : n40209;
  assign n40211 = pi19 ? n37 : n6936;
  assign n40212 = pi18 ? n37 : n40211;
  assign n40213 = pi17 ? n37 : n40212;
  assign n40214 = pi16 ? n40201 : n40213;
  assign n40215 = pi22 ? n316 : n6146;
  assign n40216 = pi21 ? n40215 : n32;
  assign n40217 = pi20 ? n40216 : n32;
  assign n40218 = pi19 ? n13371 : n40217;
  assign n40219 = pi18 ? n99 : n40218;
  assign n40220 = pi17 ? n39598 : n40219;
  assign n40221 = pi16 ? n36933 : n40220;
  assign n40222 = pi15 ? n40214 : n40221;
  assign n40223 = pi20 ? n25822 : n32;
  assign n40224 = pi19 ? n157 : n40223;
  assign n40225 = pi18 ? n39609 : n40224;
  assign n40226 = pi17 ? n34298 : n40225;
  assign n40227 = pi16 ? n36950 : n40226;
  assign n40228 = pi19 ? n20563 : n36897;
  assign n40229 = pi18 ? n31315 : n40228;
  assign n40230 = pi17 ? n32 : n40229;
  assign n40231 = pi19 ? n157 : n16507;
  assign n40232 = pi18 ? n39617 : n40231;
  assign n40233 = pi17 ? n39616 : n40232;
  assign n40234 = pi16 ? n40230 : n40233;
  assign n40235 = pi15 ? n40227 : n40234;
  assign n40236 = pi14 ? n40222 : n40235;
  assign n40237 = pi13 ? n40210 : n40236;
  assign n40238 = pi12 ? n40181 : n40237;
  assign n40239 = pi11 ? n40131 : n40238;
  assign n40240 = pi20 ? n5420 : n2747;
  assign n40241 = pi19 ? n29428 : n40240;
  assign n40242 = pi18 ? n39630 : n40241;
  assign n40243 = pi20 ? n2184 : n157;
  assign n40244 = pi19 ? n40243 : n39635;
  assign n40245 = pi19 ? n157 : n14328;
  assign n40246 = pi18 ? n40244 : n40245;
  assign n40247 = pi17 ? n40242 : n40246;
  assign n40248 = pi16 ? n35801 : n40247;
  assign n40249 = pi22 ? n30868 : n39190;
  assign n40250 = pi22 ? n39174 : n99;
  assign n40251 = pi21 ? n40249 : n40250;
  assign n40252 = pi20 ? n20563 : n40251;
  assign n40253 = pi19 ? n20563 : n40252;
  assign n40254 = pi18 ? n31315 : n40253;
  assign n40255 = pi17 ? n32 : n40254;
  assign n40256 = pi17 ? n39598 : n39648;
  assign n40257 = pi16 ? n40255 : n40256;
  assign n40258 = pi15 ? n40248 : n40257;
  assign n40259 = pi16 ? n35814 : n39660;
  assign n40260 = pi16 ? n40230 : n39666;
  assign n40261 = pi15 ? n40259 : n40260;
  assign n40262 = pi14 ? n40258 : n40261;
  assign n40263 = pi21 ? n39175 : n99;
  assign n40264 = pi20 ? n31925 : n40263;
  assign n40265 = pi19 ? n20563 : n40264;
  assign n40266 = pi18 ? n31315 : n40265;
  assign n40267 = pi17 ? n32 : n40266;
  assign n40268 = pi20 ? n99 : n3033;
  assign n40269 = pi19 ? n99 : n40268;
  assign n40270 = pi20 ? n21638 : n2181;
  assign n40271 = pi19 ? n40270 : n2191;
  assign n40272 = pi18 ? n40269 : n40271;
  assign n40273 = pi22 ? n22428 : n456;
  assign n40274 = pi22 ? n99 : n455;
  assign n40275 = pi21 ? n40273 : n40274;
  assign n40276 = pi20 ? n40275 : n16614;
  assign n40277 = pi19 ? n39682 : n40276;
  assign n40278 = pi18 ? n40277 : n39687;
  assign n40279 = pi17 ? n40272 : n40278;
  assign n40280 = pi16 ? n40267 : n40279;
  assign n40281 = pi22 ? n30868 : n39174;
  assign n40282 = pi21 ? n40281 : n99;
  assign n40283 = pi20 ? n38754 : n40282;
  assign n40284 = pi19 ? n20563 : n40283;
  assign n40285 = pi18 ? n31315 : n40284;
  assign n40286 = pi17 ? n32 : n40285;
  assign n40287 = pi16 ? n40286 : n39700;
  assign n40288 = pi15 ? n40280 : n40287;
  assign n40289 = pi21 ? n20563 : n39182;
  assign n40290 = pi20 ? n40289 : n37;
  assign n40291 = pi19 ? n20563 : n40290;
  assign n40292 = pi18 ? n31315 : n40291;
  assign n40293 = pi17 ? n32 : n40292;
  assign n40294 = pi19 ? n39711 : n3978;
  assign n40295 = pi18 ? n139 : n40294;
  assign n40296 = pi17 ? n39709 : n40295;
  assign n40297 = pi16 ? n40293 : n40296;
  assign n40298 = pi19 ? n39724 : n3321;
  assign n40299 = pi18 ? n139 : n40298;
  assign n40300 = pi17 ? n39723 : n40299;
  assign n40301 = pi16 ? n39628 : n40300;
  assign n40302 = pi15 ? n40297 : n40301;
  assign n40303 = pi14 ? n40288 : n40302;
  assign n40304 = pi13 ? n40262 : n40303;
  assign n40305 = pi19 ? n39724 : n36426;
  assign n40306 = pi18 ? n139 : n40305;
  assign n40307 = pi17 ? n11568 : n40306;
  assign n40308 = pi16 ? n39628 : n40307;
  assign n40309 = pi19 ? n26742 : n36426;
  assign n40310 = pi18 ? n39737 : n40309;
  assign n40311 = pi17 ? n39736 : n40310;
  assign n40312 = pi16 ? n39628 : n40311;
  assign n40313 = pi15 ? n40308 : n40312;
  assign n40314 = pi19 ? n20563 : n36362;
  assign n40315 = pi18 ? n31315 : n40314;
  assign n40316 = pi17 ? n32 : n40315;
  assign n40317 = pi16 ? n40316 : n39750;
  assign n40318 = pi16 ? n40316 : n39761;
  assign n40319 = pi15 ? n40317 : n40318;
  assign n40320 = pi14 ? n40313 : n40319;
  assign n40321 = pi16 ? n40316 : n39770;
  assign n40322 = pi16 ? n40230 : n39777;
  assign n40323 = pi15 ? n40321 : n40322;
  assign n40324 = pi18 ? n31938 : n35812;
  assign n40325 = pi17 ? n32 : n40324;
  assign n40326 = pi16 ? n40325 : n39783;
  assign n40327 = pi19 ? n20563 : n40149;
  assign n40328 = pi18 ? n31315 : n40327;
  assign n40329 = pi17 ? n32 : n40328;
  assign n40330 = pi19 ? n37692 : n1823;
  assign n40331 = pi18 ? n7707 : n40330;
  assign n40332 = pi17 ? n37 : n40331;
  assign n40333 = pi16 ? n40329 : n40332;
  assign n40334 = pi15 ? n40326 : n40333;
  assign n40335 = pi14 ? n40323 : n40334;
  assign n40336 = pi13 ? n40320 : n40335;
  assign n40337 = pi12 ? n40304 : n40336;
  assign n40338 = pi19 ? n38736 : n32;
  assign n40339 = pi18 ? n37 : n40338;
  assign n40340 = pi17 ? n37 : n40339;
  assign n40341 = pi16 ? n34889 : n40340;
  assign n40342 = pi23 ? n20564 : n30868;
  assign n40343 = pi22 ? n40342 : n30868;
  assign n40344 = pi21 ? n40343 : n39801;
  assign n40345 = pi20 ? n32 : n40344;
  assign n40346 = pi19 ? n32 : n40345;
  assign n40347 = pi20 ? n36885 : n37;
  assign n40348 = pi19 ? n39806 : n40347;
  assign n40349 = pi18 ? n40346 : n40348;
  assign n40350 = pi17 ? n32 : n40349;
  assign n40351 = pi21 ? n6376 : n15698;
  assign n40352 = pi20 ? n335 : n40351;
  assign n40353 = pi19 ? n40352 : n32;
  assign n40354 = pi18 ? n335 : n40353;
  assign n40355 = pi17 ? n39814 : n40354;
  assign n40356 = pi16 ? n40350 : n40355;
  assign n40357 = pi15 ? n40341 : n40356;
  assign n40358 = pi21 ? n30867 : n31200;
  assign n40359 = pi20 ? n40358 : n649;
  assign n40360 = pi19 ? n20563 : n40359;
  assign n40361 = pi18 ? n31315 : n40360;
  assign n40362 = pi17 ? n32 : n40361;
  assign n40363 = pi16 ? n40362 : n39831;
  assign n40364 = pi20 ? n40148 : n649;
  assign n40365 = pi19 ? n20563 : n40364;
  assign n40366 = pi18 ? n31315 : n40365;
  assign n40367 = pi17 ? n32 : n40366;
  assign n40368 = pi16 ? n40367 : n39840;
  assign n40369 = pi15 ? n40363 : n40368;
  assign n40370 = pi14 ? n40357 : n40369;
  assign n40371 = pi20 ? n40148 : n605;
  assign n40372 = pi19 ? n20563 : n40371;
  assign n40373 = pi18 ? n31315 : n40372;
  assign n40374 = pi17 ? n32 : n40373;
  assign n40375 = pi16 ? n40374 : n39851;
  assign n40376 = pi19 ? n20563 : n25354;
  assign n40377 = pi18 ? n31315 : n40376;
  assign n40378 = pi17 ? n32 : n40377;
  assign n40379 = pi16 ? n40378 : n39872;
  assign n40380 = pi15 ? n40375 : n40379;
  assign n40381 = pi20 ? n36929 : n37;
  assign n40382 = pi19 ? n20563 : n40381;
  assign n40383 = pi18 ? n31315 : n40382;
  assign n40384 = pi17 ? n32 : n40383;
  assign n40385 = pi16 ? n40384 : n39879;
  assign n40386 = pi23 ? n30868 : n20563;
  assign n40387 = pi23 ? n99 : n20563;
  assign n40388 = pi22 ? n40386 : n40387;
  assign n40389 = pi21 ? n36489 : n40388;
  assign n40390 = pi20 ? n40389 : n99;
  assign n40391 = pi19 ? n20563 : n40390;
  assign n40392 = pi18 ? n31315 : n40391;
  assign n40393 = pi17 ? n32 : n40392;
  assign n40394 = pi16 ? n40393 : n39893;
  assign n40395 = pi15 ? n40385 : n40394;
  assign n40396 = pi14 ? n40380 : n40395;
  assign n40397 = pi13 ? n40370 : n40396;
  assign n40398 = pi16 ? n40384 : n39908;
  assign n40399 = pi20 ? n2107 : n38823;
  assign n40400 = pi19 ? n40399 : n32;
  assign n40401 = pi18 ? n37 : n40400;
  assign n40402 = pi17 ? n37 : n40401;
  assign n40403 = pi16 ? n40316 : n40402;
  assign n40404 = pi15 ? n40398 : n40403;
  assign n40405 = pi21 ? n30868 : n37809;
  assign n40406 = pi20 ? n40405 : n99;
  assign n40407 = pi19 ? n30868 : n40406;
  assign n40408 = pi18 ? n37808 : n40407;
  assign n40409 = pi17 ? n32 : n40408;
  assign n40410 = pi21 ? n3445 : n882;
  assign n40411 = pi20 ? n685 : n40410;
  assign n40412 = pi19 ? n40411 : n32;
  assign n40413 = pi18 ? n99 : n40412;
  assign n40414 = pi17 ? n99 : n40413;
  assign n40415 = pi16 ? n40409 : n40414;
  assign n40416 = pi21 ? n30868 : n37810;
  assign n40417 = pi20 ? n40416 : n99;
  assign n40418 = pi19 ? n30868 : n40417;
  assign n40419 = pi18 ? n37808 : n40418;
  assign n40420 = pi17 ? n32 : n40419;
  assign n40421 = pi20 ? n7754 : n37820;
  assign n40422 = pi19 ? n40421 : n32;
  assign n40423 = pi18 ? n99 : n40422;
  assign n40424 = pi17 ? n99 : n40423;
  assign n40425 = pi16 ? n40420 : n40424;
  assign n40426 = pi15 ? n40415 : n40425;
  assign n40427 = pi14 ? n40404 : n40426;
  assign n40428 = pi23 ? n139 : n33792;
  assign n40429 = pi22 ? n40428 : n139;
  assign n40430 = pi21 ? n40429 : n139;
  assign n40431 = pi20 ? n33792 : n40430;
  assign n40432 = pi19 ? n39941 : n40431;
  assign n40433 = pi18 ? n37841 : n40432;
  assign n40434 = pi17 ? n32 : n40433;
  assign n40435 = pi21 ? n5113 : n20952;
  assign n40436 = pi20 ? n685 : n40435;
  assign n40437 = pi19 ? n40436 : n32;
  assign n40438 = pi18 ? n685 : n40437;
  assign n40439 = pi17 ? n38876 : n40438;
  assign n40440 = pi16 ? n40434 : n40439;
  assign n40441 = pi22 ? n36781 : n363;
  assign n40442 = pi21 ? n40441 : n363;
  assign n40443 = pi20 ? n39953 : n40442;
  assign n40444 = pi19 ? n38885 : n40443;
  assign n40445 = pi18 ? n37841 : n40444;
  assign n40446 = pi17 ? n32 : n40445;
  assign n40447 = pi18 ? n685 : n33716;
  assign n40448 = pi17 ? n39963 : n40447;
  assign n40449 = pi16 ? n40446 : n40448;
  assign n40450 = pi15 ? n40440 : n40449;
  assign n40451 = pi22 ? n36781 : n335;
  assign n40452 = pi21 ? n40451 : n38905;
  assign n40453 = pi20 ? n39975 : n40452;
  assign n40454 = pi19 ? n39974 : n40453;
  assign n40455 = pi18 ? n39971 : n40454;
  assign n40456 = pi17 ? n32 : n40455;
  assign n40457 = pi20 ? n39990 : n11695;
  assign n40458 = pi19 ? n40457 : n32;
  assign n40459 = pi18 ? n39988 : n40458;
  assign n40460 = pi17 ? n39986 : n40459;
  assign n40461 = pi16 ? n40456 : n40460;
  assign n40462 = pi21 ? n36784 : n36798;
  assign n40463 = pi20 ? n32 : n40462;
  assign n40464 = pi19 ? n32 : n40463;
  assign n40465 = pi22 ? n36781 : n157;
  assign n40466 = pi21 ? n40465 : n157;
  assign n40467 = pi20 ? n36781 : n40466;
  assign n40468 = pi19 ? n40001 : n40467;
  assign n40469 = pi18 ? n40464 : n40468;
  assign n40470 = pi17 ? n32 : n40469;
  assign n40471 = pi20 ? n34537 : n6935;
  assign n40472 = pi19 ? n40471 : n32;
  assign n40473 = pi18 ? n157 : n40472;
  assign n40474 = pi17 ? n157 : n40473;
  assign n40475 = pi16 ? n40470 : n40474;
  assign n40476 = pi15 ? n40461 : n40475;
  assign n40477 = pi14 ? n40450 : n40476;
  assign n40478 = pi13 ? n40427 : n40477;
  assign n40479 = pi12 ? n40397 : n40478;
  assign n40480 = pi11 ? n40337 : n40479;
  assign n40481 = pi10 ? n40239 : n40480;
  assign n40482 = pi09 ? n40040 : n40481;
  assign n40483 = pi08 ? n40022 : n40482;
  assign n40484 = pi07 ? n39371 : n40483;
  assign n40485 = pi19 ? n37334 : n20563;
  assign n40486 = pi18 ? n32 : n40485;
  assign n40487 = pi17 ? n32 : n40486;
  assign n40488 = pi19 ? n32898 : n23648;
  assign n40489 = pi18 ? n20563 : n40488;
  assign n40490 = pi20 ? n25223 : n32;
  assign n40491 = pi19 ? n99 : n40490;
  assign n40492 = pi18 ? n30101 : n40491;
  assign n40493 = pi17 ? n40489 : n40492;
  assign n40494 = pi16 ? n40487 : n40493;
  assign n40495 = pi15 ? n32 : n40494;
  assign n40496 = pi20 ? n37926 : n20563;
  assign n40497 = pi19 ? n40496 : n20563;
  assign n40498 = pi18 ? n32 : n40497;
  assign n40499 = pi17 ? n32 : n40498;
  assign n40500 = pi19 ? n31267 : n38638;
  assign n40501 = pi18 ? n20563 : n40500;
  assign n40502 = pi22 ? n3492 : n32;
  assign n40503 = pi21 ? n99 : n40502;
  assign n40504 = pi20 ? n40503 : n32;
  assign n40505 = pi19 ? n99 : n40504;
  assign n40506 = pi18 ? n99 : n40505;
  assign n40507 = pi17 ? n40501 : n40506;
  assign n40508 = pi16 ? n40499 : n40507;
  assign n40509 = pi20 ? n40054 : n20563;
  assign n40510 = pi19 ? n40509 : n20563;
  assign n40511 = pi18 ? n32 : n40510;
  assign n40512 = pi17 ? n32 : n40511;
  assign n40513 = pi18 ? n20563 : n37588;
  assign n40514 = pi21 ? n99 : n10453;
  assign n40515 = pi20 ? n40514 : n32;
  assign n40516 = pi19 ? n99 : n40515;
  assign n40517 = pi18 ? n99 : n40516;
  assign n40518 = pi17 ? n40513 : n40517;
  assign n40519 = pi16 ? n40512 : n40518;
  assign n40520 = pi15 ? n40508 : n40519;
  assign n40521 = pi14 ? n40495 : n40520;
  assign n40522 = pi13 ? n32 : n40521;
  assign n40523 = pi12 ? n32 : n40522;
  assign n40524 = pi11 ? n32 : n40523;
  assign n40525 = pi10 ? n32 : n40524;
  assign n40526 = pi18 ? n20563 : n37054;
  assign n40527 = pi19 ? n37 : n11395;
  assign n40528 = pi18 ? n32556 : n40527;
  assign n40529 = pi17 ? n40526 : n40528;
  assign n40530 = pi16 ? n39375 : n40529;
  assign n40531 = pi20 ? n36867 : n20563;
  assign n40532 = pi19 ? n40531 : n20563;
  assign n40533 = pi18 ? n32 : n40532;
  assign n40534 = pi17 ? n32 : n40533;
  assign n40535 = pi18 ? n20563 : n31939;
  assign n40536 = pi20 ? n25593 : n32;
  assign n40537 = pi19 ? n37 : n40536;
  assign n40538 = pi18 ? n37 : n40537;
  assign n40539 = pi17 ? n40535 : n40538;
  assign n40540 = pi16 ? n40534 : n40539;
  assign n40541 = pi15 ? n40530 : n40540;
  assign n40542 = pi18 ? n20563 : n32934;
  assign n40543 = pi21 ? n37 : n33324;
  assign n40544 = pi20 ? n40543 : n32;
  assign n40545 = pi19 ? n37 : n40544;
  assign n40546 = pi18 ? n37 : n40545;
  assign n40547 = pi17 ? n40542 : n40546;
  assign n40548 = pi16 ? n40047 : n40547;
  assign n40549 = pi20 ? n28157 : n20563;
  assign n40550 = pi19 ? n40549 : n20563;
  assign n40551 = pi18 ? n32 : n40550;
  assign n40552 = pi17 ? n32 : n40551;
  assign n40553 = pi20 ? n24689 : n32;
  assign n40554 = pi19 ? n9824 : n40553;
  assign n40555 = pi18 ? n37 : n40554;
  assign n40556 = pi17 ? n40041 : n40555;
  assign n40557 = pi16 ? n40552 : n40556;
  assign n40558 = pi15 ? n40548 : n40557;
  assign n40559 = pi14 ? n40541 : n40558;
  assign n40560 = pi20 ? n3083 : n1719;
  assign n40561 = pi19 ? n40560 : n11560;
  assign n40562 = pi18 ? n32619 : n40561;
  assign n40563 = pi17 ? n39415 : n40562;
  assign n40564 = pi16 ? n37930 : n40563;
  assign n40565 = pi20 ? n3090 : n14057;
  assign n40566 = pi19 ? n37 : n40565;
  assign n40567 = pi22 ? n1196 : n32;
  assign n40568 = pi21 ? n139 : n40567;
  assign n40569 = pi20 ? n40568 : n32;
  assign n40570 = pi19 ? n9814 : n40569;
  assign n40571 = pi18 ? n40566 : n40570;
  assign n40572 = pi17 ? n40048 : n40571;
  assign n40573 = pi16 ? n38985 : n40572;
  assign n40574 = pi15 ? n40564 : n40573;
  assign n40575 = pi18 ? n39073 : n37;
  assign n40576 = pi20 ? n37 : n13179;
  assign n40577 = pi19 ? n37 : n40576;
  assign n40578 = pi21 ? n37 : n1721;
  assign n40579 = pi20 ? n37 : n40578;
  assign n40580 = pi19 ? n40579 : n11560;
  assign n40581 = pi18 ? n40577 : n40580;
  assign n40582 = pi17 ? n40575 : n40581;
  assign n40583 = pi16 ? n39001 : n40582;
  assign n40584 = pi18 ? n34869 : n37;
  assign n40585 = pi17 ? n40584 : n40581;
  assign n40586 = pi16 ? n37324 : n40585;
  assign n40587 = pi15 ? n40583 : n40586;
  assign n40588 = pi14 ? n40574 : n40587;
  assign n40589 = pi13 ? n40559 : n40588;
  assign n40590 = pi21 ? n335 : n17630;
  assign n40591 = pi20 ? n40590 : n32;
  assign n40592 = pi19 ? n7676 : n40591;
  assign n40593 = pi18 ? n37 : n40592;
  assign n40594 = pi17 ? n40062 : n40593;
  assign n40595 = pi16 ? n38380 : n40594;
  assign n40596 = pi17 ? n40068 : n40101;
  assign n40597 = pi16 ? n39457 : n40596;
  assign n40598 = pi15 ? n40595 : n40597;
  assign n40599 = pi21 ? n37 : n40091;
  assign n40600 = pi20 ? n40599 : n32;
  assign n40601 = pi19 ? n37 : n40600;
  assign n40602 = pi18 ? n37 : n40601;
  assign n40603 = pi17 ? n38992 : n40602;
  assign n40604 = pi16 ? n35765 : n40603;
  assign n40605 = pi21 ? n2091 : n5003;
  assign n40606 = pi20 ? n40605 : n32;
  assign n40607 = pi19 ? n37 : n40606;
  assign n40608 = pi18 ? n37 : n40607;
  assign n40609 = pi17 ? n38369 : n40608;
  assign n40610 = pi16 ? n36216 : n40609;
  assign n40611 = pi15 ? n40604 : n40610;
  assign n40612 = pi14 ? n40598 : n40611;
  assign n40613 = pi21 ? n2091 : n3125;
  assign n40614 = pi20 ? n40613 : n32;
  assign n40615 = pi19 ? n37 : n40614;
  assign n40616 = pi18 ? n37 : n40615;
  assign n40617 = pi17 ? n39481 : n40616;
  assign n40618 = pi16 ? n36216 : n40617;
  assign n40619 = pi19 ? n37 : n13744;
  assign n40620 = pi18 ? n37 : n40619;
  assign n40621 = pi17 ? n39481 : n40620;
  assign n40622 = pi16 ? n36216 : n40621;
  assign n40623 = pi15 ? n40618 : n40622;
  assign n40624 = pi18 ? n33869 : n37;
  assign n40625 = pi17 ? n40624 : n40620;
  assign n40626 = pi16 ? n36216 : n40625;
  assign n40627 = pi17 ? n39489 : n40620;
  assign n40628 = pi16 ? n36216 : n40627;
  assign n40629 = pi15 ? n40626 : n40628;
  assign n40630 = pi14 ? n40623 : n40629;
  assign n40631 = pi13 ? n40612 : n40630;
  assign n40632 = pi12 ? n40589 : n40631;
  assign n40633 = pi21 ? n18462 : n6416;
  assign n40634 = pi20 ? n40633 : n32;
  assign n40635 = pi19 ? n14198 : n40634;
  assign n40636 = pi18 ? n37 : n40635;
  assign n40637 = pi17 ? n39494 : n40636;
  assign n40638 = pi16 ? n36216 : n40637;
  assign n40639 = pi20 ? n27058 : n32;
  assign n40640 = pi19 ? n5029 : n40639;
  assign n40641 = pi18 ? n37 : n40640;
  assign n40642 = pi17 ? n38425 : n40641;
  assign n40643 = pi16 ? n36216 : n40642;
  assign n40644 = pi15 ? n40638 : n40643;
  assign n40645 = pi19 ? n37 : n40639;
  assign n40646 = pi18 ? n37 : n40645;
  assign n40647 = pi17 ? n38425 : n40646;
  assign n40648 = pi16 ? n36216 : n40647;
  assign n40649 = pi21 ? n3392 : n2637;
  assign n40650 = pi20 ? n40649 : n32;
  assign n40651 = pi19 ? n37 : n40650;
  assign n40652 = pi18 ? n37 : n40651;
  assign n40653 = pi17 ? n38425 : n40652;
  assign n40654 = pi16 ? n36216 : n40653;
  assign n40655 = pi15 ? n40648 : n40654;
  assign n40656 = pi14 ? n40644 : n40655;
  assign n40657 = pi17 ? n37372 : n40646;
  assign n40658 = pi16 ? n36216 : n40657;
  assign n40659 = pi19 ? n19092 : n39523;
  assign n40660 = pi18 ? n37 : n40659;
  assign n40661 = pi17 ? n39497 : n40660;
  assign n40662 = pi16 ? n36216 : n40661;
  assign n40663 = pi15 ? n40658 : n40662;
  assign n40664 = pi18 ? n32899 : n37;
  assign n40665 = pi19 ? n5029 : n39523;
  assign n40666 = pi18 ? n37 : n40665;
  assign n40667 = pi17 ? n40664 : n40666;
  assign n40668 = pi16 ? n36216 : n40667;
  assign n40669 = pi21 ? n31885 : n37;
  assign n40670 = pi20 ? n20563 : n40669;
  assign n40671 = pi19 ? n40670 : n37;
  assign n40672 = pi18 ? n40671 : n37;
  assign n40673 = pi21 ? n6401 : n363;
  assign n40674 = pi20 ? n37 : n40673;
  assign n40675 = pi19 ? n40674 : n12102;
  assign n40676 = pi18 ? n37 : n40675;
  assign n40677 = pi17 ? n40672 : n40676;
  assign n40678 = pi16 ? n36216 : n40677;
  assign n40679 = pi15 ? n40668 : n40678;
  assign n40680 = pi14 ? n40663 : n40679;
  assign n40681 = pi13 ? n40656 : n40680;
  assign n40682 = pi19 ? n27443 : n7408;
  assign n40683 = pi18 ? n37 : n40682;
  assign n40684 = pi17 ? n37377 : n40683;
  assign n40685 = pi16 ? n36216 : n40684;
  assign n40686 = pi18 ? n32369 : n37;
  assign n40687 = pi17 ? n40686 : n40187;
  assign n40688 = pi16 ? n36216 : n40687;
  assign n40689 = pi15 ? n40685 : n40688;
  assign n40690 = pi19 ? n37 : n14305;
  assign n40691 = pi18 ? n37 : n40690;
  assign n40692 = pi17 ? n38449 : n40691;
  assign n40693 = pi16 ? n36216 : n40692;
  assign n40694 = pi19 ? n37 : n38533;
  assign n40695 = pi18 ? n37 : n40694;
  assign n40696 = pi17 ? n38449 : n40695;
  assign n40697 = pi16 ? n36216 : n40696;
  assign n40698 = pi15 ? n40693 : n40697;
  assign n40699 = pi14 ? n40689 : n40698;
  assign n40700 = pi19 ? n31267 : n24269;
  assign n40701 = pi20 ? n17960 : n37;
  assign n40702 = pi19 ? n40701 : n20660;
  assign n40703 = pi18 ? n40700 : n40702;
  assign n40704 = pi20 ? n20660 : n99;
  assign n40705 = pi19 ? n40704 : n99;
  assign n40706 = pi20 ? n2749 : n181;
  assign n40707 = pi23 ? n99 : n31328;
  assign n40708 = pi22 ? n40707 : n747;
  assign n40709 = pi21 ? n40708 : n32;
  assign n40710 = pi20 ? n40709 : n32;
  assign n40711 = pi19 ? n40706 : n40710;
  assign n40712 = pi18 ? n40705 : n40711;
  assign n40713 = pi17 ? n40703 : n40712;
  assign n40714 = pi16 ? n36216 : n40713;
  assign n40715 = pi18 ? n31939 : n99;
  assign n40716 = pi19 ? n7845 : n157;
  assign n40717 = pi19 ? n157 : n6899;
  assign n40718 = pi18 ? n40716 : n40717;
  assign n40719 = pi17 ? n40715 : n40718;
  assign n40720 = pi16 ? n36216 : n40719;
  assign n40721 = pi15 ? n40714 : n40720;
  assign n40722 = pi19 ? n31280 : n26407;
  assign n40723 = pi18 ? n40722 : n99;
  assign n40724 = pi19 ? n19134 : n157;
  assign n40725 = pi22 ? n157 : n3318;
  assign n40726 = pi21 ? n40725 : n32;
  assign n40727 = pi20 ? n40726 : n32;
  assign n40728 = pi19 ? n157 : n40727;
  assign n40729 = pi18 ? n40724 : n40728;
  assign n40730 = pi17 ? n40723 : n40729;
  assign n40731 = pi16 ? n36216 : n40730;
  assign n40732 = pi19 ? n38574 : n29428;
  assign n40733 = pi18 ? n40732 : n99;
  assign n40734 = pi21 ? n32572 : n32;
  assign n40735 = pi20 ? n40734 : n32;
  assign n40736 = pi19 ? n12525 : n40735;
  assign n40737 = pi18 ? n40724 : n40736;
  assign n40738 = pi17 ? n40733 : n40737;
  assign n40739 = pi16 ? n36216 : n40738;
  assign n40740 = pi15 ? n40731 : n40739;
  assign n40741 = pi14 ? n40721 : n40740;
  assign n40742 = pi13 ? n40699 : n40741;
  assign n40743 = pi12 ? n40681 : n40742;
  assign n40744 = pi11 ? n40632 : n40743;
  assign n40745 = pi20 ? n30096 : n3869;
  assign n40746 = pi19 ? n40745 : n99;
  assign n40747 = pi18 ? n40746 : n99;
  assign n40748 = pi22 ? n157 : n3338;
  assign n40749 = pi21 ? n40748 : n32;
  assign n40750 = pi20 ? n40749 : n32;
  assign n40751 = pi19 ? n157 : n40750;
  assign n40752 = pi18 ? n40724 : n40751;
  assign n40753 = pi17 ? n40747 : n40752;
  assign n40754 = pi16 ? n36216 : n40753;
  assign n40755 = pi21 ? n36516 : n37;
  assign n40756 = pi21 ? n2168 : n99;
  assign n40757 = pi20 ? n40755 : n40756;
  assign n40758 = pi19 ? n40757 : n99;
  assign n40759 = pi18 ? n40758 : n99;
  assign n40760 = pi20 ? n19201 : n219;
  assign n40761 = pi19 ? n28194 : n40760;
  assign n40762 = pi21 ? n777 : n204;
  assign n40763 = pi20 ? n40762 : n20978;
  assign n40764 = pi19 ? n40763 : n6936;
  assign n40765 = pi18 ? n40761 : n40764;
  assign n40766 = pi17 ? n40759 : n40765;
  assign n40767 = pi16 ? n36216 : n40766;
  assign n40768 = pi15 ? n40754 : n40767;
  assign n40769 = pi20 ? n7745 : n14844;
  assign n40770 = pi19 ? n40769 : n99;
  assign n40771 = pi18 ? n32934 : n40770;
  assign n40772 = pi20 ? n22965 : n219;
  assign n40773 = pi19 ? n99 : n40772;
  assign n40774 = pi21 ? n3759 : n2402;
  assign n40775 = pi20 ? n40774 : n316;
  assign n40776 = pi19 ? n40775 : n6936;
  assign n40777 = pi18 ? n40773 : n40776;
  assign n40778 = pi17 ? n40771 : n40777;
  assign n40779 = pi16 ? n36923 : n40778;
  assign n40780 = pi19 ? n37 : n21611;
  assign n40781 = pi18 ? n37 : n40780;
  assign n40782 = pi22 ? n99 : n37602;
  assign n40783 = pi21 ? n99 : n40782;
  assign n40784 = pi20 ? n40783 : n316;
  assign n40785 = pi19 ? n40784 : n6936;
  assign n40786 = pi18 ? n99 : n40785;
  assign n40787 = pi17 ? n40781 : n40786;
  assign n40788 = pi16 ? n36216 : n40787;
  assign n40789 = pi15 ? n40779 : n40788;
  assign n40790 = pi14 ? n40768 : n40789;
  assign n40791 = pi21 ? n20563 : n30868;
  assign n40792 = pi20 ? n20563 : n40791;
  assign n40793 = pi19 ? n20563 : n40792;
  assign n40794 = pi18 ? n31315 : n40793;
  assign n40795 = pi17 ? n32 : n40794;
  assign n40796 = pi20 ? n40755 : n37;
  assign n40797 = pi19 ? n40796 : n37;
  assign n40798 = pi18 ? n40797 : n37;
  assign n40799 = pi21 ? n37 : n3711;
  assign n40800 = pi20 ? n37 : n40799;
  assign n40801 = pi21 ? n19292 : n316;
  assign n40802 = pi20 ? n40801 : n1583;
  assign n40803 = pi19 ? n40800 : n40802;
  assign n40804 = pi20 ? n21732 : n2383;
  assign n40805 = pi19 ? n40804 : n6936;
  assign n40806 = pi18 ? n40803 : n40805;
  assign n40807 = pi17 ? n40798 : n40806;
  assign n40808 = pi16 ? n40795 : n40807;
  assign n40809 = pi22 ? n39190 : n37;
  assign n40810 = pi21 ? n40809 : n37;
  assign n40811 = pi20 ? n40810 : n37;
  assign n40812 = pi19 ? n40811 : n37;
  assign n40813 = pi18 ? n40812 : n15029;
  assign n40814 = pi20 ? n2872 : n204;
  assign n40815 = pi20 ? n27675 : n32;
  assign n40816 = pi19 ? n40814 : n40815;
  assign n40817 = pi18 ? n139 : n40816;
  assign n40818 = pi17 ? n40813 : n40817;
  assign n40819 = pi16 ? n40795 : n40818;
  assign n40820 = pi15 ? n40808 : n40819;
  assign n40821 = pi19 ? n40814 : n3978;
  assign n40822 = pi18 ? n139 : n40821;
  assign n40823 = pi17 ? n18075 : n40822;
  assign n40824 = pi16 ? n36227 : n40823;
  assign n40825 = pi20 ? n9354 : n37;
  assign n40826 = pi19 ? n40825 : n9795;
  assign n40827 = pi18 ? n37 : n40826;
  assign n40828 = pi19 ? n40814 : n3177;
  assign n40829 = pi18 ? n139 : n40828;
  assign n40830 = pi17 ? n40827 : n40829;
  assign n40831 = pi16 ? n36216 : n40830;
  assign n40832 = pi15 ? n40824 : n40831;
  assign n40833 = pi14 ? n40820 : n40832;
  assign n40834 = pi13 ? n40790 : n40833;
  assign n40835 = pi19 ? n40825 : n139;
  assign n40836 = pi18 ? n37 : n40835;
  assign n40837 = pi19 ? n16473 : n3177;
  assign n40838 = pi18 ? n139 : n40837;
  assign n40839 = pi17 ? n40836 : n40838;
  assign n40840 = pi16 ? n36216 : n40839;
  assign n40841 = pi19 ? n37 : n1800;
  assign n40842 = pi18 ? n37 : n40841;
  assign n40843 = pi19 ? n16473 : n3304;
  assign n40844 = pi18 ? n139 : n40843;
  assign n40845 = pi17 ? n40842 : n40844;
  assign n40846 = pi16 ? n36216 : n40845;
  assign n40847 = pi15 ? n40840 : n40846;
  assign n40848 = pi19 ? n37 : n947;
  assign n40849 = pi18 ? n37 : n40848;
  assign n40850 = pi20 ? n2318 : n26482;
  assign n40851 = pi19 ? n36541 : n40850;
  assign n40852 = pi20 ? n1026 : n11808;
  assign n40853 = pi19 ? n40852 : n6418;
  assign n40854 = pi18 ? n40851 : n40853;
  assign n40855 = pi17 ? n40849 : n40854;
  assign n40856 = pi16 ? n39086 : n40855;
  assign n40857 = pi20 ? n3924 : n820;
  assign n40858 = pi19 ? n377 : n40857;
  assign n40859 = pi18 ? n37 : n40858;
  assign n40860 = pi21 ? n820 : n335;
  assign n40861 = pi20 ? n939 : n40860;
  assign n40862 = pi21 ? n297 : n569;
  assign n40863 = pi20 ? n3083 : n40862;
  assign n40864 = pi19 ? n40861 : n40863;
  assign n40865 = pi19 ? n13532 : n4117;
  assign n40866 = pi18 ? n40864 : n40865;
  assign n40867 = pi17 ? n40859 : n40866;
  assign n40868 = pi16 ? n36227 : n40867;
  assign n40869 = pi15 ? n40856 : n40868;
  assign n40870 = pi14 ? n40847 : n40869;
  assign n40871 = pi21 ? n574 : n335;
  assign n40872 = pi20 ? n40871 : n642;
  assign n40873 = pi19 ? n37 : n40872;
  assign n40874 = pi18 ? n37 : n40873;
  assign n40875 = pi21 ? n570 : n6361;
  assign n40876 = pi20 ? n604 : n40875;
  assign n40877 = pi21 ? n233 : n570;
  assign n40878 = pi20 ? n40877 : n30657;
  assign n40879 = pi19 ? n40876 : n40878;
  assign n40880 = pi19 ? n30698 : n5831;
  assign n40881 = pi18 ? n40879 : n40880;
  assign n40882 = pi17 ? n40874 : n40881;
  assign n40883 = pi16 ? n36227 : n40882;
  assign n40884 = pi19 ? n39774 : n10012;
  assign n40885 = pi18 ? n37 : n40884;
  assign n40886 = pi17 ? n37 : n40885;
  assign n40887 = pi16 ? n36923 : n40886;
  assign n40888 = pi15 ? n40883 : n40887;
  assign n40889 = pi20 ? n2094 : n8927;
  assign n40890 = pi20 ? n6358 : n38469;
  assign n40891 = pi19 ? n40889 : n40890;
  assign n40892 = pi19 ? n37685 : n2654;
  assign n40893 = pi18 ? n40891 : n40892;
  assign n40894 = pi17 ? n37 : n40893;
  assign n40895 = pi16 ? n36235 : n40894;
  assign n40896 = pi19 ? n6355 : n38470;
  assign n40897 = pi22 ? n233 : n2299;
  assign n40898 = pi21 ? n233 : n40897;
  assign n40899 = pi20 ? n233 : n40898;
  assign n40900 = pi19 ? n40899 : n1823;
  assign n40901 = pi18 ? n40896 : n40900;
  assign n40902 = pi17 ? n37 : n40901;
  assign n40903 = pi16 ? n36227 : n40902;
  assign n40904 = pi15 ? n40895 : n40903;
  assign n40905 = pi14 ? n40888 : n40904;
  assign n40906 = pi13 ? n40870 : n40905;
  assign n40907 = pi12 ? n40834 : n40906;
  assign n40908 = pi22 ? n30865 : n30868;
  assign n40909 = pi21 ? n40908 : n30868;
  assign n40910 = pi20 ? n32 : n40909;
  assign n40911 = pi19 ? n32 : n40910;
  assign n40912 = pi22 ? n40386 : n30868;
  assign n40913 = pi22 ? n30868 : n40386;
  assign n40914 = pi21 ? n40912 : n40913;
  assign n40915 = pi21 ? n30868 : n39801;
  assign n40916 = pi20 ? n40914 : n40915;
  assign n40917 = pi22 ? n20563 : n40386;
  assign n40918 = pi21 ? n40917 : n30868;
  assign n40919 = pi21 ? n31924 : n29133;
  assign n40920 = pi20 ? n40918 : n40919;
  assign n40921 = pi19 ? n40916 : n40920;
  assign n40922 = pi18 ? n40911 : n40921;
  assign n40923 = pi17 ? n32 : n40922;
  assign n40924 = pi19 ? n639 : n7685;
  assign n40925 = pi21 ? n335 : n19438;
  assign n40926 = pi20 ? n335 : n40925;
  assign n40927 = pi19 ? n40926 : n32;
  assign n40928 = pi18 ? n40924 : n40927;
  assign n40929 = pi17 ? n37 : n40928;
  assign n40930 = pi16 ? n40923 : n40929;
  assign n40931 = pi21 ? n40343 : n30868;
  assign n40932 = pi20 ? n32 : n40931;
  assign n40933 = pi19 ? n32 : n40932;
  assign n40934 = pi20 ? n30868 : n33821;
  assign n40935 = pi19 ? n30868 : n40934;
  assign n40936 = pi18 ? n40933 : n40935;
  assign n40937 = pi17 ? n32 : n40936;
  assign n40938 = pi19 ? n33666 : n18408;
  assign n40939 = pi18 ? n37 : n40938;
  assign n40940 = pi20 ? n3292 : n610;
  assign n40941 = pi20 ? n31723 : n335;
  assign n40942 = pi19 ? n40940 : n40941;
  assign n40943 = pi21 ? n335 : n23543;
  assign n40944 = pi20 ? n335 : n40943;
  assign n40945 = pi19 ? n40944 : n32;
  assign n40946 = pi18 ? n40942 : n40945;
  assign n40947 = pi17 ? n40939 : n40946;
  assign n40948 = pi16 ? n40937 : n40947;
  assign n40949 = pi15 ? n40930 : n40948;
  assign n40950 = pi22 ? n30865 : n33792;
  assign n40951 = pi21 ? n40950 : n33792;
  assign n40952 = pi20 ? n32 : n40951;
  assign n40953 = pi19 ? n32 : n40952;
  assign n40954 = pi22 ? n36615 : n20563;
  assign n40955 = pi22 ? n33792 : n36615;
  assign n40956 = pi21 ? n40954 : n40955;
  assign n40957 = pi22 ? n33792 : n20563;
  assign n40958 = pi21 ? n33792 : n40957;
  assign n40959 = pi20 ? n40956 : n40958;
  assign n40960 = pi22 ? n20563 : n36615;
  assign n40961 = pi21 ? n40960 : n20563;
  assign n40962 = pi20 ? n40961 : n33821;
  assign n40963 = pi19 ? n40959 : n40962;
  assign n40964 = pi18 ? n40953 : n40963;
  assign n40965 = pi17 ? n32 : n40964;
  assign n40966 = pi20 ? n581 : n37;
  assign n40967 = pi19 ? n40966 : n14166;
  assign n40968 = pi18 ? n9856 : n40967;
  assign n40969 = pi20 ? n7591 : n610;
  assign n40970 = pi19 ? n40969 : n40941;
  assign n40971 = pi21 ? n233 : n8946;
  assign n40972 = pi20 ? n13527 : n40971;
  assign n40973 = pi19 ? n40972 : n32;
  assign n40974 = pi18 ? n40970 : n40973;
  assign n40975 = pi17 ? n40968 : n40974;
  assign n40976 = pi16 ? n40965 : n40975;
  assign n40977 = pi18 ? n31315 : n33823;
  assign n40978 = pi17 ? n32 : n40977;
  assign n40979 = pi20 ? n5766 : n605;
  assign n40980 = pi19 ? n40979 : n335;
  assign n40981 = pi18 ? n40980 : n335;
  assign n40982 = pi17 ? n40981 : n39850;
  assign n40983 = pi16 ? n40978 : n40982;
  assign n40984 = pi15 ? n40976 : n40983;
  assign n40985 = pi14 ? n40949 : n40984;
  assign n40986 = pi22 ? n20563 : n36659;
  assign n40987 = pi21 ? n40986 : n37;
  assign n40988 = pi20 ? n20563 : n40987;
  assign n40989 = pi19 ? n20563 : n40988;
  assign n40990 = pi18 ? n31315 : n40989;
  assign n40991 = pi17 ? n32 : n40990;
  assign n40992 = pi19 ? n19092 : n7731;
  assign n40993 = pi21 ? n5015 : n2091;
  assign n40994 = pi21 ? n18411 : n22919;
  assign n40995 = pi20 ? n40993 : n40994;
  assign n40996 = pi19 ? n40995 : n32;
  assign n40997 = pi18 ? n40992 : n40996;
  assign n40998 = pi17 ? n37 : n40997;
  assign n40999 = pi16 ? n40991 : n40998;
  assign n41000 = pi18 ? n31315 : n39432;
  assign n41001 = pi17 ? n32 : n41000;
  assign n41002 = pi21 ? n24222 : n696;
  assign n41003 = pi20 ? n37 : n41002;
  assign n41004 = pi19 ? n41003 : n32;
  assign n41005 = pi18 ? n7732 : n41004;
  assign n41006 = pi17 ? n37 : n41005;
  assign n41007 = pi16 ? n41001 : n41006;
  assign n41008 = pi15 ? n40999 : n41007;
  assign n41009 = pi19 ? n37 : n23903;
  assign n41010 = pi18 ? n37 : n41009;
  assign n41011 = pi20 ? n15173 : n7730;
  assign n41012 = pi19 ? n23917 : n41011;
  assign n41013 = pi20 ? n19084 : n15729;
  assign n41014 = pi19 ? n41013 : n32;
  assign n41015 = pi18 ? n41012 : n41014;
  assign n41016 = pi17 ? n41010 : n41015;
  assign n41017 = pi16 ? n39086 : n41016;
  assign n41018 = pi21 ? n36489 : n30843;
  assign n41019 = pi20 ? n38754 : n41018;
  assign n41020 = pi19 ? n20563 : n41019;
  assign n41021 = pi18 ? n31315 : n41020;
  assign n41022 = pi17 ? n32 : n41021;
  assign n41023 = pi19 ? n37 : n37510;
  assign n41024 = pi18 ? n37 : n41023;
  assign n41025 = pi20 ? n9660 : n363;
  assign n41026 = pi19 ? n41025 : n23917;
  assign n41027 = pi20 ? n363 : n39875;
  assign n41028 = pi19 ? n41027 : n32;
  assign n41029 = pi18 ? n41026 : n41028;
  assign n41030 = pi17 ? n41024 : n41029;
  assign n41031 = pi16 ? n41022 : n41030;
  assign n41032 = pi15 ? n41017 : n41031;
  assign n41033 = pi14 ? n41008 : n41032;
  assign n41034 = pi13 ? n40985 : n41033;
  assign n41035 = pi19 ? n37 : n363;
  assign n41036 = pi20 ? n10496 : n15173;
  assign n41037 = pi19 ? n41036 : n37;
  assign n41038 = pi18 ? n41035 : n41037;
  assign n41039 = pi19 ? n5029 : n35670;
  assign n41040 = pi20 ? n2729 : n39889;
  assign n41041 = pi19 ? n41040 : n32;
  assign n41042 = pi18 ? n41039 : n41041;
  assign n41043 = pi17 ? n41038 : n41042;
  assign n41044 = pi16 ? n39086 : n41043;
  assign n41045 = pi20 ? n37 : n38823;
  assign n41046 = pi19 ? n41045 : n32;
  assign n41047 = pi18 ? n37 : n41046;
  assign n41048 = pi17 ? n37 : n41047;
  assign n41049 = pi16 ? n39086 : n41048;
  assign n41050 = pi15 ? n41044 : n41049;
  assign n41051 = pi20 ? n30868 : n38250;
  assign n41052 = pi19 ? n30868 : n41051;
  assign n41053 = pi18 ? n37808 : n41052;
  assign n41054 = pi17 ? n32 : n41053;
  assign n41055 = pi20 ? n99 : n35686;
  assign n41056 = pi19 ? n41055 : n99;
  assign n41057 = pi20 ? n26891 : n37797;
  assign n41058 = pi19 ? n41057 : n32;
  assign n41059 = pi18 ? n41056 : n41058;
  assign n41060 = pi17 ? n99 : n41059;
  assign n41061 = pi16 ? n41054 : n41060;
  assign n41062 = pi19 ? n30868 : n39317;
  assign n41063 = pi18 ? n37808 : n41062;
  assign n41064 = pi17 ? n32 : n41063;
  assign n41065 = pi21 ? n4247 : n99;
  assign n41066 = pi20 ? n139 : n41065;
  assign n41067 = pi20 ? n30766 : n35686;
  assign n41068 = pi19 ? n41066 : n41067;
  assign n41069 = pi18 ? n22703 : n41068;
  assign n41070 = pi20 ? n99 : n23162;
  assign n41071 = pi20 ? n41065 : n32787;
  assign n41072 = pi19 ? n41070 : n41071;
  assign n41073 = pi20 ? n26891 : n14723;
  assign n41074 = pi19 ? n41073 : n32;
  assign n41075 = pi18 ? n41072 : n41074;
  assign n41076 = pi17 ? n41069 : n41075;
  assign n41077 = pi16 ? n41064 : n41076;
  assign n41078 = pi15 ? n41061 : n41077;
  assign n41079 = pi14 ? n41050 : n41078;
  assign n41080 = pi22 ? n37251 : n36798;
  assign n41081 = pi21 ? n41080 : n36798;
  assign n41082 = pi20 ? n32 : n41081;
  assign n41083 = pi19 ? n32 : n41082;
  assign n41084 = pi21 ? n36659 : n37253;
  assign n41085 = pi20 ? n36659 : n41084;
  assign n41086 = pi19 ? n36659 : n41085;
  assign n41087 = pi18 ? n41083 : n41086;
  assign n41088 = pi17 ? n32 : n41087;
  assign n41089 = pi20 ? n139 : n34368;
  assign n41090 = pi21 ? n335 : n685;
  assign n41091 = pi20 ? n335 : n41090;
  assign n41092 = pi19 ? n41089 : n41091;
  assign n41093 = pi18 ? n41092 : n685;
  assign n41094 = pi18 ? n685 : n37856;
  assign n41095 = pi17 ? n41093 : n41094;
  assign n41096 = pi16 ? n41088 : n41095;
  assign n41097 = pi23 ? n33793 : n36659;
  assign n41098 = pi22 ? n41097 : n36798;
  assign n41099 = pi21 ? n41098 : n36798;
  assign n41100 = pi20 ? n32 : n41099;
  assign n41101 = pi19 ? n32 : n41100;
  assign n41102 = pi20 ? n36659 : n39975;
  assign n41103 = pi19 ? n36659 : n41102;
  assign n41104 = pi18 ? n41101 : n41103;
  assign n41105 = pi17 ? n32 : n41104;
  assign n41106 = pi21 ? n40451 : n335;
  assign n41107 = pi20 ? n41106 : n335;
  assign n41108 = pi19 ? n41107 : n41091;
  assign n41109 = pi18 ? n41108 : n685;
  assign n41110 = pi22 ? n685 : n10784;
  assign n41111 = pi21 ? n41110 : n32;
  assign n41112 = pi20 ? n685 : n41111;
  assign n41113 = pi19 ? n41112 : n32;
  assign n41114 = pi18 ? n685 : n41113;
  assign n41115 = pi17 ? n41109 : n41114;
  assign n41116 = pi16 ? n41105 : n41115;
  assign n41117 = pi15 ? n41096 : n41116;
  assign n41118 = pi22 ? n37276 : n36659;
  assign n41119 = pi21 ? n41118 : n36781;
  assign n41120 = pi20 ? n36798 : n41119;
  assign n41121 = pi19 ? n36798 : n41120;
  assign n41122 = pi18 ? n39971 : n41121;
  assign n41123 = pi17 ? n32 : n41122;
  assign n41124 = pi21 ? n40451 : n157;
  assign n41125 = pi20 ? n41124 : n157;
  assign n41126 = pi19 ? n41125 : n157;
  assign n41127 = pi18 ? n41126 : n157;
  assign n41128 = pi22 ? n2244 : n759;
  assign n41129 = pi21 ? n41128 : n32;
  assign n41130 = pi20 ? n157 : n41129;
  assign n41131 = pi19 ? n41130 : n32;
  assign n41132 = pi18 ? n157 : n41131;
  assign n41133 = pi17 ? n41127 : n41132;
  assign n41134 = pi16 ? n41123 : n41133;
  assign n41135 = pi20 ? n36798 : n36781;
  assign n41136 = pi19 ? n36798 : n41135;
  assign n41137 = pi18 ? n40464 : n41136;
  assign n41138 = pi17 ? n32 : n41137;
  assign n41139 = pi22 ? n36781 : n204;
  assign n41140 = pi21 ? n41139 : n157;
  assign n41141 = pi20 ? n41140 : n157;
  assign n41142 = pi19 ? n41141 : n157;
  assign n41143 = pi18 ? n41142 : n157;
  assign n41144 = pi21 ? n7137 : n32;
  assign n41145 = pi20 ? n157 : n41144;
  assign n41146 = pi19 ? n41145 : n32;
  assign n41147 = pi18 ? n157 : n41146;
  assign n41148 = pi17 ? n41143 : n41147;
  assign n41149 = pi16 ? n41138 : n41148;
  assign n41150 = pi15 ? n41134 : n41149;
  assign n41151 = pi14 ? n41117 : n41150;
  assign n41152 = pi13 ? n41079 : n41151;
  assign n41153 = pi12 ? n41034 : n41152;
  assign n41154 = pi11 ? n40907 : n41153;
  assign n41155 = pi10 ? n40744 : n41154;
  assign n41156 = pi09 ? n40525 : n41155;
  assign n41157 = pi19 ? n38377 : n20563;
  assign n41158 = pi18 ? n32 : n41157;
  assign n41159 = pi17 ? n32 : n41158;
  assign n41160 = pi19 ? n31926 : n38638;
  assign n41161 = pi18 ? n20563 : n41160;
  assign n41162 = pi21 ? n99 : n32300;
  assign n41163 = pi20 ? n41162 : n32;
  assign n41164 = pi19 ? n99 : n41163;
  assign n41165 = pi18 ? n99 : n41164;
  assign n41166 = pi17 ? n41161 : n41165;
  assign n41167 = pi16 ? n41159 : n41166;
  assign n41168 = pi19 ? n39454 : n20563;
  assign n41169 = pi18 ? n32 : n41168;
  assign n41170 = pi17 ? n32 : n41169;
  assign n41171 = pi16 ? n41170 : n40518;
  assign n41172 = pi15 ? n41167 : n41171;
  assign n41173 = pi14 ? n40495 : n41172;
  assign n41174 = pi13 ? n32 : n41173;
  assign n41175 = pi12 ? n32 : n41174;
  assign n41176 = pi11 ? n32 : n41175;
  assign n41177 = pi10 ? n32 : n41176;
  assign n41178 = pi18 ? n20563 : n32377;
  assign n41179 = pi17 ? n41178 : n40528;
  assign n41180 = pi16 ? n40025 : n41179;
  assign n41181 = pi19 ? n30118 : n20563;
  assign n41182 = pi18 ? n32 : n41181;
  assign n41183 = pi17 ? n32 : n41182;
  assign n41184 = pi16 ? n41183 : n40539;
  assign n41185 = pi15 ? n41180 : n41184;
  assign n41186 = pi17 ? n40526 : n40546;
  assign n41187 = pi16 ? n40534 : n41186;
  assign n41188 = pi17 ? n40542 : n40555;
  assign n41189 = pi16 ? n38959 : n41188;
  assign n41190 = pi15 ? n41187 : n41189;
  assign n41191 = pi14 ? n41185 : n41190;
  assign n41192 = pi18 ? n34865 : n32934;
  assign n41193 = pi20 ? n25631 : n32;
  assign n41194 = pi19 ? n40560 : n41193;
  assign n41195 = pi18 ? n32619 : n41194;
  assign n41196 = pi17 ? n41192 : n41195;
  assign n41197 = pi16 ? n40047 : n41196;
  assign n41198 = pi18 ? n20563 : n37;
  assign n41199 = pi19 ? n9814 : n41193;
  assign n41200 = pi18 ? n40566 : n41199;
  assign n41201 = pi17 ? n41198 : n41200;
  assign n41202 = pi16 ? n39399 : n41201;
  assign n41203 = pi15 ? n41197 : n41202;
  assign n41204 = pi19 ? n40579 : n12397;
  assign n41205 = pi18 ? n40577 : n41204;
  assign n41206 = pi17 ? n39415 : n41205;
  assign n41207 = pi16 ? n38985 : n41206;
  assign n41208 = pi20 ? n25655 : n32;
  assign n41209 = pi19 ? n40579 : n41208;
  assign n41210 = pi18 ? n40577 : n41209;
  assign n41211 = pi17 ? n40584 : n41210;
  assign n41212 = pi16 ? n40058 : n41211;
  assign n41213 = pi15 ? n41207 : n41212;
  assign n41214 = pi14 ? n41203 : n41213;
  assign n41215 = pi13 ? n41191 : n41214;
  assign n41216 = pi20 ? n26551 : n32;
  assign n41217 = pi19 ? n7676 : n41216;
  assign n41218 = pi18 ? n37 : n41217;
  assign n41219 = pi17 ? n39440 : n41218;
  assign n41220 = pi16 ? n37959 : n41219;
  assign n41221 = pi22 ? n10730 : n32;
  assign n41222 = pi21 ? n335 : n41221;
  assign n41223 = pi20 ? n41222 : n32;
  assign n41224 = pi19 ? n37 : n41223;
  assign n41225 = pi18 ? n37 : n41224;
  assign n41226 = pi17 ? n39440 : n41225;
  assign n41227 = pi16 ? n39001 : n41226;
  assign n41228 = pi15 ? n41220 : n41227;
  assign n41229 = pi18 ? n40228 : n37;
  assign n41230 = pi21 ? n37 : n5783;
  assign n41231 = pi20 ? n41230 : n32;
  assign n41232 = pi19 ? n37 : n41231;
  assign n41233 = pi18 ? n37 : n41232;
  assign n41234 = pi17 ? n41229 : n41233;
  assign n41235 = pi16 ? n39001 : n41234;
  assign n41236 = pi18 ? n40314 : n37;
  assign n41237 = pi21 ? n2091 : n6381;
  assign n41238 = pi20 ? n41237 : n32;
  assign n41239 = pi19 ? n37 : n41238;
  assign n41240 = pi18 ? n37 : n41239;
  assign n41241 = pi17 ? n41236 : n41240;
  assign n41242 = pi16 ? n36216 : n41241;
  assign n41243 = pi15 ? n41235 : n41242;
  assign n41244 = pi14 ? n41228 : n41243;
  assign n41245 = pi21 ? n2091 : n32959;
  assign n41246 = pi20 ? n41245 : n32;
  assign n41247 = pi19 ? n37 : n41246;
  assign n41248 = pi18 ? n37 : n41247;
  assign n41249 = pi17 ? n39481 : n41248;
  assign n41250 = pi16 ? n36216 : n41249;
  assign n41251 = pi21 ? n233 : n26163;
  assign n41252 = pi20 ? n41251 : n32;
  assign n41253 = pi19 ? n37 : n41252;
  assign n41254 = pi18 ? n37 : n41253;
  assign n41255 = pi17 ? n40099 : n41254;
  assign n41256 = pi16 ? n36216 : n41255;
  assign n41257 = pi15 ? n41250 : n41256;
  assign n41258 = pi21 ? n233 : n5813;
  assign n41259 = pi20 ? n41258 : n32;
  assign n41260 = pi19 ? n37 : n41259;
  assign n41261 = pi18 ? n37 : n41260;
  assign n41262 = pi17 ? n39481 : n41261;
  assign n41263 = pi16 ? n36216 : n41262;
  assign n41264 = pi17 ? n38389 : n40620;
  assign n41265 = pi16 ? n36216 : n41264;
  assign n41266 = pi15 ? n41263 : n41265;
  assign n41267 = pi14 ? n41257 : n41266;
  assign n41268 = pi13 ? n41244 : n41267;
  assign n41269 = pi12 ? n41215 : n41268;
  assign n41270 = pi21 ? n35611 : n6416;
  assign n41271 = pi20 ? n41270 : n32;
  assign n41272 = pi19 ? n37 : n41271;
  assign n41273 = pi18 ? n37 : n41272;
  assign n41274 = pi17 ? n39489 : n41273;
  assign n41275 = pi16 ? n36216 : n41274;
  assign n41276 = pi17 ? n39489 : n40641;
  assign n41277 = pi16 ? n36216 : n41276;
  assign n41278 = pi15 ? n41275 : n41277;
  assign n41279 = pi17 ? n39489 : n40646;
  assign n41280 = pi16 ? n36216 : n41279;
  assign n41281 = pi15 ? n41280 : n40654;
  assign n41282 = pi14 ? n41278 : n41281;
  assign n41283 = pi18 ? n32315 : n37;
  assign n41284 = pi17 ? n41283 : n40660;
  assign n41285 = pi16 ? n36216 : n41284;
  assign n41286 = pi15 ? n40658 : n41285;
  assign n41287 = pi18 ? n33916 : n37;
  assign n41288 = pi17 ? n41287 : n40666;
  assign n41289 = pi16 ? n36216 : n41288;
  assign n41290 = pi19 ? n40674 : n12888;
  assign n41291 = pi18 ? n37 : n41290;
  assign n41292 = pi17 ? n37372 : n41291;
  assign n41293 = pi16 ? n36216 : n41292;
  assign n41294 = pi15 ? n41289 : n41293;
  assign n41295 = pi14 ? n41286 : n41294;
  assign n41296 = pi13 ? n41282 : n41295;
  assign n41297 = pi20 ? n27076 : n32;
  assign n41298 = pi19 ? n27443 : n41297;
  assign n41299 = pi18 ? n37 : n41298;
  assign n41300 = pi17 ? n40120 : n41299;
  assign n41301 = pi16 ? n36216 : n41300;
  assign n41302 = pi19 ? n37 : n14724;
  assign n41303 = pi18 ? n37 : n41302;
  assign n41304 = pi17 ? n40120 : n41303;
  assign n41305 = pi16 ? n36216 : n41304;
  assign n41306 = pi15 ? n41301 : n41305;
  assign n41307 = pi19 ? n37 : n15330;
  assign n41308 = pi18 ? n37 : n41307;
  assign n41309 = pi17 ? n40686 : n41308;
  assign n41310 = pi16 ? n36216 : n41309;
  assign n41311 = pi21 ? n20977 : n1009;
  assign n41312 = pi20 ? n41311 : n32;
  assign n41313 = pi19 ? n37 : n41312;
  assign n41314 = pi18 ? n37 : n41313;
  assign n41315 = pi17 ? n40686 : n41314;
  assign n41316 = pi16 ? n36216 : n41315;
  assign n41317 = pi15 ? n41310 : n41316;
  assign n41318 = pi14 ? n41306 : n41317;
  assign n41319 = pi20 ? n37 : n18499;
  assign n41320 = pi19 ? n36897 : n41319;
  assign n41321 = pi20 ? n18500 : n22666;
  assign n41322 = pi21 ? n2746 : n2168;
  assign n41323 = pi19 ? n41321 : n41322;
  assign n41324 = pi18 ? n41320 : n41323;
  assign n41325 = pi20 ? n41322 : n99;
  assign n41326 = pi19 ? n41325 : n99;
  assign n41327 = pi20 ? n99 : n2178;
  assign n41328 = pi21 ? n32579 : n32;
  assign n41329 = pi20 ? n41328 : n32;
  assign n41330 = pi19 ? n41327 : n41329;
  assign n41331 = pi18 ? n41326 : n41330;
  assign n41332 = pi17 ? n41324 : n41331;
  assign n41333 = pi16 ? n36216 : n41332;
  assign n41334 = pi19 ? n40381 : n37;
  assign n41335 = pi18 ? n41334 : n99;
  assign n41336 = pi21 ? n8119 : n32;
  assign n41337 = pi20 ? n41336 : n32;
  assign n41338 = pi19 ? n157 : n41337;
  assign n41339 = pi18 ? n40716 : n41338;
  assign n41340 = pi17 ? n41335 : n41339;
  assign n41341 = pi16 ? n36216 : n41340;
  assign n41342 = pi15 ? n41333 : n41341;
  assign n41343 = pi19 ? n35317 : n26407;
  assign n41344 = pi18 ? n41343 : n99;
  assign n41345 = pi19 ? n157 : n6134;
  assign n41346 = pi18 ? n40724 : n41345;
  assign n41347 = pi17 ? n41344 : n41346;
  assign n41348 = pi16 ? n36216 : n41347;
  assign n41349 = pi20 ? n33821 : n5077;
  assign n41350 = pi19 ? n41349 : n29428;
  assign n41351 = pi18 ? n41350 : n99;
  assign n41352 = pi21 ? n33058 : n32;
  assign n41353 = pi20 ? n41352 : n32;
  assign n41354 = pi19 ? n12525 : n41353;
  assign n41355 = pi18 ? n40724 : n41354;
  assign n41356 = pi17 ? n41351 : n41355;
  assign n41357 = pi16 ? n36216 : n41356;
  assign n41358 = pi15 ? n41348 : n41357;
  assign n41359 = pi14 ? n41342 : n41358;
  assign n41360 = pi13 ? n41318 : n41359;
  assign n41361 = pi12 ? n41296 : n41360;
  assign n41362 = pi11 ? n41269 : n41361;
  assign n41363 = pi20 ? n33821 : n3032;
  assign n41364 = pi19 ? n41363 : n99;
  assign n41365 = pi18 ? n41364 : n99;
  assign n41366 = pi23 ? n15293 : n624;
  assign n41367 = pi22 ? n157 : n41366;
  assign n41368 = pi21 ? n41367 : n32;
  assign n41369 = pi20 ? n41368 : n32;
  assign n41370 = pi19 ? n157 : n41369;
  assign n41371 = pi18 ? n40724 : n41370;
  assign n41372 = pi17 ? n41365 : n41371;
  assign n41373 = pi16 ? n36216 : n41372;
  assign n41374 = pi22 ? n30868 : n30195;
  assign n41375 = pi21 ? n41374 : n37;
  assign n41376 = pi20 ? n41375 : n23686;
  assign n41377 = pi19 ? n41376 : n99;
  assign n41378 = pi18 ? n41377 : n99;
  assign n41379 = pi17 ? n41378 : n40765;
  assign n41380 = pi16 ? n36216 : n41379;
  assign n41381 = pi15 ? n41373 : n41380;
  assign n41382 = pi18 ? n32924 : n40770;
  assign n41383 = pi20 ? n41144 : n32;
  assign n41384 = pi19 ? n40775 : n41383;
  assign n41385 = pi18 ? n40773 : n41384;
  assign n41386 = pi17 ? n41382 : n41385;
  assign n41387 = pi16 ? n36216 : n41386;
  assign n41388 = pi18 ? n31300 : n40780;
  assign n41389 = pi17 ? n41388 : n40786;
  assign n41390 = pi16 ? n36216 : n41389;
  assign n41391 = pi15 ? n41387 : n41390;
  assign n41392 = pi14 ? n41381 : n41391;
  assign n41393 = pi22 ? n30868 : n30869;
  assign n41394 = pi21 ? n41393 : n37;
  assign n41395 = pi20 ? n41394 : n37;
  assign n41396 = pi19 ? n41395 : n37;
  assign n41397 = pi18 ? n41396 : n37;
  assign n41398 = pi17 ? n41397 : n40806;
  assign n41399 = pi16 ? n40795 : n41398;
  assign n41400 = pi22 ? n39190 : n30867;
  assign n41401 = pi21 ? n41400 : n37;
  assign n41402 = pi20 ? n41401 : n37;
  assign n41403 = pi19 ? n41402 : n37;
  assign n41404 = pi18 ? n41403 : n15029;
  assign n41405 = pi20 ? n28084 : n32;
  assign n41406 = pi19 ? n40814 : n41405;
  assign n41407 = pi18 ? n139 : n41406;
  assign n41408 = pi17 ? n41404 : n41407;
  assign n41409 = pi16 ? n40795 : n41408;
  assign n41410 = pi15 ? n41399 : n41409;
  assign n41411 = pi18 ? n32934 : n9766;
  assign n41412 = pi19 ? n40814 : n13837;
  assign n41413 = pi18 ? n139 : n41412;
  assign n41414 = pi17 ? n41411 : n41413;
  assign n41415 = pi16 ? n36923 : n41414;
  assign n41416 = pi18 ? n32934 : n40826;
  assign n41417 = pi21 ? n25285 : n32;
  assign n41418 = pi20 ? n41417 : n32;
  assign n41419 = pi19 ? n40814 : n41418;
  assign n41420 = pi18 ? n139 : n41419;
  assign n41421 = pi17 ? n41416 : n41420;
  assign n41422 = pi16 ? n36216 : n41421;
  assign n41423 = pi15 ? n41415 : n41422;
  assign n41424 = pi14 ? n41410 : n41423;
  assign n41425 = pi13 ? n41392 : n41424;
  assign n41426 = pi18 ? n32934 : n40835;
  assign n41427 = pi17 ? n41426 : n40838;
  assign n41428 = pi16 ? n36216 : n41427;
  assign n41429 = pi18 ? n33966 : n40841;
  assign n41430 = pi17 ? n41429 : n40844;
  assign n41431 = pi16 ? n36216 : n41430;
  assign n41432 = pi15 ? n41428 : n41431;
  assign n41433 = pi16 ? n40176 : n40855;
  assign n41434 = pi19 ? n13532 : n6418;
  assign n41435 = pi18 ? n40864 : n41434;
  assign n41436 = pi17 ? n40859 : n41435;
  assign n41437 = pi16 ? n40176 : n41436;
  assign n41438 = pi15 ? n41433 : n41437;
  assign n41439 = pi14 ? n41432 : n41438;
  assign n41440 = pi16 ? n40176 : n40882;
  assign n41441 = pi19 ? n39774 : n5831;
  assign n41442 = pi18 ? n37 : n41441;
  assign n41443 = pi17 ? n36919 : n41442;
  assign n41444 = pi16 ? n36216 : n41443;
  assign n41445 = pi15 ? n41440 : n41444;
  assign n41446 = pi16 ? n40193 : n40894;
  assign n41447 = pi22 ? n233 : n27667;
  assign n41448 = pi21 ? n233 : n41447;
  assign n41449 = pi20 ? n233 : n41448;
  assign n41450 = pi19 ? n41449 : n2654;
  assign n41451 = pi18 ? n40896 : n41450;
  assign n41452 = pi17 ? n37 : n41451;
  assign n41453 = pi16 ? n36923 : n41452;
  assign n41454 = pi15 ? n41446 : n41453;
  assign n41455 = pi14 ? n41445 : n41454;
  assign n41456 = pi13 ? n41439 : n41455;
  assign n41457 = pi12 ? n41425 : n41456;
  assign n41458 = pi23 ? n34196 : n20563;
  assign n41459 = pi22 ? n41458 : n30868;
  assign n41460 = pi21 ? n41459 : n30868;
  assign n41461 = pi20 ? n32 : n41460;
  assign n41462 = pi19 ? n32 : n41461;
  assign n41463 = pi21 ? n30868 : n40913;
  assign n41464 = pi20 ? n40918 : n31266;
  assign n41465 = pi19 ? n41463 : n41464;
  assign n41466 = pi18 ? n41462 : n41465;
  assign n41467 = pi17 ? n32 : n41466;
  assign n41468 = pi19 ? n12661 : n1823;
  assign n41469 = pi18 ? n40924 : n41468;
  assign n41470 = pi17 ? n37 : n41469;
  assign n41471 = pi16 ? n41467 : n41470;
  assign n41472 = pi20 ? n30868 : n35316;
  assign n41473 = pi19 ? n30868 : n41472;
  assign n41474 = pi18 ? n37808 : n41473;
  assign n41475 = pi17 ? n32 : n41474;
  assign n41476 = pi19 ? n12661 : n32;
  assign n41477 = pi18 ? n40942 : n41476;
  assign n41478 = pi17 ? n40939 : n41477;
  assign n41479 = pi16 ? n41475 : n41478;
  assign n41480 = pi15 ? n41471 : n41479;
  assign n41481 = pi23 ? n33793 : n20563;
  assign n41482 = pi22 ? n41481 : n33792;
  assign n41483 = pi21 ? n41482 : n33792;
  assign n41484 = pi20 ? n32 : n41483;
  assign n41485 = pi19 ? n32 : n41484;
  assign n41486 = pi21 ? n40957 : n40955;
  assign n41487 = pi21 ? n33792 : n40955;
  assign n41488 = pi20 ? n41486 : n41487;
  assign n41489 = pi22 ? n20563 : n37173;
  assign n41490 = pi21 ? n40960 : n41489;
  assign n41491 = pi20 ? n41490 : n35316;
  assign n41492 = pi19 ? n41488 : n41491;
  assign n41493 = pi18 ? n41485 : n41492;
  assign n41494 = pi17 ? n32 : n41493;
  assign n41495 = pi20 ? n13527 : n24109;
  assign n41496 = pi19 ? n41495 : n32;
  assign n41497 = pi18 ? n40970 : n41496;
  assign n41498 = pi17 ? n40968 : n41497;
  assign n41499 = pi16 ? n41494 : n41498;
  assign n41500 = pi18 ? n36655 : n335;
  assign n41501 = pi20 ? n335 : n24109;
  assign n41502 = pi19 ? n41501 : n32;
  assign n41503 = pi18 ? n335 : n41502;
  assign n41504 = pi17 ? n41500 : n41503;
  assign n41505 = pi16 ? n39075 : n41504;
  assign n41506 = pi15 ? n41499 : n41505;
  assign n41507 = pi14 ? n41480 : n41506;
  assign n41508 = pi21 ? n40986 : n31200;
  assign n41509 = pi20 ? n20563 : n41508;
  assign n41510 = pi19 ? n20563 : n41509;
  assign n41511 = pi18 ? n31315 : n41510;
  assign n41512 = pi17 ? n32 : n41511;
  assign n41513 = pi21 ? n18411 : n1423;
  assign n41514 = pi20 ? n40993 : n41513;
  assign n41515 = pi19 ? n41514 : n32;
  assign n41516 = pi18 ? n40992 : n41515;
  assign n41517 = pi17 ? n37 : n41516;
  assign n41518 = pi16 ? n41512 : n41517;
  assign n41519 = pi21 ? n24222 : n1423;
  assign n41520 = pi20 ? n37 : n41519;
  assign n41521 = pi19 ? n41520 : n32;
  assign n41522 = pi18 ? n7732 : n41521;
  assign n41523 = pi17 ? n37 : n41522;
  assign n41524 = pi16 ? n40176 : n41523;
  assign n41525 = pi15 ? n41518 : n41524;
  assign n41526 = pi21 ? n685 : n2230;
  assign n41527 = pi20 ? n19084 : n41526;
  assign n41528 = pi19 ? n41527 : n32;
  assign n41529 = pi18 ? n41012 : n41528;
  assign n41530 = pi17 ? n41010 : n41529;
  assign n41531 = pi16 ? n40176 : n41530;
  assign n41532 = pi21 ? n36489 : n41400;
  assign n41533 = pi20 ? n38754 : n41532;
  assign n41534 = pi19 ? n20563 : n41533;
  assign n41535 = pi18 ? n31315 : n41534;
  assign n41536 = pi17 ? n32 : n41535;
  assign n41537 = pi20 ? n363 : n41526;
  assign n41538 = pi19 ? n41537 : n32;
  assign n41539 = pi18 ? n41026 : n41538;
  assign n41540 = pi17 ? n41024 : n41539;
  assign n41541 = pi16 ? n41536 : n41540;
  assign n41542 = pi15 ? n41531 : n41541;
  assign n41543 = pi14 ? n41525 : n41542;
  assign n41544 = pi13 ? n41507 : n41543;
  assign n41545 = pi16 ? n40176 : n41043;
  assign n41546 = pi20 ? n37 : n39889;
  assign n41547 = pi19 ? n41546 : n32;
  assign n41548 = pi18 ? n37 : n41547;
  assign n41549 = pi17 ? n37 : n41548;
  assign n41550 = pi16 ? n40176 : n41549;
  assign n41551 = pi15 ? n41545 : n41550;
  assign n41552 = pi21 ? n30868 : n37240;
  assign n41553 = pi20 ? n30868 : n41552;
  assign n41554 = pi19 ? n30868 : n41553;
  assign n41555 = pi18 ? n37808 : n41554;
  assign n41556 = pi17 ? n32 : n41555;
  assign n41557 = pi22 ? n11681 : n32;
  assign n41558 = pi21 ? n685 : n41557;
  assign n41559 = pi20 ? n26891 : n41558;
  assign n41560 = pi19 ? n41559 : n32;
  assign n41561 = pi18 ? n41056 : n41560;
  assign n41562 = pi17 ? n99 : n41561;
  assign n41563 = pi16 ? n41556 : n41562;
  assign n41564 = pi22 ? n30868 : n37240;
  assign n41565 = pi21 ? n30868 : n41564;
  assign n41566 = pi20 ? n30868 : n41565;
  assign n41567 = pi19 ? n30868 : n41566;
  assign n41568 = pi18 ? n37808 : n41567;
  assign n41569 = pi17 ? n32 : n41568;
  assign n41570 = pi21 ? n685 : n5370;
  assign n41571 = pi20 ? n26891 : n41570;
  assign n41572 = pi19 ? n41571 : n32;
  assign n41573 = pi18 ? n41072 : n41572;
  assign n41574 = pi17 ? n41069 : n41573;
  assign n41575 = pi16 ? n41569 : n41574;
  assign n41576 = pi15 ? n41563 : n41575;
  assign n41577 = pi14 ? n41551 : n41576;
  assign n41578 = pi21 ? n36659 : n33792;
  assign n41579 = pi20 ? n36659 : n41578;
  assign n41580 = pi19 ? n36659 : n41579;
  assign n41581 = pi18 ? n41083 : n41580;
  assign n41582 = pi17 ? n32 : n41581;
  assign n41583 = pi20 ? n40430 : n34368;
  assign n41584 = pi19 ? n41583 : n41091;
  assign n41585 = pi18 ? n41584 : n685;
  assign n41586 = pi18 ? n685 : n36745;
  assign n41587 = pi17 ? n41585 : n41586;
  assign n41588 = pi16 ? n41582 : n41587;
  assign n41589 = pi18 ? n38899 : n41103;
  assign n41590 = pi17 ? n32 : n41589;
  assign n41591 = pi22 ? n36781 : n39976;
  assign n41592 = pi21 ? n41591 : n335;
  assign n41593 = pi20 ? n41592 : n335;
  assign n41594 = pi19 ? n41593 : n41091;
  assign n41595 = pi18 ? n41594 : n685;
  assign n41596 = pi18 ? n685 : n34771;
  assign n41597 = pi17 ? n41595 : n41596;
  assign n41598 = pi16 ? n41590 : n41597;
  assign n41599 = pi15 ? n41588 : n41598;
  assign n41600 = pi22 ? n36831 : n36798;
  assign n41601 = pi21 ? n41600 : n36798;
  assign n41602 = pi20 ? n32 : n41601;
  assign n41603 = pi19 ? n32 : n41602;
  assign n41604 = pi18 ? n41603 : n41121;
  assign n41605 = pi17 ? n32 : n41604;
  assign n41606 = pi21 ? n41591 : n157;
  assign n41607 = pi20 ? n41606 : n157;
  assign n41608 = pi19 ? n41607 : n157;
  assign n41609 = pi18 ? n41608 : n157;
  assign n41610 = pi22 ? n18448 : n1475;
  assign n41611 = pi21 ? n41610 : n32;
  assign n41612 = pi20 ? n157 : n41611;
  assign n41613 = pi19 ? n41612 : n32;
  assign n41614 = pi18 ? n157 : n41613;
  assign n41615 = pi17 ? n41609 : n41614;
  assign n41616 = pi16 ? n41605 : n41615;
  assign n41617 = pi20 ? n157 : n13398;
  assign n41618 = pi19 ? n41617 : n32;
  assign n41619 = pi18 ? n157 : n41618;
  assign n41620 = pi17 ? n41143 : n41619;
  assign n41621 = pi16 ? n41138 : n41620;
  assign n41622 = pi15 ? n41616 : n41621;
  assign n41623 = pi14 ? n41599 : n41622;
  assign n41624 = pi13 ? n41577 : n41623;
  assign n41625 = pi12 ? n41544 : n41624;
  assign n41626 = pi11 ? n41457 : n41625;
  assign n41627 = pi10 ? n41362 : n41626;
  assign n41628 = pi09 ? n41177 : n41627;
  assign n41629 = pi08 ? n41156 : n41628;
  assign n41630 = pi19 ? n37934 : n20563;
  assign n41631 = pi18 ? n32 : n41630;
  assign n41632 = pi17 ? n32 : n41631;
  assign n41633 = pi18 ? n20563 : n32295;
  assign n41634 = pi19 ? n37 : n33275;
  assign n41635 = pi20 ? n105 : n32;
  assign n41636 = pi19 ? n7776 : n41635;
  assign n41637 = pi18 ? n41634 : n41636;
  assign n41638 = pi17 ? n41633 : n41637;
  assign n41639 = pi16 ? n41632 : n41638;
  assign n41640 = pi15 ? n32 : n41639;
  assign n41641 = pi19 ? n37956 : n20563;
  assign n41642 = pi18 ? n32 : n41641;
  assign n41643 = pi17 ? n32 : n41642;
  assign n41644 = pi18 ? n20563 : n34358;
  assign n41645 = pi21 ? n99 : n4575;
  assign n41646 = pi20 ? n41645 : n32;
  assign n41647 = pi19 ? n99 : n41646;
  assign n41648 = pi18 ? n26408 : n41647;
  assign n41649 = pi17 ? n41644 : n41648;
  assign n41650 = pi16 ? n41643 : n41649;
  assign n41651 = pi19 ? n31221 : n35209;
  assign n41652 = pi18 ? n20563 : n41651;
  assign n41653 = pi21 ? n99 : n303;
  assign n41654 = pi20 ? n41653 : n32;
  assign n41655 = pi19 ? n99 : n41654;
  assign n41656 = pi18 ? n99 : n41655;
  assign n41657 = pi17 ? n41652 : n41656;
  assign n41658 = pi16 ? n41643 : n41657;
  assign n41659 = pi15 ? n41650 : n41658;
  assign n41660 = pi14 ? n41640 : n41659;
  assign n41661 = pi13 ? n32 : n41660;
  assign n41662 = pi12 ? n32 : n41661;
  assign n41663 = pi11 ? n32 : n41662;
  assign n41664 = pi10 ? n32 : n41663;
  assign n41665 = pi22 ? n11889 : n587;
  assign n41666 = pi21 ? n37 : n41665;
  assign n41667 = pi20 ? n41666 : n32;
  assign n41668 = pi19 ? n37 : n41667;
  assign n41669 = pi18 ? n37 : n41668;
  assign n41670 = pi17 ? n41644 : n41669;
  assign n41671 = pi16 ? n40487 : n41670;
  assign n41672 = pi18 ? n20563 : n32899;
  assign n41673 = pi22 ? n583 : n5631;
  assign n41674 = pi21 ? n37 : n41673;
  assign n41675 = pi20 ? n41674 : n32;
  assign n41676 = pi19 ? n37 : n41675;
  assign n41677 = pi18 ? n37 : n41676;
  assign n41678 = pi17 ? n41672 : n41677;
  assign n41679 = pi16 ? n41159 : n41678;
  assign n41680 = pi15 ? n41671 : n41679;
  assign n41681 = pi20 ? n38981 : n20563;
  assign n41682 = pi19 ? n41681 : n20563;
  assign n41683 = pi18 ? n32 : n41682;
  assign n41684 = pi17 ? n32 : n41683;
  assign n41685 = pi18 ? n20563 : n32349;
  assign n41686 = pi21 ? n37 : n35288;
  assign n41687 = pi20 ? n41686 : n32;
  assign n41688 = pi19 ? n37 : n41687;
  assign n41689 = pi18 ? n37 : n41688;
  assign n41690 = pi17 ? n41685 : n41689;
  assign n41691 = pi16 ? n41684 : n41690;
  assign n41692 = pi18 ? n20563 : n32369;
  assign n41693 = pi19 ? n9824 : n40536;
  assign n41694 = pi18 ? n37 : n41693;
  assign n41695 = pi17 ? n41692 : n41694;
  assign n41696 = pi16 ? n39375 : n41695;
  assign n41697 = pi15 ? n41691 : n41696;
  assign n41698 = pi14 ? n41680 : n41697;
  assign n41699 = pi18 ? n20563 : n37649;
  assign n41700 = pi20 ? n3083 : n3096;
  assign n41701 = pi21 ? n139 : n3894;
  assign n41702 = pi20 ? n41701 : n32;
  assign n41703 = pi19 ? n41700 : n41702;
  assign n41704 = pi18 ? n36537 : n41703;
  assign n41705 = pi17 ? n41699 : n41704;
  assign n41706 = pi16 ? n40534 : n41705;
  assign n41707 = pi20 ? n37955 : n20563;
  assign n41708 = pi19 ? n41707 : n20563;
  assign n41709 = pi18 ? n32 : n41708;
  assign n41710 = pi17 ? n32 : n41709;
  assign n41711 = pi20 ? n939 : n947;
  assign n41712 = pi19 ? n37 : n41711;
  assign n41713 = pi19 ? n15004 : n41702;
  assign n41714 = pi18 ? n41712 : n41713;
  assign n41715 = pi17 ? n40535 : n41714;
  assign n41716 = pi16 ? n41710 : n41715;
  assign n41717 = pi15 ? n41706 : n41716;
  assign n41718 = pi19 ? n9814 : n12397;
  assign n41719 = pi18 ? n37 : n41718;
  assign n41720 = pi17 ? n40526 : n41719;
  assign n41721 = pi16 ? n39399 : n41720;
  assign n41722 = pi18 ? n20563 : n32924;
  assign n41723 = pi20 ? n25266 : n32;
  assign n41724 = pi19 ? n9814 : n41723;
  assign n41725 = pi18 ? n37 : n41724;
  assign n41726 = pi17 ? n41722 : n41725;
  assign n41727 = pi16 ? n40552 : n41726;
  assign n41728 = pi15 ? n41721 : n41727;
  assign n41729 = pi14 ? n41717 : n41728;
  assign n41730 = pi13 ? n41698 : n41729;
  assign n41731 = pi17 ? n40542 : n41218;
  assign n41732 = pi16 ? n37930 : n41731;
  assign n41733 = pi21 ? n335 : n5783;
  assign n41734 = pi20 ? n41733 : n32;
  assign n41735 = pi19 ? n37 : n41734;
  assign n41736 = pi18 ? n37 : n41735;
  assign n41737 = pi17 ? n41198 : n41736;
  assign n41738 = pi16 ? n38985 : n41737;
  assign n41739 = pi15 ? n41732 : n41738;
  assign n41740 = pi17 ? n39415 : n41233;
  assign n41741 = pi16 ? n39001 : n41740;
  assign n41742 = pi17 ? n40584 : n41240;
  assign n41743 = pi16 ? n37324 : n41742;
  assign n41744 = pi15 ? n41741 : n41743;
  assign n41745 = pi14 ? n41739 : n41744;
  assign n41746 = pi18 ? n39626 : n37;
  assign n41747 = pi21 ? n233 : n6381;
  assign n41748 = pi20 ? n41747 : n32;
  assign n41749 = pi19 ? n37 : n41748;
  assign n41750 = pi18 ? n37 : n41749;
  assign n41751 = pi17 ? n41746 : n41750;
  assign n41752 = pi16 ? n38380 : n41751;
  assign n41753 = pi18 ? n34295 : n37;
  assign n41754 = pi19 ? n37 : n14675;
  assign n41755 = pi18 ? n37 : n41754;
  assign n41756 = pi17 ? n41753 : n41755;
  assign n41757 = pi16 ? n39457 : n41756;
  assign n41758 = pi15 ? n41752 : n41757;
  assign n41759 = pi18 ? n39585 : n37;
  assign n41760 = pi17 ? n41759 : n41755;
  assign n41761 = pi16 ? n35765 : n41760;
  assign n41762 = pi17 ? n41236 : n41755;
  assign n41763 = pi16 ? n36216 : n41762;
  assign n41764 = pi15 ? n41761 : n41763;
  assign n41765 = pi14 ? n41758 : n41764;
  assign n41766 = pi13 ? n41745 : n41765;
  assign n41767 = pi12 ? n41730 : n41766;
  assign n41768 = pi20 ? n24745 : n32;
  assign n41769 = pi19 ? n37 : n41768;
  assign n41770 = pi18 ? n37 : n41769;
  assign n41771 = pi17 ? n39468 : n41770;
  assign n41772 = pi16 ? n36216 : n41771;
  assign n41773 = pi21 ? n363 : n20889;
  assign n41774 = pi20 ? n41773 : n32;
  assign n41775 = pi19 ? n5029 : n41774;
  assign n41776 = pi18 ? n37 : n41775;
  assign n41777 = pi17 ? n39468 : n41776;
  assign n41778 = pi16 ? n36216 : n41777;
  assign n41779 = pi15 ? n41772 : n41778;
  assign n41780 = pi20 ? n27977 : n32;
  assign n41781 = pi19 ? n37 : n41780;
  assign n41782 = pi18 ? n37 : n41781;
  assign n41783 = pi17 ? n39468 : n41782;
  assign n41784 = pi16 ? n36216 : n41783;
  assign n41785 = pi14 ? n41779 : n41784;
  assign n41786 = pi21 ? n363 : n3319;
  assign n41787 = pi20 ? n41786 : n32;
  assign n41788 = pi19 ? n37 : n41787;
  assign n41789 = pi18 ? n37 : n41788;
  assign n41790 = pi17 ? n39476 : n41789;
  assign n41791 = pi16 ? n36216 : n41790;
  assign n41792 = pi21 ? n363 : n3339;
  assign n41793 = pi20 ? n41792 : n32;
  assign n41794 = pi19 ? n37 : n41793;
  assign n41795 = pi18 ? n37 : n41794;
  assign n41796 = pi17 ? n39481 : n41795;
  assign n41797 = pi16 ? n36216 : n41796;
  assign n41798 = pi15 ? n41791 : n41797;
  assign n41799 = pi18 ? n33858 : n37;
  assign n41800 = pi21 ? n363 : n5829;
  assign n41801 = pi20 ? n41800 : n32;
  assign n41802 = pi19 ? n5029 : n41801;
  assign n41803 = pi18 ? n37 : n41802;
  assign n41804 = pi17 ? n41799 : n41803;
  assign n41805 = pi16 ? n36216 : n41804;
  assign n41806 = pi19 ? n7731 : n40639;
  assign n41807 = pi18 ? n37 : n41806;
  assign n41808 = pi17 ? n38389 : n41807;
  assign n41809 = pi16 ? n36216 : n41808;
  assign n41810 = pi15 ? n41805 : n41809;
  assign n41811 = pi14 ? n41798 : n41810;
  assign n41812 = pi13 ? n41785 : n41811;
  assign n41813 = pi18 ? n34921 : n37;
  assign n41814 = pi19 ? n37 : n41297;
  assign n41815 = pi18 ? n37 : n41814;
  assign n41816 = pi17 ? n41813 : n41815;
  assign n41817 = pi16 ? n36216 : n41816;
  assign n41818 = pi17 ? n39489 : n41303;
  assign n41819 = pi16 ? n36216 : n41818;
  assign n41820 = pi15 ? n41817 : n41819;
  assign n41821 = pi17 ? n38425 : n41308;
  assign n41822 = pi16 ? n36216 : n41821;
  assign n41823 = pi22 ? n37 : n1457;
  assign n41824 = pi21 ? n41823 : n1009;
  assign n41825 = pi20 ? n41824 : n32;
  assign n41826 = pi19 ? n37 : n41825;
  assign n41827 = pi18 ? n37 : n41826;
  assign n41828 = pi17 ? n38425 : n41827;
  assign n41829 = pi16 ? n36216 : n41828;
  assign n41830 = pi15 ? n41822 : n41829;
  assign n41831 = pi14 ? n41820 : n41830;
  assign n41832 = pi19 ? n31221 : n23648;
  assign n41833 = pi20 ? n5077 : n3039;
  assign n41834 = pi19 ? n41833 : n99;
  assign n41835 = pi18 ? n41832 : n41834;
  assign n41836 = pi20 ? n25357 : n32;
  assign n41837 = pi19 ? n99 : n41836;
  assign n41838 = pi18 ? n99 : n41837;
  assign n41839 = pi17 ? n41835 : n41838;
  assign n41840 = pi16 ? n36216 : n41839;
  assign n41841 = pi18 ? n33299 : n99;
  assign n41842 = pi19 ? n157 : n12509;
  assign n41843 = pi18 ? n40716 : n41842;
  assign n41844 = pi17 ? n41841 : n41843;
  assign n41845 = pi16 ? n36216 : n41844;
  assign n41846 = pi15 ? n41840 : n41845;
  assign n41847 = pi19 ? n32314 : n26407;
  assign n41848 = pi18 ? n41847 : n99;
  assign n41849 = pi18 ? n40724 : n41842;
  assign n41850 = pi17 ? n41848 : n41849;
  assign n41851 = pi16 ? n36216 : n41850;
  assign n41852 = pi19 ? n32898 : n26407;
  assign n41853 = pi18 ? n41852 : n99;
  assign n41854 = pi19 ? n6542 : n157;
  assign n41855 = pi19 ? n9035 : n12509;
  assign n41856 = pi18 ? n41854 : n41855;
  assign n41857 = pi17 ? n41853 : n41856;
  assign n41858 = pi16 ? n36216 : n41857;
  assign n41859 = pi15 ? n41851 : n41858;
  assign n41860 = pi14 ? n41846 : n41859;
  assign n41861 = pi13 ? n41831 : n41860;
  assign n41862 = pi12 ? n41812 : n41861;
  assign n41863 = pi11 ? n41767 : n41862;
  assign n41864 = pi20 ? n20563 : n40810;
  assign n41865 = pi19 ? n41864 : n18853;
  assign n41866 = pi18 ? n41865 : n99;
  assign n41867 = pi18 ? n41854 : n41842;
  assign n41868 = pi17 ? n41866 : n41867;
  assign n41869 = pi16 ? n36216 : n41868;
  assign n41870 = pi22 ? n40386 : n30869;
  assign n41871 = pi21 ? n41870 : n37;
  assign n41872 = pi20 ? n20563 : n41871;
  assign n41873 = pi19 ? n41872 : n28235;
  assign n41874 = pi18 ? n41873 : n99;
  assign n41875 = pi22 ? n99 : n456;
  assign n41876 = pi21 ? n37 : n41875;
  assign n41877 = pi20 ? n99 : n41876;
  assign n41878 = pi21 ? n777 : n1027;
  assign n41879 = pi21 ? n10021 : n99;
  assign n41880 = pi20 ? n41878 : n41879;
  assign n41881 = pi19 ? n41877 : n41880;
  assign n41882 = pi21 ? n99 : n204;
  assign n41883 = pi21 ? n2409 : n316;
  assign n41884 = pi20 ? n41882 : n41883;
  assign n41885 = pi19 ? n41884 : n13399;
  assign n41886 = pi18 ? n41881 : n41885;
  assign n41887 = pi17 ? n41874 : n41886;
  assign n41888 = pi16 ? n36216 : n41887;
  assign n41889 = pi15 ? n41869 : n41888;
  assign n41890 = pi18 ? n32899 : n40770;
  assign n41891 = pi21 ? n99 : n41875;
  assign n41892 = pi20 ? n99 : n41891;
  assign n41893 = pi21 ? n3759 : n316;
  assign n41894 = pi21 ? n204 : n99;
  assign n41895 = pi20 ? n41893 : n41894;
  assign n41896 = pi19 ? n41892 : n41895;
  assign n41897 = pi22 ? n37602 : n316;
  assign n41898 = pi21 ? n41897 : n316;
  assign n41899 = pi20 ? n19201 : n41898;
  assign n41900 = pi19 ? n41899 : n13399;
  assign n41901 = pi18 ? n41896 : n41900;
  assign n41902 = pi17 ? n41890 : n41901;
  assign n41903 = pi16 ? n36216 : n41902;
  assign n41904 = pi18 ? n35300 : n40780;
  assign n41905 = pi20 ? n22941 : n316;
  assign n41906 = pi19 ? n41905 : n13399;
  assign n41907 = pi18 ? n99 : n41906;
  assign n41908 = pi17 ? n41904 : n41907;
  assign n41909 = pi16 ? n36216 : n41908;
  assign n41910 = pi15 ? n41903 : n41909;
  assign n41911 = pi14 ? n41889 : n41910;
  assign n41912 = pi21 ? n39801 : n36489;
  assign n41913 = pi21 ? n40281 : n37;
  assign n41914 = pi20 ? n41912 : n41913;
  assign n41915 = pi19 ? n41914 : n37;
  assign n41916 = pi18 ? n41915 : n37;
  assign n41917 = pi21 ? n37 : n19286;
  assign n41918 = pi20 ? n37 : n41917;
  assign n41919 = pi21 ? n19292 : n392;
  assign n41920 = pi20 ? n41919 : n5329;
  assign n41921 = pi19 ? n41918 : n41920;
  assign n41922 = pi22 ? n456 : n1784;
  assign n41923 = pi21 ? n37 : n41922;
  assign n41924 = pi20 ? n41923 : n1027;
  assign n41925 = pi19 ? n41924 : n14328;
  assign n41926 = pi18 ? n41921 : n41925;
  assign n41927 = pi17 ? n41916 : n41926;
  assign n41928 = pi16 ? n40795 : n41927;
  assign n41929 = pi19 ? n38755 : n37;
  assign n41930 = pi18 ? n41929 : n15029;
  assign n41931 = pi19 ? n2317 : n9464;
  assign n41932 = pi18 ? n139 : n41931;
  assign n41933 = pi17 ? n41930 : n41932;
  assign n41934 = pi16 ? n40795 : n41933;
  assign n41935 = pi15 ? n41928 : n41934;
  assign n41936 = pi18 ? n32349 : n9766;
  assign n41937 = pi19 ? n2317 : n13467;
  assign n41938 = pi18 ? n139 : n41937;
  assign n41939 = pi17 ? n41936 : n41938;
  assign n41940 = pi16 ? n36216 : n41939;
  assign n41941 = pi18 ? n32349 : n14115;
  assign n41942 = pi19 ? n2317 : n3978;
  assign n41943 = pi18 ? n139 : n41942;
  assign n41944 = pi17 ? n41941 : n41943;
  assign n41945 = pi16 ? n36216 : n41944;
  assign n41946 = pi15 ? n41940 : n41945;
  assign n41947 = pi14 ? n41935 : n41946;
  assign n41948 = pi13 ? n41911 : n41947;
  assign n41949 = pi18 ? n32349 : n11567;
  assign n41950 = pi17 ? n41949 : n40838;
  assign n41951 = pi16 ? n36216 : n41950;
  assign n41952 = pi19 ? n37 : n2831;
  assign n41953 = pi18 ? n32349 : n41952;
  assign n41954 = pi17 ? n41953 : n40844;
  assign n41955 = pi16 ? n36216 : n41954;
  assign n41956 = pi15 ? n41951 : n41955;
  assign n41957 = pi19 ? n37 : n3645;
  assign n41958 = pi18 ? n32369 : n41957;
  assign n41959 = pi20 ? n2830 : n3096;
  assign n41960 = pi19 ? n23771 : n41959;
  assign n41961 = pi20 ? n139 : n38714;
  assign n41962 = pi19 ? n41961 : n4111;
  assign n41963 = pi18 ? n41960 : n41962;
  assign n41964 = pi17 ? n41958 : n41963;
  assign n41965 = pi16 ? n36216 : n41964;
  assign n41966 = pi20 ? n8742 : n577;
  assign n41967 = pi19 ? n41966 : n7676;
  assign n41968 = pi18 ? n41967 : n41434;
  assign n41969 = pi17 ? n40686 : n41968;
  assign n41970 = pi16 ? n36216 : n41969;
  assign n41971 = pi15 ? n41965 : n41970;
  assign n41972 = pi14 ? n41956 : n41971;
  assign n41973 = pi19 ? n37 : n17483;
  assign n41974 = pi18 ? n32369 : n41973;
  assign n41975 = pi20 ? n604 : n649;
  assign n41976 = pi20 ? n639 : n649;
  assign n41977 = pi19 ? n41975 : n41976;
  assign n41978 = pi19 ? n30698 : n4117;
  assign n41979 = pi18 ? n41977 : n41978;
  assign n41980 = pi17 ? n41974 : n41979;
  assign n41981 = pi16 ? n36216 : n41980;
  assign n41982 = pi22 ? n316 : n685;
  assign n41983 = pi21 ? n233 : n41982;
  assign n41984 = pi20 ? n13527 : n41983;
  assign n41985 = pi19 ? n41984 : n5831;
  assign n41986 = pi18 ? n37 : n41985;
  assign n41987 = pi17 ? n39039 : n41986;
  assign n41988 = pi16 ? n36216 : n41987;
  assign n41989 = pi15 ? n41981 : n41988;
  assign n41990 = pi19 ? n8928 : n6359;
  assign n41991 = pi19 ? n37685 : n10012;
  assign n41992 = pi18 ? n41990 : n41991;
  assign n41993 = pi17 ? n40141 : n41992;
  assign n41994 = pi16 ? n36216 : n41993;
  assign n41995 = pi19 ? n2095 : n37;
  assign n41996 = pi20 ? n233 : n28750;
  assign n41997 = pi19 ? n41996 : n2654;
  assign n41998 = pi18 ? n41995 : n41997;
  assign n41999 = pi17 ? n38449 : n41998;
  assign n42000 = pi16 ? n36216 : n41999;
  assign n42001 = pi15 ? n41994 : n42000;
  assign n42002 = pi14 ? n41989 : n42001;
  assign n42003 = pi13 ? n41972 : n42002;
  assign n42004 = pi12 ? n41948 : n42003;
  assign n42005 = pi21 ? n39801 : n30868;
  assign n42006 = pi21 ? n36489 : n20563;
  assign n42007 = pi20 ? n42005 : n42006;
  assign n42008 = pi19 ? n30868 : n42007;
  assign n42009 = pi18 ? n37808 : n42008;
  assign n42010 = pi17 ? n32 : n42009;
  assign n42011 = pi18 ? n35330 : n41468;
  assign n42012 = pi17 ? n37386 : n42011;
  assign n42013 = pi16 ? n42010 : n42012;
  assign n42014 = pi20 ? n30868 : n20563;
  assign n42015 = pi19 ? n30868 : n42014;
  assign n42016 = pi18 ? n40911 : n42015;
  assign n42017 = pi17 ? n32 : n42016;
  assign n42018 = pi19 ? n37 : n18408;
  assign n42019 = pi18 ? n31939 : n42018;
  assign n42020 = pi19 ? n17204 : n2073;
  assign n42021 = pi18 ? n42020 : n41476;
  assign n42022 = pi17 ? n42019 : n42021;
  assign n42023 = pi16 ? n42017 : n42022;
  assign n42024 = pi15 ? n42013 : n42023;
  assign n42025 = pi19 ? n31280 : n335;
  assign n42026 = pi20 ? n647 : n649;
  assign n42027 = pi19 ? n42026 : n14166;
  assign n42028 = pi18 ? n42025 : n42027;
  assign n42029 = pi20 ? n604 : n610;
  assign n42030 = pi19 ? n42029 : n2073;
  assign n42031 = pi18 ? n42030 : n41496;
  assign n42032 = pi17 ? n42028 : n42031;
  assign n42033 = pi16 ? n36216 : n42032;
  assign n42034 = pi20 ? n31220 : n5766;
  assign n42035 = pi19 ? n42034 : n335;
  assign n42036 = pi18 ? n42035 : n335;
  assign n42037 = pi21 ? n6376 : n665;
  assign n42038 = pi20 ? n335 : n42037;
  assign n42039 = pi19 ? n42038 : n32;
  assign n42040 = pi18 ? n335 : n42039;
  assign n42041 = pi17 ? n42036 : n42040;
  assign n42042 = pi16 ? n36216 : n42041;
  assign n42043 = pi15 ? n42033 : n42042;
  assign n42044 = pi14 ? n42024 : n42043;
  assign n42045 = pi21 ? n20563 : n37231;
  assign n42046 = pi20 ? n42045 : n37;
  assign n42047 = pi19 ? n42046 : n37;
  assign n42048 = pi18 ? n42047 : n37;
  assign n42049 = pi21 ? n2721 : n1423;
  assign n42050 = pi20 ? n363 : n42049;
  assign n42051 = pi19 ? n42050 : n32;
  assign n42052 = pi18 ? n7731 : n42051;
  assign n42053 = pi17 ? n42048 : n42052;
  assign n42054 = pi16 ? n36216 : n42053;
  assign n42055 = pi20 ? n37 : n31485;
  assign n42056 = pi19 ? n42055 : n32;
  assign n42057 = pi18 ? n7732 : n42056;
  assign n42058 = pi17 ? n38449 : n42057;
  assign n42059 = pi16 ? n36216 : n42058;
  assign n42060 = pi15 ? n42054 : n42059;
  assign n42061 = pi18 ? n32377 : n41009;
  assign n42062 = pi20 ? n22881 : n7730;
  assign n42063 = pi19 ? n23917 : n42062;
  assign n42064 = pi18 ? n42063 : n41538;
  assign n42065 = pi17 ? n42061 : n42064;
  assign n42066 = pi16 ? n36216 : n42065;
  assign n42067 = pi19 ? n37 : n34751;
  assign n42068 = pi18 ? n32377 : n42067;
  assign n42069 = pi19 ? n39867 : n23917;
  assign n42070 = pi18 ? n42069 : n41538;
  assign n42071 = pi17 ? n42068 : n42070;
  assign n42072 = pi16 ? n36216 : n42071;
  assign n42073 = pi15 ? n42066 : n42072;
  assign n42074 = pi14 ? n42060 : n42073;
  assign n42075 = pi13 ? n42044 : n42074;
  assign n42076 = pi20 ? n31266 : n7332;
  assign n42077 = pi19 ? n42076 : n363;
  assign n42078 = pi20 ? n363 : n29356;
  assign n42079 = pi19 ? n42078 : n3393;
  assign n42080 = pi18 ? n42077 : n42079;
  assign n42081 = pi20 ? n24865 : n3393;
  assign n42082 = pi20 ? n7730 : n15173;
  assign n42083 = pi19 ? n42081 : n42082;
  assign n42084 = pi20 ? n37 : n39875;
  assign n42085 = pi19 ? n42084 : n32;
  assign n42086 = pi18 ? n42083 : n42085;
  assign n42087 = pi17 ? n42080 : n42086;
  assign n42088 = pi16 ? n36216 : n42087;
  assign n42089 = pi18 ? n36363 : n37;
  assign n42090 = pi17 ? n42089 : n41548;
  assign n42091 = pi16 ? n36216 : n42090;
  assign n42092 = pi15 ? n42088 : n42091;
  assign n42093 = pi18 ? n37808 : n30868;
  assign n42094 = pi17 ? n32 : n42093;
  assign n42095 = pi19 ? n40406 : n99;
  assign n42096 = pi19 ? n99 : n32788;
  assign n42097 = pi18 ? n42095 : n42096;
  assign n42098 = pi21 ? n4538 : n722;
  assign n42099 = pi20 ? n42098 : n32788;
  assign n42100 = pi19 ? n42099 : n34788;
  assign n42101 = pi20 ? n26891 : n38823;
  assign n42102 = pi19 ? n42101 : n32;
  assign n42103 = pi18 ? n42100 : n42102;
  assign n42104 = pi17 ? n42097 : n42103;
  assign n42105 = pi16 ? n42094 : n42104;
  assign n42106 = pi23 ? n33792 : n30868;
  assign n42107 = pi22 ? n30868 : n42106;
  assign n42108 = pi21 ? n30868 : n42107;
  assign n42109 = pi23 ? n30868 : n33792;
  assign n42110 = pi22 ? n30868 : n42109;
  assign n42111 = pi21 ? n42110 : n30868;
  assign n42112 = pi20 ? n42111 : n42106;
  assign n42113 = pi19 ? n42108 : n42112;
  assign n42114 = pi18 ? n37808 : n42113;
  assign n42115 = pi17 ? n32 : n42114;
  assign n42116 = pi22 ? n42106 : n33792;
  assign n42117 = pi21 ? n42116 : n33792;
  assign n42118 = pi20 ? n42117 : n139;
  assign n42119 = pi19 ? n42118 : n139;
  assign n42120 = pi21 ? n20605 : n20228;
  assign n42121 = pi21 ? n363 : n20228;
  assign n42122 = pi20 ? n42120 : n42121;
  assign n42123 = pi19 ? n139 : n42122;
  assign n42124 = pi18 ? n42119 : n42123;
  assign n42125 = pi20 ? n42121 : n363;
  assign n42126 = pi19 ? n42125 : n34221;
  assign n42127 = pi18 ? n42126 : n41074;
  assign n42128 = pi17 ? n42124 : n42127;
  assign n42129 = pi16 ? n42115 : n42128;
  assign n42130 = pi15 ? n42105 : n42129;
  assign n42131 = pi14 ? n42092 : n42130;
  assign n42132 = pi23 ? n33793 : n36798;
  assign n42133 = pi22 ? n42132 : n36798;
  assign n42134 = pi21 ? n42133 : n36798;
  assign n42135 = pi20 ? n32 : n42134;
  assign n42136 = pi19 ? n32 : n42135;
  assign n42137 = pi18 ? n42136 : n41580;
  assign n42138 = pi17 ? n32 : n42137;
  assign n42139 = pi20 ? n33792 : n34368;
  assign n42140 = pi19 ? n42139 : n41091;
  assign n42141 = pi18 ? n42140 : n685;
  assign n42142 = pi17 ? n42141 : n41586;
  assign n42143 = pi16 ? n42138 : n42142;
  assign n42144 = pi18 ? n39971 : n41103;
  assign n42145 = pi17 ? n32 : n42144;
  assign n42146 = pi22 ? n36781 : n36659;
  assign n42147 = pi21 ? n42146 : n36781;
  assign n42148 = pi22 ? n36801 : n36781;
  assign n42149 = pi21 ? n42148 : n335;
  assign n42150 = pi20 ? n42147 : n42149;
  assign n42151 = pi19 ? n42150 : n41091;
  assign n42152 = pi18 ? n42151 : n685;
  assign n42153 = pi17 ? n42152 : n41596;
  assign n42154 = pi16 ? n42145 : n42153;
  assign n42155 = pi15 ? n42143 : n42154;
  assign n42156 = pi20 ? n36798 : n39975;
  assign n42157 = pi19 ? n36798 : n42156;
  assign n42158 = pi18 ? n38899 : n42157;
  assign n42159 = pi17 ? n32 : n42158;
  assign n42160 = pi22 ? n3935 : n157;
  assign n42161 = pi21 ? n42148 : n42160;
  assign n42162 = pi20 ? n42147 : n42161;
  assign n42163 = pi19 ? n42162 : n157;
  assign n42164 = pi18 ? n42163 : n157;
  assign n42165 = pi20 ? n157 : n12508;
  assign n42166 = pi19 ? n42165 : n32;
  assign n42167 = pi18 ? n157 : n42166;
  assign n42168 = pi17 ? n42164 : n42167;
  assign n42169 = pi16 ? n42159 : n42168;
  assign n42170 = pi21 ? n36781 : n36798;
  assign n42171 = pi23 ? n36798 : n363;
  assign n42172 = pi23 ? n36798 : n204;
  assign n42173 = pi22 ? n42171 : n42172;
  assign n42174 = pi21 ? n42173 : n157;
  assign n42175 = pi20 ? n42170 : n42174;
  assign n42176 = pi19 ? n42175 : n157;
  assign n42177 = pi18 ? n42176 : n157;
  assign n42178 = pi22 ? n15294 : n316;
  assign n42179 = pi21 ? n42178 : n32;
  assign n42180 = pi20 ? n157 : n42179;
  assign n42181 = pi19 ? n42180 : n32;
  assign n42182 = pi18 ? n157 : n42181;
  assign n42183 = pi17 ? n42177 : n42182;
  assign n42184 = pi16 ? n41138 : n42183;
  assign n42185 = pi15 ? n42169 : n42184;
  assign n42186 = pi14 ? n42155 : n42185;
  assign n42187 = pi13 ? n42131 : n42186;
  assign n42188 = pi12 ? n42075 : n42187;
  assign n42189 = pi11 ? n42004 : n42188;
  assign n42190 = pi10 ? n41863 : n42189;
  assign n42191 = pi09 ? n41664 : n42190;
  assign n42192 = pi20 ? n30117 : n20563;
  assign n42193 = pi19 ? n32 : n42192;
  assign n42194 = pi18 ? n32 : n42193;
  assign n42195 = pi17 ? n32 : n42194;
  assign n42196 = pi18 ? n20563 : n32877;
  assign n42197 = pi17 ? n42196 : n41637;
  assign n42198 = pi16 ? n42195 : n42197;
  assign n42199 = pi15 ? n32 : n42198;
  assign n42200 = pi19 ? n32 : n38315;
  assign n42201 = pi18 ? n32 : n42200;
  assign n42202 = pi17 ? n32 : n42201;
  assign n42203 = pi18 ? n20563 : n32315;
  assign n42204 = pi17 ? n42203 : n41648;
  assign n42205 = pi16 ? n42202 : n42204;
  assign n42206 = pi19 ? n40055 : n20563;
  assign n42207 = pi18 ? n32 : n42206;
  assign n42208 = pi17 ? n32 : n42207;
  assign n42209 = pi16 ? n42208 : n41657;
  assign n42210 = pi15 ? n42205 : n42209;
  assign n42211 = pi14 ? n42199 : n42210;
  assign n42212 = pi13 ? n32 : n42211;
  assign n42213 = pi12 ? n32 : n42212;
  assign n42214 = pi11 ? n32 : n42213;
  assign n42215 = pi10 ? n32 : n42214;
  assign n42216 = pi18 ? n20563 : n35855;
  assign n42217 = pi22 ? n583 : n587;
  assign n42218 = pi21 ? n37 : n42217;
  assign n42219 = pi20 ? n42218 : n32;
  assign n42220 = pi19 ? n37 : n42219;
  assign n42221 = pi18 ? n37 : n42220;
  assign n42222 = pi17 ? n42216 : n42221;
  assign n42223 = pi16 ? n41632 : n42222;
  assign n42224 = pi18 ? n20563 : n33906;
  assign n42225 = pi17 ? n42224 : n41677;
  assign n42226 = pi16 ? n41159 : n42225;
  assign n42227 = pi15 ? n42223 : n42226;
  assign n42228 = pi18 ? n20563 : n33924;
  assign n42229 = pi17 ? n42228 : n41689;
  assign n42230 = pi16 ? n41170 : n42229;
  assign n42231 = pi16 ? n40025 : n41695;
  assign n42232 = pi15 ? n42230 : n42231;
  assign n42233 = pi14 ? n42227 : n42232;
  assign n42234 = pi18 ? n20563 : n36363;
  assign n42235 = pi19 ? n41700 : n13185;
  assign n42236 = pi18 ? n36537 : n42235;
  assign n42237 = pi17 ? n42234 : n42236;
  assign n42238 = pi16 ? n41183 : n42237;
  assign n42239 = pi19 ? n31264 : n20563;
  assign n42240 = pi18 ? n32 : n42239;
  assign n42241 = pi17 ? n32 : n42240;
  assign n42242 = pi19 ? n15004 : n13185;
  assign n42243 = pi18 ? n41712 : n42242;
  assign n42244 = pi17 ? n40535 : n42243;
  assign n42245 = pi16 ? n42241 : n42244;
  assign n42246 = pi15 ? n42238 : n42245;
  assign n42247 = pi19 ? n9814 : n13185;
  assign n42248 = pi18 ? n37 : n42247;
  assign n42249 = pi17 ? n40535 : n42248;
  assign n42250 = pi16 ? n41710 : n42249;
  assign n42251 = pi18 ? n20563 : n33950;
  assign n42252 = pi20 ? n26118 : n32;
  assign n42253 = pi19 ? n9814 : n42252;
  assign n42254 = pi18 ? n37 : n42253;
  assign n42255 = pi17 ? n42251 : n42254;
  assign n42256 = pi16 ? n38959 : n42255;
  assign n42257 = pi15 ? n42250 : n42256;
  assign n42258 = pi14 ? n42246 : n42257;
  assign n42259 = pi13 ? n42233 : n42258;
  assign n42260 = pi20 ? n627 : n32;
  assign n42261 = pi19 ? n7676 : n42260;
  assign n42262 = pi18 ? n37 : n42261;
  assign n42263 = pi17 ? n40542 : n42262;
  assign n42264 = pi16 ? n40047 : n42263;
  assign n42265 = pi19 ? n40347 : n37;
  assign n42266 = pi18 ? n20563 : n42265;
  assign n42267 = pi21 ? n335 : n18927;
  assign n42268 = pi20 ? n42267 : n32;
  assign n42269 = pi19 ? n37 : n42268;
  assign n42270 = pi18 ? n37 : n42269;
  assign n42271 = pi17 ? n42266 : n42270;
  assign n42272 = pi16 ? n39399 : n42271;
  assign n42273 = pi15 ? n42264 : n42272;
  assign n42274 = pi21 ? n37 : n6990;
  assign n42275 = pi20 ? n42274 : n32;
  assign n42276 = pi19 ? n37 : n42275;
  assign n42277 = pi18 ? n37 : n42276;
  assign n42278 = pi17 ? n41192 : n42277;
  assign n42279 = pi16 ? n38985 : n42278;
  assign n42280 = pi21 ? n2091 : n7009;
  assign n42281 = pi20 ? n42280 : n32;
  assign n42282 = pi19 ? n37 : n42281;
  assign n42283 = pi18 ? n37 : n42282;
  assign n42284 = pi17 ? n40584 : n42283;
  assign n42285 = pi16 ? n40058 : n42284;
  assign n42286 = pi15 ? n42279 : n42285;
  assign n42287 = pi14 ? n42273 : n42286;
  assign n42288 = pi21 ? n233 : n7009;
  assign n42289 = pi20 ? n42288 : n32;
  assign n42290 = pi19 ? n37 : n42289;
  assign n42291 = pi18 ? n37 : n42290;
  assign n42292 = pi17 ? n41753 : n42291;
  assign n42293 = pi16 ? n37959 : n42292;
  assign n42294 = pi18 ? n35799 : n37;
  assign n42295 = pi17 ? n42294 : n41755;
  assign n42296 = pi16 ? n39001 : n42295;
  assign n42297 = pi15 ? n42293 : n42296;
  assign n42298 = pi17 ? n39440 : n41755;
  assign n42299 = pi16 ? n39001 : n42298;
  assign n42300 = pi16 ? n36216 : n41756;
  assign n42301 = pi15 ? n42299 : n42300;
  assign n42302 = pi14 ? n42297 : n42301;
  assign n42303 = pi13 ? n42287 : n42302;
  assign n42304 = pi12 ? n42259 : n42303;
  assign n42305 = pi17 ? n38369 : n41770;
  assign n42306 = pi16 ? n36216 : n42305;
  assign n42307 = pi21 ? n363 : n6406;
  assign n42308 = pi20 ? n42307 : n32;
  assign n42309 = pi19 ? n5029 : n42308;
  assign n42310 = pi18 ? n37 : n42309;
  assign n42311 = pi17 ? n38369 : n42310;
  assign n42312 = pi16 ? n36216 : n42311;
  assign n42313 = pi15 ? n42306 : n42312;
  assign n42314 = pi21 ? n3392 : n748;
  assign n42315 = pi20 ? n42314 : n32;
  assign n42316 = pi19 ? n37 : n42315;
  assign n42317 = pi18 ? n37 : n42316;
  assign n42318 = pi17 ? n38369 : n42317;
  assign n42319 = pi16 ? n36216 : n42318;
  assign n42320 = pi17 ? n38369 : n41782;
  assign n42321 = pi16 ? n36216 : n42320;
  assign n42322 = pi15 ? n42319 : n42321;
  assign n42323 = pi14 ? n42313 : n42322;
  assign n42324 = pi17 ? n39481 : n41789;
  assign n42325 = pi16 ? n36216 : n42324;
  assign n42326 = pi18 ? n32288 : n37;
  assign n42327 = pi21 ? n363 : n6416;
  assign n42328 = pi20 ? n42327 : n32;
  assign n42329 = pi19 ? n37 : n42328;
  assign n42330 = pi18 ? n37 : n42329;
  assign n42331 = pi17 ? n42326 : n42330;
  assign n42332 = pi16 ? n36216 : n42331;
  assign n42333 = pi15 ? n42325 : n42332;
  assign n42334 = pi21 ? n363 : n760;
  assign n42335 = pi20 ? n42334 : n32;
  assign n42336 = pi19 ? n5029 : n42335;
  assign n42337 = pi18 ? n37 : n42336;
  assign n42338 = pi17 ? n40099 : n42337;
  assign n42339 = pi16 ? n36216 : n42338;
  assign n42340 = pi19 ? n7731 : n42335;
  assign n42341 = pi18 ? n37 : n42340;
  assign n42342 = pi17 ? n39476 : n42341;
  assign n42343 = pi16 ? n36216 : n42342;
  assign n42344 = pi15 ? n42339 : n42343;
  assign n42345 = pi14 ? n42333 : n42344;
  assign n42346 = pi13 ? n42323 : n42345;
  assign n42347 = pi20 ? n28002 : n32;
  assign n42348 = pi19 ? n37 : n42347;
  assign n42349 = pi18 ? n37 : n42348;
  assign n42350 = pi17 ? n38389 : n42349;
  assign n42351 = pi16 ? n36216 : n42350;
  assign n42352 = pi20 ? n37797 : n32;
  assign n42353 = pi19 ? n37 : n42352;
  assign n42354 = pi18 ? n37 : n42353;
  assign n42355 = pi17 ? n38389 : n42354;
  assign n42356 = pi16 ? n36216 : n42355;
  assign n42357 = pi15 ? n42351 : n42356;
  assign n42358 = pi19 ? n34246 : n37;
  assign n42359 = pi18 ? n42358 : n37;
  assign n42360 = pi19 ? n37 : n9756;
  assign n42361 = pi18 ? n37 : n42360;
  assign n42362 = pi17 ? n42359 : n42361;
  assign n42363 = pi16 ? n36216 : n42362;
  assign n42364 = pi21 ? n244 : n928;
  assign n42365 = pi20 ? n42364 : n32;
  assign n42366 = pi19 ? n37 : n42365;
  assign n42367 = pi18 ? n37 : n42366;
  assign n42368 = pi17 ? n39489 : n42367;
  assign n42369 = pi16 ? n36216 : n42368;
  assign n42370 = pi15 ? n42363 : n42369;
  assign n42371 = pi14 ? n42357 : n42370;
  assign n42372 = pi19 ? n34920 : n23648;
  assign n42373 = pi18 ? n42372 : n41834;
  assign n42374 = pi21 ? n157 : n1009;
  assign n42375 = pi20 ? n42374 : n32;
  assign n42376 = pi19 ? n99 : n42375;
  assign n42377 = pi18 ? n99 : n42376;
  assign n42378 = pi17 ? n42373 : n42377;
  assign n42379 = pi16 ? n36216 : n42378;
  assign n42380 = pi19 ? n157 : n12920;
  assign n42381 = pi18 ? n40716 : n42380;
  assign n42382 = pi17 ? n41841 : n42381;
  assign n42383 = pi16 ? n36216 : n42382;
  assign n42384 = pi15 ? n42379 : n42383;
  assign n42385 = pi19 ? n32294 : n26407;
  assign n42386 = pi18 ? n42385 : n99;
  assign n42387 = pi17 ? n42386 : n41849;
  assign n42388 = pi16 ? n36216 : n42387;
  assign n42389 = pi19 ? n35776 : n26407;
  assign n42390 = pi18 ? n42389 : n99;
  assign n42391 = pi17 ? n42390 : n41856;
  assign n42392 = pi16 ? n36216 : n42391;
  assign n42393 = pi15 ? n42388 : n42392;
  assign n42394 = pi14 ? n42384 : n42393;
  assign n42395 = pi13 ? n42371 : n42394;
  assign n42396 = pi12 ? n42346 : n42395;
  assign n42397 = pi11 ? n42304 : n42396;
  assign n42398 = pi20 ? n20563 : n41401;
  assign n42399 = pi19 ? n42398 : n18853;
  assign n42400 = pi18 ? n42399 : n99;
  assign n42401 = pi17 ? n42400 : n41867;
  assign n42402 = pi16 ? n36216 : n42401;
  assign n42403 = pi21 ? n39191 : n39182;
  assign n42404 = pi20 ? n20563 : n42403;
  assign n42405 = pi19 ? n42404 : n28235;
  assign n42406 = pi18 ? n42405 : n99;
  assign n42407 = pi17 ? n42406 : n41886;
  assign n42408 = pi16 ? n36216 : n42407;
  assign n42409 = pi15 ? n42402 : n42408;
  assign n42410 = pi18 ? n33916 : n40770;
  assign n42411 = pi17 ? n42410 : n41901;
  assign n42412 = pi16 ? n36216 : n42411;
  assign n42413 = pi18 ? n33916 : n40780;
  assign n42414 = pi17 ? n42413 : n41907;
  assign n42415 = pi16 ? n36216 : n42414;
  assign n42416 = pi15 ? n42412 : n42415;
  assign n42417 = pi14 ? n42409 : n42416;
  assign n42418 = pi21 ? n30868 : n37;
  assign n42419 = pi20 ? n41912 : n42418;
  assign n42420 = pi19 ? n42419 : n37;
  assign n42421 = pi18 ? n42420 : n37;
  assign n42422 = pi20 ? n37 : n2644;
  assign n42423 = pi21 ? n1056 : n3258;
  assign n42424 = pi20 ? n42423 : n5329;
  assign n42425 = pi19 ? n42422 : n42424;
  assign n42426 = pi22 ? n204 : n7262;
  assign n42427 = pi21 ? n42426 : n32;
  assign n42428 = pi20 ? n42427 : n32;
  assign n42429 = pi19 ? n41924 : n42428;
  assign n42430 = pi18 ? n42425 : n42429;
  assign n42431 = pi17 ? n42421 : n42430;
  assign n42432 = pi16 ? n40795 : n42431;
  assign n42433 = pi21 ? n30870 : n37;
  assign n42434 = pi20 ? n38754 : n42433;
  assign n42435 = pi19 ? n42434 : n37;
  assign n42436 = pi18 ? n42435 : n15029;
  assign n42437 = pi22 ? n5061 : n2192;
  assign n42438 = pi21 ? n42437 : n32;
  assign n42439 = pi20 ? n42438 : n32;
  assign n42440 = pi19 ? n2317 : n42439;
  assign n42441 = pi18 ? n139 : n42440;
  assign n42442 = pi17 ? n42436 : n42441;
  assign n42443 = pi16 ? n40795 : n42442;
  assign n42444 = pi15 ? n42432 : n42443;
  assign n42445 = pi18 ? n32899 : n9766;
  assign n42446 = pi19 ? n2317 : n13430;
  assign n42447 = pi18 ? n139 : n42446;
  assign n42448 = pi17 ? n42445 : n42447;
  assign n42449 = pi16 ? n36216 : n42448;
  assign n42450 = pi18 ? n32899 : n14115;
  assign n42451 = pi19 ? n2317 : n14353;
  assign n42452 = pi18 ? n139 : n42451;
  assign n42453 = pi17 ? n42450 : n42452;
  assign n42454 = pi16 ? n36216 : n42453;
  assign n42455 = pi15 ? n42449 : n42454;
  assign n42456 = pi14 ? n42444 : n42455;
  assign n42457 = pi13 ? n42417 : n42456;
  assign n42458 = pi18 ? n32899 : n11567;
  assign n42459 = pi19 ? n16473 : n4082;
  assign n42460 = pi18 ? n139 : n42459;
  assign n42461 = pi17 ? n42458 : n42460;
  assign n42462 = pi16 ? n36216 : n42461;
  assign n42463 = pi18 ? n35300 : n41952;
  assign n42464 = pi17 ? n42463 : n42460;
  assign n42465 = pi16 ? n36216 : n42464;
  assign n42466 = pi15 ? n42462 : n42465;
  assign n42467 = pi18 ? n35300 : n41957;
  assign n42468 = pi19 ? n41961 : n7043;
  assign n42469 = pi18 ? n41960 : n42468;
  assign n42470 = pi17 ? n42467 : n42469;
  assign n42471 = pi16 ? n36216 : n42470;
  assign n42472 = pi19 ? n7685 : n7676;
  assign n42473 = pi19 ? n13532 : n7043;
  assign n42474 = pi18 ? n42472 : n42473;
  assign n42475 = pi17 ? n38443 : n42474;
  assign n42476 = pi16 ? n36216 : n42475;
  assign n42477 = pi15 ? n42471 : n42476;
  assign n42478 = pi14 ? n42466 : n42477;
  assign n42479 = pi18 ? n35300 : n41973;
  assign n42480 = pi19 ? n30698 : n7050;
  assign n42481 = pi18 ? n41977 : n42480;
  assign n42482 = pi17 ? n42479 : n42481;
  assign n42483 = pi16 ? n36216 : n42482;
  assign n42484 = pi19 ? n41984 : n7050;
  assign n42485 = pi18 ? n37 : n42484;
  assign n42486 = pi17 ? n40664 : n42485;
  assign n42487 = pi16 ? n36216 : n42486;
  assign n42488 = pi15 ? n42483 : n42487;
  assign n42489 = pi17 ? n37377 : n41992;
  assign n42490 = pi16 ? n36216 : n42489;
  assign n42491 = pi19 ? n41996 : n10012;
  assign n42492 = pi18 ? n41995 : n42491;
  assign n42493 = pi17 ? n37377 : n42492;
  assign n42494 = pi16 ? n36216 : n42493;
  assign n42495 = pi15 ? n42490 : n42494;
  assign n42496 = pi14 ? n42488 : n42495;
  assign n42497 = pi13 ? n42478 : n42496;
  assign n42498 = pi12 ? n42457 : n42497;
  assign n42499 = pi18 ? n40933 : n42008;
  assign n42500 = pi17 ? n32 : n42499;
  assign n42501 = pi19 ? n12661 : n2654;
  assign n42502 = pi18 ? n35330 : n42501;
  assign n42503 = pi17 ? n38455 : n42502;
  assign n42504 = pi16 ? n42500 : n42503;
  assign n42505 = pi18 ? n36363 : n42018;
  assign n42506 = pi17 ? n42505 : n42021;
  assign n42507 = pi16 ? n42017 : n42506;
  assign n42508 = pi15 ? n42504 : n42507;
  assign n42509 = pi19 ? n36362 : n335;
  assign n42510 = pi18 ? n42509 : n42027;
  assign n42511 = pi20 ? n13527 : n25118;
  assign n42512 = pi19 ? n42511 : n32;
  assign n42513 = pi18 ? n42030 : n42512;
  assign n42514 = pi17 ? n42510 : n42513;
  assign n42515 = pi16 ? n36216 : n42514;
  assign n42516 = pi20 ? n34919 : n649;
  assign n42517 = pi19 ? n42516 : n335;
  assign n42518 = pi18 ? n42517 : n335;
  assign n42519 = pi21 ? n6376 : n17509;
  assign n42520 = pi20 ? n335 : n42519;
  assign n42521 = pi19 ? n42520 : n32;
  assign n42522 = pi18 ? n335 : n42521;
  assign n42523 = pi17 ? n42518 : n42522;
  assign n42524 = pi16 ? n36216 : n42523;
  assign n42525 = pi15 ? n42515 : n42524;
  assign n42526 = pi14 ? n42508 : n42525;
  assign n42527 = pi22 ? n36659 : n30195;
  assign n42528 = pi21 ? n20563 : n42527;
  assign n42529 = pi20 ? n42528 : n37;
  assign n42530 = pi19 ? n42529 : n37;
  assign n42531 = pi18 ? n42530 : n37;
  assign n42532 = pi21 ? n2721 : n2147;
  assign n42533 = pi20 ? n363 : n42532;
  assign n42534 = pi19 ? n42533 : n32;
  assign n42535 = pi18 ? n7731 : n42534;
  assign n42536 = pi17 ? n42531 : n42535;
  assign n42537 = pi16 ? n36216 : n42536;
  assign n42538 = pi21 ? n30843 : n2981;
  assign n42539 = pi20 ? n31925 : n42538;
  assign n42540 = pi19 ? n42539 : n37;
  assign n42541 = pi18 ? n42540 : n37;
  assign n42542 = pi20 ? n37 : n28783;
  assign n42543 = pi19 ? n42542 : n32;
  assign n42544 = pi18 ? n7732 : n42543;
  assign n42545 = pi17 ? n42541 : n42544;
  assign n42546 = pi16 ? n36216 : n42545;
  assign n42547 = pi15 ? n42537 : n42546;
  assign n42548 = pi21 ? n30843 : n3668;
  assign n42549 = pi20 ? n31925 : n42548;
  assign n42550 = pi19 ? n42549 : n37;
  assign n42551 = pi18 ? n42550 : n41009;
  assign n42552 = pi21 ? n685 : n10325;
  assign n42553 = pi20 ? n363 : n42552;
  assign n42554 = pi19 ? n42553 : n32;
  assign n42555 = pi18 ? n42063 : n42554;
  assign n42556 = pi17 ? n42551 : n42555;
  assign n42557 = pi16 ? n36216 : n42556;
  assign n42558 = pi18 ? n42550 : n42067;
  assign n42559 = pi17 ? n42558 : n42070;
  assign n42560 = pi16 ? n36216 : n42559;
  assign n42561 = pi15 ? n42557 : n42560;
  assign n42562 = pi14 ? n42547 : n42561;
  assign n42563 = pi13 ? n42526 : n42562;
  assign n42564 = pi21 ? n30843 : n574;
  assign n42565 = pi20 ? n31925 : n42564;
  assign n42566 = pi19 ? n42565 : n363;
  assign n42567 = pi18 ? n42566 : n42079;
  assign n42568 = pi20 ? n37 : n41526;
  assign n42569 = pi19 ? n42568 : n32;
  assign n42570 = pi18 ? n42083 : n42569;
  assign n42571 = pi17 ? n42567 : n42570;
  assign n42572 = pi16 ? n36216 : n42571;
  assign n42573 = pi17 ? n37377 : n41548;
  assign n42574 = pi16 ? n36216 : n42573;
  assign n42575 = pi15 ? n42572 : n42574;
  assign n42576 = pi20 ? n30868 : n99;
  assign n42577 = pi19 ? n42576 : n99;
  assign n42578 = pi18 ? n42577 : n42096;
  assign n42579 = pi17 ? n42578 : n42103;
  assign n42580 = pi16 ? n42094 : n42579;
  assign n42581 = pi22 ? n36781 : n38271;
  assign n42582 = pi21 ? n37252 : n42581;
  assign n42583 = pi20 ? n32 : n42582;
  assign n42584 = pi19 ? n32 : n42583;
  assign n42585 = pi18 ? n42584 : n33792;
  assign n42586 = pi17 ? n32 : n42585;
  assign n42587 = pi21 ? n36762 : n139;
  assign n42588 = pi20 ? n33792 : n42587;
  assign n42589 = pi19 ? n42588 : n139;
  assign n42590 = pi18 ? n42589 : n42123;
  assign n42591 = pi18 ? n42126 : n41058;
  assign n42592 = pi17 ? n42590 : n42591;
  assign n42593 = pi16 ? n42586 : n42592;
  assign n42594 = pi15 ? n42580 : n42593;
  assign n42595 = pi14 ? n42575 : n42594;
  assign n42596 = pi21 ? n36762 : n335;
  assign n42597 = pi20 ? n33792 : n42596;
  assign n42598 = pi19 ? n42597 : n41091;
  assign n42599 = pi18 ? n42598 : n685;
  assign n42600 = pi18 ? n685 : n37822;
  assign n42601 = pi17 ? n42599 : n42600;
  assign n42602 = pi16 ? n42138 : n42601;
  assign n42603 = pi21 ? n36781 : n335;
  assign n42604 = pi20 ? n42147 : n42603;
  assign n42605 = pi19 ? n42604 : n41091;
  assign n42606 = pi18 ? n42605 : n685;
  assign n42607 = pi20 ? n685 : n13793;
  assign n42608 = pi19 ? n42607 : n32;
  assign n42609 = pi18 ? n685 : n42608;
  assign n42610 = pi17 ? n42606 : n42609;
  assign n42611 = pi16 ? n42145 : n42610;
  assign n42612 = pi15 ? n42602 : n42611;
  assign n42613 = pi21 ? n36781 : n36837;
  assign n42614 = pi20 ? n42147 : n42613;
  assign n42615 = pi19 ? n42614 : n157;
  assign n42616 = pi18 ? n42615 : n157;
  assign n42617 = pi20 ? n157 : n12919;
  assign n42618 = pi19 ? n42617 : n32;
  assign n42619 = pi18 ? n157 : n42618;
  assign n42620 = pi17 ? n42616 : n42619;
  assign n42621 = pi16 ? n42159 : n42620;
  assign n42622 = pi22 ? n36798 : n42172;
  assign n42623 = pi21 ? n42622 : n157;
  assign n42624 = pi20 ? n42170 : n42623;
  assign n42625 = pi19 ? n42624 : n157;
  assign n42626 = pi18 ? n42625 : n157;
  assign n42627 = pi22 ? n18448 : n316;
  assign n42628 = pi21 ? n42627 : n32;
  assign n42629 = pi20 ? n157 : n42628;
  assign n42630 = pi19 ? n42629 : n32;
  assign n42631 = pi18 ? n157 : n42630;
  assign n42632 = pi17 ? n42626 : n42631;
  assign n42633 = pi16 ? n41138 : n42632;
  assign n42634 = pi15 ? n42621 : n42633;
  assign n42635 = pi14 ? n42612 : n42634;
  assign n42636 = pi13 ? n42595 : n42635;
  assign n42637 = pi12 ? n42563 : n42636;
  assign n42638 = pi11 ? n42498 : n42637;
  assign n42639 = pi10 ? n42397 : n42638;
  assign n42640 = pi09 ? n42215 : n42639;
  assign n42641 = pi08 ? n42191 : n42640;
  assign n42642 = pi07 ? n41629 : n42641;
  assign n42643 = pi06 ? n40484 : n42642;
  assign n42644 = pi19 ? n32 : n40044;
  assign n42645 = pi18 ? n32 : n42644;
  assign n42646 = pi17 ? n32 : n42645;
  assign n42647 = pi18 ? n20563 : n34295;
  assign n42648 = pi20 ? n121 : n32;
  assign n42649 = pi19 ? n6489 : n42648;
  assign n42650 = pi18 ? n34262 : n42649;
  assign n42651 = pi17 ? n42647 : n42650;
  assign n42652 = pi16 ? n42646 : n42651;
  assign n42653 = pi15 ? n32 : n42652;
  assign n42654 = pi19 ? n32 : n39396;
  assign n42655 = pi18 ? n32 : n42654;
  assign n42656 = pi17 ? n32 : n42655;
  assign n42657 = pi18 ? n20563 : n33260;
  assign n42658 = pi20 ? n142 : n32;
  assign n42659 = pi19 ? n22400 : n42658;
  assign n42660 = pi18 ? n26408 : n42659;
  assign n42661 = pi17 ? n42657 : n42660;
  assign n42662 = pi16 ? n42656 : n42661;
  assign n42663 = pi18 ? n20563 : n33285;
  assign n42664 = pi20 ? n37 : n3871;
  assign n42665 = pi20 ? n2973 : n39676;
  assign n42666 = pi19 ? n42664 : n42665;
  assign n42667 = pi20 ? n14526 : n23671;
  assign n42668 = pi21 ? n2156 : n141;
  assign n42669 = pi20 ? n42668 : n32;
  assign n42670 = pi19 ? n42667 : n42669;
  assign n42671 = pi18 ? n42666 : n42670;
  assign n42672 = pi17 ? n42663 : n42671;
  assign n42673 = pi16 ? n42656 : n42672;
  assign n42674 = pi15 ? n42662 : n42673;
  assign n42675 = pi14 ? n42653 : n42674;
  assign n42676 = pi13 ? n32 : n42675;
  assign n42677 = pi12 ? n32 : n42676;
  assign n42678 = pi11 ? n32 : n42677;
  assign n42679 = pi10 ? n32 : n42678;
  assign n42680 = pi19 ? n32 : n40549;
  assign n42681 = pi18 ? n32 : n42680;
  assign n42682 = pi17 ? n32 : n42681;
  assign n42683 = pi19 ? n37 : n13051;
  assign n42684 = pi18 ? n37 : n42683;
  assign n42685 = pi17 ? n42663 : n42684;
  assign n42686 = pi16 ? n42682 : n42685;
  assign n42687 = pi19 ? n36868 : n20563;
  assign n42688 = pi18 ? n32 : n42687;
  assign n42689 = pi17 ? n32 : n42688;
  assign n42690 = pi18 ? n20563 : n33299;
  assign n42691 = pi22 ? n139 : n1370;
  assign n42692 = pi21 ? n37 : n42691;
  assign n42693 = pi20 ? n42692 : n32;
  assign n42694 = pi19 ? n37 : n42693;
  assign n42695 = pi18 ? n37 : n42694;
  assign n42696 = pi17 ? n42690 : n42695;
  assign n42697 = pi16 ? n42689 : n42696;
  assign n42698 = pi15 ? n42686 : n42697;
  assign n42699 = pi19 ? n38998 : n20563;
  assign n42700 = pi18 ? n32 : n42699;
  assign n42701 = pi17 ? n32 : n42700;
  assign n42702 = pi22 ? n139 : n1378;
  assign n42703 = pi21 ? n37 : n42702;
  assign n42704 = pi20 ? n42703 : n32;
  assign n42705 = pi19 ? n37 : n42704;
  assign n42706 = pi18 ? n37 : n42705;
  assign n42707 = pi17 ? n41633 : n42706;
  assign n42708 = pi16 ? n42701 : n42707;
  assign n42709 = pi22 ? n139 : n5631;
  assign n42710 = pi21 ? n139 : n42709;
  assign n42711 = pi20 ? n42710 : n32;
  assign n42712 = pi19 ? n3086 : n42711;
  assign n42713 = pi18 ? n12371 : n42712;
  assign n42714 = pi17 ? n41633 : n42713;
  assign n42715 = pi16 ? n42701 : n42714;
  assign n42716 = pi15 ? n42708 : n42715;
  assign n42717 = pi14 ? n42698 : n42716;
  assign n42718 = pi19 ? n139 : n13636;
  assign n42719 = pi18 ? n9766 : n42718;
  assign n42720 = pi17 ? n41633 : n42719;
  assign n42721 = pi16 ? n41159 : n42720;
  assign n42722 = pi20 ? n3096 : n942;
  assign n42723 = pi19 ? n42722 : n13185;
  assign n42724 = pi18 ? n37 : n42723;
  assign n42725 = pi17 ? n41644 : n42724;
  assign n42726 = pi16 ? n41170 : n42725;
  assign n42727 = pi15 ? n42721 : n42726;
  assign n42728 = pi21 ? n335 : n4736;
  assign n42729 = pi20 ? n42728 : n32;
  assign n42730 = pi19 ? n577 : n42729;
  assign n42731 = pi18 ? n37 : n42730;
  assign n42732 = pi17 ? n41672 : n42731;
  assign n42733 = pi16 ? n40512 : n42732;
  assign n42734 = pi19 ? n577 : n42260;
  assign n42735 = pi18 ? n37 : n42734;
  assign n42736 = pi17 ? n41672 : n42735;
  assign n42737 = pi16 ? n39375 : n42736;
  assign n42738 = pi15 ? n42733 : n42737;
  assign n42739 = pi14 ? n42727 : n42738;
  assign n42740 = pi13 ? n42717 : n42739;
  assign n42741 = pi19 ? n37 : n42260;
  assign n42742 = pi18 ? n37 : n42741;
  assign n42743 = pi17 ? n42234 : n42742;
  assign n42744 = pi16 ? n40534 : n42743;
  assign n42745 = pi21 ? n37 : n18927;
  assign n42746 = pi20 ? n42745 : n32;
  assign n42747 = pi19 ? n37 : n42746;
  assign n42748 = pi18 ? n37 : n42747;
  assign n42749 = pi17 ? n41178 : n42748;
  assign n42750 = pi16 ? n41710 : n42749;
  assign n42751 = pi15 ? n42744 : n42750;
  assign n42752 = pi18 ? n37448 : n42269;
  assign n42753 = pi17 ? n40535 : n42752;
  assign n42754 = pi16 ? n39399 : n42753;
  assign n42755 = pi20 ? n27017 : n32;
  assign n42756 = pi19 ? n7685 : n42755;
  assign n42757 = pi18 ? n37448 : n42756;
  assign n42758 = pi17 ? n41722 : n42757;
  assign n42759 = pi16 ? n40552 : n42758;
  assign n42760 = pi15 ? n42754 : n42759;
  assign n42761 = pi14 ? n42751 : n42760;
  assign n42762 = pi19 ? n37 : n42755;
  assign n42763 = pi18 ? n37 : n42762;
  assign n42764 = pi17 ? n39415 : n42763;
  assign n42765 = pi16 ? n37930 : n42764;
  assign n42766 = pi19 ? n37 : n12818;
  assign n42767 = pi18 ? n37 : n42766;
  assign n42768 = pi17 ? n41198 : n42767;
  assign n42769 = pi16 ? n38985 : n42768;
  assign n42770 = pi15 ? n42765 : n42769;
  assign n42771 = pi20 ? n647 : n604;
  assign n42772 = pi19 ? n37 : n42771;
  assign n42773 = pi19 ? n11632 : n13258;
  assign n42774 = pi18 ? n42772 : n42773;
  assign n42775 = pi17 ? n41198 : n42774;
  assign n42776 = pi16 ? n39001 : n42775;
  assign n42777 = pi20 ? n30408 : n32;
  assign n42778 = pi19 ? n37 : n42777;
  assign n42779 = pi18 ? n37 : n42778;
  assign n42780 = pi17 ? n39415 : n42779;
  assign n42781 = pi16 ? n37324 : n42780;
  assign n42782 = pi15 ? n42776 : n42781;
  assign n42783 = pi14 ? n42770 : n42782;
  assign n42784 = pi13 ? n42761 : n42783;
  assign n42785 = pi12 ? n42740 : n42784;
  assign n42786 = pi21 ? n37 : n8486;
  assign n42787 = pi20 ? n42786 : n32;
  assign n42788 = pi19 ? n37 : n42787;
  assign n42789 = pi18 ? n37 : n42788;
  assign n42790 = pi17 ? n40584 : n42789;
  assign n42791 = pi16 ? n38380 : n42790;
  assign n42792 = pi20 ? n28913 : n32;
  assign n42793 = pi19 ? n37 : n42792;
  assign n42794 = pi18 ? n37 : n42793;
  assign n42795 = pi17 ? n40575 : n42794;
  assign n42796 = pi16 ? n38380 : n42795;
  assign n42797 = pi15 ? n42791 : n42796;
  assign n42798 = pi17 ? n40584 : n42794;
  assign n42799 = pi16 ? n34860 : n42798;
  assign n42800 = pi21 ? n5015 : n21387;
  assign n42801 = pi20 ? n42800 : n32;
  assign n42802 = pi19 ? n37 : n42801;
  assign n42803 = pi18 ? n41009 : n42802;
  assign n42804 = pi17 ? n39440 : n42803;
  assign n42805 = pi16 ? n35765 : n42804;
  assign n42806 = pi15 ? n42799 : n42805;
  assign n42807 = pi14 ? n42797 : n42806;
  assign n42808 = pi21 ? n363 : n32959;
  assign n42809 = pi20 ? n42808 : n32;
  assign n42810 = pi19 ? n5029 : n42809;
  assign n42811 = pi18 ? n37 : n42810;
  assign n42812 = pi17 ? n39448 : n42811;
  assign n42813 = pi16 ? n36216 : n42812;
  assign n42814 = pi19 ? n37 : n14699;
  assign n42815 = pi18 ? n37 : n42814;
  assign n42816 = pi17 ? n41753 : n42815;
  assign n42817 = pi16 ? n36216 : n42816;
  assign n42818 = pi15 ? n42813 : n42817;
  assign n42819 = pi17 ? n40068 : n42349;
  assign n42820 = pi16 ? n36216 : n42819;
  assign n42821 = pi21 ? n9657 : n2106;
  assign n42822 = pi20 ? n13310 : n42821;
  assign n42823 = pi19 ? n42822 : n42347;
  assign n42824 = pi18 ? n15175 : n42823;
  assign n42825 = pi17 ? n41746 : n42824;
  assign n42826 = pi16 ? n36216 : n42825;
  assign n42827 = pi15 ? n42820 : n42826;
  assign n42828 = pi14 ? n42818 : n42827;
  assign n42829 = pi13 ? n42807 : n42828;
  assign n42830 = pi17 ? n38369 : n42349;
  assign n42831 = pi16 ? n36216 : n42830;
  assign n42832 = pi21 ? n381 : n882;
  assign n42833 = pi20 ? n42832 : n32;
  assign n42834 = pi19 ? n37 : n42833;
  assign n42835 = pi18 ? n37 : n42834;
  assign n42836 = pi17 ? n38369 : n42835;
  assign n42837 = pi16 ? n36216 : n42836;
  assign n42838 = pi15 ? n42831 : n42837;
  assign n42839 = pi21 ? n244 : n882;
  assign n42840 = pi20 ? n42839 : n32;
  assign n42841 = pi19 ? n37 : n42840;
  assign n42842 = pi18 ? n37 : n42841;
  assign n42843 = pi17 ? n38369 : n42842;
  assign n42844 = pi16 ? n36216 : n42843;
  assign n42845 = pi19 ? n37 : n17013;
  assign n42846 = pi19 ? n7746 : n42365;
  assign n42847 = pi18 ? n42845 : n42846;
  assign n42848 = pi17 ? n39463 : n42847;
  assign n42849 = pi16 ? n36216 : n42848;
  assign n42850 = pi15 ? n42844 : n42849;
  assign n42851 = pi14 ? n42838 : n42850;
  assign n42852 = pi18 ? n32275 : n21612;
  assign n42853 = pi21 ? n7429 : n1009;
  assign n42854 = pi20 ? n42853 : n32;
  assign n42855 = pi19 ? n99 : n42854;
  assign n42856 = pi18 ? n99 : n42855;
  assign n42857 = pi17 ? n42852 : n42856;
  assign n42858 = pi16 ? n36216 : n42857;
  assign n42859 = pi22 ? n316 : n18448;
  assign n42860 = pi21 ? n42859 : n1009;
  assign n42861 = pi20 ? n42860 : n32;
  assign n42862 = pi19 ? n157 : n42861;
  assign n42863 = pi18 ? n17340 : n42862;
  assign n42864 = pi17 ? n42852 : n42863;
  assign n42865 = pi16 ? n36216 : n42864;
  assign n42866 = pi15 ? n42858 : n42865;
  assign n42867 = pi18 ? n33285 : n21612;
  assign n42868 = pi20 ? n17337 : n10532;
  assign n42869 = pi19 ? n99 : n42868;
  assign n42870 = pi19 ? n157 : n13399;
  assign n42871 = pi18 ? n42869 : n42870;
  assign n42872 = pi17 ? n42867 : n42871;
  assign n42873 = pi16 ? n36216 : n42872;
  assign n42874 = pi19 ? n38638 : n99;
  assign n42875 = pi18 ? n34891 : n42874;
  assign n42876 = pi18 ? n99 : n41842;
  assign n42877 = pi17 ? n42875 : n42876;
  assign n42878 = pi16 ? n36216 : n42877;
  assign n42879 = pi15 ? n42873 : n42878;
  assign n42880 = pi14 ? n42866 : n42879;
  assign n42881 = pi13 ? n42851 : n42880;
  assign n42882 = pi12 ? n42829 : n42881;
  assign n42883 = pi11 ? n42785 : n42882;
  assign n42884 = pi18 ? n38549 : n19774;
  assign n42885 = pi21 ? n99 : n3759;
  assign n42886 = pi20 ? n42885 : n204;
  assign n42887 = pi19 ? n42886 : n13399;
  assign n42888 = pi18 ? n99 : n42887;
  assign n42889 = pi17 ? n42884 : n42888;
  assign n42890 = pi16 ? n36216 : n42889;
  assign n42891 = pi21 ? n40809 : n2957;
  assign n42892 = pi20 ? n42891 : n3042;
  assign n42893 = pi19 ? n20563 : n42892;
  assign n42894 = pi18 ? n42893 : n99;
  assign n42895 = pi20 ? n24957 : n36505;
  assign n42896 = pi19 ? n99 : n42895;
  assign n42897 = pi19 ? n38631 : n13399;
  assign n42898 = pi18 ? n42896 : n42897;
  assign n42899 = pi17 ? n42894 : n42898;
  assign n42900 = pi16 ? n36216 : n42899;
  assign n42901 = pi15 ? n42890 : n42900;
  assign n42902 = pi18 ? n33858 : n30851;
  assign n42903 = pi20 ? n24957 : n99;
  assign n42904 = pi19 ? n21611 : n42903;
  assign n42905 = pi18 ? n42904 : n42897;
  assign n42906 = pi17 ? n42902 : n42905;
  assign n42907 = pi16 ? n36216 : n42906;
  assign n42908 = pi20 ? n1912 : n1019;
  assign n42909 = pi19 ? n42908 : n13399;
  assign n42910 = pi18 ? n37 : n42909;
  assign n42911 = pi17 ? n39476 : n42910;
  assign n42912 = pi16 ? n36216 : n42911;
  assign n42913 = pi15 ? n42907 : n42912;
  assign n42914 = pi14 ? n42901 : n42913;
  assign n42915 = pi20 ? n20563 : n38754;
  assign n42916 = pi19 ? n42915 : n32933;
  assign n42917 = pi18 ? n42916 : n37;
  assign n42918 = pi19 ? n37 : n39745;
  assign n42919 = pi19 ? n22775 : n14754;
  assign n42920 = pi18 ? n42918 : n42919;
  assign n42921 = pi17 ? n42917 : n42920;
  assign n42922 = pi16 ? n36216 : n42921;
  assign n42923 = pi18 ? n33869 : n15029;
  assign n42924 = pi19 ? n1017 : n15408;
  assign n42925 = pi18 ? n139 : n42924;
  assign n42926 = pi17 ? n42923 : n42925;
  assign n42927 = pi16 ? n36216 : n42926;
  assign n42928 = pi15 ? n42922 : n42927;
  assign n42929 = pi18 ? n32877 : n14115;
  assign n42930 = pi19 ? n1017 : n13430;
  assign n42931 = pi18 ? n139 : n42930;
  assign n42932 = pi17 ? n42929 : n42931;
  assign n42933 = pi16 ? n36216 : n42932;
  assign n42934 = pi18 ? n33299 : n9815;
  assign n42935 = pi19 ? n1017 : n14353;
  assign n42936 = pi18 ? n139 : n42935;
  assign n42937 = pi17 ? n42934 : n42936;
  assign n42938 = pi16 ? n36216 : n42937;
  assign n42939 = pi15 ? n42933 : n42938;
  assign n42940 = pi14 ? n42928 : n42939;
  assign n42941 = pi13 ? n42914 : n42940;
  assign n42942 = pi18 ? n33299 : n14115;
  assign n42943 = pi19 ? n1017 : n7036;
  assign n42944 = pi18 ? n139 : n42943;
  assign n42945 = pi17 ? n42942 : n42944;
  assign n42946 = pi16 ? n36216 : n42945;
  assign n42947 = pi21 ? n3668 : n139;
  assign n42948 = pi20 ? n992 : n42947;
  assign n42949 = pi19 ? n139 : n42948;
  assign n42950 = pi18 ? n42358 : n42949;
  assign n42951 = pi20 ? n5273 : n1026;
  assign n42952 = pi20 ? n6568 : n6172;
  assign n42953 = pi19 ? n42951 : n42952;
  assign n42954 = pi21 ? n2863 : n139;
  assign n42955 = pi20 ? n42954 : n1016;
  assign n42956 = pi19 ? n42955 : n7036;
  assign n42957 = pi18 ? n42953 : n42956;
  assign n42958 = pi17 ? n42950 : n42957;
  assign n42959 = pi16 ? n36216 : n42958;
  assign n42960 = pi15 ? n42946 : n42959;
  assign n42961 = pi19 ? n6373 : n28290;
  assign n42962 = pi20 ? n577 : n13527;
  assign n42963 = pi19 ? n42962 : n7725;
  assign n42964 = pi18 ? n42961 : n42963;
  assign n42965 = pi17 ? n38425 : n42964;
  assign n42966 = pi16 ? n36216 : n42965;
  assign n42967 = pi20 ? n25947 : n2092;
  assign n42968 = pi19 ? n7685 : n42967;
  assign n42969 = pi18 ? n42968 : n42963;
  assign n42970 = pi17 ? n39489 : n42969;
  assign n42971 = pi16 ? n36216 : n42970;
  assign n42972 = pi15 ? n42966 : n42971;
  assign n42973 = pi14 ? n42960 : n42972;
  assign n42974 = pi20 ? n233 : n6389;
  assign n42975 = pi19 ? n2095 : n42974;
  assign n42976 = pi20 ? n31760 : n25978;
  assign n42977 = pi19 ? n42976 : n3211;
  assign n42978 = pi18 ? n42975 : n42977;
  assign n42979 = pi17 ? n39489 : n42978;
  assign n42980 = pi16 ? n36216 : n42979;
  assign n42981 = pi21 ? n4891 : n2048;
  assign n42982 = pi20 ? n2049 : n42981;
  assign n42983 = pi19 ? n2095 : n42982;
  assign n42984 = pi19 ? n13337 : n3211;
  assign n42985 = pi18 ? n42983 : n42984;
  assign n42986 = pi17 ? n41813 : n42985;
  assign n42987 = pi16 ? n36216 : n42986;
  assign n42988 = pi15 ? n42980 : n42987;
  assign n42989 = pi20 ? n26846 : n21124;
  assign n42990 = pi19 ? n37 : n42989;
  assign n42991 = pi21 ? n1920 : n233;
  assign n42992 = pi20 ? n42991 : n233;
  assign n42993 = pi19 ? n42992 : n5831;
  assign n42994 = pi18 ? n42990 : n42993;
  assign n42995 = pi17 ? n41283 : n42994;
  assign n42996 = pi16 ? n36216 : n42995;
  assign n42997 = pi20 ? n33430 : n21124;
  assign n42998 = pi19 ? n37 : n42997;
  assign n42999 = pi19 ? n42992 : n10012;
  assign n43000 = pi18 ? n42998 : n42999;
  assign n43001 = pi17 ? n37372 : n43000;
  assign n43002 = pi16 ? n36216 : n43001;
  assign n43003 = pi15 ? n42996 : n43002;
  assign n43004 = pi14 ? n42988 : n43003;
  assign n43005 = pi13 ? n42973 : n43004;
  assign n43006 = pi12 ? n42941 : n43005;
  assign n43007 = pi21 ? n40908 : n20563;
  assign n43008 = pi20 ? n32 : n43007;
  assign n43009 = pi19 ? n32 : n43008;
  assign n43010 = pi21 ? n30868 : n20563;
  assign n43011 = pi20 ? n43010 : n20563;
  assign n43012 = pi19 ? n43011 : n20563;
  assign n43013 = pi18 ? n43009 : n43012;
  assign n43014 = pi17 ? n32 : n43013;
  assign n43015 = pi20 ? n2094 : n25965;
  assign n43016 = pi19 ? n43015 : n2654;
  assign n43017 = pi18 ? n41973 : n43016;
  assign n43018 = pi17 ? n37372 : n43017;
  assign n43019 = pi16 ? n43014 : n43018;
  assign n43020 = pi18 ? n34358 : n15082;
  assign n43021 = pi21 ? n335 : n25977;
  assign n43022 = pi20 ? n335 : n43021;
  assign n43023 = pi19 ? n43022 : n32;
  assign n43024 = pi18 ? n335 : n43023;
  assign n43025 = pi17 ? n43020 : n43024;
  assign n43026 = pi16 ? n43014 : n43025;
  assign n43027 = pi15 ? n43019 : n43026;
  assign n43028 = pi18 ? n34358 : n335;
  assign n43029 = pi21 ? n335 : n1389;
  assign n43030 = pi20 ? n335 : n43029;
  assign n43031 = pi19 ? n43030 : n32;
  assign n43032 = pi18 ? n335 : n43031;
  assign n43033 = pi17 ? n43028 : n43032;
  assign n43034 = pi16 ? n36216 : n43033;
  assign n43035 = pi20 ? n37 : n32055;
  assign n43036 = pi19 ? n43035 : n32;
  assign n43037 = pi18 ? n37 : n43036;
  assign n43038 = pi17 ? n37372 : n43037;
  assign n43039 = pi16 ? n36216 : n43038;
  assign n43040 = pi15 ? n43034 : n43039;
  assign n43041 = pi14 ? n43027 : n43040;
  assign n43042 = pi18 ? n35855 : n35637;
  assign n43043 = pi18 ? n363 : n32057;
  assign n43044 = pi17 ? n43042 : n43043;
  assign n43045 = pi16 ? n36216 : n43044;
  assign n43046 = pi21 ? n3392 : n2200;
  assign n43047 = pi20 ? n363 : n43046;
  assign n43048 = pi19 ? n43047 : n32;
  assign n43049 = pi18 ? n363 : n43048;
  assign n43050 = pi17 ? n43042 : n43049;
  assign n43051 = pi16 ? n36216 : n43050;
  assign n43052 = pi15 ? n43045 : n43051;
  assign n43053 = pi20 ? n19106 : n37;
  assign n43054 = pi19 ? n23917 : n43053;
  assign n43055 = pi20 ? n2107 : n2782;
  assign n43056 = pi19 ? n43055 : n32;
  assign n43057 = pi18 ? n43054 : n43056;
  assign n43058 = pi17 ? n39494 : n43057;
  assign n43059 = pi16 ? n36216 : n43058;
  assign n43060 = pi19 ? n37510 : n42062;
  assign n43061 = pi18 ? n35855 : n43060;
  assign n43062 = pi21 ? n3392 : n19958;
  assign n43063 = pi20 ? n43062 : n29421;
  assign n43064 = pi19 ? n363 : n43063;
  assign n43065 = pi20 ? n27520 : n41526;
  assign n43066 = pi19 ? n43065 : n32;
  assign n43067 = pi18 ? n43064 : n43066;
  assign n43068 = pi17 ? n43061 : n43067;
  assign n43069 = pi16 ? n36216 : n43068;
  assign n43070 = pi15 ? n43059 : n43069;
  assign n43071 = pi14 ? n43052 : n43070;
  assign n43072 = pi13 ? n43041 : n43071;
  assign n43073 = pi20 ? n16188 : n27520;
  assign n43074 = pi19 ? n35854 : n43073;
  assign n43075 = pi20 ? n22881 : n37;
  assign n43076 = pi19 ? n43075 : n36692;
  assign n43077 = pi18 ? n43074 : n43076;
  assign n43078 = pi20 ? n26890 : n10496;
  assign n43079 = pi19 ? n363 : n43078;
  assign n43080 = pi20 ? n21803 : n41526;
  assign n43081 = pi19 ? n43080 : n32;
  assign n43082 = pi18 ? n43079 : n43081;
  assign n43083 = pi17 ? n43077 : n43082;
  assign n43084 = pi16 ? n36216 : n43083;
  assign n43085 = pi22 ? n30867 : n112;
  assign n43086 = pi21 ? n43085 : n33758;
  assign n43087 = pi20 ? n43086 : n363;
  assign n43088 = pi19 ? n32314 : n43087;
  assign n43089 = pi22 ? n2160 : n363;
  assign n43090 = pi21 ? n10490 : n43089;
  assign n43091 = pi22 ? n7326 : n2160;
  assign n43092 = pi21 ? n7367 : n43091;
  assign n43093 = pi20 ? n43090 : n43092;
  assign n43094 = pi22 ? n363 : n112;
  assign n43095 = pi21 ? n43094 : n363;
  assign n43096 = pi21 ? n363 : n10488;
  assign n43097 = pi20 ? n43095 : n43096;
  assign n43098 = pi19 ? n43093 : n43097;
  assign n43099 = pi18 ? n43088 : n43098;
  assign n43100 = pi22 ? n5011 : n2160;
  assign n43101 = pi21 ? n363 : n43100;
  assign n43102 = pi21 ? n363 : n43089;
  assign n43103 = pi20 ? n43101 : n43102;
  assign n43104 = pi20 ? n685 : n363;
  assign n43105 = pi19 ? n43103 : n43104;
  assign n43106 = pi21 ? n43089 : n11208;
  assign n43107 = pi21 ? n2721 : n3523;
  assign n43108 = pi20 ? n43106 : n43107;
  assign n43109 = pi19 ? n43108 : n32;
  assign n43110 = pi18 ? n43105 : n43109;
  assign n43111 = pi17 ? n43099 : n43110;
  assign n43112 = pi16 ? n36216 : n43111;
  assign n43113 = pi15 ? n43084 : n43112;
  assign n43114 = pi18 ? n39318 : n99;
  assign n43115 = pi20 ? n30766 : n26891;
  assign n43116 = pi19 ? n43115 : n363;
  assign n43117 = pi20 ? n23150 : n38823;
  assign n43118 = pi19 ? n43117 : n32;
  assign n43119 = pi18 ? n43116 : n43118;
  assign n43120 = pi17 ? n43114 : n43119;
  assign n43121 = pi16 ? n42094 : n43120;
  assign n43122 = pi20 ? n36781 : n33792;
  assign n43123 = pi19 ? n43122 : n33792;
  assign n43124 = pi18 ? n37264 : n43123;
  assign n43125 = pi17 ? n32 : n43124;
  assign n43126 = pi19 ? n33792 : n139;
  assign n43127 = pi20 ? n139 : n685;
  assign n43128 = pi19 ? n139 : n43127;
  assign n43129 = pi18 ? n43126 : n43128;
  assign n43130 = pi20 ? n685 : n33780;
  assign n43131 = pi19 ? n43130 : n36772;
  assign n43132 = pi20 ? n685 : n14262;
  assign n43133 = pi19 ? n43132 : n32;
  assign n43134 = pi18 ? n43131 : n43133;
  assign n43135 = pi17 ? n43129 : n43134;
  assign n43136 = pi16 ? n43125 : n43135;
  assign n43137 = pi15 ? n43121 : n43136;
  assign n43138 = pi14 ? n43113 : n43137;
  assign n43139 = pi20 ? n36798 : n36659;
  assign n43140 = pi19 ? n43139 : n36659;
  assign n43141 = pi18 ? n41101 : n43140;
  assign n43142 = pi17 ? n32 : n43141;
  assign n43143 = pi19 ? n41579 : n41089;
  assign n43144 = pi22 ? n685 : n139;
  assign n43145 = pi21 ? n139 : n43144;
  assign n43146 = pi22 ? n139 : n685;
  assign n43147 = pi21 ? n139 : n43146;
  assign n43148 = pi20 ? n43145 : n43147;
  assign n43149 = pi19 ? n139 : n43148;
  assign n43150 = pi18 ? n43143 : n43149;
  assign n43151 = pi21 ? n43144 : n43146;
  assign n43152 = pi21 ? n685 : n43146;
  assign n43153 = pi20 ? n43151 : n43152;
  assign n43154 = pi20 ? n685 : n7829;
  assign n43155 = pi19 ? n43153 : n43154;
  assign n43156 = pi20 ? n27551 : n14723;
  assign n43157 = pi19 ? n43156 : n32;
  assign n43158 = pi18 ? n43155 : n43157;
  assign n43159 = pi17 ? n43150 : n43158;
  assign n43160 = pi16 ? n43142 : n43159;
  assign n43161 = pi22 ? n39996 : n36798;
  assign n43162 = pi21 ? n43161 : n36798;
  assign n43163 = pi20 ? n32 : n43162;
  assign n43164 = pi19 ? n32 : n43163;
  assign n43165 = pi18 ? n43164 : n43140;
  assign n43166 = pi17 ? n32 : n43165;
  assign n43167 = pi19 ? n41102 : n41107;
  assign n43168 = pi21 ? n335 : n1091;
  assign n43169 = pi20 ? n43168 : n316;
  assign n43170 = pi19 ? n43169 : n316;
  assign n43171 = pi18 ? n43167 : n43170;
  assign n43172 = pi20 ? n316 : n34537;
  assign n43173 = pi19 ? n316 : n43172;
  assign n43174 = pi20 ? n316 : n1010;
  assign n43175 = pi19 ? n43174 : n32;
  assign n43176 = pi18 ? n43173 : n43175;
  assign n43177 = pi17 ? n43171 : n43176;
  assign n43178 = pi16 ? n43166 : n43177;
  assign n43179 = pi15 ? n43160 : n43178;
  assign n43180 = pi21 ? n39997 : n36781;
  assign n43181 = pi20 ? n32 : n43180;
  assign n43182 = pi19 ? n32 : n43181;
  assign n43183 = pi19 ? n41135 : n36781;
  assign n43184 = pi18 ? n43182 : n43183;
  assign n43185 = pi17 ? n32 : n43184;
  assign n43186 = pi20 ? n36781 : n39975;
  assign n43187 = pi19 ? n43186 : n41125;
  assign n43188 = pi18 ? n43187 : n157;
  assign n43189 = pi17 ? n43188 : n42619;
  assign n43190 = pi16 ? n43185 : n43189;
  assign n43191 = pi23 ? n36782 : n36798;
  assign n43192 = pi22 ? n43191 : n36798;
  assign n43193 = pi21 ? n43192 : n36781;
  assign n43194 = pi20 ? n32 : n43193;
  assign n43195 = pi19 ? n32 : n43194;
  assign n43196 = pi18 ? n43195 : n43183;
  assign n43197 = pi17 ? n32 : n43196;
  assign n43198 = pi25 ? n203 : n32;
  assign n43199 = pi23 ? n36781 : n43198;
  assign n43200 = pi22 ? n36781 : n43199;
  assign n43201 = pi21 ? n43200 : n36798;
  assign n43202 = pi20 ? n36781 : n43201;
  assign n43203 = pi22 ? n36798 : n363;
  assign n43204 = pi21 ? n43203 : n157;
  assign n43205 = pi20 ? n43204 : n157;
  assign n43206 = pi19 ? n43202 : n43205;
  assign n43207 = pi18 ? n43206 : n157;
  assign n43208 = pi17 ? n43207 : n42619;
  assign n43209 = pi16 ? n43197 : n43208;
  assign n43210 = pi15 ? n43190 : n43209;
  assign n43211 = pi14 ? n43179 : n43210;
  assign n43212 = pi13 ? n43138 : n43211;
  assign n43213 = pi12 ? n43072 : n43212;
  assign n43214 = pi11 ? n43006 : n43213;
  assign n43215 = pi10 ? n42883 : n43214;
  assign n43216 = pi09 ? n42679 : n43215;
  assign n43217 = pi19 ? n32 : n40509;
  assign n43218 = pi18 ? n32 : n43217;
  assign n43219 = pi17 ? n32 : n43218;
  assign n43220 = pi16 ? n43219 : n42651;
  assign n43221 = pi15 ? n32 : n43220;
  assign n43222 = pi19 ? n32 : n40531;
  assign n43223 = pi18 ? n32 : n43222;
  assign n43224 = pi17 ? n32 : n43223;
  assign n43225 = pi16 ? n43224 : n42661;
  assign n43226 = pi19 ? n32 : n41707;
  assign n43227 = pi18 ? n32 : n43226;
  assign n43228 = pi17 ? n32 : n43227;
  assign n43229 = pi20 ? n37 : n3033;
  assign n43230 = pi20 ? n2973 : n21638;
  assign n43231 = pi19 ? n43229 : n43230;
  assign n43232 = pi20 ? n14524 : n2176;
  assign n43233 = pi22 ? n112 : n140;
  assign n43234 = pi21 ? n37 : n43233;
  assign n43235 = pi20 ? n43234 : n32;
  assign n43236 = pi19 ? n43232 : n43235;
  assign n43237 = pi18 ? n43231 : n43236;
  assign n43238 = pi17 ? n42663 : n43237;
  assign n43239 = pi16 ? n43228 : n43238;
  assign n43240 = pi15 ? n43225 : n43239;
  assign n43241 = pi14 ? n43221 : n43240;
  assign n43242 = pi13 ? n32 : n43241;
  assign n43243 = pi12 ? n32 : n43242;
  assign n43244 = pi11 ? n32 : n43243;
  assign n43245 = pi10 ? n32 : n43244;
  assign n43246 = pi20 ? n38997 : n20563;
  assign n43247 = pi19 ? n32 : n43246;
  assign n43248 = pi18 ? n32 : n43247;
  assign n43249 = pi17 ? n32 : n43248;
  assign n43250 = pi18 ? n20563 : n32288;
  assign n43251 = pi17 ? n43250 : n42684;
  assign n43252 = pi16 ? n43249 : n43251;
  assign n43253 = pi20 ? n31263 : n20563;
  assign n43254 = pi19 ? n32 : n43253;
  assign n43255 = pi18 ? n32 : n43254;
  assign n43256 = pi17 ? n32 : n43255;
  assign n43257 = pi18 ? n20563 : n38549;
  assign n43258 = pi17 ? n43257 : n42695;
  assign n43259 = pi16 ? n43256 : n43258;
  assign n43260 = pi15 ? n43252 : n43259;
  assign n43261 = pi19 ? n32 : n20563;
  assign n43262 = pi18 ? n32 : n43261;
  assign n43263 = pi17 ? n32 : n43262;
  assign n43264 = pi18 ? n20563 : n42358;
  assign n43265 = pi17 ? n43264 : n42706;
  assign n43266 = pi16 ? n43263 : n43265;
  assign n43267 = pi16 ? n41632 : n42714;
  assign n43268 = pi15 ? n43266 : n43267;
  assign n43269 = pi14 ? n43260 : n43268;
  assign n43270 = pi19 ? n139 : n14108;
  assign n43271 = pi18 ? n9766 : n43270;
  assign n43272 = pi17 ? n42196 : n43271;
  assign n43273 = pi16 ? n42689 : n43272;
  assign n43274 = pi19 ? n42722 : n14108;
  assign n43275 = pi18 ? n37 : n43274;
  assign n43276 = pi17 ? n41644 : n43275;
  assign n43277 = pi16 ? n41170 : n43276;
  assign n43278 = pi15 ? n43273 : n43277;
  assign n43279 = pi18 ? n20563 : n37029;
  assign n43280 = pi21 ? n335 : n13102;
  assign n43281 = pi20 ? n43280 : n32;
  assign n43282 = pi19 ? n577 : n43281;
  assign n43283 = pi18 ? n37 : n43282;
  assign n43284 = pi17 ? n43279 : n43283;
  assign n43285 = pi16 ? n41170 : n43284;
  assign n43286 = pi20 ? n28355 : n32;
  assign n43287 = pi19 ? n577 : n43286;
  assign n43288 = pi18 ? n37 : n43287;
  assign n43289 = pi17 ? n41672 : n43288;
  assign n43290 = pi16 ? n40025 : n43289;
  assign n43291 = pi15 ? n43285 : n43290;
  assign n43292 = pi14 ? n43278 : n43291;
  assign n43293 = pi13 ? n43269 : n43292;
  assign n43294 = pi18 ? n20563 : n35300;
  assign n43295 = pi19 ? n37 : n43286;
  assign n43296 = pi18 ? n37 : n43295;
  assign n43297 = pi17 ? n43294 : n43296;
  assign n43298 = pi16 ? n41183 : n43297;
  assign n43299 = pi21 ? n37 : n8260;
  assign n43300 = pi20 ? n43299 : n32;
  assign n43301 = pi19 ? n37 : n43300;
  assign n43302 = pi18 ? n37 : n43301;
  assign n43303 = pi17 ? n41178 : n43302;
  assign n43304 = pi16 ? n42241 : n43303;
  assign n43305 = pi15 ? n43298 : n43304;
  assign n43306 = pi21 ? n335 : n8260;
  assign n43307 = pi20 ? n43306 : n32;
  assign n43308 = pi19 ? n37 : n43307;
  assign n43309 = pi18 ? n37448 : n43308;
  assign n43310 = pi17 ? n42234 : n43309;
  assign n43311 = pi16 ? n41710 : n43310;
  assign n43312 = pi18 ? n20563 : n33976;
  assign n43313 = pi19 ? n7685 : n23550;
  assign n43314 = pi18 ? n37448 : n43313;
  assign n43315 = pi17 ? n43312 : n43314;
  assign n43316 = pi16 ? n38959 : n43315;
  assign n43317 = pi15 ? n43311 : n43316;
  assign n43318 = pi14 ? n43305 : n43317;
  assign n43319 = pi18 ? n34247 : n31300;
  assign n43320 = pi19 ? n37 : n23550;
  assign n43321 = pi18 ? n37 : n43320;
  assign n43322 = pi17 ? n43319 : n43321;
  assign n43323 = pi16 ? n40047 : n43322;
  assign n43324 = pi17 ? n40542 : n42767;
  assign n43325 = pi16 ? n39399 : n43324;
  assign n43326 = pi15 ? n43323 : n43325;
  assign n43327 = pi17 ? n40542 : n42774;
  assign n43328 = pi16 ? n38985 : n43327;
  assign n43329 = pi16 ? n40058 : n42780;
  assign n43330 = pi15 ? n43328 : n43329;
  assign n43331 = pi14 ? n43326 : n43330;
  assign n43332 = pi13 ? n43318 : n43331;
  assign n43333 = pi12 ? n43293 : n43332;
  assign n43334 = pi17 ? n40575 : n42789;
  assign n43335 = pi16 ? n37959 : n43334;
  assign n43336 = pi21 ? n37 : n35928;
  assign n43337 = pi20 ? n43336 : n32;
  assign n43338 = pi19 ? n37 : n43337;
  assign n43339 = pi18 ? n37 : n43338;
  assign n43340 = pi17 ? n39415 : n43339;
  assign n43341 = pi16 ? n37959 : n43340;
  assign n43342 = pi15 ? n43335 : n43341;
  assign n43343 = pi18 ? n40191 : n37;
  assign n43344 = pi23 ? n363 : n778;
  assign n43345 = pi22 ? n43344 : n32;
  assign n43346 = pi21 ? n37 : n43345;
  assign n43347 = pi20 ? n43346 : n32;
  assign n43348 = pi19 ? n37 : n43347;
  assign n43349 = pi18 ? n37 : n43348;
  assign n43350 = pi17 ? n43343 : n43349;
  assign n43351 = pi16 ? n37959 : n43350;
  assign n43352 = pi22 ? n21501 : n32;
  assign n43353 = pi21 ? n5015 : n43352;
  assign n43354 = pi20 ? n43353 : n32;
  assign n43355 = pi19 ? n37 : n43354;
  assign n43356 = pi18 ? n41009 : n43355;
  assign n43357 = pi17 ? n39433 : n43356;
  assign n43358 = pi16 ? n39001 : n43357;
  assign n43359 = pi15 ? n43351 : n43358;
  assign n43360 = pi14 ? n43342 : n43359;
  assign n43361 = pi21 ? n363 : n21387;
  assign n43362 = pi20 ? n43361 : n32;
  assign n43363 = pi19 ? n5029 : n43362;
  assign n43364 = pi18 ? n37 : n43363;
  assign n43365 = pi17 ? n41753 : n43364;
  assign n43366 = pi16 ? n37337 : n43365;
  assign n43367 = pi19 ? n20563 : n36886;
  assign n43368 = pi18 ? n43367 : n37;
  assign n43369 = pi19 ? n37 : n15198;
  assign n43370 = pi18 ? n37 : n43369;
  assign n43371 = pi17 ? n43368 : n43370;
  assign n43372 = pi16 ? n37337 : n43371;
  assign n43373 = pi15 ? n43366 : n43372;
  assign n43374 = pi17 ? n39440 : n43370;
  assign n43375 = pi16 ? n36163 : n43374;
  assign n43376 = pi19 ? n42822 : n15198;
  assign n43377 = pi18 ? n15175 : n43376;
  assign n43378 = pi17 ? n40062 : n43377;
  assign n43379 = pi16 ? n34860 : n43378;
  assign n43380 = pi15 ? n43375 : n43379;
  assign n43381 = pi14 ? n43373 : n43380;
  assign n43382 = pi13 ? n43360 : n43381;
  assign n43383 = pi17 ? n38992 : n42815;
  assign n43384 = pi16 ? n36216 : n43383;
  assign n43385 = pi21 ? n381 : n2320;
  assign n43386 = pi20 ? n43385 : n32;
  assign n43387 = pi19 ? n37 : n43386;
  assign n43388 = pi18 ? n37 : n43387;
  assign n43389 = pi17 ? n38992 : n43388;
  assign n43390 = pi16 ? n36216 : n43389;
  assign n43391 = pi15 ? n43384 : n43390;
  assign n43392 = pi17 ? n38992 : n42842;
  assign n43393 = pi16 ? n36216 : n43392;
  assign n43394 = pi19 ? n7746 : n42840;
  assign n43395 = pi18 ? n42845 : n43394;
  assign n43396 = pi17 ? n38992 : n43395;
  assign n43397 = pi16 ? n36216 : n43396;
  assign n43398 = pi15 ? n43393 : n43397;
  assign n43399 = pi14 ? n43391 : n43398;
  assign n43400 = pi18 ? n32872 : n21612;
  assign n43401 = pi21 ? n7429 : n928;
  assign n43402 = pi20 ? n43401 : n32;
  assign n43403 = pi19 ? n99 : n43402;
  assign n43404 = pi18 ? n99 : n43403;
  assign n43405 = pi17 ? n43400 : n43404;
  assign n43406 = pi16 ? n36216 : n43405;
  assign n43407 = pi18 ? n40314 : n21612;
  assign n43408 = pi21 ? n42859 : n928;
  assign n43409 = pi20 ? n43408 : n32;
  assign n43410 = pi19 ? n157 : n43409;
  assign n43411 = pi18 ? n17340 : n43410;
  assign n43412 = pi17 ? n43407 : n43411;
  assign n43413 = pi16 ? n36216 : n43412;
  assign n43414 = pi15 ? n43406 : n43413;
  assign n43415 = pi18 ? n33847 : n21612;
  assign n43416 = pi19 ? n157 : n14305;
  assign n43417 = pi18 ? n42869 : n43416;
  assign n43418 = pi17 ? n43415 : n43417;
  assign n43419 = pi16 ? n36216 : n43418;
  assign n43420 = pi18 ? n32275 : n42874;
  assign n43421 = pi18 ? n99 : n42380;
  assign n43422 = pi17 ? n43420 : n43421;
  assign n43423 = pi16 ? n36216 : n43422;
  assign n43424 = pi15 ? n43419 : n43423;
  assign n43425 = pi14 ? n43414 : n43424;
  assign n43426 = pi13 ? n43399 : n43425;
  assign n43427 = pi12 ? n43382 : n43426;
  assign n43428 = pi11 ? n43333 : n43427;
  assign n43429 = pi18 ? n33285 : n19774;
  assign n43430 = pi19 ? n42886 : n14305;
  assign n43431 = pi18 ? n99 : n43430;
  assign n43432 = pi17 ? n43429 : n43431;
  assign n43433 = pi16 ? n36216 : n43432;
  assign n43434 = pi21 ? n41400 : n2957;
  assign n43435 = pi20 ? n43434 : n14844;
  assign n43436 = pi19 ? n20563 : n43435;
  assign n43437 = pi18 ? n43436 : n99;
  assign n43438 = pi19 ? n38631 : n14305;
  assign n43439 = pi18 ? n42896 : n43438;
  assign n43440 = pi17 ? n43437 : n43439;
  assign n43441 = pi16 ? n36216 : n43440;
  assign n43442 = pi15 ? n43433 : n43441;
  assign n43443 = pi18 ? n34891 : n30851;
  assign n43444 = pi18 ? n42904 : n43438;
  assign n43445 = pi17 ? n43443 : n43444;
  assign n43446 = pi16 ? n36216 : n43445;
  assign n43447 = pi18 ? n34899 : n37;
  assign n43448 = pi19 ? n42908 : n14305;
  assign n43449 = pi18 ? n37 : n43448;
  assign n43450 = pi17 ? n43447 : n43449;
  assign n43451 = pi16 ? n36216 : n43450;
  assign n43452 = pi15 ? n43446 : n43451;
  assign n43453 = pi14 ? n43442 : n43452;
  assign n43454 = pi19 ? n42915 : n40811;
  assign n43455 = pi18 ? n43454 : n37;
  assign n43456 = pi17 ? n43455 : n42920;
  assign n43457 = pi16 ? n36216 : n43456;
  assign n43458 = pi18 ? n33285 : n15029;
  assign n43459 = pi21 ? n10410 : n32;
  assign n43460 = pi20 ? n43459 : n32;
  assign n43461 = pi19 ? n1017 : n43460;
  assign n43462 = pi18 ? n139 : n43461;
  assign n43463 = pi17 ? n43458 : n43462;
  assign n43464 = pi16 ? n36216 : n43463;
  assign n43465 = pi15 ? n43457 : n43464;
  assign n43466 = pi18 ? n33858 : n14115;
  assign n43467 = pi19 ? n1017 : n14328;
  assign n43468 = pi18 ? n139 : n43467;
  assign n43469 = pi17 ? n43466 : n43468;
  assign n43470 = pi16 ? n36216 : n43469;
  assign n43471 = pi18 ? n33858 : n9815;
  assign n43472 = pi20 ? n19549 : n32;
  assign n43473 = pi19 ? n1017 : n43472;
  assign n43474 = pi18 ? n139 : n43473;
  assign n43475 = pi17 ? n43471 : n43474;
  assign n43476 = pi16 ? n36216 : n43475;
  assign n43477 = pi15 ? n43470 : n43476;
  assign n43478 = pi14 ? n43465 : n43477;
  assign n43479 = pi13 ? n43453 : n43478;
  assign n43480 = pi19 ? n1017 : n4853;
  assign n43481 = pi18 ? n139 : n43480;
  assign n43482 = pi17 ? n42942 : n43481;
  assign n43483 = pi16 ? n36216 : n43482;
  assign n43484 = pi18 ? n38549 : n42949;
  assign n43485 = pi19 ? n42955 : n15447;
  assign n43486 = pi18 ? n42953 : n43485;
  assign n43487 = pi17 ? n43484 : n43486;
  assign n43488 = pi16 ? n36216 : n43487;
  assign n43489 = pi15 ? n43483 : n43488;
  assign n43490 = pi19 ? n42962 : n8296;
  assign n43491 = pi18 ? n42961 : n43490;
  assign n43492 = pi17 ? n40624 : n43491;
  assign n43493 = pi16 ? n36216 : n43492;
  assign n43494 = pi19 ? n42962 : n9483;
  assign n43495 = pi18 ? n42968 : n43494;
  assign n43496 = pi17 ? n40624 : n43495;
  assign n43497 = pi16 ? n36216 : n43496;
  assign n43498 = pi15 ? n43493 : n43497;
  assign n43499 = pi14 ? n43489 : n43498;
  assign n43500 = pi19 ? n42976 : n4009;
  assign n43501 = pi18 ? n42975 : n43500;
  assign n43502 = pi17 ? n40624 : n43501;
  assign n43503 = pi16 ? n36216 : n43502;
  assign n43504 = pi17 ? n38389 : n42985;
  assign n43505 = pi16 ? n36216 : n43504;
  assign n43506 = pi15 ? n43503 : n43505;
  assign n43507 = pi19 ? n42992 : n7050;
  assign n43508 = pi18 ? n42990 : n43507;
  assign n43509 = pi17 ? n42359 : n43508;
  assign n43510 = pi16 ? n36216 : n43509;
  assign n43511 = pi17 ? n41283 : n43000;
  assign n43512 = pi16 ? n36216 : n43511;
  assign n43513 = pi15 ? n43510 : n43512;
  assign n43514 = pi14 ? n43506 : n43513;
  assign n43515 = pi13 ? n43499 : n43514;
  assign n43516 = pi12 ? n43479 : n43515;
  assign n43517 = pi17 ? n41283 : n43017;
  assign n43518 = pi16 ? n43014 : n43517;
  assign n43519 = pi18 ? n32315 : n15082;
  assign n43520 = pi19 ? n43022 : n1823;
  assign n43521 = pi18 ? n335 : n43520;
  assign n43522 = pi17 ? n43519 : n43521;
  assign n43523 = pi16 ? n43014 : n43522;
  assign n43524 = pi15 ? n43518 : n43523;
  assign n43525 = pi18 ? n32315 : n335;
  assign n43526 = pi19 ? n12637 : n32;
  assign n43527 = pi18 ? n335 : n43526;
  assign n43528 = pi17 ? n43525 : n43527;
  assign n43529 = pi16 ? n36216 : n43528;
  assign n43530 = pi20 ? n37 : n28769;
  assign n43531 = pi19 ? n43530 : n32;
  assign n43532 = pi18 ? n37 : n43531;
  assign n43533 = pi17 ? n41283 : n43532;
  assign n43534 = pi16 ? n36216 : n43533;
  assign n43535 = pi15 ? n43529 : n43534;
  assign n43536 = pi14 ? n43524 : n43535;
  assign n43537 = pi18 ? n32877 : n35637;
  assign n43538 = pi20 ? n363 : n28769;
  assign n43539 = pi19 ? n43538 : n32;
  assign n43540 = pi18 ? n363 : n43539;
  assign n43541 = pi17 ? n43537 : n43540;
  assign n43542 = pi16 ? n36216 : n43541;
  assign n43543 = pi22 ? n40386 : n30195;
  assign n43544 = pi21 ? n20563 : n43543;
  assign n43545 = pi20 ? n20563 : n43544;
  assign n43546 = pi19 ? n43545 : n37;
  assign n43547 = pi18 ? n43546 : n35637;
  assign n43548 = pi21 ? n3392 : n2147;
  assign n43549 = pi20 ? n363 : n43548;
  assign n43550 = pi19 ? n43549 : n32;
  assign n43551 = pi18 ? n363 : n43550;
  assign n43552 = pi17 ? n43547 : n43551;
  assign n43553 = pi16 ? n36216 : n43552;
  assign n43554 = pi15 ? n43542 : n43553;
  assign n43555 = pi22 ? n36615 : n30195;
  assign n43556 = pi21 ? n20563 : n43555;
  assign n43557 = pi20 ? n20563 : n43556;
  assign n43558 = pi19 ? n43557 : n37;
  assign n43559 = pi18 ? n43558 : n37;
  assign n43560 = pi17 ? n43559 : n43057;
  assign n43561 = pi16 ? n36216 : n43560;
  assign n43562 = pi18 ? n43558 : n43060;
  assign n43563 = pi20 ? n27520 : n42552;
  assign n43564 = pi19 ? n43563 : n32;
  assign n43565 = pi18 ? n43064 : n43564;
  assign n43566 = pi17 ? n43562 : n43565;
  assign n43567 = pi16 ? n36216 : n43566;
  assign n43568 = pi15 ? n43561 : n43567;
  assign n43569 = pi14 ? n43554 : n43568;
  assign n43570 = pi13 ? n43536 : n43569;
  assign n43571 = pi23 ? n36659 : n20563;
  assign n43572 = pi22 ? n43571 : n30195;
  assign n43573 = pi21 ? n20563 : n43572;
  assign n43574 = pi20 ? n20563 : n43573;
  assign n43575 = pi19 ? n43574 : n43073;
  assign n43576 = pi18 ? n43575 : n43076;
  assign n43577 = pi17 ? n43576 : n43082;
  assign n43578 = pi16 ? n36216 : n43577;
  assign n43579 = pi23 ? n20563 : n99;
  assign n43580 = pi22 ? n20563 : n43579;
  assign n43581 = pi21 ? n43580 : n33758;
  assign n43582 = pi20 ? n43581 : n363;
  assign n43583 = pi19 ? n20563 : n43582;
  assign n43584 = pi21 ? n32817 : n31833;
  assign n43585 = pi22 ? n4543 : n4537;
  assign n43586 = pi21 ? n722 : n43585;
  assign n43587 = pi20 ? n43584 : n43586;
  assign n43588 = pi21 ? n363 : n31833;
  assign n43589 = pi20 ? n23150 : n43588;
  assign n43590 = pi19 ? n43587 : n43589;
  assign n43591 = pi18 ? n43583 : n43590;
  assign n43592 = pi21 ? n363 : n4538;
  assign n43593 = pi20 ? n43592 : n23162;
  assign n43594 = pi19 ? n43593 : n43104;
  assign n43595 = pi22 ? n4537 : n685;
  assign n43596 = pi21 ? n722 : n43595;
  assign n43597 = pi20 ? n43596 : n43107;
  assign n43598 = pi19 ? n43597 : n32;
  assign n43599 = pi18 ? n43594 : n43598;
  assign n43600 = pi17 ? n43591 : n43599;
  assign n43601 = pi16 ? n36216 : n43600;
  assign n43602 = pi15 ? n43578 : n43601;
  assign n43603 = pi20 ? n30868 : n40416;
  assign n43604 = pi19 ? n43603 : n99;
  assign n43605 = pi18 ? n43604 : n99;
  assign n43606 = pi17 ? n43605 : n43119;
  assign n43607 = pi16 ? n42094 : n43606;
  assign n43608 = pi21 ? n36763 : n139;
  assign n43609 = pi20 ? n43608 : n139;
  assign n43610 = pi19 ? n33792 : n43609;
  assign n43611 = pi18 ? n43610 : n43128;
  assign n43612 = pi20 ? n685 : n14698;
  assign n43613 = pi19 ? n43612 : n32;
  assign n43614 = pi18 ? n43131 : n43613;
  assign n43615 = pi17 ? n43611 : n43614;
  assign n43616 = pi16 ? n43125 : n43615;
  assign n43617 = pi15 ? n43607 : n43616;
  assign n43618 = pi14 ? n43602 : n43617;
  assign n43619 = pi20 ? n43608 : n34368;
  assign n43620 = pi19 ? n41579 : n43619;
  assign n43621 = pi18 ? n43620 : n43149;
  assign n43622 = pi20 ? n27551 : n37797;
  assign n43623 = pi19 ? n43622 : n32;
  assign n43624 = pi18 ? n43155 : n43623;
  assign n43625 = pi17 ? n43621 : n43624;
  assign n43626 = pi16 ? n43142 : n43625;
  assign n43627 = pi22 ? n36781 : n36801;
  assign n43628 = pi21 ? n43627 : n335;
  assign n43629 = pi20 ? n43628 : n335;
  assign n43630 = pi19 ? n41102 : n43629;
  assign n43631 = pi18 ? n43630 : n43170;
  assign n43632 = pi18 ? n43173 : n30497;
  assign n43633 = pi17 ? n43631 : n43632;
  assign n43634 = pi16 ? n43166 : n43633;
  assign n43635 = pi15 ? n43626 : n43634;
  assign n43636 = pi23 ? n36798 : n335;
  assign n43637 = pi22 ? n36781 : n43636;
  assign n43638 = pi21 ? n43637 : n157;
  assign n43639 = pi20 ? n43638 : n157;
  assign n43640 = pi19 ? n43186 : n43639;
  assign n43641 = pi18 ? n43640 : n157;
  assign n43642 = pi17 ? n43641 : n42619;
  assign n43643 = pi16 ? n43185 : n43642;
  assign n43644 = pi22 ? n36798 : n42171;
  assign n43645 = pi21 ? n43644 : n157;
  assign n43646 = pi20 ? n43645 : n157;
  assign n43647 = pi19 ? n43202 : n43646;
  assign n43648 = pi18 ? n43647 : n157;
  assign n43649 = pi21 ? n42627 : n1009;
  assign n43650 = pi20 ? n157 : n43649;
  assign n43651 = pi19 ? n43650 : n32;
  assign n43652 = pi18 ? n157 : n43651;
  assign n43653 = pi17 ? n43648 : n43652;
  assign n43654 = pi16 ? n43197 : n43653;
  assign n43655 = pi15 ? n43643 : n43654;
  assign n43656 = pi14 ? n43635 : n43655;
  assign n43657 = pi13 ? n43618 : n43656;
  assign n43658 = pi12 ? n43570 : n43657;
  assign n43659 = pi11 ? n43516 : n43658;
  assign n43660 = pi10 ? n43428 : n43659;
  assign n43661 = pi09 ? n43245 : n43660;
  assign n43662 = pi08 ? n43216 : n43661;
  assign n43663 = pi18 ? n32 : n31265;
  assign n43664 = pi17 ? n32 : n43663;
  assign n43665 = pi18 ? n20563 : n34258;
  assign n43666 = pi20 ? n27252 : n32;
  assign n43667 = pi19 ? n5121 : n43666;
  assign n43668 = pi18 ? n34262 : n43667;
  assign n43669 = pi17 ? n43665 : n43668;
  assign n43670 = pi16 ? n43664 : n43669;
  assign n43671 = pi15 ? n32 : n43670;
  assign n43672 = pi20 ? n32 : n20563;
  assign n43673 = pi19 ? n32 : n43672;
  assign n43674 = pi18 ? n32 : n43673;
  assign n43675 = pi17 ? n32 : n43674;
  assign n43676 = pi18 ? n20563 : n33245;
  assign n43677 = pi21 ? n99 : n19759;
  assign n43678 = pi20 ? n43677 : n32;
  assign n43679 = pi19 ? n99 : n43678;
  assign n43680 = pi18 ? n26408 : n43679;
  assign n43681 = pi17 ? n43676 : n43680;
  assign n43682 = pi16 ? n43675 : n43681;
  assign n43683 = pi19 ? n32 : n40496;
  assign n43684 = pi18 ? n32 : n43683;
  assign n43685 = pi17 ? n32 : n43684;
  assign n43686 = pi22 ? n37 : n18038;
  assign n43687 = pi21 ? n37 : n43686;
  assign n43688 = pi20 ? n43687 : n32;
  assign n43689 = pi19 ? n37 : n43688;
  assign n43690 = pi18 ? n37 : n43689;
  assign n43691 = pi17 ? n42657 : n43690;
  assign n43692 = pi16 ? n43685 : n43691;
  assign n43693 = pi15 ? n43682 : n43692;
  assign n43694 = pi14 ? n43671 : n43693;
  assign n43695 = pi13 ? n32 : n43694;
  assign n43696 = pi12 ? n32 : n43695;
  assign n43697 = pi11 ? n32 : n43696;
  assign n43698 = pi10 ? n32 : n43697;
  assign n43699 = pi21 ? n37 : n2027;
  assign n43700 = pi20 ? n43699 : n32;
  assign n43701 = pi19 ? n37 : n43700;
  assign n43702 = pi18 ? n37 : n43701;
  assign n43703 = pi17 ? n42657 : n43702;
  assign n43704 = pi16 ? n43685 : n43703;
  assign n43705 = pi22 ? n139 : n8198;
  assign n43706 = pi21 ? n37 : n43705;
  assign n43707 = pi20 ? n43706 : n32;
  assign n43708 = pi19 ? n37 : n43707;
  assign n43709 = pi18 ? n37 : n43708;
  assign n43710 = pi17 ? n42647 : n43709;
  assign n43711 = pi16 ? n42656 : n43710;
  assign n43712 = pi15 ? n43704 : n43711;
  assign n43713 = pi22 ? n139 : n1159;
  assign n43714 = pi21 ? n297 : n43713;
  assign n43715 = pi20 ? n43714 : n32;
  assign n43716 = pi19 ? n37 : n43715;
  assign n43717 = pi18 ? n37 : n43716;
  assign n43718 = pi17 ? n42663 : n43717;
  assign n43719 = pi16 ? n42682 : n43718;
  assign n43720 = pi22 ? n139 : n3146;
  assign n43721 = pi21 ? n139 : n43720;
  assign n43722 = pi20 ? n43721 : n32;
  assign n43723 = pi19 ? n3554 : n43722;
  assign n43724 = pi18 ? n18083 : n43723;
  assign n43725 = pi17 ? n42663 : n43724;
  assign n43726 = pi16 ? n42682 : n43725;
  assign n43727 = pi15 ? n43719 : n43726;
  assign n43728 = pi14 ? n43712 : n43727;
  assign n43729 = pi19 ? n139 : n43722;
  assign n43730 = pi18 ? n13193 : n43729;
  assign n43731 = pi17 ? n42657 : n43730;
  assign n43732 = pi16 ? n42195 : n43731;
  assign n43733 = pi22 ? n139 : n23361;
  assign n43734 = pi21 ? n139 : n43733;
  assign n43735 = pi20 ? n43734 : n32;
  assign n43736 = pi19 ? n3096 : n43735;
  assign n43737 = pi18 ? n13110 : n43736;
  assign n43738 = pi17 ? n42690 : n43737;
  assign n43739 = pi16 ? n41643 : n43738;
  assign n43740 = pi15 ? n43732 : n43739;
  assign n43741 = pi21 ? n335 : n43733;
  assign n43742 = pi20 ? n43741 : n32;
  assign n43743 = pi19 ? n577 : n43742;
  assign n43744 = pi18 ? n13110 : n43743;
  assign n43745 = pi17 ? n42690 : n43744;
  assign n43746 = pi16 ? n42701 : n43745;
  assign n43747 = pi23 ? n6960 : n32;
  assign n43748 = pi22 ? n335 : n43747;
  assign n43749 = pi21 ? n335 : n43748;
  assign n43750 = pi20 ? n43749 : n32;
  assign n43751 = pi19 ? n577 : n43750;
  assign n43752 = pi18 ? n14149 : n43751;
  assign n43753 = pi17 ? n42690 : n43752;
  assign n43754 = pi16 ? n42701 : n43753;
  assign n43755 = pi15 ? n43746 : n43754;
  assign n43756 = pi14 ? n43740 : n43755;
  assign n43757 = pi13 ? n43728 : n43756;
  assign n43758 = pi19 ? n37 : n43750;
  assign n43759 = pi18 ? n37 : n43758;
  assign n43760 = pi17 ? n42663 : n43759;
  assign n43761 = pi16 ? n41159 : n43760;
  assign n43762 = pi21 ? n37 : n20800;
  assign n43763 = pi20 ? n43762 : n32;
  assign n43764 = pi19 ? n37 : n43763;
  assign n43765 = pi18 ? n37 : n43764;
  assign n43766 = pi17 ? n42203 : n43765;
  assign n43767 = pi16 ? n41170 : n43766;
  assign n43768 = pi15 ? n43761 : n43767;
  assign n43769 = pi19 ? n6373 : n43286;
  assign n43770 = pi18 ? n37 : n43769;
  assign n43771 = pi17 ? n41644 : n43770;
  assign n43772 = pi16 ? n40512 : n43771;
  assign n43773 = pi19 ? n7685 : n24093;
  assign n43774 = pi18 ? n37 : n43773;
  assign n43775 = pi17 ? n41685 : n43774;
  assign n43776 = pi16 ? n39375 : n43775;
  assign n43777 = pi15 ? n43772 : n43776;
  assign n43778 = pi14 ? n43768 : n43777;
  assign n43779 = pi19 ? n37 : n24093;
  assign n43780 = pi18 ? n37 : n43779;
  assign n43781 = pi17 ? n41178 : n43780;
  assign n43782 = pi16 ? n40534 : n43781;
  assign n43783 = pi21 ? n569 : n665;
  assign n43784 = pi20 ? n43783 : n32;
  assign n43785 = pi19 ? n37 : n43784;
  assign n43786 = pi18 ? n37 : n43785;
  assign n43787 = pi17 ? n41178 : n43786;
  assign n43788 = pi16 ? n41710 : n43787;
  assign n43789 = pi15 ? n43782 : n43788;
  assign n43790 = pi19 ? n17224 : n24093;
  assign n43791 = pi18 ? n37 : n43790;
  assign n43792 = pi17 ? n41178 : n43791;
  assign n43793 = pi16 ? n39399 : n43792;
  assign n43794 = pi20 ? n1424 : n32;
  assign n43795 = pi19 ? n37 : n43794;
  assign n43796 = pi18 ? n37 : n43795;
  assign n43797 = pi17 ? n41178 : n43796;
  assign n43798 = pi16 ? n40552 : n43797;
  assign n43799 = pi15 ? n43793 : n43798;
  assign n43800 = pi14 ? n43789 : n43799;
  assign n43801 = pi13 ? n43778 : n43800;
  assign n43802 = pi12 ? n43757 : n43801;
  assign n43803 = pi20 ? n28420 : n32;
  assign n43804 = pi19 ? n37 : n43803;
  assign n43805 = pi18 ? n37 : n43804;
  assign n43806 = pi17 ? n40535 : n43805;
  assign n43807 = pi16 ? n37930 : n43806;
  assign n43808 = pi22 ? n3944 : n688;
  assign n43809 = pi21 ? n37 : n43808;
  assign n43810 = pi20 ? n43809 : n32;
  assign n43811 = pi19 ? n37 : n43810;
  assign n43812 = pi18 ? n37 : n43811;
  assign n43813 = pi17 ? n40535 : n43812;
  assign n43814 = pi16 ? n37930 : n43813;
  assign n43815 = pi15 ? n43807 : n43814;
  assign n43816 = pi22 ? n5061 : n688;
  assign n43817 = pi21 ? n37 : n43816;
  assign n43818 = pi20 ? n43817 : n32;
  assign n43819 = pi19 ? n37 : n43818;
  assign n43820 = pi18 ? n37 : n43819;
  assign n43821 = pi17 ? n41722 : n43820;
  assign n43822 = pi16 ? n37930 : n43821;
  assign n43823 = pi21 ? n5015 : n8486;
  assign n43824 = pi20 ? n43823 : n32;
  assign n43825 = pi19 ? n37 : n43824;
  assign n43826 = pi18 ? n41009 : n43825;
  assign n43827 = pi17 ? n41198 : n43826;
  assign n43828 = pi16 ? n38985 : n43827;
  assign n43829 = pi15 ? n43822 : n43828;
  assign n43830 = pi14 ? n43815 : n43829;
  assign n43831 = pi19 ? n6403 : n14693;
  assign n43832 = pi18 ? n37 : n43831;
  assign n43833 = pi17 ? n41192 : n43832;
  assign n43834 = pi16 ? n36871 : n43833;
  assign n43835 = pi17 ? n41198 : n43370;
  assign n43836 = pi16 ? n36871 : n43835;
  assign n43837 = pi15 ? n43834 : n43836;
  assign n43838 = pi20 ? n15173 : n5013;
  assign n43839 = pi19 ? n37 : n43838;
  assign n43840 = pi19 ? n18192 : n15198;
  assign n43841 = pi18 ? n43839 : n43840;
  assign n43842 = pi17 ? n41198 : n43841;
  assign n43843 = pi16 ? n37959 : n43842;
  assign n43844 = pi15 ? n43836 : n43843;
  assign n43845 = pi14 ? n43837 : n43844;
  assign n43846 = pi13 ? n43830 : n43845;
  assign n43847 = pi18 ? n38951 : n37;
  assign n43848 = pi17 ? n43847 : n43370;
  assign n43849 = pi16 ? n37324 : n43848;
  assign n43850 = pi17 ? n43343 : n43388;
  assign n43851 = pi16 ? n37324 : n43850;
  assign n43852 = pi15 ? n43849 : n43851;
  assign n43853 = pi21 ? n6433 : n2320;
  assign n43854 = pi20 ? n43853 : n32;
  assign n43855 = pi19 ? n37 : n43854;
  assign n43856 = pi18 ? n37 : n43855;
  assign n43857 = pi17 ? n43847 : n43856;
  assign n43858 = pi16 ? n39457 : n43857;
  assign n43859 = pi21 ? n777 : n882;
  assign n43860 = pi20 ? n43859 : n32;
  assign n43861 = pi19 ? n99 : n43860;
  assign n43862 = pi18 ? n19774 : n43861;
  assign n43863 = pi17 ? n40584 : n43862;
  assign n43864 = pi16 ? n36163 : n43863;
  assign n43865 = pi15 ? n43858 : n43864;
  assign n43866 = pi14 ? n43852 : n43865;
  assign n43867 = pi18 ? n33245 : n19774;
  assign n43868 = pi17 ? n43867 : n43404;
  assign n43869 = pi16 ? n34860 : n43868;
  assign n43870 = pi18 ? n34258 : n21612;
  assign n43871 = pi19 ? n157 : n43402;
  assign n43872 = pi18 ? n17340 : n43871;
  assign n43873 = pi17 ? n43870 : n43872;
  assign n43874 = pi16 ? n34860 : n43873;
  assign n43875 = pi15 ? n43869 : n43874;
  assign n43876 = pi18 ? n33245 : n21612;
  assign n43877 = pi21 ? n164 : n3013;
  assign n43878 = pi20 ? n43877 : n787;
  assign n43879 = pi19 ? n43878 : n6532;
  assign n43880 = pi18 ? n43879 : n43416;
  assign n43881 = pi17 ? n43876 : n43880;
  assign n43882 = pi16 ? n35765 : n43881;
  assign n43883 = pi20 ? n3039 : n14844;
  assign n43884 = pi19 ? n43883 : n99;
  assign n43885 = pi18 ? n35799 : n43884;
  assign n43886 = pi20 ? n169 : n776;
  assign n43887 = pi19 ? n99 : n43886;
  assign n43888 = pi21 ? n3562 : n2678;
  assign n43889 = pi20 ? n43888 : n32;
  assign n43890 = pi19 ? n157 : n43889;
  assign n43891 = pi18 ? n43887 : n43890;
  assign n43892 = pi17 ? n43885 : n43891;
  assign n43893 = pi16 ? n36216 : n43892;
  assign n43894 = pi15 ? n43882 : n43893;
  assign n43895 = pi14 ? n43875 : n43894;
  assign n43896 = pi13 ? n43866 : n43895;
  assign n43897 = pi12 ? n43846 : n43896;
  assign n43898 = pi11 ? n43802 : n43897;
  assign n43899 = pi18 ? n34295 : n19774;
  assign n43900 = pi22 ? n3961 : n99;
  assign n43901 = pi21 ? n43900 : n99;
  assign n43902 = pi20 ? n43901 : n19201;
  assign n43903 = pi19 ? n99 : n43902;
  assign n43904 = pi20 ? n3759 : n204;
  assign n43905 = pi21 ? n316 : n2700;
  assign n43906 = pi20 ? n43905 : n32;
  assign n43907 = pi19 ? n43904 : n43906;
  assign n43908 = pi18 ? n43903 : n43907;
  assign n43909 = pi17 ? n43899 : n43908;
  assign n43910 = pi16 ? n36216 : n43909;
  assign n43911 = pi20 ? n39192 : n37;
  assign n43912 = pi19 ? n20563 : n43911;
  assign n43913 = pi18 ? n43912 : n21612;
  assign n43914 = pi21 ? n17375 : n99;
  assign n43915 = pi20 ? n99 : n43914;
  assign n43916 = pi19 ? n99 : n43915;
  assign n43917 = pi19 ? n38631 : n43906;
  assign n43918 = pi18 ? n43916 : n43917;
  assign n43919 = pi17 ? n43913 : n43918;
  assign n43920 = pi16 ? n36216 : n43919;
  assign n43921 = pi15 ? n43910 : n43920;
  assign n43922 = pi18 ? n34295 : n30851;
  assign n43923 = pi18 ? n21612 : n43438;
  assign n43924 = pi17 ? n43922 : n43923;
  assign n43925 = pi16 ? n36216 : n43924;
  assign n43926 = pi20 ? n947 : n3096;
  assign n43927 = pi19 ? n37 : n43926;
  assign n43928 = pi20 ? n13147 : n204;
  assign n43929 = pi19 ? n43928 : n15383;
  assign n43930 = pi18 ? n43927 : n43929;
  assign n43931 = pi17 ? n41753 : n43930;
  assign n43932 = pi16 ? n36216 : n43931;
  assign n43933 = pi15 ? n43925 : n43932;
  assign n43934 = pi14 ? n43921 : n43933;
  assign n43935 = pi21 ? n20563 : n39801;
  assign n43936 = pi20 ? n43935 : n39183;
  assign n43937 = pi19 ? n20563 : n43936;
  assign n43938 = pi18 ? n43937 : n37;
  assign n43939 = pi21 ? n1711 : n37;
  assign n43940 = pi20 ? n43939 : n204;
  assign n43941 = pi19 ? n43940 : n14754;
  assign n43942 = pi18 ? n10652 : n43941;
  assign n43943 = pi17 ? n43938 : n43942;
  assign n43944 = pi16 ? n36216 : n43943;
  assign n43945 = pi22 ? n39190 : n30195;
  assign n43946 = pi21 ? n20563 : n43945;
  assign n43947 = pi20 ? n43946 : n39183;
  assign n43948 = pi19 ? n20563 : n43947;
  assign n43949 = pi18 ? n43948 : n15029;
  assign n43950 = pi19 ? n12589 : n14754;
  assign n43951 = pi18 ? n139 : n43950;
  assign n43952 = pi17 ? n43949 : n43951;
  assign n43953 = pi16 ? n36216 : n43952;
  assign n43954 = pi15 ? n43944 : n43953;
  assign n43955 = pi18 ? n39447 : n14115;
  assign n43956 = pi22 ? n204 : n19327;
  assign n43957 = pi21 ? n43956 : n32;
  assign n43958 = pi20 ? n43957 : n32;
  assign n43959 = pi19 ? n12589 : n43958;
  assign n43960 = pi18 ? n139 : n43959;
  assign n43961 = pi17 ? n43955 : n43960;
  assign n43962 = pi16 ? n36216 : n43961;
  assign n43963 = pi18 ? n39447 : n9796;
  assign n43964 = pi19 ? n12589 : n43472;
  assign n43965 = pi18 ? n139 : n43964;
  assign n43966 = pi17 ? n43963 : n43965;
  assign n43967 = pi16 ? n36216 : n43966;
  assign n43968 = pi15 ? n43962 : n43967;
  assign n43969 = pi14 ? n43954 : n43968;
  assign n43970 = pi13 ? n43934 : n43969;
  assign n43971 = pi19 ? n31363 : n9795;
  assign n43972 = pi18 ? n33260 : n43971;
  assign n43973 = pi17 ? n43972 : n43965;
  assign n43974 = pi16 ? n36216 : n43973;
  assign n43975 = pi19 ? n139 : n26471;
  assign n43976 = pi18 ? n33260 : n43975;
  assign n43977 = pi22 ? n37 : n918;
  assign n43978 = pi21 ? n139 : n43977;
  assign n43979 = pi20 ? n43978 : n947;
  assign n43980 = pi19 ? n139 : n43979;
  assign n43981 = pi23 ? n233 : n4882;
  assign n43982 = pi22 ? n43981 : n688;
  assign n43983 = pi21 ? n43982 : n32;
  assign n43984 = pi20 ? n43983 : n32;
  assign n43985 = pi19 ? n9769 : n43984;
  assign n43986 = pi18 ? n43980 : n43985;
  assign n43987 = pi17 ? n43976 : n43986;
  assign n43988 = pi16 ? n36216 : n43987;
  assign n43989 = pi15 ? n43974 : n43988;
  assign n43990 = pi19 ? n6373 : n37;
  assign n43991 = pi18 ? n43990 : n43490;
  assign n43992 = pi17 ? n38992 : n43991;
  assign n43993 = pi16 ? n36216 : n43992;
  assign n43994 = pi20 ? n8927 : n3410;
  assign n43995 = pi19 ? n7685 : n43994;
  assign n43996 = pi20 ? n30674 : n13527;
  assign n43997 = pi19 ? n43996 : n9483;
  assign n43998 = pi18 ? n43995 : n43997;
  assign n43999 = pi17 ? n38992 : n43998;
  assign n44000 = pi16 ? n36216 : n43999;
  assign n44001 = pi15 ? n43993 : n44000;
  assign n44002 = pi14 ? n43989 : n44001;
  assign n44003 = pi20 ? n233 : n26846;
  assign n44004 = pi19 ? n2095 : n44003;
  assign n44005 = pi21 ? n3409 : n335;
  assign n44006 = pi20 ? n44005 : n15465;
  assign n44007 = pi19 ? n44006 : n4009;
  assign n44008 = pi18 ? n44004 : n44007;
  assign n44009 = pi17 ? n38992 : n44008;
  assign n44010 = pi16 ? n36216 : n44009;
  assign n44011 = pi20 ? n5023 : n7705;
  assign n44012 = pi19 ? n2095 : n44011;
  assign n44013 = pi20 ? n21160 : n233;
  assign n44014 = pi19 ? n44013 : n3211;
  assign n44015 = pi18 ? n44012 : n44014;
  assign n44016 = pi17 ? n38369 : n44015;
  assign n44017 = pi16 ? n36216 : n44016;
  assign n44018 = pi15 ? n44010 : n44017;
  assign n44019 = pi21 ? n37 : n6361;
  assign n44020 = pi20 ? n44019 : n37;
  assign n44021 = pi19 ? n37 : n44020;
  assign n44022 = pi21 ? n24208 : n32;
  assign n44023 = pi20 ? n44022 : n32;
  assign n44024 = pi19 ? n6391 : n44023;
  assign n44025 = pi18 ? n44021 : n44024;
  assign n44026 = pi17 ? n38369 : n44025;
  assign n44027 = pi16 ? n36216 : n44026;
  assign n44028 = pi23 ? n2120 : n316;
  assign n44029 = pi22 ? n44028 : n32;
  assign n44030 = pi21 ? n44029 : n32;
  assign n44031 = pi20 ? n44030 : n32;
  assign n44032 = pi19 ? n6391 : n44031;
  assign n44033 = pi18 ? n44021 : n44032;
  assign n44034 = pi17 ? n39481 : n44033;
  assign n44035 = pi16 ? n36216 : n44034;
  assign n44036 = pi15 ? n44027 : n44035;
  assign n44037 = pi14 ? n44018 : n44036;
  assign n44038 = pi13 ? n44002 : n44037;
  assign n44039 = pi12 ? n43970 : n44038;
  assign n44040 = pi19 ? n6391 : n7833;
  assign n44041 = pi18 ? n41973 : n44040;
  assign n44042 = pi17 ? n42326 : n44041;
  assign n44043 = pi16 ? n43014 : n44042;
  assign n44044 = pi18 ? n32288 : n15082;
  assign n44045 = pi19 ? n13528 : n1823;
  assign n44046 = pi18 ? n335 : n44045;
  assign n44047 = pi17 ? n44044 : n44046;
  assign n44048 = pi16 ? n36216 : n44047;
  assign n44049 = pi15 ? n44043 : n44048;
  assign n44050 = pi18 ? n32288 : n335;
  assign n44051 = pi21 ? n335 : n18411;
  assign n44052 = pi20 ? n335 : n44051;
  assign n44053 = pi19 ? n44052 : n32;
  assign n44054 = pi18 ? n335 : n44053;
  assign n44055 = pi17 ? n44050 : n44054;
  assign n44056 = pi16 ? n36216 : n44055;
  assign n44057 = pi20 ? n40987 : n37;
  assign n44058 = pi19 ? n20563 : n44057;
  assign n44059 = pi18 ? n44058 : n37;
  assign n44060 = pi20 ? n37 : n25199;
  assign n44061 = pi19 ? n44060 : n32;
  assign n44062 = pi18 ? n37 : n44061;
  assign n44063 = pi17 ? n44059 : n44062;
  assign n44064 = pi16 ? n36216 : n44063;
  assign n44065 = pi15 ? n44056 : n44064;
  assign n44066 = pi14 ? n44049 : n44065;
  assign n44067 = pi20 ? n35316 : n14530;
  assign n44068 = pi19 ? n20563 : n44067;
  assign n44069 = pi18 ? n44068 : n35637;
  assign n44070 = pi17 ? n44069 : n43540;
  assign n44071 = pi16 ? n36216 : n44070;
  assign n44072 = pi22 ? n14245 : n363;
  assign n44073 = pi21 ? n44072 : n5113;
  assign n44074 = pi20 ? n363 : n44073;
  assign n44075 = pi19 ? n44074 : n32;
  assign n44076 = pi18 ? n363 : n44075;
  assign n44077 = pi17 ? n44069 : n44076;
  assign n44078 = pi16 ? n36216 : n44077;
  assign n44079 = pi15 ? n44071 : n44078;
  assign n44080 = pi20 ? n35316 : n13179;
  assign n44081 = pi19 ? n20563 : n44080;
  assign n44082 = pi18 ? n44081 : n37;
  assign n44083 = pi20 ? n2107 : n37;
  assign n44084 = pi19 ? n23917 : n44083;
  assign n44085 = pi20 ? n2107 : n42552;
  assign n44086 = pi19 ? n44085 : n32;
  assign n44087 = pi18 ? n44084 : n44086;
  assign n44088 = pi17 ? n44082 : n44087;
  assign n44089 = pi16 ? n36216 : n44088;
  assign n44090 = pi18 ? n44081 : n42063;
  assign n44091 = pi20 ? n29741 : n685;
  assign n44092 = pi19 ? n363 : n44091;
  assign n44093 = pi20 ? n18194 : n42552;
  assign n44094 = pi19 ? n44093 : n32;
  assign n44095 = pi18 ? n44092 : n44094;
  assign n44096 = pi17 ? n44090 : n44095;
  assign n44097 = pi16 ? n36216 : n44096;
  assign n44098 = pi15 ? n44089 : n44097;
  assign n44099 = pi14 ? n44079 : n44098;
  assign n44100 = pi13 ? n44066 : n44099;
  assign n44101 = pi22 ? n36781 : n37;
  assign n44102 = pi21 ? n20563 : n44101;
  assign n44103 = pi21 ? n574 : n5015;
  assign n44104 = pi20 ? n44102 : n44103;
  assign n44105 = pi19 ? n20563 : n44104;
  assign n44106 = pi18 ? n44105 : n43076;
  assign n44107 = pi20 ? n685 : n29741;
  assign n44108 = pi19 ? n363 : n44107;
  assign n44109 = pi20 ? n26891 : n42552;
  assign n44110 = pi19 ? n44109 : n32;
  assign n44111 = pi18 ? n44108 : n44110;
  assign n44112 = pi17 ? n44106 : n44111;
  assign n44113 = pi16 ? n36216 : n44112;
  assign n44114 = pi22 ? n36781 : n99;
  assign n44115 = pi21 ? n30868 : n44114;
  assign n44116 = pi22 ? n22116 : n99;
  assign n44117 = pi21 ? n44116 : n22549;
  assign n44118 = pi20 ? n44115 : n44117;
  assign n44119 = pi19 ? n30868 : n44118;
  assign n44120 = pi20 ? n23162 : n29686;
  assign n44121 = pi19 ? n44120 : n363;
  assign n44122 = pi18 ? n44119 : n44121;
  assign n44123 = pi19 ? n363 : n43104;
  assign n44124 = pi22 ? n363 : n3944;
  assign n44125 = pi21 ? n44124 : n5178;
  assign n44126 = pi20 ? n23162 : n44125;
  assign n44127 = pi19 ? n44126 : n32;
  assign n44128 = pi18 ? n44123 : n44127;
  assign n44129 = pi17 ? n44122 : n44128;
  assign n44130 = pi16 ? n42094 : n44129;
  assign n44131 = pi15 ? n44113 : n44130;
  assign n44132 = pi18 ? n39917 : n99;
  assign n44133 = pi20 ? n363 : n38823;
  assign n44134 = pi19 ? n44133 : n32;
  assign n44135 = pi18 ? n43116 : n44134;
  assign n44136 = pi17 ? n44132 : n44135;
  assign n44137 = pi16 ? n42094 : n44136;
  assign n44138 = pi21 ? n36784 : n36781;
  assign n44139 = pi20 ? n32 : n44138;
  assign n44140 = pi19 ? n32 : n44139;
  assign n44141 = pi18 ? n44140 : n43123;
  assign n44142 = pi17 ? n32 : n44141;
  assign n44143 = pi22 ? n33792 : n40428;
  assign n44144 = pi21 ? n33792 : n44143;
  assign n44145 = pi20 ? n44144 : n139;
  assign n44146 = pi19 ? n33792 : n44145;
  assign n44147 = pi18 ? n44146 : n43128;
  assign n44148 = pi21 ? n43144 : n685;
  assign n44149 = pi21 ? n43146 : n685;
  assign n44150 = pi20 ? n44148 : n44149;
  assign n44151 = pi19 ? n685 : n44150;
  assign n44152 = pi20 ? n685 : n38823;
  assign n44153 = pi19 ? n44152 : n32;
  assign n44154 = pi18 ? n44151 : n44153;
  assign n44155 = pi17 ? n44147 : n44154;
  assign n44156 = pi16 ? n44142 : n44155;
  assign n44157 = pi15 ? n44137 : n44156;
  assign n44158 = pi14 ? n44131 : n44157;
  assign n44159 = pi18 ? n41603 : n43140;
  assign n44160 = pi17 ? n32 : n44159;
  assign n44161 = pi20 ? n44144 : n34368;
  assign n44162 = pi19 ? n41579 : n44161;
  assign n44163 = pi23 ? n685 : n139;
  assign n44164 = pi22 ? n139 : n44163;
  assign n44165 = pi21 ? n44164 : n139;
  assign n44166 = pi20 ? n139 : n44165;
  assign n44167 = pi19 ? n139 : n44166;
  assign n44168 = pi18 ? n44162 : n44167;
  assign n44169 = pi22 ? n3472 : n139;
  assign n44170 = pi21 ? n258 : n44169;
  assign n44171 = pi22 ? n3472 : n157;
  assign n44172 = pi21 ? n258 : n44171;
  assign n44173 = pi20 ? n44170 : n44172;
  assign n44174 = pi21 ? n43144 : n157;
  assign n44175 = pi21 ? n20460 : n248;
  assign n44176 = pi20 ? n44174 : n44175;
  assign n44177 = pi19 ? n44173 : n44176;
  assign n44178 = pi20 ? n873 : n14713;
  assign n44179 = pi19 ? n44178 : n32;
  assign n44180 = pi18 ? n44177 : n44179;
  assign n44181 = pi17 ? n44168 : n44180;
  assign n44182 = pi16 ? n44160 : n44181;
  assign n44183 = pi20 ? n42147 : n41106;
  assign n44184 = pi19 ? n41102 : n44183;
  assign n44185 = pi20 ? n335 : n3707;
  assign n44186 = pi19 ? n44185 : n316;
  assign n44187 = pi18 ? n44184 : n44186;
  assign n44188 = pi17 ? n44187 : n43632;
  assign n44189 = pi16 ? n44160 : n44188;
  assign n44190 = pi15 ? n44182 : n44189;
  assign n44191 = pi21 ? n42146 : n36798;
  assign n44192 = pi22 ? n36798 : n335;
  assign n44193 = pi21 ? n44192 : n157;
  assign n44194 = pi20 ? n44191 : n44193;
  assign n44195 = pi19 ? n43186 : n44194;
  assign n44196 = pi18 ? n44195 : n157;
  assign n44197 = pi20 ? n157 : n27095;
  assign n44198 = pi19 ? n44197 : n32;
  assign n44199 = pi18 ? n157 : n44198;
  assign n44200 = pi17 ? n44196 : n44199;
  assign n44201 = pi16 ? n43185 : n44200;
  assign n44202 = pi22 ? n36783 : n36798;
  assign n44203 = pi21 ? n44202 : n36781;
  assign n44204 = pi20 ? n32 : n44203;
  assign n44205 = pi19 ? n32 : n44204;
  assign n44206 = pi18 ? n44205 : n43183;
  assign n44207 = pi17 ? n32 : n44206;
  assign n44208 = pi20 ? n36781 : n42170;
  assign n44209 = pi21 ? n38901 : n36798;
  assign n44210 = pi20 ? n44209 : n43204;
  assign n44211 = pi19 ? n44208 : n44210;
  assign n44212 = pi18 ? n44211 : n157;
  assign n44213 = pi17 ? n44212 : n43652;
  assign n44214 = pi16 ? n44207 : n44213;
  assign n44215 = pi15 ? n44201 : n44214;
  assign n44216 = pi14 ? n44190 : n44215;
  assign n44217 = pi13 ? n44158 : n44216;
  assign n44218 = pi12 ? n44100 : n44217;
  assign n44219 = pi11 ? n44039 : n44218;
  assign n44220 = pi10 ? n43898 : n44219;
  assign n44221 = pi09 ? n43698 : n44220;
  assign n44222 = pi18 ? n32 : n37335;
  assign n44223 = pi17 ? n32 : n44222;
  assign n44224 = pi16 ? n44223 : n43669;
  assign n44225 = pi15 ? n32 : n44224;
  assign n44226 = pi18 ? n32 : n30119;
  assign n44227 = pi17 ? n32 : n44226;
  assign n44228 = pi19 ? n99 : n43666;
  assign n44229 = pi18 ? n26408 : n44228;
  assign n44230 = pi17 ? n43676 : n44229;
  assign n44231 = pi16 ? n44227 : n44230;
  assign n44232 = pi16 ? n44227 : n43691;
  assign n44233 = pi15 ? n44231 : n44232;
  assign n44234 = pi14 ? n44225 : n44233;
  assign n44235 = pi13 ? n32 : n44234;
  assign n44236 = pi12 ? n32 : n44235;
  assign n44237 = pi11 ? n32 : n44236;
  assign n44238 = pi10 ? n32 : n44237;
  assign n44239 = pi22 ? n37 : n8174;
  assign n44240 = pi21 ? n37 : n44239;
  assign n44241 = pi20 ? n44240 : n32;
  assign n44242 = pi19 ? n37 : n44241;
  assign n44243 = pi18 ? n37 : n44242;
  assign n44244 = pi17 ? n42657 : n44243;
  assign n44245 = pi16 ? n43664 : n44244;
  assign n44246 = pi19 ? n32 : n39372;
  assign n44247 = pi18 ? n32 : n44246;
  assign n44248 = pi17 ? n32 : n44247;
  assign n44249 = pi18 ? n20563 : n33828;
  assign n44250 = pi23 ? n139 : n5630;
  assign n44251 = pi22 ? n139 : n44250;
  assign n44252 = pi21 ? n37 : n44251;
  assign n44253 = pi20 ? n44252 : n32;
  assign n44254 = pi19 ? n37 : n44253;
  assign n44255 = pi18 ? n37 : n44254;
  assign n44256 = pi17 ? n44249 : n44255;
  assign n44257 = pi16 ? n44248 : n44256;
  assign n44258 = pi15 ? n44245 : n44257;
  assign n44259 = pi21 ? n297 : n28259;
  assign n44260 = pi20 ? n44259 : n32;
  assign n44261 = pi19 ? n37 : n44260;
  assign n44262 = pi18 ? n37 : n44261;
  assign n44263 = pi17 ? n42663 : n44262;
  assign n44264 = pi16 ? n43228 : n44263;
  assign n44265 = pi21 ? n139 : n12243;
  assign n44266 = pi20 ? n44265 : n32;
  assign n44267 = pi19 ? n3554 : n44266;
  assign n44268 = pi18 ? n18083 : n44267;
  assign n44269 = pi17 ? n43250 : n44268;
  assign n44270 = pi16 ? n43249 : n44269;
  assign n44271 = pi15 ? n44264 : n44270;
  assign n44272 = pi14 ? n44258 : n44271;
  assign n44273 = pi19 ? n32 : n38947;
  assign n44274 = pi18 ? n32 : n44273;
  assign n44275 = pi17 ? n32 : n44274;
  assign n44276 = pi19 ? n139 : n15621;
  assign n44277 = pi18 ? n13193 : n44276;
  assign n44278 = pi17 ? n42657 : n44277;
  assign n44279 = pi16 ? n44275 : n44278;
  assign n44280 = pi18 ? n20563 : n33858;
  assign n44281 = pi19 ? n3096 : n15621;
  assign n44282 = pi18 ? n13110 : n44281;
  assign n44283 = pi17 ? n44280 : n44282;
  assign n44284 = pi16 ? n42202 : n44283;
  assign n44285 = pi15 ? n44279 : n44284;
  assign n44286 = pi21 ? n335 : n20300;
  assign n44287 = pi20 ? n44286 : n32;
  assign n44288 = pi19 ? n577 : n44287;
  assign n44289 = pi18 ? n13110 : n44288;
  assign n44290 = pi17 ? n42690 : n44289;
  assign n44291 = pi16 ? n43263 : n44290;
  assign n44292 = pi20 ? n29288 : n32;
  assign n44293 = pi19 ? n577 : n44292;
  assign n44294 = pi18 ? n14149 : n44293;
  assign n44295 = pi17 ? n42690 : n44294;
  assign n44296 = pi16 ? n41632 : n44295;
  assign n44297 = pi15 ? n44291 : n44296;
  assign n44298 = pi14 ? n44285 : n44297;
  assign n44299 = pi13 ? n44272 : n44298;
  assign n44300 = pi19 ? n37 : n44292;
  assign n44301 = pi18 ? n37 : n44300;
  assign n44302 = pi17 ? n42663 : n44301;
  assign n44303 = pi16 ? n42689 : n44302;
  assign n44304 = pi21 ? n37 : n7658;
  assign n44305 = pi20 ? n44304 : n32;
  assign n44306 = pi19 ? n37 : n44305;
  assign n44307 = pi18 ? n37 : n44306;
  assign n44308 = pi17 ? n43264 : n44307;
  assign n44309 = pi16 ? n41170 : n44308;
  assign n44310 = pi15 ? n44303 : n44309;
  assign n44311 = pi21 ? n335 : n7658;
  assign n44312 = pi20 ? n44311 : n32;
  assign n44313 = pi19 ? n6373 : n44312;
  assign n44314 = pi18 ? n37 : n44313;
  assign n44315 = pi17 ? n42203 : n44314;
  assign n44316 = pi16 ? n41170 : n44315;
  assign n44317 = pi20 ? n11857 : n32;
  assign n44318 = pi19 ? n7685 : n44317;
  assign n44319 = pi18 ? n37 : n44318;
  assign n44320 = pi17 ? n43294 : n44319;
  assign n44321 = pi16 ? n40025 : n44320;
  assign n44322 = pi15 ? n44316 : n44321;
  assign n44323 = pi14 ? n44310 : n44322;
  assign n44324 = pi16 ? n41183 : n43781;
  assign n44325 = pi16 ? n42241 : n43787;
  assign n44326 = pi15 ? n44324 : n44325;
  assign n44327 = pi17 ? n41692 : n43791;
  assign n44328 = pi16 ? n41710 : n44327;
  assign n44329 = pi17 ? n41692 : n43796;
  assign n44330 = pi16 ? n38959 : n44329;
  assign n44331 = pi15 ? n44328 : n44330;
  assign n44332 = pi14 ? n44326 : n44331;
  assign n44333 = pi13 ? n44323 : n44332;
  assign n44334 = pi12 ? n44299 : n44333;
  assign n44335 = pi18 ? n20563 : n35318;
  assign n44336 = pi17 ? n44335 : n43805;
  assign n44337 = pi16 ? n40047 : n44336;
  assign n44338 = pi22 ? n35912 : n688;
  assign n44339 = pi21 ? n37 : n44338;
  assign n44340 = pi20 ? n44339 : n32;
  assign n44341 = pi19 ? n37 : n44340;
  assign n44342 = pi18 ? n37 : n44341;
  assign n44343 = pi17 ? n44335 : n44342;
  assign n44344 = pi16 ? n40047 : n44343;
  assign n44345 = pi15 ? n44337 : n44344;
  assign n44346 = pi22 ? n11680 : n688;
  assign n44347 = pi21 ? n37 : n44346;
  assign n44348 = pi20 ? n44347 : n32;
  assign n44349 = pi19 ? n37 : n44348;
  assign n44350 = pi18 ? n37 : n44349;
  assign n44351 = pi17 ? n41722 : n44350;
  assign n44352 = pi16 ? n40047 : n44351;
  assign n44353 = pi17 ? n40542 : n43826;
  assign n44354 = pi16 ? n39399 : n44353;
  assign n44355 = pi15 ? n44352 : n44354;
  assign n44356 = pi14 ? n44345 : n44355;
  assign n44357 = pi17 ? n41722 : n43832;
  assign n44358 = pi16 ? n38331 : n44357;
  assign n44359 = pi18 ? n20563 : n31300;
  assign n44360 = pi17 ? n44359 : n43370;
  assign n44361 = pi16 ? n38331 : n44360;
  assign n44362 = pi15 ? n44358 : n44361;
  assign n44363 = pi18 ? n15175 : n43840;
  assign n44364 = pi17 ? n41198 : n44363;
  assign n44365 = pi16 ? n37930 : n44364;
  assign n44366 = pi15 ? n44361 : n44365;
  assign n44367 = pi14 ? n44362 : n44366;
  assign n44368 = pi13 ? n44356 : n44367;
  assign n44369 = pi17 ? n43343 : n43370;
  assign n44370 = pi16 ? n37937 : n44369;
  assign n44371 = pi17 ? n40048 : n43388;
  assign n44372 = pi16 ? n37937 : n44371;
  assign n44373 = pi15 ? n44370 : n44372;
  assign n44374 = pi17 ? n40041 : n43856;
  assign n44375 = pi16 ? n37937 : n44374;
  assign n44376 = pi18 ? n36931 : n37;
  assign n44377 = pi20 ? n30461 : n32;
  assign n44378 = pi19 ? n99 : n44377;
  assign n44379 = pi18 ? n19774 : n44378;
  assign n44380 = pi17 ? n44376 : n44379;
  assign n44381 = pi16 ? n36871 : n44380;
  assign n44382 = pi15 ? n44375 : n44381;
  assign n44383 = pi14 ? n44373 : n44382;
  assign n44384 = pi18 ? n39432 : n19774;
  assign n44385 = pi21 ? n7429 : n882;
  assign n44386 = pi20 ? n44385 : n32;
  assign n44387 = pi19 ? n99 : n44386;
  assign n44388 = pi18 ? n99 : n44387;
  assign n44389 = pi17 ? n44384 : n44388;
  assign n44390 = pi16 ? n37959 : n44389;
  assign n44391 = pi16 ? n37959 : n43873;
  assign n44392 = pi15 ? n44390 : n44391;
  assign n44393 = pi18 ? n33823 : n21612;
  assign n44394 = pi19 ? n157 : n15330;
  assign n44395 = pi18 ? n43879 : n44394;
  assign n44396 = pi17 ? n44393 : n44395;
  assign n44397 = pi16 ? n37337 : n44396;
  assign n44398 = pi18 ? n33823 : n43884;
  assign n44399 = pi20 ? n27095 : n32;
  assign n44400 = pi19 ? n157 : n44399;
  assign n44401 = pi18 ? n43887 : n44400;
  assign n44402 = pi17 ? n44398 : n44401;
  assign n44403 = pi16 ? n38380 : n44402;
  assign n44404 = pi15 ? n44397 : n44403;
  assign n44405 = pi14 ? n44392 : n44404;
  assign n44406 = pi13 ? n44383 : n44405;
  assign n44407 = pi12 ? n44368 : n44406;
  assign n44408 = pi11 ? n44334 : n44407;
  assign n44409 = pi19 ? n43904 : n15330;
  assign n44410 = pi18 ? n43903 : n44409;
  assign n44411 = pi17 ? n43899 : n44410;
  assign n44412 = pi16 ? n39457 : n44411;
  assign n44413 = pi20 ? n39192 : n31298;
  assign n44414 = pi19 ? n20563 : n44413;
  assign n44415 = pi18 ? n44414 : n21612;
  assign n44416 = pi19 ? n38631 : n15330;
  assign n44417 = pi18 ? n43916 : n44416;
  assign n44418 = pi17 ? n44415 : n44417;
  assign n44419 = pi16 ? n39457 : n44418;
  assign n44420 = pi15 ? n44412 : n44419;
  assign n44421 = pi18 ? n33245 : n30851;
  assign n44422 = pi18 ? n21612 : n44416;
  assign n44423 = pi17 ? n44421 : n44422;
  assign n44424 = pi16 ? n36163 : n44423;
  assign n44425 = pi20 ? n2889 : n32;
  assign n44426 = pi19 ? n43928 : n44425;
  assign n44427 = pi18 ? n43927 : n44426;
  assign n44428 = pi17 ? n40062 : n44427;
  assign n44429 = pi16 ? n34860 : n44428;
  assign n44430 = pi15 ? n44424 : n44429;
  assign n44431 = pi14 ? n44420 : n44430;
  assign n44432 = pi19 ? n43940 : n15383;
  assign n44433 = pi18 ? n10652 : n44432;
  assign n44434 = pi17 ? n43938 : n44433;
  assign n44435 = pi16 ? n35765 : n44434;
  assign n44436 = pi20 ? n20563 : n39183;
  assign n44437 = pi19 ? n20563 : n44436;
  assign n44438 = pi18 ? n44437 : n15029;
  assign n44439 = pi17 ? n44438 : n43951;
  assign n44440 = pi16 ? n35765 : n44439;
  assign n44441 = pi15 ? n44435 : n44440;
  assign n44442 = pi18 ? n34295 : n14115;
  assign n44443 = pi21 ? n36058 : n32;
  assign n44444 = pi20 ? n44443 : n32;
  assign n44445 = pi19 ? n12589 : n44444;
  assign n44446 = pi18 ? n139 : n44445;
  assign n44447 = pi17 ? n44442 : n44446;
  assign n44448 = pi16 ? n36216 : n44447;
  assign n44449 = pi18 ? n34295 : n9796;
  assign n44450 = pi19 ? n12589 : n6272;
  assign n44451 = pi18 ? n139 : n44450;
  assign n44452 = pi17 ? n44449 : n44451;
  assign n44453 = pi16 ? n36216 : n44452;
  assign n44454 = pi15 ? n44448 : n44453;
  assign n44455 = pi14 ? n44441 : n44454;
  assign n44456 = pi13 ? n44431 : n44455;
  assign n44457 = pi18 ? n39626 : n43971;
  assign n44458 = pi19 ? n12589 : n10336;
  assign n44459 = pi18 ? n139 : n44458;
  assign n44460 = pi17 ? n44457 : n44459;
  assign n44461 = pi16 ? n36216 : n44460;
  assign n44462 = pi18 ? n34295 : n43975;
  assign n44463 = pi20 ? n30562 : n947;
  assign n44464 = pi19 ? n139 : n44463;
  assign n44465 = pi19 ? n9769 : n16520;
  assign n44466 = pi18 ? n44464 : n44465;
  assign n44467 = pi17 ? n44462 : n44466;
  assign n44468 = pi16 ? n36216 : n44467;
  assign n44469 = pi15 ? n44461 : n44468;
  assign n44470 = pi19 ? n42962 : n9964;
  assign n44471 = pi18 ? n43990 : n44470;
  assign n44472 = pi17 ? n39448 : n44471;
  assign n44473 = pi16 ? n36216 : n44472;
  assign n44474 = pi19 ? n43996 : n8296;
  assign n44475 = pi18 ? n43995 : n44474;
  assign n44476 = pi17 ? n39448 : n44475;
  assign n44477 = pi16 ? n36216 : n44476;
  assign n44478 = pi15 ? n44473 : n44477;
  assign n44479 = pi14 ? n44469 : n44478;
  assign n44480 = pi19 ? n44006 : n12150;
  assign n44481 = pi18 ? n44004 : n44480;
  assign n44482 = pi17 ? n39448 : n44481;
  assign n44483 = pi16 ? n36216 : n44482;
  assign n44484 = pi19 ? n44013 : n4009;
  assign n44485 = pi18 ? n44012 : n44484;
  assign n44486 = pi17 ? n39448 : n44485;
  assign n44487 = pi16 ? n36216 : n44486;
  assign n44488 = pi15 ? n44483 : n44487;
  assign n44489 = pi19 ? n6391 : n4103;
  assign n44490 = pi18 ? n44021 : n44489;
  assign n44491 = pi17 ? n38992 : n44490;
  assign n44492 = pi16 ? n36216 : n44491;
  assign n44493 = pi19 ? n6391 : n3341;
  assign n44494 = pi18 ? n44021 : n44493;
  assign n44495 = pi17 ? n39468 : n44494;
  assign n44496 = pi16 ? n36216 : n44495;
  assign n44497 = pi15 ? n44492 : n44496;
  assign n44498 = pi14 ? n44488 : n44497;
  assign n44499 = pi13 ? n44479 : n44498;
  assign n44500 = pi12 ? n44456 : n44499;
  assign n44501 = pi19 ? n6391 : n2639;
  assign n44502 = pi18 ? n41973 : n44501;
  assign n44503 = pi17 ? n39468 : n44502;
  assign n44504 = pi16 ? n43014 : n44503;
  assign n44505 = pi18 ? n32872 : n15082;
  assign n44506 = pi19 ? n13528 : n2654;
  assign n44507 = pi18 ? n335 : n44506;
  assign n44508 = pi17 ? n44505 : n44507;
  assign n44509 = pi16 ? n36216 : n44508;
  assign n44510 = pi15 ? n44504 : n44509;
  assign n44511 = pi18 ? n32872 : n335;
  assign n44512 = pi19 ? n44052 : n2702;
  assign n44513 = pi18 ? n335 : n44512;
  assign n44514 = pi17 ? n44511 : n44513;
  assign n44515 = pi16 ? n36216 : n44514;
  assign n44516 = pi21 ? n40986 : n30843;
  assign n44517 = pi20 ? n44516 : n37;
  assign n44518 = pi19 ? n20563 : n44517;
  assign n44519 = pi18 ? n44518 : n37;
  assign n44520 = pi19 ? n44060 : n1823;
  assign n44521 = pi18 ? n37 : n44520;
  assign n44522 = pi17 ? n44519 : n44521;
  assign n44523 = pi16 ? n36216 : n44522;
  assign n44524 = pi15 ? n44515 : n44523;
  assign n44525 = pi14 ? n44510 : n44524;
  assign n44526 = pi20 ? n31266 : n14530;
  assign n44527 = pi19 ? n20563 : n44526;
  assign n44528 = pi18 ? n44527 : n35637;
  assign n44529 = pi17 ? n44528 : n43540;
  assign n44530 = pi16 ? n36216 : n44529;
  assign n44531 = pi20 ? n31925 : n14530;
  assign n44532 = pi19 ? n20563 : n44531;
  assign n44533 = pi18 ? n44532 : n35637;
  assign n44534 = pi17 ? n44533 : n44076;
  assign n44535 = pi16 ? n36216 : n44534;
  assign n44536 = pi15 ? n44530 : n44535;
  assign n44537 = pi20 ? n31925 : n13179;
  assign n44538 = pi19 ? n20563 : n44537;
  assign n44539 = pi18 ? n44538 : n37;
  assign n44540 = pi20 ? n2107 : n18233;
  assign n44541 = pi19 ? n44540 : n32;
  assign n44542 = pi18 ? n44084 : n44541;
  assign n44543 = pi17 ? n44539 : n44542;
  assign n44544 = pi16 ? n36216 : n44543;
  assign n44545 = pi18 ? n44538 : n42063;
  assign n44546 = pi17 ? n44545 : n44095;
  assign n44547 = pi16 ? n36216 : n44546;
  assign n44548 = pi15 ? n44544 : n44547;
  assign n44549 = pi14 ? n44536 : n44548;
  assign n44550 = pi13 ? n44525 : n44549;
  assign n44551 = pi22 ? n36781 : n30195;
  assign n44552 = pi21 ? n20563 : n44551;
  assign n44553 = pi20 ? n44552 : n44103;
  assign n44554 = pi19 ? n20563 : n44553;
  assign n44555 = pi18 ? n44554 : n43076;
  assign n44556 = pi20 ? n26891 : n41526;
  assign n44557 = pi19 ? n44556 : n32;
  assign n44558 = pi18 ? n44108 : n44557;
  assign n44559 = pi17 ? n44555 : n44558;
  assign n44560 = pi16 ? n36216 : n44559;
  assign n44561 = pi22 ? n36781 : n37809;
  assign n44562 = pi21 ? n30868 : n44561;
  assign n44563 = pi23 ? n36781 : n99;
  assign n44564 = pi22 ? n44563 : n99;
  assign n44565 = pi21 ? n44564 : n22549;
  assign n44566 = pi20 ? n44562 : n44565;
  assign n44567 = pi19 ? n30868 : n44566;
  assign n44568 = pi18 ? n44567 : n44121;
  assign n44569 = pi21 ? n44124 : n3494;
  assign n44570 = pi20 ? n23162 : n44569;
  assign n44571 = pi19 ? n44570 : n32;
  assign n44572 = pi18 ? n44123 : n44571;
  assign n44573 = pi17 ? n44568 : n44572;
  assign n44574 = pi16 ? n42094 : n44573;
  assign n44575 = pi15 ? n44560 : n44574;
  assign n44576 = pi18 ? n40407 : n99;
  assign n44577 = pi20 ? n363 : n39889;
  assign n44578 = pi19 ? n44577 : n32;
  assign n44579 = pi18 ? n43116 : n44578;
  assign n44580 = pi17 ? n44576 : n44579;
  assign n44581 = pi16 ? n42094 : n44580;
  assign n44582 = pi20 ? n33792 : n43608;
  assign n44583 = pi19 ? n33792 : n44582;
  assign n44584 = pi18 ? n44583 : n43128;
  assign n44585 = pi17 ? n44584 : n44154;
  assign n44586 = pi16 ? n43125 : n44585;
  assign n44587 = pi15 ? n44581 : n44586;
  assign n44588 = pi14 ? n44575 : n44587;
  assign n44589 = pi18 ? n39971 : n43140;
  assign n44590 = pi17 ? n32 : n44589;
  assign n44591 = pi21 ? n36763 : n335;
  assign n44592 = pi20 ? n33792 : n44591;
  assign n44593 = pi19 ? n41579 : n44592;
  assign n44594 = pi18 ? n44593 : n139;
  assign n44595 = pi21 ? n4638 : n248;
  assign n44596 = pi20 ? n44174 : n44595;
  assign n44597 = pi19 ? n44173 : n44596;
  assign n44598 = pi18 ? n44597 : n44179;
  assign n44599 = pi17 ? n44594 : n44598;
  assign n44600 = pi16 ? n44590 : n44599;
  assign n44601 = pi20 ? n42147 : n43628;
  assign n44602 = pi19 ? n41102 : n44601;
  assign n44603 = pi18 ? n44602 : n44186;
  assign n44604 = pi17 ? n44603 : n43632;
  assign n44605 = pi16 ? n44590 : n44604;
  assign n44606 = pi15 ? n44600 : n44605;
  assign n44607 = pi18 ? n44140 : n43183;
  assign n44608 = pi17 ? n32 : n44607;
  assign n44609 = pi22 ? n36798 : n43636;
  assign n44610 = pi21 ? n44609 : n157;
  assign n44611 = pi20 ? n44191 : n44610;
  assign n44612 = pi19 ? n43186 : n44611;
  assign n44613 = pi18 ? n44612 : n157;
  assign n44614 = pi17 ? n44613 : n44199;
  assign n44615 = pi16 ? n44608 : n44614;
  assign n44616 = pi20 ? n44209 : n43645;
  assign n44617 = pi19 ? n44208 : n44616;
  assign n44618 = pi18 ? n44617 : n157;
  assign n44619 = pi21 ? n42627 : n928;
  assign n44620 = pi20 ? n157 : n44619;
  assign n44621 = pi19 ? n44620 : n32;
  assign n44622 = pi18 ? n157 : n44621;
  assign n44623 = pi17 ? n44618 : n44622;
  assign n44624 = pi16 ? n44207 : n44623;
  assign n44625 = pi15 ? n44615 : n44624;
  assign n44626 = pi14 ? n44606 : n44625;
  assign n44627 = pi13 ? n44588 : n44626;
  assign n44628 = pi12 ? n44550 : n44627;
  assign n44629 = pi11 ? n44500 : n44628;
  assign n44630 = pi10 ? n44408 : n44629;
  assign n44631 = pi09 ? n44238 : n44630;
  assign n44632 = pi08 ? n44221 : n44631;
  assign n44633 = pi07 ? n43662 : n44632;
  assign n44634 = pi18 ? n32 : n40056;
  assign n44635 = pi17 ? n32 : n44634;
  assign n44636 = pi19 ? n31267 : n35209;
  assign n44637 = pi20 ? n99 : n32;
  assign n44638 = pi19 ? n99 : n44637;
  assign n44639 = pi18 ? n44636 : n44638;
  assign n44640 = pi17 ? n20563 : n44639;
  assign n44641 = pi16 ? n44635 : n44640;
  assign n44642 = pi15 ? n32 : n44641;
  assign n44643 = pi18 ? n32 : n38999;
  assign n44644 = pi17 ? n32 : n44643;
  assign n44645 = pi19 ? n31280 : n17013;
  assign n44646 = pi20 ? n16008 : n181;
  assign n44647 = pi20 ? n1650 : n32;
  assign n44648 = pi19 ? n44646 : n44647;
  assign n44649 = pi18 ? n44645 : n44648;
  assign n44650 = pi17 ? n20563 : n44649;
  assign n44651 = pi16 ? n44644 : n44650;
  assign n44652 = pi18 ? n32 : n37322;
  assign n44653 = pi17 ? n32 : n44652;
  assign n44654 = pi20 ? n3096 : n32;
  assign n44655 = pi19 ? n37 : n44654;
  assign n44656 = pi18 ? n37 : n44655;
  assign n44657 = pi17 ? n20563 : n44656;
  assign n44658 = pi16 ? n44653 : n44657;
  assign n44659 = pi15 ? n44651 : n44658;
  assign n44660 = pi14 ? n44642 : n44659;
  assign n44661 = pi13 ? n32 : n44660;
  assign n44662 = pi12 ? n32 : n44661;
  assign n44663 = pi11 ? n32 : n44662;
  assign n44664 = pi10 ? n32 : n44663;
  assign n44665 = pi20 ? n3299 : n32;
  assign n44666 = pi19 ? n37 : n44665;
  assign n44667 = pi18 ? n37 : n44666;
  assign n44668 = pi17 ? n20563 : n44667;
  assign n44669 = pi16 ? n43664 : n44668;
  assign n44670 = pi18 ? n32 : n31315;
  assign n44671 = pi17 ? n32 : n44670;
  assign n44672 = pi22 ? n139 : n5011;
  assign n44673 = pi21 ? n139 : n44672;
  assign n44674 = pi20 ? n44673 : n32;
  assign n44675 = pi19 ? n13125 : n44674;
  assign n44676 = pi18 ? n32924 : n44675;
  assign n44677 = pi17 ? n20563 : n44676;
  assign n44678 = pi16 ? n44671 : n44677;
  assign n44679 = pi15 ? n44669 : n44678;
  assign n44680 = pi18 ? n20563 : n34869;
  assign n44681 = pi20 ? n29210 : n32;
  assign n44682 = pi19 ? n37 : n44681;
  assign n44683 = pi18 ? n37 : n44682;
  assign n44684 = pi17 ? n44680 : n44683;
  assign n44685 = pi16 ? n43685 : n44684;
  assign n44686 = pi19 ? n32 : n41681;
  assign n44687 = pi18 ? n32 : n44686;
  assign n44688 = pi17 ? n32 : n44687;
  assign n44689 = pi20 ? n28260 : n32;
  assign n44690 = pi19 ? n22792 : n44689;
  assign n44691 = pi18 ? n34582 : n44690;
  assign n44692 = pi17 ? n43676 : n44691;
  assign n44693 = pi16 ? n44688 : n44692;
  assign n44694 = pi15 ? n44685 : n44693;
  assign n44695 = pi14 ? n44679 : n44694;
  assign n44696 = pi18 ? n11567 : n44276;
  assign n44697 = pi17 ? n20563 : n44696;
  assign n44698 = pi16 ? n44688 : n44697;
  assign n44699 = pi19 ? n37 : n10621;
  assign n44700 = pi20 ? n28301 : n32;
  assign n44701 = pi19 ? n139 : n44700;
  assign n44702 = pi18 ? n44699 : n44701;
  assign n44703 = pi17 ? n44680 : n44702;
  assign n44704 = pi16 ? n42682 : n44703;
  assign n44705 = pi15 ? n44698 : n44704;
  assign n44706 = pi20 ? n8742 : n14573;
  assign n44707 = pi19 ? n37 : n44706;
  assign n44708 = pi20 ? n1704 : n37;
  assign n44709 = pi22 ? n335 : n6069;
  assign n44710 = pi21 ? n297 : n44709;
  assign n44711 = pi20 ? n44710 : n32;
  assign n44712 = pi19 ? n44708 : n44711;
  assign n44713 = pi18 ? n44707 : n44712;
  assign n44714 = pi17 ? n42657 : n44713;
  assign n44715 = pi16 ? n42682 : n44714;
  assign n44716 = pi21 ? n37 : n22278;
  assign n44717 = pi20 ? n44716 : n32;
  assign n44718 = pi19 ? n37 : n44717;
  assign n44719 = pi18 ? n37 : n44718;
  assign n44720 = pi17 ? n42657 : n44719;
  assign n44721 = pi16 ? n42682 : n44720;
  assign n44722 = pi15 ? n44715 : n44721;
  assign n44723 = pi14 ? n44705 : n44722;
  assign n44724 = pi13 ? n44695 : n44723;
  assign n44725 = pi22 ? n37 : n6077;
  assign n44726 = pi21 ? n37 : n44725;
  assign n44727 = pi20 ? n44726 : n32;
  assign n44728 = pi19 ? n37 : n44727;
  assign n44729 = pi18 ? n37 : n44728;
  assign n44730 = pi17 ? n42647 : n44729;
  assign n44731 = pi16 ? n42195 : n44730;
  assign n44732 = pi18 ? n20563 : n32275;
  assign n44733 = pi17 ? n44732 : n44719;
  assign n44734 = pi16 ? n41643 : n44733;
  assign n44735 = pi15 ? n44731 : n44734;
  assign n44736 = pi21 ? n569 : n7658;
  assign n44737 = pi20 ? n44736 : n32;
  assign n44738 = pi19 ? n37 : n44737;
  assign n44739 = pi18 ? n37 : n44738;
  assign n44740 = pi17 ? n42663 : n44739;
  assign n44741 = pi16 ? n42701 : n44740;
  assign n44742 = pi20 ? n3299 : n13273;
  assign n44743 = pi19 ? n37 : n44742;
  assign n44744 = pi19 ? n14394 : n44312;
  assign n44745 = pi18 ? n44743 : n44744;
  assign n44746 = pi17 ? n42690 : n44745;
  assign n44747 = pi16 ? n42701 : n44746;
  assign n44748 = pi15 ? n44741 : n44747;
  assign n44749 = pi14 ? n44735 : n44748;
  assign n44750 = pi19 ? n32876 : n30097;
  assign n44751 = pi18 ? n20563 : n44750;
  assign n44752 = pi19 ? n37 : n44317;
  assign n44753 = pi18 ? n37 : n44752;
  assign n44754 = pi17 ? n44751 : n44753;
  assign n44755 = pi16 ? n41159 : n44754;
  assign n44756 = pi21 ? n569 : n15100;
  assign n44757 = pi20 ? n44756 : n32;
  assign n44758 = pi19 ? n37 : n44757;
  assign n44759 = pi18 ? n37 : n44758;
  assign n44760 = pi17 ? n42690 : n44759;
  assign n44761 = pi16 ? n41170 : n44760;
  assign n44762 = pi15 ? n44755 : n44761;
  assign n44763 = pi21 ? n584 : n41110;
  assign n44764 = pi20 ? n44763 : n32;
  assign n44765 = pi19 ? n33694 : n44764;
  assign n44766 = pi18 ? n37 : n44765;
  assign n44767 = pi17 ? n41633 : n44766;
  assign n44768 = pi16 ? n40512 : n44767;
  assign n44769 = pi20 ? n2140 : n32;
  assign n44770 = pi19 ? n37 : n44769;
  assign n44771 = pi18 ? n37 : n44770;
  assign n44772 = pi17 ? n41633 : n44771;
  assign n44773 = pi16 ? n39375 : n44772;
  assign n44774 = pi15 ? n44768 : n44773;
  assign n44775 = pi14 ? n44762 : n44774;
  assign n44776 = pi13 ? n44749 : n44775;
  assign n44777 = pi12 ? n44724 : n44776;
  assign n44778 = pi20 ? n1409 : n32;
  assign n44779 = pi19 ? n37 : n44778;
  assign n44780 = pi18 ? n37 : n44779;
  assign n44781 = pi17 ? n43294 : n44780;
  assign n44782 = pi16 ? n40534 : n44781;
  assign n44783 = pi21 ? n3392 : n1408;
  assign n44784 = pi20 ? n44783 : n32;
  assign n44785 = pi19 ? n37 : n44784;
  assign n44786 = pi18 ? n37 : n44785;
  assign n44787 = pi17 ? n41672 : n44786;
  assign n44788 = pi16 ? n40534 : n44787;
  assign n44789 = pi15 ? n44782 : n44788;
  assign n44790 = pi21 ? n3392 : n34942;
  assign n44791 = pi20 ? n44790 : n32;
  assign n44792 = pi19 ? n37 : n44791;
  assign n44793 = pi18 ? n37 : n44792;
  assign n44794 = pi17 ? n41672 : n44793;
  assign n44795 = pi16 ? n40534 : n44794;
  assign n44796 = pi19 ? n35667 : n44791;
  assign n44797 = pi18 ? n37 : n44796;
  assign n44798 = pi17 ? n42228 : n44797;
  assign n44799 = pi16 ? n38950 : n44798;
  assign n44800 = pi15 ? n44795 : n44799;
  assign n44801 = pi14 ? n44789 : n44800;
  assign n44802 = pi19 ? n19092 : n15723;
  assign n44803 = pi18 ? n37 : n44802;
  assign n44804 = pi17 ? n41685 : n44803;
  assign n44805 = pi16 ? n38959 : n44804;
  assign n44806 = pi19 ? n37 : n15723;
  assign n44807 = pi18 ? n37 : n44806;
  assign n44808 = pi17 ? n41685 : n44807;
  assign n44809 = pi16 ? n38959 : n44808;
  assign n44810 = pi15 ? n44805 : n44809;
  assign n44811 = pi19 ? n37 : n15736;
  assign n44812 = pi18 ? n37 : n44811;
  assign n44813 = pi17 ? n41178 : n44812;
  assign n44814 = pi16 ? n38959 : n44813;
  assign n44815 = pi16 ? n40047 : n44813;
  assign n44816 = pi15 ? n44814 : n44815;
  assign n44817 = pi14 ? n44810 : n44816;
  assign n44818 = pi13 ? n44801 : n44817;
  assign n44819 = pi21 ? n6433 : n3523;
  assign n44820 = pi20 ? n44819 : n32;
  assign n44821 = pi19 ? n37 : n44820;
  assign n44822 = pi18 ? n37 : n44821;
  assign n44823 = pi17 ? n41178 : n44822;
  assign n44824 = pi16 ? n38318 : n44823;
  assign n44825 = pi17 ? n41178 : n43388;
  assign n44826 = pi16 ? n38318 : n44825;
  assign n44827 = pi19 ? n30097 : n21611;
  assign n44828 = pi18 ? n20563 : n44827;
  assign n44829 = pi22 ? n19177 : n316;
  assign n44830 = pi21 ? n44829 : n2320;
  assign n44831 = pi20 ? n44830 : n32;
  assign n44832 = pi19 ? n99 : n44831;
  assign n44833 = pi18 ? n99 : n44832;
  assign n44834 = pi17 ? n44828 : n44833;
  assign n44835 = pi16 ? n38331 : n44834;
  assign n44836 = pi15 ? n44826 : n44835;
  assign n44837 = pi14 ? n44824 : n44836;
  assign n44838 = pi18 ? n20563 : n31281;
  assign n44839 = pi18 ? n99 : n43861;
  assign n44840 = pi17 ? n44838 : n44839;
  assign n44841 = pi16 ? n38985 : n44840;
  assign n44842 = pi18 ? n20563 : n36403;
  assign n44843 = pi19 ? n19134 : n44399;
  assign n44844 = pi18 ? n26668 : n44843;
  assign n44845 = pi17 ? n44842 : n44844;
  assign n44846 = pi16 ? n38985 : n44845;
  assign n44847 = pi15 ? n44841 : n44846;
  assign n44848 = pi20 ? n32286 : n14844;
  assign n44849 = pi21 ? n99 : n3013;
  assign n44850 = pi20 ? n99 : n44849;
  assign n44851 = pi19 ? n44848 : n44850;
  assign n44852 = pi18 ? n20563 : n44851;
  assign n44853 = pi20 ? n10532 : n157;
  assign n44854 = pi19 ? n10527 : n44853;
  assign n44855 = pi19 ? n6532 : n15288;
  assign n44856 = pi18 ? n44854 : n44855;
  assign n44857 = pi17 ? n44852 : n44856;
  assign n44858 = pi16 ? n38985 : n44857;
  assign n44859 = pi20 ? n160 : n6508;
  assign n44860 = pi19 ? n99 : n44859;
  assign n44861 = pi20 ? n2243 : n10021;
  assign n44862 = pi21 ? n3562 : n2578;
  assign n44863 = pi20 ? n44862 : n32;
  assign n44864 = pi19 ? n44861 : n44863;
  assign n44865 = pi18 ? n44860 : n44864;
  assign n44866 = pi17 ? n44828 : n44865;
  assign n44867 = pi16 ? n40058 : n44866;
  assign n44868 = pi15 ? n44858 : n44867;
  assign n44869 = pi14 ? n44847 : n44868;
  assign n44870 = pi13 ? n44837 : n44869;
  assign n44871 = pi12 ? n44818 : n44870;
  assign n44872 = pi11 ? n44777 : n44871;
  assign n44873 = pi21 ? n41875 : n99;
  assign n44874 = pi20 ? n44873 : n3760;
  assign n44875 = pi19 ? n99 : n44874;
  assign n44876 = pi20 ? n41882 : n2383;
  assign n44877 = pi20 ? n3737 : n32;
  assign n44878 = pi19 ? n44876 : n44877;
  assign n44879 = pi18 ? n44875 : n44878;
  assign n44880 = pi17 ? n41192 : n44879;
  assign n44881 = pi16 ? n37937 : n44880;
  assign n44882 = pi20 ? n31903 : n14844;
  assign n44883 = pi19 ? n44882 : n3050;
  assign n44884 = pi18 ? n20563 : n44883;
  assign n44885 = pi19 ? n99 : n21611;
  assign n44886 = pi20 ? n99 : n2383;
  assign n44887 = pi19 ? n44886 : n44877;
  assign n44888 = pi18 ? n44885 : n44887;
  assign n44889 = pi17 ? n44884 : n44888;
  assign n44890 = pi16 ? n37937 : n44889;
  assign n44891 = pi15 ? n44881 : n44890;
  assign n44892 = pi20 ? n37 : n941;
  assign n44893 = pi19 ? n37 : n44892;
  assign n44894 = pi21 ? n20098 : n1027;
  assign n44895 = pi20 ? n139 : n44894;
  assign n44896 = pi19 ? n44895 : n44877;
  assign n44897 = pi18 ? n44893 : n44896;
  assign n44898 = pi17 ? n41198 : n44897;
  assign n44899 = pi16 ? n39001 : n44898;
  assign n44900 = pi20 ? n297 : n992;
  assign n44901 = pi19 ? n37 : n44900;
  assign n44902 = pi20 ? n992 : n2316;
  assign n44903 = pi21 ? n25463 : n2700;
  assign n44904 = pi20 ? n44903 : n32;
  assign n44905 = pi19 ? n44902 : n44904;
  assign n44906 = pi18 ? n44901 : n44905;
  assign n44907 = pi17 ? n44359 : n44906;
  assign n44908 = pi16 ? n37324 : n44907;
  assign n44909 = pi15 ? n44899 : n44908;
  assign n44910 = pi14 ? n44891 : n44909;
  assign n44911 = pi19 ? n20563 : n42915;
  assign n44912 = pi18 ? n44911 : n37;
  assign n44913 = pi21 ? n25463 : n1009;
  assign n44914 = pi20 ? n44913 : n32;
  assign n44915 = pi19 ? n2317 : n44914;
  assign n44916 = pi18 ? n8766 : n44915;
  assign n44917 = pi17 ? n44912 : n44916;
  assign n44918 = pi16 ? n37337 : n44917;
  assign n44919 = pi18 ? n34258 : n16093;
  assign n44920 = pi20 ? n139 : n6172;
  assign n44921 = pi22 ? n204 : n27692;
  assign n44922 = pi21 ? n44921 : n20952;
  assign n44923 = pi20 ? n44922 : n32;
  assign n44924 = pi19 ? n44920 : n44923;
  assign n44925 = pi18 ? n139 : n44924;
  assign n44926 = pi17 ? n44919 : n44925;
  assign n44927 = pi16 ? n37337 : n44926;
  assign n44928 = pi15 ? n44918 : n44927;
  assign n44929 = pi19 ? n32933 : n9765;
  assign n44930 = pi18 ? n34865 : n44929;
  assign n44931 = pi19 ? n36541 : n16507;
  assign n44932 = pi18 ? n139 : n44931;
  assign n44933 = pi17 ? n44930 : n44932;
  assign n44934 = pi16 ? n38380 : n44933;
  assign n44935 = pi19 ? n32933 : n14962;
  assign n44936 = pi18 ? n34865 : n44935;
  assign n44937 = pi19 ? n1017 : n6272;
  assign n44938 = pi18 ? n139 : n44937;
  assign n44939 = pi17 ? n44936 : n44938;
  assign n44940 = pi16 ? n38380 : n44939;
  assign n44941 = pi15 ? n44934 : n44940;
  assign n44942 = pi14 ? n44928 : n44941;
  assign n44943 = pi13 ? n44910 : n44942;
  assign n44944 = pi20 ? n942 : n947;
  assign n44945 = pi19 ? n9765 : n44944;
  assign n44946 = pi18 ? n34258 : n44945;
  assign n44947 = pi19 ? n139 : n9442;
  assign n44948 = pi18 ? n139 : n44947;
  assign n44949 = pi17 ? n44946 : n44948;
  assign n44950 = pi16 ? n39457 : n44949;
  assign n44951 = pi20 ? n376 : n947;
  assign n44952 = pi19 ? n44951 : n139;
  assign n44953 = pi18 ? n34258 : n44952;
  assign n44954 = pi19 ? n139 : n16520;
  assign n44955 = pi18 ? n139 : n44954;
  assign n44956 = pi17 ? n44953 : n44955;
  assign n44957 = pi16 ? n39457 : n44956;
  assign n44958 = pi15 ? n44950 : n44957;
  assign n44959 = pi19 ? n19405 : n16520;
  assign n44960 = pi18 ? n10682 : n44959;
  assign n44961 = pi17 ? n40041 : n44960;
  assign n44962 = pi16 ? n36163 : n44961;
  assign n44963 = pi20 ? n577 : n30674;
  assign n44964 = pi19 ? n37 : n44963;
  assign n44965 = pi20 ? n26002 : n233;
  assign n44966 = pi19 ? n44965 : n9964;
  assign n44967 = pi18 ? n44964 : n44966;
  assign n44968 = pi17 ? n40041 : n44967;
  assign n44969 = pi16 ? n36163 : n44968;
  assign n44970 = pi15 ? n44962 : n44969;
  assign n44971 = pi14 ? n44958 : n44970;
  assign n44972 = pi20 ? n31811 : n233;
  assign n44973 = pi19 ? n37 : n44972;
  assign n44974 = pi20 ? n233 : n6376;
  assign n44975 = pi19 ? n44974 : n8296;
  assign n44976 = pi18 ? n44973 : n44975;
  assign n44977 = pi17 ? n39415 : n44976;
  assign n44978 = pi16 ? n36216 : n44977;
  assign n44979 = pi19 ? n233 : n4009;
  assign n44980 = pi18 ? n28724 : n44979;
  assign n44981 = pi17 ? n39415 : n44980;
  assign n44982 = pi16 ? n36216 : n44981;
  assign n44983 = pi15 ? n44978 : n44982;
  assign n44984 = pi20 ? n26846 : n233;
  assign n44985 = pi19 ? n37 : n44984;
  assign n44986 = pi19 ? n7981 : n4009;
  assign n44987 = pi18 ? n44985 : n44986;
  assign n44988 = pi17 ? n40584 : n44987;
  assign n44989 = pi16 ? n36216 : n44988;
  assign n44990 = pi18 ? n37808 : n42015;
  assign n44991 = pi17 ? n32 : n44990;
  assign n44992 = pi23 ? n233 : n20004;
  assign n44993 = pi22 ? n44992 : n32;
  assign n44994 = pi21 ? n44993 : n32;
  assign n44995 = pi20 ? n44994 : n32;
  assign n44996 = pi19 ? n32703 : n44995;
  assign n44997 = pi18 ? n15161 : n44996;
  assign n44998 = pi17 ? n39440 : n44997;
  assign n44999 = pi16 ? n44991 : n44998;
  assign n45000 = pi15 ? n44989 : n44999;
  assign n45001 = pi14 ? n44983 : n45000;
  assign n45002 = pi13 ? n44971 : n45001;
  assign n45003 = pi12 ? n44943 : n45002;
  assign n45004 = pi22 ? n37804 : n33792;
  assign n45005 = pi21 ? n45004 : n33792;
  assign n45006 = pi20 ? n32 : n45005;
  assign n45007 = pi19 ? n32 : n45006;
  assign n45008 = pi22 ? n36615 : n33792;
  assign n45009 = pi21 ? n33792 : n45008;
  assign n45010 = pi21 ? n40955 : n33792;
  assign n45011 = pi20 ? n45009 : n45010;
  assign n45012 = pi19 ? n33792 : n45011;
  assign n45013 = pi18 ? n45007 : n45012;
  assign n45014 = pi17 ? n32 : n45013;
  assign n45015 = pi21 ? n40957 : n40960;
  assign n45016 = pi22 ? n20563 : n33792;
  assign n45017 = pi21 ? n40957 : n45016;
  assign n45018 = pi20 ? n45015 : n45017;
  assign n45019 = pi20 ? n45009 : n30096;
  assign n45020 = pi19 ? n45018 : n45019;
  assign n45021 = pi18 ? n45020 : n37;
  assign n45022 = pi20 ? n647 : n233;
  assign n45023 = pi19 ? n45022 : n2639;
  assign n45024 = pi18 ? n25114 : n45023;
  assign n45025 = pi17 ? n45021 : n45024;
  assign n45026 = pi16 ? n45014 : n45025;
  assign n45027 = pi18 ? n33245 : n16147;
  assign n45028 = pi20 ? n335 : n6376;
  assign n45029 = pi19 ? n45028 : n2654;
  assign n45030 = pi18 ? n335 : n45029;
  assign n45031 = pi17 ? n45027 : n45030;
  assign n45032 = pi16 ? n36216 : n45031;
  assign n45033 = pi15 ? n45026 : n45032;
  assign n45034 = pi19 ? n37 : n29400;
  assign n45035 = pi21 ? n6401 : n2721;
  assign n45036 = pi20 ? n37 : n45035;
  assign n45037 = pi19 ? n45036 : n2702;
  assign n45038 = pi18 ? n45034 : n45037;
  assign n45039 = pi17 ? n40584 : n45038;
  assign n45040 = pi16 ? n36216 : n45039;
  assign n45041 = pi21 ? n2106 : n6461;
  assign n45042 = pi20 ? n37 : n45041;
  assign n45043 = pi19 ? n45042 : n2702;
  assign n45044 = pi18 ? n45034 : n45043;
  assign n45045 = pi17 ? n40584 : n45044;
  assign n45046 = pi16 ? n36216 : n45045;
  assign n45047 = pi15 ? n45040 : n45046;
  assign n45048 = pi14 ? n45033 : n45047;
  assign n45049 = pi22 ? n40386 : n20563;
  assign n45050 = pi21 ? n45049 : n37;
  assign n45051 = pi20 ? n20563 : n45050;
  assign n45052 = pi19 ? n20563 : n45051;
  assign n45053 = pi20 ? n363 : n27501;
  assign n45054 = pi19 ? n23302 : n45053;
  assign n45055 = pi18 ? n45052 : n45054;
  assign n45056 = pi19 ? n24880 : n39867;
  assign n45057 = pi20 ? n22881 : n25199;
  assign n45058 = pi19 ? n45057 : n1823;
  assign n45059 = pi18 ? n45056 : n45058;
  assign n45060 = pi17 ? n45055 : n45059;
  assign n45061 = pi16 ? n36216 : n45060;
  assign n45062 = pi20 ? n16008 : n14887;
  assign n45063 = pi19 ? n45062 : n43075;
  assign n45064 = pi18 ? n45052 : n45063;
  assign n45065 = pi19 ? n37 : n43075;
  assign n45066 = pi21 ? n3392 : n685;
  assign n45067 = pi20 ? n22881 : n45066;
  assign n45068 = pi19 ? n45067 : n32;
  assign n45069 = pi18 ? n45065 : n45068;
  assign n45070 = pi17 ? n45064 : n45069;
  assign n45071 = pi16 ? n36216 : n45070;
  assign n45072 = pi15 ? n45061 : n45071;
  assign n45073 = pi21 ? n40954 : n29133;
  assign n45074 = pi20 ? n20563 : n45073;
  assign n45075 = pi19 ? n20563 : n45074;
  assign n45076 = pi18 ? n45075 : n19855;
  assign n45077 = pi21 ? n685 : n5113;
  assign n45078 = pi20 ? n363 : n45077;
  assign n45079 = pi19 ? n45078 : n32;
  assign n45080 = pi18 ? n24881 : n45079;
  assign n45081 = pi17 ? n45076 : n45080;
  assign n45082 = pi16 ? n36216 : n45081;
  assign n45083 = pi19 ? n39867 : n30805;
  assign n45084 = pi20 ? n24220 : n2782;
  assign n45085 = pi19 ? n45084 : n32;
  assign n45086 = pi18 ? n45083 : n45085;
  assign n45087 = pi17 ? n45076 : n45086;
  assign n45088 = pi16 ? n36216 : n45087;
  assign n45089 = pi15 ? n45082 : n45088;
  assign n45090 = pi14 ? n45072 : n45089;
  assign n45091 = pi13 ? n45048 : n45090;
  assign n45092 = pi22 ? n43571 : n20563;
  assign n45093 = pi21 ? n45092 : n29133;
  assign n45094 = pi20 ? n20563 : n45093;
  assign n45095 = pi19 ? n20563 : n45094;
  assign n45096 = pi20 ? n3292 : n37;
  assign n45097 = pi20 ? n7730 : n685;
  assign n45098 = pi19 ? n45096 : n45097;
  assign n45099 = pi18 ? n45095 : n45098;
  assign n45100 = pi19 ? n685 : n35660;
  assign n45101 = pi20 ? n685 : n42552;
  assign n45102 = pi19 ? n45101 : n32;
  assign n45103 = pi18 ? n45100 : n45102;
  assign n45104 = pi17 ? n45099 : n45103;
  assign n45105 = pi16 ? n36216 : n45104;
  assign n45106 = pi23 ? n36659 : n30868;
  assign n45107 = pi22 ? n45106 : n30868;
  assign n45108 = pi21 ? n45107 : n39926;
  assign n45109 = pi20 ? n30868 : n45108;
  assign n45110 = pi19 ? n30868 : n45109;
  assign n45111 = pi21 ? n22113 : n99;
  assign n45112 = pi20 ? n45111 : n23150;
  assign n45113 = pi19 ? n45112 : n363;
  assign n45114 = pi18 ? n45110 : n45113;
  assign n45115 = pi19 ? n28767 : n35660;
  assign n45116 = pi21 ? n14255 : n26377;
  assign n45117 = pi20 ? n26891 : n45116;
  assign n45118 = pi19 ? n45117 : n32;
  assign n45119 = pi18 ? n45115 : n45118;
  assign n45120 = pi17 ? n45114 : n45119;
  assign n45121 = pi16 ? n42094 : n45120;
  assign n45122 = pi15 ? n45105 : n45121;
  assign n45123 = pi20 ? n30868 : n39927;
  assign n45124 = pi19 ? n30868 : n45123;
  assign n45125 = pi18 ? n45124 : n99;
  assign n45126 = pi21 ? n722 : n685;
  assign n45127 = pi20 ? n99 : n45126;
  assign n45128 = pi19 ? n45127 : n685;
  assign n45129 = pi21 ? n14255 : n8486;
  assign n45130 = pi20 ? n363 : n45129;
  assign n45131 = pi19 ? n45130 : n32;
  assign n45132 = pi18 ? n45128 : n45131;
  assign n45133 = pi17 ? n45125 : n45132;
  assign n45134 = pi16 ? n42094 : n45133;
  assign n45135 = pi23 ? n32 : n36781;
  assign n45136 = pi22 ? n45135 : n36781;
  assign n45137 = pi21 ? n45136 : n36781;
  assign n45138 = pi20 ? n32 : n45137;
  assign n45139 = pi19 ? n32 : n45138;
  assign n45140 = pi21 ? n39972 : n36798;
  assign n45141 = pi20 ? n45140 : n36798;
  assign n45142 = pi22 ? n36798 : n33792;
  assign n45143 = pi21 ? n36798 : n45142;
  assign n45144 = pi20 ? n45143 : n33792;
  assign n45145 = pi19 ? n45141 : n45144;
  assign n45146 = pi18 ? n45139 : n45145;
  assign n45147 = pi17 ? n32 : n45146;
  assign n45148 = pi18 ? n33792 : n139;
  assign n45149 = pi21 ? n43146 : n43144;
  assign n45150 = pi20 ? n45149 : n44149;
  assign n45151 = pi20 ? n44149 : n28516;
  assign n45152 = pi19 ? n45150 : n45151;
  assign n45153 = pi20 ? n685 : n15754;
  assign n45154 = pi19 ? n45153 : n32;
  assign n45155 = pi18 ? n45152 : n45154;
  assign n45156 = pi17 ? n45148 : n45155;
  assign n45157 = pi16 ? n45147 : n45156;
  assign n45158 = pi15 ? n45134 : n45157;
  assign n45159 = pi14 ? n45122 : n45158;
  assign n45160 = pi23 ? n32 : n36798;
  assign n45161 = pi22 ? n45160 : n36798;
  assign n45162 = pi21 ? n45161 : n36798;
  assign n45163 = pi20 ? n32 : n45162;
  assign n45164 = pi19 ? n32 : n45163;
  assign n45165 = pi20 ? n45143 : n36659;
  assign n45166 = pi19 ? n36798 : n45165;
  assign n45167 = pi18 ? n45164 : n45166;
  assign n45168 = pi17 ? n32 : n45167;
  assign n45169 = pi19 ? n41089 : n335;
  assign n45170 = pi18 ? n41580 : n45169;
  assign n45171 = pi21 ? n157 : n1785;
  assign n45172 = pi20 ? n45171 : n316;
  assign n45173 = pi19 ? n139 : n45172;
  assign n45174 = pi21 ? n6132 : n2320;
  assign n45175 = pi20 ? n157 : n45174;
  assign n45176 = pi19 ? n45175 : n32;
  assign n45177 = pi18 ? n45173 : n45176;
  assign n45178 = pi17 ? n45170 : n45177;
  assign n45179 = pi16 ? n45168 : n45178;
  assign n45180 = pi20 ? n36781 : n36659;
  assign n45181 = pi19 ? n36781 : n45180;
  assign n45182 = pi18 ? n45139 : n45181;
  assign n45183 = pi17 ? n32 : n45182;
  assign n45184 = pi19 ? n41107 : n335;
  assign n45185 = pi18 ? n41103 : n45184;
  assign n45186 = pi21 ? n3693 : n1091;
  assign n45187 = pi20 ? n45186 : n34537;
  assign n45188 = pi20 ? n7435 : n34538;
  assign n45189 = pi19 ? n45187 : n45188;
  assign n45190 = pi20 ? n17390 : n2330;
  assign n45191 = pi19 ? n45190 : n32;
  assign n45192 = pi18 ? n45189 : n45191;
  assign n45193 = pi17 ? n45185 : n45192;
  assign n45194 = pi16 ? n45183 : n45193;
  assign n45195 = pi15 ? n45179 : n45194;
  assign n45196 = pi18 ? n45164 : n41136;
  assign n45197 = pi17 ? n32 : n45196;
  assign n45198 = pi19 ? n36781 : n44208;
  assign n45199 = pi21 ? n44192 : n36837;
  assign n45200 = pi20 ? n45199 : n157;
  assign n45201 = pi19 ? n45200 : n157;
  assign n45202 = pi18 ? n45198 : n45201;
  assign n45203 = pi23 ? n15293 : n233;
  assign n45204 = pi22 ? n157 : n45203;
  assign n45205 = pi21 ? n45204 : n928;
  assign n45206 = pi20 ? n157 : n45205;
  assign n45207 = pi19 ? n45206 : n32;
  assign n45208 = pi18 ? n157 : n45207;
  assign n45209 = pi17 ? n45202 : n45208;
  assign n45210 = pi16 ? n45197 : n45209;
  assign n45211 = pi22 ? n32 : n36783;
  assign n45212 = pi21 ? n45211 : n36781;
  assign n45213 = pi20 ? n32 : n45212;
  assign n45214 = pi19 ? n32 : n45213;
  assign n45215 = pi18 ? n45214 : n36781;
  assign n45216 = pi17 ? n32 : n45215;
  assign n45217 = pi21 ? n43203 : n5054;
  assign n45218 = pi20 ? n45217 : n157;
  assign n45219 = pi19 ? n45218 : n157;
  assign n45220 = pi18 ? n45198 : n45219;
  assign n45221 = pi17 ? n45220 : n44199;
  assign n45222 = pi16 ? n45216 : n45221;
  assign n45223 = pi15 ? n45210 : n45222;
  assign n45224 = pi14 ? n45195 : n45223;
  assign n45225 = pi13 ? n45159 : n45224;
  assign n45226 = pi12 ? n45091 : n45225;
  assign n45227 = pi11 ? n45003 : n45226;
  assign n45228 = pi10 ? n44872 : n45227;
  assign n45229 = pi09 ? n44664 : n45228;
  assign n45230 = pi16 ? n32 : n44640;
  assign n45231 = pi15 ? n32 : n45230;
  assign n45232 = pi18 ? n32 : n38983;
  assign n45233 = pi17 ? n32 : n45232;
  assign n45234 = pi16 ? n45233 : n44650;
  assign n45235 = pi15 ? n45234 : n44658;
  assign n45236 = pi14 ? n45231 : n45235;
  assign n45237 = pi13 ? n32 : n45236;
  assign n45238 = pi12 ? n32 : n45237;
  assign n45239 = pi11 ? n32 : n45238;
  assign n45240 = pi10 ? n32 : n45239;
  assign n45241 = pi16 ? n44223 : n44668;
  assign n45242 = pi18 ? n32 : n38378;
  assign n45243 = pi17 ? n32 : n45242;
  assign n45244 = pi16 ? n45243 : n44677;
  assign n45245 = pi15 ? n45241 : n45244;
  assign n45246 = pi18 ? n20563 : n36931;
  assign n45247 = pi17 ? n45246 : n44683;
  assign n45248 = pi16 ? n43664 : n45247;
  assign n45249 = pi19 ? n22792 : n16100;
  assign n45250 = pi18 ? n34582 : n45249;
  assign n45251 = pi17 ? n43676 : n45250;
  assign n45252 = pi16 ? n43664 : n45251;
  assign n45253 = pi15 ? n45248 : n45252;
  assign n45254 = pi14 ? n45245 : n45253;
  assign n45255 = pi19 ? n139 : n16100;
  assign n45256 = pi18 ? n11567 : n45255;
  assign n45257 = pi17 ? n20563 : n45256;
  assign n45258 = pi16 ? n44671 : n45257;
  assign n45259 = pi19 ? n139 : n14954;
  assign n45260 = pi18 ? n44699 : n45259;
  assign n45261 = pi17 ? n44680 : n45260;
  assign n45262 = pi16 ? n43224 : n45261;
  assign n45263 = pi15 ? n45258 : n45262;
  assign n45264 = pi19 ? n37 : n13124;
  assign n45265 = pi20 ? n31082 : n37;
  assign n45266 = pi22 ? n335 : n6833;
  assign n45267 = pi21 ? n297 : n45266;
  assign n45268 = pi20 ? n45267 : n32;
  assign n45269 = pi19 ? n45265 : n45268;
  assign n45270 = pi18 ? n45264 : n45269;
  assign n45271 = pi17 ? n42657 : n45270;
  assign n45272 = pi16 ? n43228 : n45271;
  assign n45273 = pi21 ? n37 : n2061;
  assign n45274 = pi20 ? n45273 : n32;
  assign n45275 = pi19 ? n37 : n45274;
  assign n45276 = pi18 ? n37 : n45275;
  assign n45277 = pi17 ? n42657 : n45276;
  assign n45278 = pi16 ? n43249 : n45277;
  assign n45279 = pi15 ? n45272 : n45278;
  assign n45280 = pi14 ? n45263 : n45279;
  assign n45281 = pi13 ? n45254 : n45280;
  assign n45282 = pi21 ? n37 : n17755;
  assign n45283 = pi20 ? n45282 : n32;
  assign n45284 = pi19 ? n37 : n45283;
  assign n45285 = pi18 ? n37 : n45284;
  assign n45286 = pi17 ? n42647 : n45285;
  assign n45287 = pi16 ? n44275 : n45286;
  assign n45288 = pi21 ? n37 : n9900;
  assign n45289 = pi20 ? n45288 : n32;
  assign n45290 = pi19 ? n37 : n45289;
  assign n45291 = pi18 ? n37 : n45290;
  assign n45292 = pi17 ? n44732 : n45291;
  assign n45293 = pi16 ? n42202 : n45292;
  assign n45294 = pi15 ? n45287 : n45293;
  assign n45295 = pi21 ? n569 : n8869;
  assign n45296 = pi20 ? n45295 : n32;
  assign n45297 = pi19 ? n37 : n45296;
  assign n45298 = pi18 ? n37 : n45297;
  assign n45299 = pi17 ? n42663 : n45298;
  assign n45300 = pi16 ? n43263 : n45299;
  assign n45301 = pi22 ? n335 : n10768;
  assign n45302 = pi21 ? n335 : n45301;
  assign n45303 = pi20 ? n45302 : n32;
  assign n45304 = pi19 ? n14394 : n45303;
  assign n45305 = pi18 ? n44743 : n45304;
  assign n45306 = pi17 ? n43257 : n45305;
  assign n45307 = pi16 ? n41632 : n45306;
  assign n45308 = pi15 ? n45300 : n45307;
  assign n45309 = pi14 ? n45294 : n45308;
  assign n45310 = pi22 ? n233 : n10768;
  assign n45311 = pi21 ? n335 : n45310;
  assign n45312 = pi20 ? n45311 : n32;
  assign n45313 = pi19 ? n37 : n45312;
  assign n45314 = pi18 ? n37 : n45313;
  assign n45315 = pi17 ? n42663 : n45314;
  assign n45316 = pi16 ? n42689 : n45315;
  assign n45317 = pi15 ? n45316 : n44761;
  assign n45318 = pi22 ? n685 : n730;
  assign n45319 = pi21 ? n37 : n45318;
  assign n45320 = pi20 ? n45319 : n32;
  assign n45321 = pi19 ? n37 : n45320;
  assign n45322 = pi18 ? n37 : n45321;
  assign n45323 = pi17 ? n42196 : n45322;
  assign n45324 = pi16 ? n41170 : n45323;
  assign n45325 = pi16 ? n40025 : n44772;
  assign n45326 = pi15 ? n45324 : n45325;
  assign n45327 = pi14 ? n45317 : n45326;
  assign n45328 = pi13 ? n45309 : n45327;
  assign n45329 = pi12 ? n45281 : n45328;
  assign n45330 = pi20 ? n30972 : n32;
  assign n45331 = pi19 ? n37 : n45330;
  assign n45332 = pi18 ? n37 : n45331;
  assign n45333 = pi17 ? n43279 : n45332;
  assign n45334 = pi16 ? n41183 : n45333;
  assign n45335 = pi19 ? n40198 : n37;
  assign n45336 = pi18 ? n20563 : n45335;
  assign n45337 = pi17 ? n45336 : n44786;
  assign n45338 = pi16 ? n41183 : n45337;
  assign n45339 = pi15 ? n45334 : n45338;
  assign n45340 = pi17 ? n43279 : n44793;
  assign n45341 = pi16 ? n41684 : n45340;
  assign n45342 = pi17 ? n41672 : n44797;
  assign n45343 = pi16 ? n40512 : n45342;
  assign n45344 = pi15 ? n45341 : n45343;
  assign n45345 = pi14 ? n45339 : n45344;
  assign n45346 = pi21 ? n363 : n13687;
  assign n45347 = pi20 ? n45346 : n32;
  assign n45348 = pi19 ? n19092 : n45347;
  assign n45349 = pi18 ? n37 : n45348;
  assign n45350 = pi17 ? n41685 : n45349;
  assign n45351 = pi16 ? n39375 : n45350;
  assign n45352 = pi21 ? n363 : n22919;
  assign n45353 = pi20 ? n45352 : n32;
  assign n45354 = pi19 ? n37 : n45353;
  assign n45355 = pi18 ? n37 : n45354;
  assign n45356 = pi17 ? n41685 : n45355;
  assign n45357 = pi16 ? n39375 : n45356;
  assign n45358 = pi15 ? n45351 : n45357;
  assign n45359 = pi18 ? n20563 : n34949;
  assign n45360 = pi21 ? n2106 : n22919;
  assign n45361 = pi20 ? n45360 : n32;
  assign n45362 = pi19 ? n37 : n45361;
  assign n45363 = pi18 ? n37 : n45362;
  assign n45364 = pi17 ? n45359 : n45363;
  assign n45365 = pi16 ? n39375 : n45364;
  assign n45366 = pi19 ? n43246 : n20563;
  assign n45367 = pi18 ? n32 : n45366;
  assign n45368 = pi17 ? n32 : n45367;
  assign n45369 = pi17 ? n45359 : n44812;
  assign n45370 = pi16 ? n45368 : n45369;
  assign n45371 = pi15 ? n45365 : n45370;
  assign n45372 = pi14 ? n45358 : n45371;
  assign n45373 = pi13 ? n45345 : n45372;
  assign n45374 = pi17 ? n41692 : n44822;
  assign n45375 = pi16 ? n38950 : n45374;
  assign n45376 = pi21 ? n381 : n3523;
  assign n45377 = pi20 ? n45376 : n32;
  assign n45378 = pi19 ? n37 : n45377;
  assign n45379 = pi18 ? n37 : n45378;
  assign n45380 = pi17 ? n41178 : n45379;
  assign n45381 = pi16 ? n38950 : n45380;
  assign n45382 = pi19 ? n40149 : n21611;
  assign n45383 = pi18 ? n20563 : n45382;
  assign n45384 = pi21 ? n44829 : n3523;
  assign n45385 = pi20 ? n45384 : n32;
  assign n45386 = pi19 ? n99 : n45385;
  assign n45387 = pi18 ? n99 : n45386;
  assign n45388 = pi17 ? n45383 : n45387;
  assign n45389 = pi16 ? n38959 : n45388;
  assign n45390 = pi15 ? n45381 : n45389;
  assign n45391 = pi14 ? n45375 : n45390;
  assign n45392 = pi19 ? n42192 : n20563;
  assign n45393 = pi18 ? n32 : n45392;
  assign n45394 = pi17 ? n32 : n45393;
  assign n45395 = pi19 ? n35317 : n99;
  assign n45396 = pi18 ? n20563 : n45395;
  assign n45397 = pi18 ? n99 : n44378;
  assign n45398 = pi17 ? n45396 : n45397;
  assign n45399 = pi16 ? n45394 : n45398;
  assign n45400 = pi20 ? n28024 : n32;
  assign n45401 = pi19 ? n19134 : n45400;
  assign n45402 = pi18 ? n26668 : n45401;
  assign n45403 = pi17 ? n44842 : n45402;
  assign n45404 = pi16 ? n45394 : n45403;
  assign n45405 = pi15 ? n45399 : n45404;
  assign n45406 = pi20 ? n31220 : n14844;
  assign n45407 = pi19 ? n45406 : n44850;
  assign n45408 = pi18 ? n20563 : n45407;
  assign n45409 = pi19 ? n6532 : n15788;
  assign n45410 = pi18 ? n44854 : n45409;
  assign n45411 = pi17 ? n45408 : n45410;
  assign n45412 = pi16 ? n45394 : n45411;
  assign n45413 = pi19 ? n43253 : n20563;
  assign n45414 = pi18 ? n32 : n45413;
  assign n45415 = pi17 ? n32 : n45414;
  assign n45416 = pi21 ? n3562 : n3339;
  assign n45417 = pi20 ? n45416 : n32;
  assign n45418 = pi19 ? n44861 : n45417;
  assign n45419 = pi18 ? n44860 : n45418;
  assign n45420 = pi17 ? n44828 : n45419;
  assign n45421 = pi16 ? n45415 : n45420;
  assign n45422 = pi15 ? n45412 : n45421;
  assign n45423 = pi14 ? n45405 : n45422;
  assign n45424 = pi13 ? n45391 : n45423;
  assign n45425 = pi12 ? n45373 : n45424;
  assign n45426 = pi11 ? n45329 : n45425;
  assign n45427 = pi21 ? n1027 : n882;
  assign n45428 = pi20 ? n45427 : n32;
  assign n45429 = pi19 ? n44876 : n45428;
  assign n45430 = pi18 ? n44875 : n45429;
  assign n45431 = pi17 ? n41722 : n45430;
  assign n45432 = pi16 ? n38331 : n45431;
  assign n45433 = pi19 ? n44848 : n3050;
  assign n45434 = pi18 ? n20563 : n45433;
  assign n45435 = pi19 ? n44886 : n45428;
  assign n45436 = pi18 ? n44885 : n45435;
  assign n45437 = pi17 ? n45434 : n45436;
  assign n45438 = pi16 ? n38331 : n45437;
  assign n45439 = pi15 ? n45432 : n45438;
  assign n45440 = pi17 ? n44359 : n44897;
  assign n45441 = pi16 ? n38331 : n45440;
  assign n45442 = pi19 ? n44902 : n18375;
  assign n45443 = pi18 ? n44901 : n45442;
  assign n45444 = pi17 ? n41722 : n45443;
  assign n45445 = pi16 ? n37930 : n45444;
  assign n45446 = pi15 ? n45441 : n45445;
  assign n45447 = pi14 ? n45439 : n45446;
  assign n45448 = pi19 ? n2317 : n18375;
  assign n45449 = pi18 ? n8766 : n45448;
  assign n45450 = pi17 ? n44912 : n45449;
  assign n45451 = pi16 ? n38985 : n45450;
  assign n45452 = pi19 ? n33965 : n9814;
  assign n45453 = pi18 ? n34865 : n45452;
  assign n45454 = pi21 ? n3763 : n20952;
  assign n45455 = pi20 ? n45454 : n32;
  assign n45456 = pi19 ? n44920 : n45455;
  assign n45457 = pi18 ? n139 : n45456;
  assign n45458 = pi17 ? n45453 : n45457;
  assign n45459 = pi16 ? n38985 : n45458;
  assign n45460 = pi15 ? n45451 : n45459;
  assign n45461 = pi18 ? n20563 : n44929;
  assign n45462 = pi19 ? n36541 : n16477;
  assign n45463 = pi18 ? n139 : n45462;
  assign n45464 = pi17 ? n45461 : n45463;
  assign n45465 = pi16 ? n36871 : n45464;
  assign n45466 = pi18 ? n20563 : n44935;
  assign n45467 = pi19 ? n1017 : n7639;
  assign n45468 = pi18 ? n139 : n45467;
  assign n45469 = pi17 ? n45466 : n45468;
  assign n45470 = pi16 ? n36871 : n45469;
  assign n45471 = pi15 ? n45465 : n45470;
  assign n45472 = pi14 ? n45460 : n45471;
  assign n45473 = pi13 ? n45447 : n45472;
  assign n45474 = pi19 ? n139 : n17511;
  assign n45475 = pi18 ? n139 : n45474;
  assign n45476 = pi17 ? n44946 : n45475;
  assign n45477 = pi16 ? n37959 : n45476;
  assign n45478 = pi18 ? n34247 : n20723;
  assign n45479 = pi19 ? n139 : n16945;
  assign n45480 = pi18 ? n139 : n45479;
  assign n45481 = pi17 ? n45478 : n45480;
  assign n45482 = pi16 ? n37959 : n45481;
  assign n45483 = pi15 ? n45477 : n45482;
  assign n45484 = pi19 ? n19405 : n16945;
  assign n45485 = pi18 ? n10682 : n45484;
  assign n45486 = pi17 ? n41198 : n45485;
  assign n45487 = pi16 ? n39001 : n45486;
  assign n45488 = pi17 ? n41198 : n44967;
  assign n45489 = pi16 ? n39001 : n45488;
  assign n45490 = pi15 ? n45487 : n45489;
  assign n45491 = pi14 ? n45483 : n45490;
  assign n45492 = pi19 ? n44974 : n9457;
  assign n45493 = pi18 ? n44973 : n45492;
  assign n45494 = pi17 ? n39415 : n45493;
  assign n45495 = pi16 ? n37324 : n45494;
  assign n45496 = pi19 ? n233 : n5668;
  assign n45497 = pi18 ? n28724 : n45496;
  assign n45498 = pi17 ? n40048 : n45497;
  assign n45499 = pi16 ? n37324 : n45498;
  assign n45500 = pi15 ? n45495 : n45499;
  assign n45501 = pi16 ? n37337 : n44988;
  assign n45502 = pi21 ? n37332 : n30868;
  assign n45503 = pi20 ? n32 : n45502;
  assign n45504 = pi19 ? n32 : n45503;
  assign n45505 = pi18 ? n45504 : n42015;
  assign n45506 = pi17 ? n32 : n45505;
  assign n45507 = pi18 ? n35777 : n37;
  assign n45508 = pi19 ? n32703 : n4103;
  assign n45509 = pi18 ? n15161 : n45508;
  assign n45510 = pi17 ? n45507 : n45509;
  assign n45511 = pi16 ? n45506 : n45510;
  assign n45512 = pi15 ? n45501 : n45511;
  assign n45513 = pi14 ? n45500 : n45512;
  assign n45514 = pi13 ? n45491 : n45513;
  assign n45515 = pi12 ? n45473 : n45514;
  assign n45516 = pi23 ? n32 : n33793;
  assign n45517 = pi22 ? n45516 : n33792;
  assign n45518 = pi21 ? n45517 : n33792;
  assign n45519 = pi20 ? n32 : n45518;
  assign n45520 = pi19 ? n32 : n45519;
  assign n45521 = pi20 ? n33792 : n45010;
  assign n45522 = pi19 ? n33792 : n45521;
  assign n45523 = pi18 ? n45520 : n45522;
  assign n45524 = pi17 ? n32 : n45523;
  assign n45525 = pi21 ? n40955 : n40960;
  assign n45526 = pi22 ? n33792 : n37173;
  assign n45527 = pi21 ? n45526 : n45016;
  assign n45528 = pi20 ? n45525 : n45527;
  assign n45529 = pi22 ? n37173 : n30867;
  assign n45530 = pi21 ? n45529 : n37;
  assign n45531 = pi20 ? n33792 : n45530;
  assign n45532 = pi19 ? n45528 : n45531;
  assign n45533 = pi18 ? n45532 : n37;
  assign n45534 = pi19 ? n45022 : n4117;
  assign n45535 = pi18 ? n25114 : n45534;
  assign n45536 = pi17 ? n45533 : n45535;
  assign n45537 = pi16 ? n45524 : n45536;
  assign n45538 = pi18 ? n40199 : n16147;
  assign n45539 = pi19 ? n45028 : n10012;
  assign n45540 = pi18 ? n335 : n45539;
  assign n45541 = pi17 ? n45538 : n45540;
  assign n45542 = pi16 ? n35765 : n45541;
  assign n45543 = pi15 ? n45537 : n45542;
  assign n45544 = pi19 ? n45036 : n2654;
  assign n45545 = pi18 ? n45034 : n45544;
  assign n45546 = pi17 ? n40575 : n45545;
  assign n45547 = pi16 ? n35765 : n45546;
  assign n45548 = pi17 ? n40575 : n45044;
  assign n45549 = pi16 ? n35765 : n45548;
  assign n45550 = pi15 ? n45547 : n45549;
  assign n45551 = pi14 ? n45543 : n45550;
  assign n45552 = pi21 ? n45049 : n31200;
  assign n45553 = pi20 ? n20563 : n45552;
  assign n45554 = pi19 ? n20563 : n45553;
  assign n45555 = pi19 ? n37 : n45053;
  assign n45556 = pi18 ? n45554 : n45555;
  assign n45557 = pi19 ? n45057 : n2702;
  assign n45558 = pi18 ? n45056 : n45557;
  assign n45559 = pi17 ? n45556 : n45558;
  assign n45560 = pi16 ? n34860 : n45559;
  assign n45561 = pi21 ? n45049 : n30867;
  assign n45562 = pi20 ? n20563 : n45561;
  assign n45563 = pi19 ? n20563 : n45562;
  assign n45564 = pi19 ? n24263 : n43075;
  assign n45565 = pi18 ? n45563 : n45564;
  assign n45566 = pi19 ? n45067 : n2702;
  assign n45567 = pi18 ? n45065 : n45566;
  assign n45568 = pi17 ? n45565 : n45567;
  assign n45569 = pi16 ? n34860 : n45568;
  assign n45570 = pi15 ? n45560 : n45569;
  assign n45571 = pi21 ? n40954 : n31294;
  assign n45572 = pi20 ? n20563 : n45571;
  assign n45573 = pi19 ? n20563 : n45572;
  assign n45574 = pi18 ? n45573 : n37;
  assign n45575 = pi19 ? n45078 : n1823;
  assign n45576 = pi18 ? n24881 : n45575;
  assign n45577 = pi17 ? n45574 : n45576;
  assign n45578 = pi16 ? n38380 : n45577;
  assign n45579 = pi23 ? n685 : n13482;
  assign n45580 = pi22 ? n685 : n45579;
  assign n45581 = pi21 ? n685 : n45580;
  assign n45582 = pi20 ? n24220 : n45581;
  assign n45583 = pi19 ? n45582 : n32;
  assign n45584 = pi18 ? n45083 : n45583;
  assign n45585 = pi17 ? n45574 : n45584;
  assign n45586 = pi16 ? n38380 : n45585;
  assign n45587 = pi15 ? n45578 : n45586;
  assign n45588 = pi14 ? n45570 : n45587;
  assign n45589 = pi13 ? n45551 : n45588;
  assign n45590 = pi21 ? n45092 : n31294;
  assign n45591 = pi20 ? n20563 : n45590;
  assign n45592 = pi19 ? n20563 : n45591;
  assign n45593 = pi19 ? n37 : n45097;
  assign n45594 = pi18 ? n45592 : n45593;
  assign n45595 = pi17 ? n45594 : n45103;
  assign n45596 = pi16 ? n38380 : n45595;
  assign n45597 = pi23 ? n32 : n30868;
  assign n45598 = pi22 ? n32 : n45597;
  assign n45599 = pi21 ? n45598 : n30868;
  assign n45600 = pi20 ? n32 : n45599;
  assign n45601 = pi19 ? n32 : n45600;
  assign n45602 = pi18 ? n45601 : n30868;
  assign n45603 = pi17 ? n32 : n45602;
  assign n45604 = pi21 ? n45107 : n41564;
  assign n45605 = pi20 ? n30868 : n45604;
  assign n45606 = pi19 ? n30868 : n45605;
  assign n45607 = pi23 ? n99 : n36781;
  assign n45608 = pi22 ? n45607 : n99;
  assign n45609 = pi21 ? n45608 : n99;
  assign n45610 = pi20 ? n45609 : n23150;
  assign n45611 = pi19 ? n45610 : n363;
  assign n45612 = pi18 ? n45606 : n45611;
  assign n45613 = pi21 ? n14255 : n1423;
  assign n45614 = pi20 ? n26891 : n45613;
  assign n45615 = pi19 ? n45614 : n32;
  assign n45616 = pi18 ? n45115 : n45615;
  assign n45617 = pi17 ? n45612 : n45616;
  assign n45618 = pi16 ? n45603 : n45617;
  assign n45619 = pi15 ? n45596 : n45618;
  assign n45620 = pi22 ? n32 : n37804;
  assign n45621 = pi21 ? n45620 : n30868;
  assign n45622 = pi20 ? n32 : n45621;
  assign n45623 = pi19 ? n32 : n45622;
  assign n45624 = pi18 ? n45623 : n30868;
  assign n45625 = pi17 ? n32 : n45624;
  assign n45626 = pi19 ? n30868 : n43603;
  assign n45627 = pi18 ? n45626 : n99;
  assign n45628 = pi21 ? n14255 : n2230;
  assign n45629 = pi20 ? n363 : n45628;
  assign n45630 = pi19 ? n45629 : n32;
  assign n45631 = pi18 ? n45128 : n45630;
  assign n45632 = pi17 ? n45627 : n45631;
  assign n45633 = pi16 ? n45625 : n45632;
  assign n45634 = pi23 ? n32 : n36782;
  assign n45635 = pi22 ? n32 : n45634;
  assign n45636 = pi21 ? n45635 : n36781;
  assign n45637 = pi20 ? n32 : n45636;
  assign n45638 = pi19 ? n32 : n45637;
  assign n45639 = pi18 ? n45638 : n45145;
  assign n45640 = pi17 ? n32 : n45639;
  assign n45641 = pi20 ? n40430 : n139;
  assign n45642 = pi19 ? n45641 : n139;
  assign n45643 = pi18 ? n33792 : n45642;
  assign n45644 = pi21 ? n6461 : n37547;
  assign n45645 = pi20 ? n685 : n45644;
  assign n45646 = pi19 ? n45645 : n32;
  assign n45647 = pi18 ? n45152 : n45646;
  assign n45648 = pi17 ? n45643 : n45647;
  assign n45649 = pi16 ? n45640 : n45648;
  assign n45650 = pi15 ? n45633 : n45649;
  assign n45651 = pi14 ? n45619 : n45650;
  assign n45652 = pi23 ? n32 : n36830;
  assign n45653 = pi22 ? n32 : n45652;
  assign n45654 = pi21 ? n45653 : n36798;
  assign n45655 = pi20 ? n32 : n45654;
  assign n45656 = pi19 ? n32 : n45655;
  assign n45657 = pi18 ? n45656 : n45166;
  assign n45658 = pi17 ? n32 : n45657;
  assign n45659 = pi19 ? n41583 : n335;
  assign n45660 = pi18 ? n41580 : n45659;
  assign n45661 = pi17 ? n45660 : n45177;
  assign n45662 = pi16 ? n45658 : n45661;
  assign n45663 = pi21 ? n32 : n45136;
  assign n45664 = pi20 ? n32 : n45663;
  assign n45665 = pi19 ? n32 : n45664;
  assign n45666 = pi18 ? n45665 : n45181;
  assign n45667 = pi17 ? n32 : n45666;
  assign n45668 = pi16 ? n45667 : n45193;
  assign n45669 = pi15 ? n45662 : n45668;
  assign n45670 = pi21 ? n32 : n45161;
  assign n45671 = pi20 ? n32 : n45670;
  assign n45672 = pi19 ? n32 : n45671;
  assign n45673 = pi18 ? n45672 : n41136;
  assign n45674 = pi17 ? n32 : n45673;
  assign n45675 = pi23 ? n335 : n36798;
  assign n45676 = pi22 ? n36798 : n45675;
  assign n45677 = pi21 ? n45676 : n36837;
  assign n45678 = pi20 ? n45677 : n157;
  assign n45679 = pi19 ? n45678 : n157;
  assign n45680 = pi18 ? n45198 : n45679;
  assign n45681 = pi22 ? n157 : n1457;
  assign n45682 = pi21 ? n45681 : n882;
  assign n45683 = pi20 ? n157 : n45682;
  assign n45684 = pi19 ? n45683 : n32;
  assign n45685 = pi18 ? n157 : n45684;
  assign n45686 = pi17 ? n45680 : n45685;
  assign n45687 = pi16 ? n45674 : n45686;
  assign n45688 = pi18 ? n45665 : n36781;
  assign n45689 = pi17 ? n32 : n45688;
  assign n45690 = pi21 ? n36798 : n5054;
  assign n45691 = pi20 ? n45690 : n157;
  assign n45692 = pi19 ? n45691 : n157;
  assign n45693 = pi18 ? n45198 : n45692;
  assign n45694 = pi20 ? n157 : n28024;
  assign n45695 = pi19 ? n45694 : n32;
  assign n45696 = pi18 ? n157 : n45695;
  assign n45697 = pi17 ? n45693 : n45696;
  assign n45698 = pi16 ? n45689 : n45697;
  assign n45699 = pi15 ? n45687 : n45698;
  assign n45700 = pi14 ? n45669 : n45699;
  assign n45701 = pi13 ? n45651 : n45700;
  assign n45702 = pi12 ? n45589 : n45701;
  assign n45703 = pi11 ? n45515 : n45702;
  assign n45704 = pi10 ? n45426 : n45703;
  assign n45705 = pi09 ? n45240 : n45704;
  assign n45706 = pi08 ? n45229 : n45705;
  assign n45707 = pi18 ? n40045 : n20563;
  assign n45708 = pi20 ? n5077 : n14844;
  assign n45709 = pi19 ? n32294 : n45708;
  assign n45710 = pi19 ? n99 : n14836;
  assign n45711 = pi18 ? n45709 : n45710;
  assign n45712 = pi17 ? n45707 : n45711;
  assign n45713 = pi16 ? n32 : n45712;
  assign n45714 = pi15 ? n32 : n45713;
  assign n45715 = pi18 ? n40550 : n20563;
  assign n45716 = pi21 ? n1698 : n820;
  assign n45717 = pi20 ? n45716 : n942;
  assign n45718 = pi20 ? n139 : n14835;
  assign n45719 = pi19 ? n45717 : n45718;
  assign n45720 = pi18 ? n32295 : n45719;
  assign n45721 = pi17 ? n45715 : n45720;
  assign n45722 = pi16 ? n32 : n45721;
  assign n45723 = pi20 ? n3096 : n14847;
  assign n45724 = pi19 ? n37 : n45723;
  assign n45725 = pi18 ? n32899 : n45724;
  assign n45726 = pi17 ? n20563 : n45725;
  assign n45727 = pi16 ? n45233 : n45726;
  assign n45728 = pi15 ? n45722 : n45727;
  assign n45729 = pi14 ? n45714 : n45728;
  assign n45730 = pi13 ? n32 : n45729;
  assign n45731 = pi12 ? n32 : n45730;
  assign n45732 = pi11 ? n32 : n45731;
  assign n45733 = pi10 ? n32 : n45732;
  assign n45734 = pi20 ? n3299 : n15978;
  assign n45735 = pi19 ? n37 : n45734;
  assign n45736 = pi18 ? n32349 : n45735;
  assign n45737 = pi17 ? n20563 : n45736;
  assign n45738 = pi16 ? n44635 : n45737;
  assign n45739 = pi18 ? n32 : n37935;
  assign n45740 = pi17 ? n32 : n45739;
  assign n45741 = pi20 ? n44673 : n15978;
  assign n45742 = pi19 ? n13125 : n45741;
  assign n45743 = pi18 ? n32899 : n45742;
  assign n45744 = pi17 ? n20563 : n45743;
  assign n45745 = pi16 ? n45740 : n45744;
  assign n45746 = pi15 ? n45738 : n45745;
  assign n45747 = pi20 ? n29210 : n2470;
  assign n45748 = pi19 ? n13148 : n45747;
  assign n45749 = pi18 ? n31939 : n45748;
  assign n45750 = pi17 ? n20563 : n45749;
  assign n45751 = pi16 ? n44653 : n45750;
  assign n45752 = pi18 ? n17061 : n45249;
  assign n45753 = pi17 ? n20563 : n45752;
  assign n45754 = pi16 ? n44223 : n45753;
  assign n45755 = pi15 ? n45751 : n45754;
  assign n45756 = pi14 ? n45746 : n45755;
  assign n45757 = pi20 ? n37 : n3922;
  assign n45758 = pi19 ? n30097 : n45757;
  assign n45759 = pi20 ? n3092 : n2512;
  assign n45760 = pi19 ? n45759 : n16100;
  assign n45761 = pi18 ? n45758 : n45760;
  assign n45762 = pi17 ? n20563 : n45761;
  assign n45763 = pi16 ? n44671 : n45762;
  assign n45764 = pi21 ? n3668 : n3073;
  assign n45765 = pi20 ? n376 : n45764;
  assign n45766 = pi21 ? n297 : n14952;
  assign n45767 = pi20 ? n45766 : n32;
  assign n45768 = pi19 ? n45765 : n45767;
  assign n45769 = pi18 ? n31939 : n45768;
  assign n45770 = pi17 ? n20563 : n45769;
  assign n45771 = pi16 ? n43675 : n45770;
  assign n45772 = pi15 ? n45763 : n45771;
  assign n45773 = pi17 ? n20563 : n45276;
  assign n45774 = pi16 ? n43685 : n45773;
  assign n45775 = pi18 ? n20563 : n35777;
  assign n45776 = pi21 ? n37 : n13253;
  assign n45777 = pi20 ? n45776 : n32;
  assign n45778 = pi19 ? n37 : n45777;
  assign n45779 = pi18 ? n37 : n45778;
  assign n45780 = pi17 ? n45775 : n45779;
  assign n45781 = pi16 ? n44688 : n45780;
  assign n45782 = pi15 ? n45774 : n45781;
  assign n45783 = pi14 ? n45772 : n45782;
  assign n45784 = pi13 ? n45756 : n45783;
  assign n45785 = pi20 ? n19934 : n32;
  assign n45786 = pi19 ? n7676 : n45785;
  assign n45787 = pi18 ? n37 : n45786;
  assign n45788 = pi17 ? n42647 : n45787;
  assign n45789 = pi16 ? n44688 : n45788;
  assign n45790 = pi22 ? n335 : n19177;
  assign n45791 = pi21 ? n37 : n45790;
  assign n45792 = pi20 ? n45791 : n32;
  assign n45793 = pi19 ? n7676 : n45792;
  assign n45794 = pi18 ? n37 : n45793;
  assign n45795 = pi17 ? n44680 : n45794;
  assign n45796 = pi16 ? n42682 : n45795;
  assign n45797 = pi15 ? n45789 : n45796;
  assign n45798 = pi19 ? n37 : n33694;
  assign n45799 = pi21 ? n583 : n4975;
  assign n45800 = pi20 ? n4951 : n45799;
  assign n45801 = pi21 ? n570 : n9900;
  assign n45802 = pi20 ? n45801 : n32;
  assign n45803 = pi19 ? n45800 : n45802;
  assign n45804 = pi18 ? n45798 : n45803;
  assign n45805 = pi17 ? n42657 : n45804;
  assign n45806 = pi16 ? n42682 : n45805;
  assign n45807 = pi21 ? n583 : n4938;
  assign n45808 = pi20 ? n4951 : n45807;
  assign n45809 = pi22 ? n335 : n1150;
  assign n45810 = pi21 ? n570 : n45809;
  assign n45811 = pi20 ? n45810 : n32;
  assign n45812 = pi19 ? n45808 : n45811;
  assign n45813 = pi18 ? n37 : n45812;
  assign n45814 = pi17 ? n42657 : n45813;
  assign n45815 = pi16 ? n42682 : n45814;
  assign n45816 = pi15 ? n45806 : n45815;
  assign n45817 = pi14 ? n45797 : n45816;
  assign n45818 = pi21 ? n570 : n45310;
  assign n45819 = pi20 ? n45818 : n32;
  assign n45820 = pi19 ? n12440 : n45819;
  assign n45821 = pi18 ? n37 : n45820;
  assign n45822 = pi17 ? n42657 : n45821;
  assign n45823 = pi16 ? n42195 : n45822;
  assign n45824 = pi20 ? n31770 : n32;
  assign n45825 = pi19 ? n37 : n45824;
  assign n45826 = pi18 ? n37 : n45825;
  assign n45827 = pi17 ? n42663 : n45826;
  assign n45828 = pi16 ? n41643 : n45827;
  assign n45829 = pi15 ? n45823 : n45828;
  assign n45830 = pi21 ? n37 : n41110;
  assign n45831 = pi20 ? n45830 : n32;
  assign n45832 = pi19 ? n37 : n45831;
  assign n45833 = pi18 ? n37 : n45832;
  assign n45834 = pi17 ? n42663 : n45833;
  assign n45835 = pi16 ? n42701 : n45834;
  assign n45836 = pi20 ? n31465 : n32;
  assign n45837 = pi19 ? n37 : n45836;
  assign n45838 = pi18 ? n37 : n45837;
  assign n45839 = pi17 ? n42663 : n45838;
  assign n45840 = pi16 ? n42701 : n45839;
  assign n45841 = pi15 ? n45835 : n45840;
  assign n45842 = pi14 ? n45829 : n45841;
  assign n45843 = pi13 ? n45817 : n45842;
  assign n45844 = pi12 ? n45784 : n45843;
  assign n45845 = pi21 ? n37 : n17284;
  assign n45846 = pi20 ? n45845 : n32;
  assign n45847 = pi19 ? n37 : n45846;
  assign n45848 = pi18 ? n37 : n45847;
  assign n45849 = pi17 ? n44732 : n45848;
  assign n45850 = pi16 ? n41159 : n45849;
  assign n45851 = pi20 ? n37 : n27484;
  assign n45852 = pi21 ? n363 : n2139;
  assign n45853 = pi20 ? n45852 : n32;
  assign n45854 = pi19 ? n45851 : n45853;
  assign n45855 = pi18 ? n6404 : n45854;
  assign n45856 = pi17 ? n42663 : n45855;
  assign n45857 = pi16 ? n41159 : n45856;
  assign n45858 = pi15 ? n45850 : n45857;
  assign n45859 = pi21 ? n363 : n2193;
  assign n45860 = pi20 ? n45859 : n32;
  assign n45861 = pi19 ? n45851 : n45860;
  assign n45862 = pi18 ? n6404 : n45861;
  assign n45863 = pi17 ? n42690 : n45862;
  assign n45864 = pi16 ? n41159 : n45863;
  assign n45865 = pi19 ? n37 : n45860;
  assign n45866 = pi18 ? n6404 : n45865;
  assign n45867 = pi17 ? n42690 : n45866;
  assign n45868 = pi16 ? n41170 : n45867;
  assign n45869 = pi15 ? n45864 : n45868;
  assign n45870 = pi14 ? n45858 : n45869;
  assign n45871 = pi20 ? n29373 : n32;
  assign n45872 = pi19 ? n37 : n45871;
  assign n45873 = pi18 ? n37 : n45872;
  assign n45874 = pi17 ? n42690 : n45873;
  assign n45875 = pi16 ? n40025 : n45874;
  assign n45876 = pi17 ? n42663 : n45873;
  assign n45877 = pi16 ? n40025 : n45876;
  assign n45878 = pi15 ? n45875 : n45877;
  assign n45879 = pi19 ? n37 : n16246;
  assign n45880 = pi18 ? n37 : n45879;
  assign n45881 = pi17 ? n41633 : n45880;
  assign n45882 = pi16 ? n40499 : n45881;
  assign n45883 = pi16 ? n41684 : n45881;
  assign n45884 = pi15 ? n45882 : n45883;
  assign n45885 = pi14 ? n45878 : n45884;
  assign n45886 = pi13 ? n45870 : n45885;
  assign n45887 = pi19 ? n37 : n12376;
  assign n45888 = pi18 ? n37 : n45887;
  assign n45889 = pi17 ? n41672 : n45888;
  assign n45890 = pi16 ? n40512 : n45889;
  assign n45891 = pi17 ? n41644 : n45888;
  assign n45892 = pi16 ? n40512 : n45891;
  assign n45893 = pi15 ? n45890 : n45892;
  assign n45894 = pi19 ? n32294 : n35209;
  assign n45895 = pi18 ? n20563 : n45894;
  assign n45896 = pi21 ? n99 : n3523;
  assign n45897 = pi20 ? n45896 : n32;
  assign n45898 = pi19 ? n99 : n45897;
  assign n45899 = pi18 ? n34567 : n45898;
  assign n45900 = pi17 ? n45895 : n45899;
  assign n45901 = pi16 ? n40512 : n45900;
  assign n45902 = pi18 ? n20563 : n38094;
  assign n45903 = pi18 ? n99 : n45898;
  assign n45904 = pi17 ? n45902 : n45903;
  assign n45905 = pi16 ? n41710 : n45904;
  assign n45906 = pi15 ? n45901 : n45905;
  assign n45907 = pi14 ? n45893 : n45906;
  assign n45908 = pi19 ? n32898 : n18853;
  assign n45909 = pi18 ? n20563 : n45908;
  assign n45910 = pi21 ? n22940 : n2320;
  assign n45911 = pi20 ? n45910 : n32;
  assign n45912 = pi19 ? n99 : n45911;
  assign n45913 = pi18 ? n99 : n45912;
  assign n45914 = pi17 ? n45909 : n45913;
  assign n45915 = pi16 ? n41710 : n45914;
  assign n45916 = pi18 ? n20563 : n37559;
  assign n45917 = pi21 ? n3562 : n31963;
  assign n45918 = pi20 ? n45917 : n32;
  assign n45919 = pi19 ? n19134 : n45918;
  assign n45920 = pi18 ? n99 : n45919;
  assign n45921 = pi17 ? n45916 : n45920;
  assign n45922 = pi16 ? n41710 : n45921;
  assign n45923 = pi15 ? n45915 : n45922;
  assign n45924 = pi19 ? n33923 : n99;
  assign n45925 = pi18 ? n20563 : n45924;
  assign n45926 = pi21 ? n157 : n3302;
  assign n45927 = pi20 ? n45926 : n32;
  assign n45928 = pi19 ? n34498 : n45927;
  assign n45929 = pi18 ? n19124 : n45928;
  assign n45930 = pi17 ? n45925 : n45929;
  assign n45931 = pi16 ? n41710 : n45930;
  assign n45932 = pi19 ? n32348 : n21611;
  assign n45933 = pi18 ? n20563 : n45932;
  assign n45934 = pi21 ? n204 : n21929;
  assign n45935 = pi20 ? n42885 : n45934;
  assign n45936 = pi21 ? n316 : n3302;
  assign n45937 = pi20 ? n45936 : n32;
  assign n45938 = pi19 ? n45935 : n45937;
  assign n45939 = pi18 ? n99 : n45938;
  assign n45940 = pi17 ? n45933 : n45939;
  assign n45941 = pi16 ? n45368 : n45940;
  assign n45942 = pi15 ? n45931 : n45941;
  assign n45943 = pi14 ? n45923 : n45942;
  assign n45944 = pi13 ? n45907 : n45943;
  assign n45945 = pi12 ? n45886 : n45944;
  assign n45946 = pi11 ? n45844 : n45945;
  assign n45947 = pi21 ? n29133 : n181;
  assign n45948 = pi20 ? n20563 : n45947;
  assign n45949 = pi20 ? n5077 : n219;
  assign n45950 = pi19 ? n45948 : n45949;
  assign n45951 = pi18 ? n20563 : n45950;
  assign n45952 = pi20 ? n42885 : n22965;
  assign n45953 = pi19 ? n45952 : n17867;
  assign n45954 = pi18 ? n99 : n45953;
  assign n45955 = pi17 ? n45951 : n45954;
  assign n45956 = pi16 ? n39399 : n45955;
  assign n45957 = pi21 ? n30843 : n99;
  assign n45958 = pi20 ? n20563 : n45957;
  assign n45959 = pi19 ? n45958 : n25381;
  assign n45960 = pi18 ? n20563 : n45959;
  assign n45961 = pi19 ? n27596 : n9756;
  assign n45962 = pi18 ? n44885 : n45961;
  assign n45963 = pi17 ? n45960 : n45962;
  assign n45964 = pi16 ? n39399 : n45963;
  assign n45965 = pi15 ? n45956 : n45964;
  assign n45966 = pi19 ? n2862 : n19691;
  assign n45967 = pi18 ? n44893 : n45966;
  assign n45968 = pi17 ? n41685 : n45967;
  assign n45969 = pi16 ? n39399 : n45968;
  assign n45970 = pi18 ? n18083 : n45448;
  assign n45971 = pi17 ? n45359 : n45970;
  assign n45972 = pi16 ? n40552 : n45971;
  assign n45973 = pi15 ? n45969 : n45972;
  assign n45974 = pi14 ? n45965 : n45973;
  assign n45975 = pi18 ? n20563 : n41929;
  assign n45976 = pi17 ? n45975 : n45449;
  assign n45977 = pi16 ? n45415 : n45976;
  assign n45978 = pi19 ? n32348 : n9814;
  assign n45979 = pi18 ? n20563 : n45978;
  assign n45980 = pi21 ? n3763 : n37639;
  assign n45981 = pi20 ? n45980 : n32;
  assign n45982 = pi19 ? n36541 : n45981;
  assign n45983 = pi18 ? n139 : n45982;
  assign n45984 = pi17 ? n45979 : n45983;
  assign n45985 = pi16 ? n45415 : n45984;
  assign n45986 = pi15 ? n45977 : n45985;
  assign n45987 = pi17 ? n45979 : n45463;
  assign n45988 = pi16 ? n45415 : n45987;
  assign n45989 = pi18 ? n20563 : n38140;
  assign n45990 = pi20 ? n21338 : n32;
  assign n45991 = pi19 ? n36541 : n45990;
  assign n45992 = pi18 ? n139 : n45991;
  assign n45993 = pi17 ? n45989 : n45992;
  assign n45994 = pi16 ? n45415 : n45993;
  assign n45995 = pi15 ? n45988 : n45994;
  assign n45996 = pi14 ? n45986 : n45995;
  assign n45997 = pi13 ? n45974 : n45996;
  assign n45998 = pi20 ? n8729 : n8731;
  assign n45999 = pi19 ? n36362 : n45998;
  assign n46000 = pi18 ? n20563 : n45999;
  assign n46001 = pi23 ? n233 : n139;
  assign n46002 = pi22 ? n46001 : n139;
  assign n46003 = pi21 ? n139 : n46002;
  assign n46004 = pi20 ? n139 : n46003;
  assign n46005 = pi19 ? n46004 : n10298;
  assign n46006 = pi18 ? n139 : n46005;
  assign n46007 = pi17 ? n46000 : n46006;
  assign n46008 = pi16 ? n38318 : n46007;
  assign n46009 = pi20 ? n34919 : n3086;
  assign n46010 = pi19 ? n46009 : n9769;
  assign n46011 = pi18 ? n20563 : n46010;
  assign n46012 = pi22 ? n6833 : n6415;
  assign n46013 = pi21 ? n46012 : n32;
  assign n46014 = pi20 ? n46013 : n32;
  assign n46015 = pi19 ? n139 : n46014;
  assign n46016 = pi18 ? n139 : n46015;
  assign n46017 = pi17 ? n46011 : n46016;
  assign n46018 = pi16 ? n38318 : n46017;
  assign n46019 = pi15 ? n46008 : n46018;
  assign n46020 = pi21 ? n335 : n4903;
  assign n46021 = pi20 ? n335 : n46020;
  assign n46022 = pi19 ? n46021 : n9432;
  assign n46023 = pi18 ? n10682 : n46022;
  assign n46024 = pi17 ? n41178 : n46023;
  assign n46025 = pi16 ? n38985 : n46024;
  assign n46026 = pi19 ? n37 : n27685;
  assign n46027 = pi19 ? n233 : n16945;
  assign n46028 = pi18 ? n46026 : n46027;
  assign n46029 = pi17 ? n41178 : n46028;
  assign n46030 = pi16 ? n38985 : n46029;
  assign n46031 = pi15 ? n46025 : n46030;
  assign n46032 = pi14 ? n46019 : n46031;
  assign n46033 = pi20 ? n649 : n233;
  assign n46034 = pi19 ? n37 : n46033;
  assign n46035 = pi20 ? n233 : n6361;
  assign n46036 = pi19 ? n46035 : n8918;
  assign n46037 = pi18 ? n46034 : n46036;
  assign n46038 = pi17 ? n44335 : n46037;
  assign n46039 = pi16 ? n40058 : n46038;
  assign n46040 = pi22 ? n40387 : n112;
  assign n46041 = pi21 ? n20563 : n46040;
  assign n46042 = pi20 ? n46041 : n2973;
  assign n46043 = pi19 ? n46042 : n37;
  assign n46044 = pi18 ? n20563 : n46043;
  assign n46045 = pi20 ? n29667 : n233;
  assign n46046 = pi19 ? n37 : n46045;
  assign n46047 = pi19 ? n233 : n15891;
  assign n46048 = pi18 ? n46046 : n46047;
  assign n46049 = pi17 ? n46044 : n46048;
  assign n46050 = pi16 ? n40058 : n46049;
  assign n46051 = pi15 ? n46039 : n46050;
  assign n46052 = pi20 ? n40919 : n37;
  assign n46053 = pi19 ? n46052 : n37;
  assign n46054 = pi18 ? n20563 : n46053;
  assign n46055 = pi20 ? n20391 : n32;
  assign n46056 = pi19 ? n7981 : n46055;
  assign n46057 = pi18 ? n16209 : n46056;
  assign n46058 = pi17 ? n46054 : n46057;
  assign n46059 = pi16 ? n37937 : n46058;
  assign n46060 = pi22 ? n32 : n30868;
  assign n46061 = pi21 ? n32 : n46060;
  assign n46062 = pi20 ? n32 : n46061;
  assign n46063 = pi19 ? n32 : n46062;
  assign n46064 = pi18 ? n46063 : n42015;
  assign n46065 = pi17 ? n32 : n46064;
  assign n46066 = pi22 ? n1070 : n14363;
  assign n46067 = pi21 ? n46066 : n32;
  assign n46068 = pi20 ? n46067 : n32;
  assign n46069 = pi19 ? n32703 : n46068;
  assign n46070 = pi18 ? n15161 : n46069;
  assign n46071 = pi17 ? n46054 : n46070;
  assign n46072 = pi16 ? n46065 : n46071;
  assign n46073 = pi15 ? n46059 : n46072;
  assign n46074 = pi14 ? n46051 : n46073;
  assign n46075 = pi13 ? n46032 : n46074;
  assign n46076 = pi12 ? n45997 : n46075;
  assign n46077 = pi21 ? n32 : n45517;
  assign n46078 = pi20 ? n32 : n46077;
  assign n46079 = pi19 ? n32 : n46078;
  assign n46080 = pi18 ? n46079 : n33792;
  assign n46081 = pi17 ? n32 : n46080;
  assign n46082 = pi21 ? n33792 : n45016;
  assign n46083 = pi20 ? n33792 : n46082;
  assign n46084 = pi18 ? n46083 : n46053;
  assign n46085 = pi20 ? n37 : n31764;
  assign n46086 = pi19 ? n37 : n46085;
  assign n46087 = pi19 ? n45022 : n6418;
  assign n46088 = pi18 ? n46086 : n46087;
  assign n46089 = pi17 ? n46084 : n46088;
  assign n46090 = pi16 ? n46081 : n46089;
  assign n46091 = pi19 ? n33846 : n335;
  assign n46092 = pi18 ? n20563 : n46091;
  assign n46093 = pi21 ? n335 : n29868;
  assign n46094 = pi20 ? n335 : n46093;
  assign n46095 = pi19 ? n46094 : n3341;
  assign n46096 = pi18 ? n335 : n46095;
  assign n46097 = pi17 ? n46092 : n46096;
  assign n46098 = pi16 ? n37337 : n46097;
  assign n46099 = pi15 ? n46090 : n46098;
  assign n46100 = pi21 ? n37 : n25347;
  assign n46101 = pi20 ? n37 : n46100;
  assign n46102 = pi19 ? n46101 : n2639;
  assign n46103 = pi18 ? n45034 : n46102;
  assign n46104 = pi17 ? n41699 : n46103;
  assign n46105 = pi16 ? n37337 : n46104;
  assign n46106 = pi23 ? n11910 : n363;
  assign n46107 = pi22 ? n46106 : n2244;
  assign n46108 = pi21 ? n37 : n46107;
  assign n46109 = pi20 ? n37 : n46108;
  assign n46110 = pi19 ? n46109 : n2654;
  assign n46111 = pi18 ? n45034 : n46110;
  assign n46112 = pi17 ? n41699 : n46111;
  assign n46113 = pi16 ? n37337 : n46112;
  assign n46114 = pi15 ? n46105 : n46113;
  assign n46115 = pi14 ? n46099 : n46114;
  assign n46116 = pi22 ? n39190 : n20563;
  assign n46117 = pi21 ? n46116 : n31885;
  assign n46118 = pi20 ? n46117 : n16008;
  assign n46119 = pi20 ? n10496 : n9660;
  assign n46120 = pi19 ? n46118 : n46119;
  assign n46121 = pi18 ? n20563 : n46120;
  assign n46122 = pi20 ? n15173 : n16188;
  assign n46123 = pi20 ? n39902 : n3392;
  assign n46124 = pi19 ? n46122 : n46123;
  assign n46125 = pi19 ? n45057 : n2654;
  assign n46126 = pi18 ? n46124 : n46125;
  assign n46127 = pi17 ? n46121 : n46126;
  assign n46128 = pi16 ? n36871 : n46127;
  assign n46129 = pi21 ? n46116 : n30195;
  assign n46130 = pi20 ? n46129 : n14887;
  assign n46131 = pi19 ? n46130 : n43075;
  assign n46132 = pi18 ? n20563 : n46131;
  assign n46133 = pi21 ? n2106 : n2768;
  assign n46134 = pi20 ? n22881 : n46133;
  assign n46135 = pi19 ? n46134 : n1823;
  assign n46136 = pi18 ? n45065 : n46135;
  assign n46137 = pi17 ? n46132 : n46136;
  assign n46138 = pi16 ? n36871 : n46137;
  assign n46139 = pi15 ? n46128 : n46138;
  assign n46140 = pi21 ? n37768 : n31924;
  assign n46141 = pi20 ? n46140 : n13613;
  assign n46142 = pi19 ? n46141 : n37;
  assign n46143 = pi18 ? n20563 : n46142;
  assign n46144 = pi17 ? n46143 : n45576;
  assign n46145 = pi16 ? n36871 : n46144;
  assign n46146 = pi19 ? n39867 : n37753;
  assign n46147 = pi21 ? n685 : n38878;
  assign n46148 = pi20 ? n24220 : n46147;
  assign n46149 = pi19 ? n46148 : n32;
  assign n46150 = pi18 ? n46146 : n46149;
  assign n46151 = pi17 ? n46143 : n46150;
  assign n46152 = pi16 ? n36871 : n46151;
  assign n46153 = pi15 ? n46145 : n46152;
  assign n46154 = pi14 ? n46139 : n46153;
  assign n46155 = pi13 ? n46115 : n46154;
  assign n46156 = pi21 ? n37784 : n31924;
  assign n46157 = pi20 ? n46156 : n3292;
  assign n46158 = pi19 ? n46157 : n45097;
  assign n46159 = pi18 ? n20563 : n46158;
  assign n46160 = pi20 ? n685 : n2782;
  assign n46161 = pi19 ? n46160 : n32;
  assign n46162 = pi18 ? n45100 : n46161;
  assign n46163 = pi17 ? n46159 : n46162;
  assign n46164 = pi16 ? n36871 : n46163;
  assign n46165 = pi23 ? n32 : n34196;
  assign n46166 = pi22 ? n46165 : n30868;
  assign n46167 = pi21 ? n32 : n46166;
  assign n46168 = pi20 ? n32 : n46167;
  assign n46169 = pi19 ? n32 : n46168;
  assign n46170 = pi18 ? n46169 : n30868;
  assign n46171 = pi17 ? n32 : n46170;
  assign n46172 = pi23 ? n30868 : n36659;
  assign n46173 = pi22 ? n46172 : n30868;
  assign n46174 = pi21 ? n46173 : n37810;
  assign n46175 = pi21 ? n4538 : n363;
  assign n46176 = pi20 ? n46174 : n46175;
  assign n46177 = pi19 ? n46176 : n34796;
  assign n46178 = pi18 ? n30868 : n46177;
  assign n46179 = pi22 ? n685 : n19696;
  assign n46180 = pi21 ? n363 : n46179;
  assign n46181 = pi20 ? n26891 : n46180;
  assign n46182 = pi19 ? n46181 : n32;
  assign n46183 = pi18 ? n45115 : n46182;
  assign n46184 = pi17 ? n46178 : n46183;
  assign n46185 = pi16 ? n46171 : n46184;
  assign n46186 = pi15 ? n46164 : n46185;
  assign n46187 = pi22 ? n45597 : n30868;
  assign n46188 = pi21 ? n32 : n46187;
  assign n46189 = pi20 ? n32 : n46188;
  assign n46190 = pi19 ? n32 : n46189;
  assign n46191 = pi18 ? n46190 : n30868;
  assign n46192 = pi17 ? n32 : n46191;
  assign n46193 = pi19 ? n39928 : n99;
  assign n46194 = pi18 ? n30868 : n46193;
  assign n46195 = pi19 ? n5086 : n685;
  assign n46196 = pi20 ? n99 : n41526;
  assign n46197 = pi19 ? n46196 : n32;
  assign n46198 = pi18 ? n46195 : n46197;
  assign n46199 = pi17 ? n46194 : n46198;
  assign n46200 = pi16 ? n46192 : n46199;
  assign n46201 = pi21 ? n32 : n45635;
  assign n46202 = pi20 ? n32 : n46201;
  assign n46203 = pi19 ? n32 : n46202;
  assign n46204 = pi20 ? n36798 : n33792;
  assign n46205 = pi19 ? n45141 : n46204;
  assign n46206 = pi18 ? n46203 : n46205;
  assign n46207 = pi17 ? n32 : n46206;
  assign n46208 = pi19 ? n44582 : n139;
  assign n46209 = pi18 ? n33792 : n46208;
  assign n46210 = pi22 ? n44163 : n139;
  assign n46211 = pi21 ? n46210 : n139;
  assign n46212 = pi22 ? n316 : n3472;
  assign n46213 = pi21 ? n316 : n46212;
  assign n46214 = pi20 ? n46211 : n46213;
  assign n46215 = pi19 ? n139 : n46214;
  assign n46216 = pi21 ? n44169 : n139;
  assign n46217 = pi21 ? n157 : n3494;
  assign n46218 = pi20 ? n46216 : n46217;
  assign n46219 = pi19 ? n46218 : n32;
  assign n46220 = pi18 ? n46215 : n46219;
  assign n46221 = pi17 ? n46209 : n46220;
  assign n46222 = pi16 ? n46207 : n46221;
  assign n46223 = pi15 ? n46200 : n46222;
  assign n46224 = pi14 ? n46186 : n46223;
  assign n46225 = pi21 ? n32 : n45653;
  assign n46226 = pi20 ? n32 : n46225;
  assign n46227 = pi19 ? n32 : n46226;
  assign n46228 = pi19 ? n36798 : n43139;
  assign n46229 = pi18 ? n46227 : n46228;
  assign n46230 = pi17 ? n32 : n46229;
  assign n46231 = pi19 ? n44592 : n335;
  assign n46232 = pi18 ? n41580 : n46231;
  assign n46233 = pi20 ? n880 : n316;
  assign n46234 = pi19 ? n139 : n46233;
  assign n46235 = pi20 ? n249 : n18285;
  assign n46236 = pi19 ? n46235 : n32;
  assign n46237 = pi18 ? n46234 : n46236;
  assign n46238 = pi17 ? n46232 : n46237;
  assign n46239 = pi16 ? n46230 : n46238;
  assign n46240 = pi18 ? n46203 : n45181;
  assign n46241 = pi17 ? n32 : n46240;
  assign n46242 = pi21 ? n42146 : n36659;
  assign n46243 = pi22 ? n36710 : n335;
  assign n46244 = pi21 ? n46243 : n335;
  assign n46245 = pi20 ? n46242 : n46244;
  assign n46246 = pi19 ? n46245 : n335;
  assign n46247 = pi18 ? n41103 : n46246;
  assign n46248 = pi21 ? n3693 : n335;
  assign n46249 = pi20 ? n46248 : n17366;
  assign n46250 = pi20 ? n157 : n3562;
  assign n46251 = pi19 ? n46249 : n46250;
  assign n46252 = pi20 ? n17390 : n3619;
  assign n46253 = pi19 ? n46252 : n32;
  assign n46254 = pi18 ? n46251 : n46253;
  assign n46255 = pi17 ? n46247 : n46254;
  assign n46256 = pi16 ? n46241 : n46255;
  assign n46257 = pi15 ? n46239 : n46256;
  assign n46258 = pi18 ? n46227 : n41136;
  assign n46259 = pi17 ? n32 : n46258;
  assign n46260 = pi22 ? n36659 : n36798;
  assign n46261 = pi21 ? n37899 : n46260;
  assign n46262 = pi22 ? n36798 : n36710;
  assign n46263 = pi21 ? n46262 : n34833;
  assign n46264 = pi20 ? n46261 : n46263;
  assign n46265 = pi19 ? n46264 : n157;
  assign n46266 = pi18 ? n45198 : n46265;
  assign n46267 = pi22 ? n157 : n18448;
  assign n46268 = pi21 ? n46267 : n882;
  assign n46269 = pi20 ? n157 : n46268;
  assign n46270 = pi19 ? n46269 : n32;
  assign n46271 = pi18 ? n157 : n46270;
  assign n46272 = pi17 ? n46266 : n46271;
  assign n46273 = pi16 ? n46259 : n46272;
  assign n46274 = pi24 ? n32 : n43198;
  assign n46275 = pi23 ? n32 : n46274;
  assign n46276 = pi22 ? n32 : n46275;
  assign n46277 = pi21 ? n32 : n46276;
  assign n46278 = pi20 ? n32 : n46277;
  assign n46279 = pi19 ? n32 : n46278;
  assign n46280 = pi22 ? n43198 : n36781;
  assign n46281 = pi21 ? n43198 : n46280;
  assign n46282 = pi20 ? n43198 : n46281;
  assign n46283 = pi22 ? n36781 : n43198;
  assign n46284 = pi21 ? n46283 : n43198;
  assign n46285 = pi20 ? n46284 : n36781;
  assign n46286 = pi19 ? n46282 : n46285;
  assign n46287 = pi18 ? n46279 : n46286;
  assign n46288 = pi17 ? n32 : n46287;
  assign n46289 = pi21 ? n38901 : n39972;
  assign n46290 = pi20 ? n46289 : n43204;
  assign n46291 = pi19 ? n46290 : n157;
  assign n46292 = pi18 ? n45198 : n46291;
  assign n46293 = pi17 ? n46292 : n45696;
  assign n46294 = pi16 ? n46288 : n46293;
  assign n46295 = pi15 ? n46273 : n46294;
  assign n46296 = pi14 ? n46257 : n46295;
  assign n46297 = pi13 ? n46224 : n46296;
  assign n46298 = pi12 ? n46155 : n46297;
  assign n46299 = pi11 ? n46076 : n46298;
  assign n46300 = pi10 ? n45946 : n46299;
  assign n46301 = pi09 ? n45733 : n46300;
  assign n46302 = pi18 ? n40532 : n20563;
  assign n46303 = pi17 ? n46302 : n45711;
  assign n46304 = pi16 ? n32 : n46303;
  assign n46305 = pi15 ? n32 : n46304;
  assign n46306 = pi21 ? n3073 : n820;
  assign n46307 = pi20 ? n46306 : n942;
  assign n46308 = pi19 ? n46307 : n45718;
  assign n46309 = pi18 ? n32295 : n46308;
  assign n46310 = pi17 ? n45715 : n46309;
  assign n46311 = pi16 ? n32 : n46310;
  assign n46312 = pi18 ? n38316 : n20563;
  assign n46313 = pi18 ? n45335 : n45724;
  assign n46314 = pi17 ? n46312 : n46313;
  assign n46315 = pi16 ? n32 : n46314;
  assign n46316 = pi15 ? n46311 : n46315;
  assign n46317 = pi14 ? n46305 : n46316;
  assign n46318 = pi13 ? n32 : n46317;
  assign n46319 = pi12 ? n32 : n46318;
  assign n46320 = pi11 ? n32 : n46319;
  assign n46321 = pi10 ? n32 : n46320;
  assign n46322 = pi18 ? n37981 : n45735;
  assign n46323 = pi17 ? n20563 : n46322;
  assign n46324 = pi16 ? n32 : n46323;
  assign n46325 = pi18 ? n32 : n37928;
  assign n46326 = pi17 ? n32 : n46325;
  assign n46327 = pi18 ? n33906 : n45742;
  assign n46328 = pi17 ? n20563 : n46327;
  assign n46329 = pi16 ? n46326 : n46328;
  assign n46330 = pi15 ? n46324 : n46329;
  assign n46331 = pi20 ? n36929 : n36885;
  assign n46332 = pi19 ? n46331 : n37;
  assign n46333 = pi18 ? n46332 : n45748;
  assign n46334 = pi17 ? n20563 : n46333;
  assign n46335 = pi16 ? n44635 : n46334;
  assign n46336 = pi19 ? n40347 : n9824;
  assign n46337 = pi20 ? n1794 : n2554;
  assign n46338 = pi19 ? n22792 : n46337;
  assign n46339 = pi18 ? n46336 : n46338;
  assign n46340 = pi17 ? n20563 : n46339;
  assign n46341 = pi16 ? n44223 : n46340;
  assign n46342 = pi15 ? n46335 : n46341;
  assign n46343 = pi14 ? n46330 : n46342;
  assign n46344 = pi19 ? n33949 : n45757;
  assign n46345 = pi18 ? n46344 : n45760;
  assign n46346 = pi17 ? n20563 : n46345;
  assign n46347 = pi16 ? n45243 : n46346;
  assign n46348 = pi18 ? n32 : n39455;
  assign n46349 = pi17 ? n32 : n46348;
  assign n46350 = pi20 ? n942 : n2679;
  assign n46351 = pi19 ? n45765 : n46350;
  assign n46352 = pi18 ? n31939 : n46351;
  assign n46353 = pi17 ? n20563 : n46352;
  assign n46354 = pi16 ? n46349 : n46353;
  assign n46355 = pi15 ? n46347 : n46354;
  assign n46356 = pi20 ? n45273 : n2679;
  assign n46357 = pi19 ? n37 : n46356;
  assign n46358 = pi18 ? n37 : n46357;
  assign n46359 = pi17 ? n20563 : n46358;
  assign n46360 = pi16 ? n43664 : n46359;
  assign n46361 = pi20 ? n13273 : n2701;
  assign n46362 = pi19 ? n37 : n46361;
  assign n46363 = pi18 ? n37 : n46362;
  assign n46364 = pi17 ? n45775 : n46363;
  assign n46365 = pi16 ? n43664 : n46364;
  assign n46366 = pi15 ? n46360 : n46365;
  assign n46367 = pi14 ? n46355 : n46366;
  assign n46368 = pi13 ? n46343 : n46367;
  assign n46369 = pi20 ? n3299 : n2701;
  assign n46370 = pi19 ? n7676 : n46369;
  assign n46371 = pi18 ? n37 : n46370;
  assign n46372 = pi17 ? n44249 : n46371;
  assign n46373 = pi16 ? n44671 : n46372;
  assign n46374 = pi22 ? n335 : n11047;
  assign n46375 = pi21 ? n37 : n46374;
  assign n46376 = pi20 ? n46375 : n1822;
  assign n46377 = pi19 ? n7676 : n46376;
  assign n46378 = pi18 ? n37 : n46377;
  assign n46379 = pi17 ? n45246 : n46378;
  assign n46380 = pi16 ? n43224 : n46379;
  assign n46381 = pi15 ? n46373 : n46380;
  assign n46382 = pi20 ? n30300 : n1822;
  assign n46383 = pi19 ? n45800 : n46382;
  assign n46384 = pi18 ? n45798 : n46383;
  assign n46385 = pi17 ? n42657 : n46384;
  assign n46386 = pi16 ? n43228 : n46385;
  assign n46387 = pi20 ? n30300 : n32;
  assign n46388 = pi19 ? n45808 : n46387;
  assign n46389 = pi18 ? n37 : n46388;
  assign n46390 = pi17 ? n42657 : n46389;
  assign n46391 = pi16 ? n43249 : n46390;
  assign n46392 = pi15 ? n46386 : n46391;
  assign n46393 = pi14 ? n46381 : n46392;
  assign n46394 = pi20 ? n25146 : n32;
  assign n46395 = pi19 ? n12440 : n46394;
  assign n46396 = pi18 ? n37 : n46395;
  assign n46397 = pi17 ? n42657 : n46396;
  assign n46398 = pi16 ? n44275 : n46397;
  assign n46399 = pi16 ? n42202 : n45827;
  assign n46400 = pi15 ? n46398 : n46399;
  assign n46401 = pi20 ? n2729 : n32;
  assign n46402 = pi19 ? n37 : n46401;
  assign n46403 = pi18 ? n37 : n46402;
  assign n46404 = pi17 ? n43250 : n46403;
  assign n46405 = pi16 ? n43263 : n46404;
  assign n46406 = pi18 ? n20563 : n34891;
  assign n46407 = pi20 ? n2107 : n32;
  assign n46408 = pi19 ? n37 : n46407;
  assign n46409 = pi18 ? n37 : n46408;
  assign n46410 = pi17 ? n46406 : n46409;
  assign n46411 = pi16 ? n41632 : n46410;
  assign n46412 = pi15 ? n46405 : n46411;
  assign n46413 = pi14 ? n46400 : n46412;
  assign n46414 = pi13 ? n46393 : n46413;
  assign n46415 = pi12 ? n46368 : n46414;
  assign n46416 = pi22 ? n5011 : n1475;
  assign n46417 = pi21 ? n37 : n46416;
  assign n46418 = pi20 ? n46417 : n32;
  assign n46419 = pi19 ? n37 : n46418;
  assign n46420 = pi18 ? n37 : n46419;
  assign n46421 = pi17 ? n44732 : n46420;
  assign n46422 = pi16 ? n42689 : n46421;
  assign n46423 = pi16 ? n42689 : n45856;
  assign n46424 = pi15 ? n46422 : n46423;
  assign n46425 = pi16 ? n41643 : n45863;
  assign n46426 = pi17 ? n44280 : n45866;
  assign n46427 = pi16 ? n41643 : n46426;
  assign n46428 = pi15 ? n46425 : n46427;
  assign n46429 = pi14 ? n46424 : n46428;
  assign n46430 = pi17 ? n43257 : n45873;
  assign n46431 = pi16 ? n40487 : n46430;
  assign n46432 = pi16 ? n40487 : n45876;
  assign n46433 = pi15 ? n46431 : n46432;
  assign n46434 = pi17 ? n43264 : n45880;
  assign n46435 = pi16 ? n40487 : n46434;
  assign n46436 = pi16 ? n41159 : n45881;
  assign n46437 = pi15 ? n46435 : n46436;
  assign n46438 = pi14 ? n46433 : n46437;
  assign n46439 = pi13 ? n46429 : n46438;
  assign n46440 = pi17 ? n42224 : n45888;
  assign n46441 = pi16 ? n41170 : n46440;
  assign n46442 = pi18 ? n20563 : n34921;
  assign n46443 = pi17 ? n46442 : n45888;
  assign n46444 = pi16 ? n41170 : n46443;
  assign n46445 = pi15 ? n46441 : n46444;
  assign n46446 = pi19 ? n43672 : n20563;
  assign n46447 = pi18 ? n32 : n46446;
  assign n46448 = pi17 ? n32 : n46447;
  assign n46449 = pi20 ? n32591 : n32;
  assign n46450 = pi19 ? n99 : n46449;
  assign n46451 = pi18 ? n34567 : n46450;
  assign n46452 = pi17 ? n45895 : n46451;
  assign n46453 = pi16 ? n46448 : n46452;
  assign n46454 = pi19 ? n35854 : n21611;
  assign n46455 = pi18 ? n20563 : n46454;
  assign n46456 = pi18 ? n99 : n46450;
  assign n46457 = pi17 ? n46455 : n46456;
  assign n46458 = pi16 ? n40499 : n46457;
  assign n46459 = pi15 ? n46453 : n46458;
  assign n46460 = pi14 ? n46445 : n46459;
  assign n46461 = pi16 ? n40499 : n45914;
  assign n46462 = pi21 ? n3562 : n1485;
  assign n46463 = pi20 ? n46462 : n32;
  assign n46464 = pi19 ? n19134 : n46463;
  assign n46465 = pi18 ? n99 : n46464;
  assign n46466 = pi17 ? n45916 : n46465;
  assign n46467 = pi16 ? n40499 : n46466;
  assign n46468 = pi15 ? n46461 : n46467;
  assign n46469 = pi19 ? n32898 : n99;
  assign n46470 = pi18 ? n20563 : n46469;
  assign n46471 = pi21 ? n157 : n2300;
  assign n46472 = pi20 ? n46471 : n32;
  assign n46473 = pi19 ? n34498 : n46472;
  assign n46474 = pi18 ? n19124 : n46473;
  assign n46475 = pi17 ? n46470 : n46474;
  assign n46476 = pi16 ? n40499 : n46475;
  assign n46477 = pi19 ? n31904 : n21611;
  assign n46478 = pi18 ? n20563 : n46477;
  assign n46479 = pi21 ? n316 : n2300;
  assign n46480 = pi20 ? n46479 : n32;
  assign n46481 = pi19 ? n45935 : n46480;
  assign n46482 = pi18 ? n99 : n46481;
  assign n46483 = pi17 ? n46478 : n46482;
  assign n46484 = pi16 ? n39375 : n46483;
  assign n46485 = pi15 ? n46476 : n46484;
  assign n46486 = pi14 ? n46468 : n46485;
  assign n46487 = pi13 ? n46460 : n46486;
  assign n46488 = pi12 ? n46439 : n46487;
  assign n46489 = pi11 ? n46415 : n46488;
  assign n46490 = pi21 ? n31924 : n181;
  assign n46491 = pi20 ? n20563 : n46490;
  assign n46492 = pi19 ? n46491 : n45949;
  assign n46493 = pi18 ? n20563 : n46492;
  assign n46494 = pi19 ? n45952 : n10595;
  assign n46495 = pi18 ? n99 : n46494;
  assign n46496 = pi17 ? n46493 : n46495;
  assign n46497 = pi16 ? n39375 : n46496;
  assign n46498 = pi21 ? n31924 : n99;
  assign n46499 = pi20 ? n20563 : n46498;
  assign n46500 = pi19 ? n46499 : n3050;
  assign n46501 = pi18 ? n20563 : n46500;
  assign n46502 = pi19 ? n27596 : n10595;
  assign n46503 = pi18 ? n44885 : n46502;
  assign n46504 = pi17 ? n46501 : n46503;
  assign n46505 = pi16 ? n39375 : n46504;
  assign n46506 = pi15 ? n46497 : n46505;
  assign n46507 = pi21 ? n204 : n6416;
  assign n46508 = pi20 ? n46507 : n32;
  assign n46509 = pi19 ? n2862 : n46508;
  assign n46510 = pi18 ? n44893 : n46509;
  assign n46511 = pi17 ? n41685 : n46510;
  assign n46512 = pi16 ? n39375 : n46511;
  assign n46513 = pi20 ? n7264 : n32;
  assign n46514 = pi19 ? n2317 : n46513;
  assign n46515 = pi18 ? n18083 : n46514;
  assign n46516 = pi17 ? n41685 : n46515;
  assign n46517 = pi16 ? n40534 : n46516;
  assign n46518 = pi15 ? n46512 : n46517;
  assign n46519 = pi14 ? n46506 : n46518;
  assign n46520 = pi19 ? n2317 : n19330;
  assign n46521 = pi18 ? n8766 : n46520;
  assign n46522 = pi17 ? n45975 : n46521;
  assign n46523 = pi16 ? n38959 : n46522;
  assign n46524 = pi19 ? n31904 : n9814;
  assign n46525 = pi18 ? n20563 : n46524;
  assign n46526 = pi22 ? n204 : n4883;
  assign n46527 = pi21 ? n46526 : n928;
  assign n46528 = pi20 ? n46527 : n32;
  assign n46529 = pi19 ? n36541 : n46528;
  assign n46530 = pi18 ? n139 : n46529;
  assign n46531 = pi17 ? n46525 : n46530;
  assign n46532 = pi16 ? n38959 : n46531;
  assign n46533 = pi15 ? n46523 : n46532;
  assign n46534 = pi21 ? n46526 : n1009;
  assign n46535 = pi20 ? n46534 : n32;
  assign n46536 = pi19 ? n36541 : n46535;
  assign n46537 = pi18 ? n139 : n46536;
  assign n46538 = pi17 ? n46525 : n46537;
  assign n46539 = pi16 ? n38959 : n46538;
  assign n46540 = pi21 ? n25463 : n32;
  assign n46541 = pi20 ? n46540 : n32;
  assign n46542 = pi19 ? n36541 : n46541;
  assign n46543 = pi18 ? n139 : n46542;
  assign n46544 = pi17 ? n45989 : n46543;
  assign n46545 = pi16 ? n38959 : n46544;
  assign n46546 = pi15 ? n46539 : n46545;
  assign n46547 = pi14 ? n46533 : n46546;
  assign n46548 = pi13 ? n46519 : n46547;
  assign n46549 = pi20 ? n3075 : n16047;
  assign n46550 = pi19 ? n31926 : n46549;
  assign n46551 = pi18 ? n20563 : n46550;
  assign n46552 = pi20 ? n33658 : n32;
  assign n46553 = pi19 ? n46004 : n46552;
  assign n46554 = pi18 ? n139 : n46553;
  assign n46555 = pi17 ? n46551 : n46554;
  assign n46556 = pi16 ? n39399 : n46555;
  assign n46557 = pi20 ? n20563 : n3086;
  assign n46558 = pi19 ? n46557 : n9769;
  assign n46559 = pi18 ? n20563 : n46558;
  assign n46560 = pi22 ? n6833 : n2121;
  assign n46561 = pi21 ? n46560 : n32;
  assign n46562 = pi20 ? n46561 : n32;
  assign n46563 = pi19 ? n139 : n46562;
  assign n46564 = pi18 ? n139 : n46563;
  assign n46565 = pi17 ? n46559 : n46564;
  assign n46566 = pi16 ? n39399 : n46565;
  assign n46567 = pi15 ? n46556 : n46566;
  assign n46568 = pi19 ? n46021 : n10298;
  assign n46569 = pi18 ? n10682 : n46568;
  assign n46570 = pi17 ? n45359 : n46569;
  assign n46571 = pi16 ? n39399 : n46570;
  assign n46572 = pi22 ? n233 : n21537;
  assign n46573 = pi21 ? n46572 : n32;
  assign n46574 = pi20 ? n46573 : n32;
  assign n46575 = pi19 ? n233 : n46574;
  assign n46576 = pi18 ? n46026 : n46575;
  assign n46577 = pi17 ? n45359 : n46576;
  assign n46578 = pi16 ? n39399 : n46577;
  assign n46579 = pi15 ? n46571 : n46578;
  assign n46580 = pi14 ? n46567 : n46579;
  assign n46581 = pi21 ? n15698 : n32;
  assign n46582 = pi20 ? n46581 : n32;
  assign n46583 = pi19 ? n46035 : n46582;
  assign n46584 = pi18 ? n46034 : n46583;
  assign n46585 = pi17 ? n41178 : n46584;
  assign n46586 = pi16 ? n38318 : n46585;
  assign n46587 = pi21 ? n20563 : n43580;
  assign n46588 = pi20 ? n46587 : n2973;
  assign n46589 = pi19 ? n46588 : n37;
  assign n46590 = pi18 ? n20563 : n46589;
  assign n46591 = pi22 ? n6365 : n18256;
  assign n46592 = pi21 ? n46591 : n32;
  assign n46593 = pi20 ? n46592 : n32;
  assign n46594 = pi19 ? n233 : n46593;
  assign n46595 = pi18 ? n46046 : n46594;
  assign n46596 = pi17 ? n46590 : n46595;
  assign n46597 = pi16 ? n40552 : n46596;
  assign n46598 = pi15 ? n46586 : n46597;
  assign n46599 = pi22 ? n37804 : n20563;
  assign n46600 = pi21 ? n46599 : n20563;
  assign n46601 = pi20 ? n46600 : n20563;
  assign n46602 = pi19 ? n46601 : n20563;
  assign n46603 = pi18 ? n32 : n46602;
  assign n46604 = pi17 ? n32 : n46603;
  assign n46605 = pi21 ? n38763 : n32;
  assign n46606 = pi20 ? n46605 : n32;
  assign n46607 = pi19 ? n7981 : n46606;
  assign n46608 = pi18 ? n16209 : n46607;
  assign n46609 = pi17 ? n41178 : n46608;
  assign n46610 = pi16 ? n46604 : n46609;
  assign n46611 = pi22 ? n37251 : n30868;
  assign n46612 = pi21 ? n46611 : n30868;
  assign n46613 = pi20 ? n46612 : n30868;
  assign n46614 = pi19 ? n46613 : n42014;
  assign n46615 = pi18 ? n32 : n46614;
  assign n46616 = pi17 ? n32 : n46615;
  assign n46617 = pi19 ? n32703 : n46055;
  assign n46618 = pi18 ? n15161 : n46617;
  assign n46619 = pi17 ? n41178 : n46618;
  assign n46620 = pi16 ? n46616 : n46619;
  assign n46621 = pi15 ? n46610 : n46620;
  assign n46622 = pi14 ? n46598 : n46621;
  assign n46623 = pi13 ? n46580 : n46622;
  assign n46624 = pi12 ? n46548 : n46623;
  assign n46625 = pi18 ? n32 : n33792;
  assign n46626 = pi17 ? n32 : n46625;
  assign n46627 = pi21 ? n37768 : n29133;
  assign n46628 = pi20 ? n46627 : n37;
  assign n46629 = pi19 ? n46628 : n37;
  assign n46630 = pi18 ? n46083 : n46629;
  assign n46631 = pi19 ? n45022 : n4103;
  assign n46632 = pi18 ? n46086 : n46631;
  assign n46633 = pi17 ? n46630 : n46632;
  assign n46634 = pi16 ? n46626 : n46633;
  assign n46635 = pi19 ? n31267 : n335;
  assign n46636 = pi18 ? n20563 : n46635;
  assign n46637 = pi23 ? n19714 : n685;
  assign n46638 = pi22 ? n335 : n46637;
  assign n46639 = pi21 ? n335 : n46638;
  assign n46640 = pi20 ? n335 : n46639;
  assign n46641 = pi19 ? n46640 : n4103;
  assign n46642 = pi18 ? n335 : n46641;
  assign n46643 = pi17 ? n46636 : n46642;
  assign n46644 = pi16 ? n37930 : n46643;
  assign n46645 = pi15 ? n46634 : n46644;
  assign n46646 = pi22 ? n363 : n8311;
  assign n46647 = pi21 ? n37 : n46646;
  assign n46648 = pi20 ? n37 : n46647;
  assign n46649 = pi19 ? n46648 : n2639;
  assign n46650 = pi18 ? n45034 : n46649;
  assign n46651 = pi17 ? n41178 : n46650;
  assign n46652 = pi16 ? n37930 : n46651;
  assign n46653 = pi22 ? n4537 : n2244;
  assign n46654 = pi21 ? n37 : n46653;
  assign n46655 = pi20 ? n37 : n46654;
  assign n46656 = pi19 ? n46655 : n2654;
  assign n46657 = pi18 ? n45034 : n46656;
  assign n46658 = pi17 ? n41178 : n46657;
  assign n46659 = pi16 ? n37930 : n46658;
  assign n46660 = pi15 ? n46652 : n46659;
  assign n46661 = pi14 ? n46645 : n46660;
  assign n46662 = pi20 ? n20563 : n16008;
  assign n46663 = pi19 ? n46662 : n46119;
  assign n46664 = pi18 ? n20563 : n46663;
  assign n46665 = pi17 ? n46664 : n46126;
  assign n46666 = pi16 ? n38331 : n46665;
  assign n46667 = pi20 ? n20563 : n14887;
  assign n46668 = pi19 ? n46667 : n43075;
  assign n46669 = pi18 ? n20563 : n46668;
  assign n46670 = pi20 ? n22881 : n38841;
  assign n46671 = pi19 ? n46670 : n2654;
  assign n46672 = pi18 ? n45065 : n46671;
  assign n46673 = pi17 ? n46669 : n46672;
  assign n46674 = pi16 ? n38331 : n46673;
  assign n46675 = pi15 ? n46666 : n46674;
  assign n46676 = pi20 ? n20563 : n13613;
  assign n46677 = pi19 ? n46676 : n37;
  assign n46678 = pi18 ? n20563 : n46677;
  assign n46679 = pi19 ? n28767 : n2654;
  assign n46680 = pi18 ? n24881 : n46679;
  assign n46681 = pi17 ? n46678 : n46680;
  assign n46682 = pi16 ? n45394 : n46681;
  assign n46683 = pi20 ? n24220 : n45077;
  assign n46684 = pi19 ? n46683 : n35482;
  assign n46685 = pi18 ? n46146 : n46684;
  assign n46686 = pi17 ? n46678 : n46685;
  assign n46687 = pi16 ? n45394 : n46686;
  assign n46688 = pi15 ? n46682 : n46687;
  assign n46689 = pi14 ? n46675 : n46688;
  assign n46690 = pi13 ? n46661 : n46689;
  assign n46691 = pi20 ? n20563 : n3292;
  assign n46692 = pi19 ? n46691 : n45097;
  assign n46693 = pi18 ? n20563 : n46692;
  assign n46694 = pi20 ? n685 : n45077;
  assign n46695 = pi19 ? n46694 : n32;
  assign n46696 = pi18 ? n45100 : n46695;
  assign n46697 = pi17 ? n46693 : n46696;
  assign n46698 = pi16 ? n45394 : n46697;
  assign n46699 = pi21 ? n46166 : n30868;
  assign n46700 = pi20 ? n46699 : n30868;
  assign n46701 = pi19 ? n46700 : n30868;
  assign n46702 = pi18 ? n32 : n46701;
  assign n46703 = pi17 ? n32 : n46702;
  assign n46704 = pi21 ? n45608 : n363;
  assign n46705 = pi20 ? n30868 : n46704;
  assign n46706 = pi19 ? n46705 : n34796;
  assign n46707 = pi18 ? n30868 : n46706;
  assign n46708 = pi20 ? n26891 : n27218;
  assign n46709 = pi19 ? n46708 : n32;
  assign n46710 = pi18 ? n45115 : n46709;
  assign n46711 = pi17 ? n46707 : n46710;
  assign n46712 = pi16 ? n46703 : n46711;
  assign n46713 = pi15 ? n46698 : n46712;
  assign n46714 = pi21 ? n46187 : n30868;
  assign n46715 = pi20 ? n46714 : n30868;
  assign n46716 = pi19 ? n46715 : n30868;
  assign n46717 = pi18 ? n32 : n46716;
  assign n46718 = pi17 ? n32 : n46717;
  assign n46719 = pi20 ? n41565 : n99;
  assign n46720 = pi19 ? n46719 : n99;
  assign n46721 = pi18 ? n30868 : n46720;
  assign n46722 = pi20 ? n99 : n42552;
  assign n46723 = pi19 ? n46722 : n32;
  assign n46724 = pi18 ? n46195 : n46723;
  assign n46725 = pi17 ? n46721 : n46724;
  assign n46726 = pi16 ? n46718 : n46725;
  assign n46727 = pi22 ? n32 : n36798;
  assign n46728 = pi21 ? n46727 : n36798;
  assign n46729 = pi20 ? n46728 : n36798;
  assign n46730 = pi19 ? n46729 : n46204;
  assign n46731 = pi18 ? n32 : n46730;
  assign n46732 = pi17 ? n32 : n46731;
  assign n46733 = pi21 ? n38867 : n139;
  assign n46734 = pi20 ? n33792 : n46733;
  assign n46735 = pi19 ? n46734 : n139;
  assign n46736 = pi18 ? n33792 : n46735;
  assign n46737 = pi20 ? n139 : n46213;
  assign n46738 = pi19 ? n139 : n46737;
  assign n46739 = pi22 ? n316 : n26376;
  assign n46740 = pi21 ? n157 : n46739;
  assign n46741 = pi20 ? n139 : n46740;
  assign n46742 = pi19 ? n46741 : n32;
  assign n46743 = pi18 ? n46738 : n46742;
  assign n46744 = pi17 ? n46736 : n46743;
  assign n46745 = pi16 ? n46732 : n46744;
  assign n46746 = pi15 ? n46726 : n46745;
  assign n46747 = pi14 ? n46713 : n46746;
  assign n46748 = pi19 ? n46729 : n43139;
  assign n46749 = pi18 ? n32 : n46748;
  assign n46750 = pi17 ? n32 : n46749;
  assign n46751 = pi21 ? n38867 : n335;
  assign n46752 = pi20 ? n33792 : n46751;
  assign n46753 = pi19 ? n46752 : n335;
  assign n46754 = pi18 ? n41580 : n46753;
  assign n46755 = pi17 ? n46754 : n46237;
  assign n46756 = pi16 ? n46750 : n46755;
  assign n46757 = pi23 ? n32 : n37273;
  assign n46758 = pi22 ? n32 : n46757;
  assign n46759 = pi21 ? n46758 : n36781;
  assign n46760 = pi20 ? n46759 : n36781;
  assign n46761 = pi19 ? n46760 : n45180;
  assign n46762 = pi18 ? n32 : n46761;
  assign n46763 = pi17 ? n32 : n46762;
  assign n46764 = pi22 ? n36659 : n335;
  assign n46765 = pi21 ? n46764 : n335;
  assign n46766 = pi20 ? n46242 : n46765;
  assign n46767 = pi19 ? n46766 : n335;
  assign n46768 = pi18 ? n41103 : n46767;
  assign n46769 = pi17 ? n46768 : n46254;
  assign n46770 = pi16 ? n46763 : n46769;
  assign n46771 = pi15 ? n46756 : n46770;
  assign n46772 = pi22 ? n32 : n45160;
  assign n46773 = pi21 ? n46772 : n36798;
  assign n46774 = pi20 ? n46773 : n36798;
  assign n46775 = pi19 ? n46774 : n41135;
  assign n46776 = pi18 ? n32 : n46775;
  assign n46777 = pi17 ? n32 : n46776;
  assign n46778 = pi22 ? n36798 : n37276;
  assign n46779 = pi21 ? n46778 : n34833;
  assign n46780 = pi20 ? n46261 : n46779;
  assign n46781 = pi19 ? n46780 : n157;
  assign n46782 = pi18 ? n45198 : n46781;
  assign n46783 = pi21 ? n46267 : n2320;
  assign n46784 = pi20 ? n157 : n46783;
  assign n46785 = pi19 ? n46784 : n32;
  assign n46786 = pi18 ? n157 : n46785;
  assign n46787 = pi17 ? n46782 : n46786;
  assign n46788 = pi16 ? n46777 : n46787;
  assign n46789 = pi23 ? n32 : n43198;
  assign n46790 = pi22 ? n32 : n46789;
  assign n46791 = pi21 ? n46790 : n43198;
  assign n46792 = pi20 ? n46791 : n46281;
  assign n46793 = pi19 ? n46792 : n46285;
  assign n46794 = pi18 ? n32 : n46793;
  assign n46795 = pi17 ? n32 : n46794;
  assign n46796 = pi23 ? n363 : n36798;
  assign n46797 = pi22 ? n36798 : n46796;
  assign n46798 = pi21 ? n46797 : n157;
  assign n46799 = pi20 ? n46289 : n46798;
  assign n46800 = pi19 ? n46799 : n157;
  assign n46801 = pi18 ? n45198 : n46800;
  assign n46802 = pi17 ? n46801 : n45696;
  assign n46803 = pi16 ? n46795 : n46802;
  assign n46804 = pi15 ? n46788 : n46803;
  assign n46805 = pi14 ? n46771 : n46804;
  assign n46806 = pi13 ? n46747 : n46805;
  assign n46807 = pi12 ? n46690 : n46806;
  assign n46808 = pi11 ? n46624 : n46807;
  assign n46809 = pi10 ? n46489 : n46808;
  assign n46810 = pi09 ? n46321 : n46809;
  assign n46811 = pi08 ? n46301 : n46810;
  assign n46812 = pi07 ? n45706 : n46811;
  assign n46813 = pi06 ? n44633 : n46812;
  assign n46814 = pi05 ? n42643 : n46813;
  assign n46815 = pi21 ? n29133 : n36249;
  assign n46816 = pi20 ? n46815 : n20563;
  assign n46817 = pi19 ? n34920 : n46816;
  assign n46818 = pi18 ? n46446 : n46817;
  assign n46819 = pi21 ? n31200 : n31924;
  assign n46820 = pi20 ? n46819 : n33964;
  assign n46821 = pi19 ? n46820 : n37;
  assign n46822 = pi20 ? n37 : n38969;
  assign n46823 = pi23 ? n3491 : n32;
  assign n46824 = pi22 ? n46823 : n32;
  assign n46825 = pi21 ? n46824 : n32;
  assign n46826 = pi20 ? n14844 : n46825;
  assign n46827 = pi19 ? n46822 : n46826;
  assign n46828 = pi18 ? n46821 : n46827;
  assign n46829 = pi17 ? n46818 : n46828;
  assign n46830 = pi16 ? n32 : n46829;
  assign n46831 = pi15 ? n32 : n46830;
  assign n46832 = pi18 ? n41708 : n20563;
  assign n46833 = pi21 ? n23269 : n32;
  assign n46834 = pi20 ? n3086 : n46833;
  assign n46835 = pi19 ? n37 : n46834;
  assign n46836 = pi18 ? n32295 : n46835;
  assign n46837 = pi17 ? n46832 : n46836;
  assign n46838 = pi16 ? n32 : n46837;
  assign n46839 = pi18 ? n38957 : n20563;
  assign n46840 = pi20 ? n8742 : n46833;
  assign n46841 = pi19 ? n37 : n46840;
  assign n46842 = pi18 ? n33299 : n46841;
  assign n46843 = pi17 ? n46839 : n46842;
  assign n46844 = pi16 ? n32 : n46843;
  assign n46845 = pi15 ? n46838 : n46844;
  assign n46846 = pi14 ? n46831 : n46845;
  assign n46847 = pi13 ? n32 : n46846;
  assign n46848 = pi12 ? n32 : n46847;
  assign n46849 = pi11 ? n32 : n46848;
  assign n46850 = pi10 ? n32 : n46849;
  assign n46851 = pi23 ? n19714 : n32;
  assign n46852 = pi22 ? n46851 : n32;
  assign n46853 = pi21 ? n46852 : n32;
  assign n46854 = pi20 ? n3086 : n46853;
  assign n46855 = pi19 ? n37 : n46854;
  assign n46856 = pi18 ? n33285 : n46855;
  assign n46857 = pi17 ? n45707 : n46856;
  assign n46858 = pi16 ? n32 : n46857;
  assign n46859 = pi18 ? n39397 : n20563;
  assign n46860 = pi20 ? n942 : n17032;
  assign n46861 = pi19 ? n12370 : n46860;
  assign n46862 = pi18 ? n32872 : n46861;
  assign n46863 = pi17 ? n46859 : n46862;
  assign n46864 = pi16 ? n32 : n46863;
  assign n46865 = pi15 ? n46858 : n46864;
  assign n46866 = pi18 ? n45392 : n20563;
  assign n46867 = pi20 ? n139 : n2470;
  assign n46868 = pi19 ? n37 : n46867;
  assign n46869 = pi18 ? n33299 : n46868;
  assign n46870 = pi17 ? n46866 : n46869;
  assign n46871 = pi16 ? n32 : n46870;
  assign n46872 = pi20 ? n3090 : n2470;
  assign n46873 = pi19 ? n37 : n46872;
  assign n46874 = pi18 ? n33869 : n46873;
  assign n46875 = pi17 ? n20563 : n46874;
  assign n46876 = pi16 ? n44635 : n46875;
  assign n46877 = pi15 ? n46871 : n46876;
  assign n46878 = pi14 ? n46865 : n46877;
  assign n46879 = pi20 ? n942 : n2554;
  assign n46880 = pi19 ? n9824 : n46879;
  assign n46881 = pi18 ? n34358 : n46880;
  assign n46882 = pi17 ? n20563 : n46881;
  assign n46883 = pi16 ? n45740 : n46882;
  assign n46884 = pi18 ? n32 : n36869;
  assign n46885 = pi17 ? n32 : n46884;
  assign n46886 = pi20 ? n577 : n2554;
  assign n46887 = pi19 ? n37 : n46886;
  assign n46888 = pi18 ? n42358 : n46887;
  assign n46889 = pi17 ? n20563 : n46888;
  assign n46890 = pi16 ? n46885 : n46889;
  assign n46891 = pi15 ? n46883 : n46890;
  assign n46892 = pi20 ? n577 : n2679;
  assign n46893 = pi19 ? n37 : n46892;
  assign n46894 = pi18 ? n34358 : n46893;
  assign n46895 = pi17 ? n20563 : n46894;
  assign n46896 = pi16 ? n44653 : n46895;
  assign n46897 = pi20 ? n649 : n2701;
  assign n46898 = pi19 ? n37 : n46897;
  assign n46899 = pi18 ? n33916 : n46898;
  assign n46900 = pi17 ? n20563 : n46899;
  assign n46901 = pi16 ? n44223 : n46900;
  assign n46902 = pi15 ? n46896 : n46901;
  assign n46903 = pi14 ? n46891 : n46902;
  assign n46904 = pi13 ? n46878 : n46903;
  assign n46905 = pi18 ? n32349 : n46898;
  assign n46906 = pi17 ? n20563 : n46905;
  assign n46907 = pi16 ? n44671 : n46906;
  assign n46908 = pi21 ? n37 : n10684;
  assign n46909 = pi20 ? n46908 : n1822;
  assign n46910 = pi19 ? n37 : n46909;
  assign n46911 = pi18 ? n37029 : n46910;
  assign n46912 = pi17 ? n20563 : n46911;
  assign n46913 = pi16 ? n43675 : n46912;
  assign n46914 = pi15 ? n46907 : n46913;
  assign n46915 = pi21 ? n569 : n10684;
  assign n46916 = pi20 ? n46915 : n1822;
  assign n46917 = pi19 ? n8802 : n46916;
  assign n46918 = pi18 ? n37 : n46917;
  assign n46919 = pi17 ? n20563 : n46918;
  assign n46920 = pi16 ? n43685 : n46919;
  assign n46921 = pi19 ? n8802 : n45824;
  assign n46922 = pi18 ? n37 : n46921;
  assign n46923 = pi17 ? n42647 : n46922;
  assign n46924 = pi16 ? n44688 : n46923;
  assign n46925 = pi15 ? n46920 : n46924;
  assign n46926 = pi14 ? n46914 : n46925;
  assign n46927 = pi20 ? n2094 : n32;
  assign n46928 = pi19 ? n37 : n46927;
  assign n46929 = pi18 ? n37 : n46928;
  assign n46930 = pi17 ? n42647 : n46929;
  assign n46931 = pi16 ? n44688 : n46930;
  assign n46932 = pi20 ? n2085 : n2679;
  assign n46933 = pi19 ? n37 : n46932;
  assign n46934 = pi18 ? n37 : n46933;
  assign n46935 = pi17 ? n20563 : n46934;
  assign n46936 = pi16 ? n42682 : n46935;
  assign n46937 = pi15 ? n46931 : n46936;
  assign n46938 = pi17 ? n20563 : n46409;
  assign n46939 = pi16 ? n42682 : n46938;
  assign n46940 = pi19 ? n37 : n18629;
  assign n46941 = pi18 ? n37 : n46940;
  assign n46942 = pi17 ? n42657 : n46941;
  assign n46943 = pi16 ? n42682 : n46942;
  assign n46944 = pi15 ? n46939 : n46943;
  assign n46945 = pi14 ? n46937 : n46944;
  assign n46946 = pi13 ? n46926 : n46945;
  assign n46947 = pi12 ? n46904 : n46946;
  assign n46948 = pi17 ? n42657 : n46409;
  assign n46949 = pi16 ? n42195 : n46948;
  assign n46950 = pi18 ? n20563 : n40314;
  assign n46951 = pi21 ? n6401 : n14255;
  assign n46952 = pi20 ? n46951 : n32;
  assign n46953 = pi19 ? n5029 : n46952;
  assign n46954 = pi18 ? n37 : n46953;
  assign n46955 = pi17 ? n46950 : n46954;
  assign n46956 = pi16 ? n43256 : n46955;
  assign n46957 = pi15 ? n46949 : n46956;
  assign n46958 = pi18 ? n20563 : n39447;
  assign n46959 = pi22 ? n37 : n705;
  assign n46960 = pi21 ? n37 : n46959;
  assign n46961 = pi20 ? n46960 : n32;
  assign n46962 = pi19 ? n37 : n46961;
  assign n46963 = pi18 ? n37 : n46962;
  assign n46964 = pi17 ? n46958 : n46963;
  assign n46965 = pi16 ? n42202 : n46964;
  assign n46966 = pi21 ? n37 : n2759;
  assign n46967 = pi20 ? n46966 : n32;
  assign n46968 = pi19 ? n37 : n46967;
  assign n46969 = pi18 ? n37 : n46968;
  assign n46970 = pi17 ? n43676 : n46969;
  assign n46971 = pi16 ? n42208 : n46970;
  assign n46972 = pi15 ? n46965 : n46971;
  assign n46973 = pi14 ? n46957 : n46972;
  assign n46974 = pi17 ? n20563 : n44771;
  assign n46975 = pi16 ? n41632 : n46974;
  assign n46976 = pi17 ? n43665 : n44771;
  assign n46977 = pi16 ? n41632 : n46976;
  assign n46978 = pi15 ? n46975 : n46977;
  assign n46979 = pi21 ? n37 : n10318;
  assign n46980 = pi20 ? n46979 : n32;
  assign n46981 = pi19 ? n37 : n46980;
  assign n46982 = pi18 ? n37 : n46981;
  assign n46983 = pi17 ? n44732 : n46982;
  assign n46984 = pi16 ? n42689 : n46983;
  assign n46985 = pi18 ? n20563 : n33847;
  assign n46986 = pi21 ? n24501 : n272;
  assign n46987 = pi20 ? n37 : n46986;
  assign n46988 = pi21 ? n272 : n6535;
  assign n46989 = pi20 ? n46988 : n32;
  assign n46990 = pi19 ? n46987 : n46989;
  assign n46991 = pi18 ? n37 : n46990;
  assign n46992 = pi17 ? n46985 : n46991;
  assign n46993 = pi16 ? n42689 : n46992;
  assign n46994 = pi15 ? n46984 : n46993;
  assign n46995 = pi14 ? n46978 : n46994;
  assign n46996 = pi13 ? n46973 : n46995;
  assign n46997 = pi19 ? n37321 : n20563;
  assign n46998 = pi18 ? n32 : n46997;
  assign n46999 = pi17 ? n32 : n46998;
  assign n47000 = pi21 ? n37 : n6535;
  assign n47001 = pi20 ? n47000 : n32;
  assign n47002 = pi19 ? n37 : n47001;
  assign n47003 = pi18 ? n37 : n47002;
  assign n47004 = pi17 ? n42657 : n47003;
  assign n47005 = pi16 ? n46999 : n47004;
  assign n47006 = pi19 ? n37 : n13111;
  assign n47007 = pi18 ? n37 : n47006;
  assign n47008 = pi17 ? n42657 : n47007;
  assign n47009 = pi16 ? n46999 : n47008;
  assign n47010 = pi15 ? n47005 : n47009;
  assign n47011 = pi20 ? n22644 : n99;
  assign n47012 = pi19 ? n47011 : n99;
  assign n47013 = pi18 ? n47012 : n46450;
  assign n47014 = pi17 ? n44732 : n47013;
  assign n47015 = pi16 ? n46999 : n47014;
  assign n47016 = pi20 ? n31220 : n21635;
  assign n47017 = pi19 ? n20563 : n47016;
  assign n47018 = pi18 ? n20563 : n47017;
  assign n47019 = pi20 ? n3869 : n99;
  assign n47020 = pi19 ? n47019 : n99;
  assign n47021 = pi18 ? n47020 : n46450;
  assign n47022 = pi17 ? n47018 : n47021;
  assign n47023 = pi16 ? n40487 : n47022;
  assign n47024 = pi15 ? n47015 : n47023;
  assign n47025 = pi14 ? n47010 : n47024;
  assign n47026 = pi20 ? n38966 : n37;
  assign n47027 = pi19 ? n20563 : n47026;
  assign n47028 = pi18 ? n20563 : n47027;
  assign n47029 = pi20 ? n99 : n9687;
  assign n47030 = pi19 ? n47029 : n16340;
  assign n47031 = pi18 ? n99 : n47030;
  assign n47032 = pi17 ? n47028 : n47031;
  assign n47033 = pi16 ? n40487 : n47032;
  assign n47034 = pi20 ? n40919 : n14844;
  assign n47035 = pi19 ? n20563 : n47034;
  assign n47036 = pi18 ? n20563 : n47035;
  assign n47037 = pi19 ? n11445 : n16325;
  assign n47038 = pi18 ? n38578 : n47037;
  assign n47039 = pi17 ? n47036 : n47038;
  assign n47040 = pi16 ? n40487 : n47039;
  assign n47041 = pi15 ? n47033 : n47040;
  assign n47042 = pi20 ? n40755 : n15964;
  assign n47043 = pi19 ? n20563 : n47042;
  assign n47044 = pi18 ? n20563 : n47043;
  assign n47045 = pi20 ? n18499 : n99;
  assign n47046 = pi20 ? n6477 : n99;
  assign n47047 = pi19 ? n47045 : n47046;
  assign n47048 = pi21 ? n775 : n5176;
  assign n47049 = pi20 ? n2238 : n47048;
  assign n47050 = pi21 ? n5176 : n2320;
  assign n47051 = pi20 ? n47050 : n32;
  assign n47052 = pi19 ? n47049 : n47051;
  assign n47053 = pi18 ? n47047 : n47052;
  assign n47054 = pi17 ? n47044 : n47053;
  assign n47055 = pi16 ? n42241 : n47054;
  assign n47056 = pi19 ? n31314 : n20563;
  assign n47057 = pi18 ? n32 : n47056;
  assign n47058 = pi17 ? n32 : n47057;
  assign n47059 = pi20 ? n30096 : n2970;
  assign n47060 = pi19 ? n20563 : n47059;
  assign n47061 = pi18 ? n20563 : n47060;
  assign n47062 = pi20 ? n30108 : n3824;
  assign n47063 = pi19 ? n47062 : n23318;
  assign n47064 = pi20 ? n99 : n19201;
  assign n47065 = pi21 ? n204 : n2320;
  assign n47066 = pi20 ? n47065 : n32;
  assign n47067 = pi19 ? n47064 : n47066;
  assign n47068 = pi18 ? n47063 : n47067;
  assign n47069 = pi17 ? n47061 : n47068;
  assign n47070 = pi16 ? n47058 : n47069;
  assign n47071 = pi15 ? n47055 : n47070;
  assign n47072 = pi14 ? n47041 : n47071;
  assign n47073 = pi13 ? n47025 : n47072;
  assign n47074 = pi12 ? n46996 : n47073;
  assign n47075 = pi11 ? n46947 : n47074;
  assign n47076 = pi19 ? n42915 : n30109;
  assign n47077 = pi18 ? n20563 : n47076;
  assign n47078 = pi21 ? n16438 : n2320;
  assign n47079 = pi20 ? n47078 : n32;
  assign n47080 = pi19 ? n99 : n47079;
  assign n47081 = pi18 ? n34285 : n47080;
  assign n47082 = pi17 ? n47077 : n47081;
  assign n47083 = pi16 ? n47058 : n47082;
  assign n47084 = pi20 ? n40755 : n38969;
  assign n47085 = pi19 ? n32876 : n47084;
  assign n47086 = pi18 ? n20563 : n47085;
  assign n47087 = pi20 ? n3884 : n2959;
  assign n47088 = pi19 ? n99 : n47087;
  assign n47089 = pi22 ? n112 : n745;
  assign n47090 = pi21 ? n47089 : n204;
  assign n47091 = pi20 ? n3042 : n47090;
  assign n47092 = pi21 ? n204 : n4101;
  assign n47093 = pi20 ? n47092 : n32;
  assign n47094 = pi19 ? n47091 : n47093;
  assign n47095 = pi18 ? n47088 : n47094;
  assign n47096 = pi17 ? n47086 : n47095;
  assign n47097 = pi16 ? n47058 : n47096;
  assign n47098 = pi15 ? n47083 : n47097;
  assign n47099 = pi21 ? n39175 : n37;
  assign n47100 = pi20 ? n47099 : n8742;
  assign n47101 = pi19 ? n32876 : n47100;
  assign n47102 = pi18 ? n20563 : n47101;
  assign n47103 = pi19 ? n28290 : n28582;
  assign n47104 = pi19 ? n1017 : n19321;
  assign n47105 = pi18 ? n47103 : n47104;
  assign n47106 = pi17 ? n47102 : n47105;
  assign n47107 = pi16 ? n47058 : n47106;
  assign n47108 = pi19 ? n32663 : n19691;
  assign n47109 = pi18 ? n37 : n47108;
  assign n47110 = pi17 ? n42196 : n47109;
  assign n47111 = pi16 ? n41684 : n47110;
  assign n47112 = pi15 ? n47107 : n47111;
  assign n47113 = pi14 ? n47098 : n47112;
  assign n47114 = pi19 ? n32294 : n20759;
  assign n47115 = pi18 ? n20563 : n47114;
  assign n47116 = pi21 ? n204 : n882;
  assign n47117 = pi20 ? n47116 : n32;
  assign n47118 = pi19 ? n12589 : n47117;
  assign n47119 = pi18 ? n17061 : n47118;
  assign n47120 = pi17 ? n47115 : n47119;
  assign n47121 = pi16 ? n41684 : n47120;
  assign n47122 = pi21 ? n1696 : n1043;
  assign n47123 = pi20 ? n37 : n47122;
  assign n47124 = pi19 ? n20563 : n47123;
  assign n47125 = pi18 ? n20563 : n47124;
  assign n47126 = pi21 ? n1721 : n297;
  assign n47127 = pi20 ? n47126 : n139;
  assign n47128 = pi19 ? n47127 : n139;
  assign n47129 = pi19 ? n12589 : n18370;
  assign n47130 = pi18 ? n47128 : n47129;
  assign n47131 = pi17 ? n47125 : n47130;
  assign n47132 = pi16 ? n41684 : n47131;
  assign n47133 = pi15 ? n47121 : n47132;
  assign n47134 = pi19 ? n19816 : n9769;
  assign n47135 = pi19 ? n12589 : n18387;
  assign n47136 = pi18 ? n47134 : n47135;
  assign n47137 = pi17 ? n42690 : n47136;
  assign n47138 = pi16 ? n41684 : n47137;
  assign n47139 = pi19 ? n16023 : n139;
  assign n47140 = pi20 ? n139 : n37159;
  assign n47141 = pi20 ? n22805 : n32;
  assign n47142 = pi19 ? n47140 : n47141;
  assign n47143 = pi18 ? n47139 : n47142;
  assign n47144 = pi17 ? n41633 : n47143;
  assign n47145 = pi16 ? n41684 : n47144;
  assign n47146 = pi15 ? n47138 : n47145;
  assign n47147 = pi14 ? n47133 : n47146;
  assign n47148 = pi13 ? n47113 : n47147;
  assign n47149 = pi20 ? n37 : n3087;
  assign n47150 = pi19 ? n32294 : n47149;
  assign n47151 = pi18 ? n20563 : n47150;
  assign n47152 = pi21 ? n335 : n139;
  assign n47153 = pi20 ? n139 : n47152;
  assign n47154 = pi19 ? n47153 : n18413;
  assign n47155 = pi18 ? n139 : n47154;
  assign n47156 = pi17 ? n47151 : n47155;
  assign n47157 = pi16 ? n41710 : n47156;
  assign n47158 = pi21 ? n20563 : n45016;
  assign n47159 = pi20 ? n20563 : n47158;
  assign n47160 = pi19 ? n47159 : n37;
  assign n47161 = pi18 ? n20563 : n47160;
  assign n47162 = pi21 ? n4973 : n2007;
  assign n47163 = pi21 ? n566 : n570;
  assign n47164 = pi20 ? n47162 : n47163;
  assign n47165 = pi19 ? n47164 : n2004;
  assign n47166 = pi20 ? n647 : n6377;
  assign n47167 = pi19 ? n47166 : n18413;
  assign n47168 = pi18 ? n47165 : n47167;
  assign n47169 = pi17 ? n47161 : n47168;
  assign n47170 = pi16 ? n41710 : n47169;
  assign n47171 = pi15 ? n47157 : n47170;
  assign n47172 = pi18 ? n20563 : n33869;
  assign n47173 = pi20 ? n3292 : n604;
  assign n47174 = pi19 ? n37 : n47173;
  assign n47175 = pi20 ? n638 : n42991;
  assign n47176 = pi19 ? n47175 : n19440;
  assign n47177 = pi18 ? n47174 : n47176;
  assign n47178 = pi17 ? n47172 : n47177;
  assign n47179 = pi16 ? n41710 : n47178;
  assign n47180 = pi20 ? n30606 : n32;
  assign n47181 = pi19 ? n13337 : n47180;
  assign n47182 = pi18 ? n6374 : n47181;
  assign n47183 = pi17 ? n41633 : n47182;
  assign n47184 = pi16 ? n41710 : n47183;
  assign n47185 = pi15 ? n47179 : n47184;
  assign n47186 = pi14 ? n47171 : n47185;
  assign n47187 = pi20 ? n30006 : n32;
  assign n47188 = pi19 ? n19358 : n47187;
  assign n47189 = pi18 ? n45798 : n47188;
  assign n47190 = pi17 ? n41644 : n47189;
  assign n47191 = pi16 ? n38950 : n47190;
  assign n47192 = pi21 ? n32 : n30868;
  assign n47193 = pi20 ? n47192 : n30868;
  assign n47194 = pi19 ? n47193 : n30868;
  assign n47195 = pi18 ? n32 : n47194;
  assign n47196 = pi17 ? n32 : n47195;
  assign n47197 = pi22 ? n43579 : n37;
  assign n47198 = pi21 ? n30868 : n47197;
  assign n47199 = pi20 ? n30868 : n47198;
  assign n47200 = pi19 ? n47199 : n37;
  assign n47201 = pi18 ? n30868 : n47200;
  assign n47202 = pi20 ? n649 : n21148;
  assign n47203 = pi19 ? n37 : n47202;
  assign n47204 = pi19 ? n5024 : n47187;
  assign n47205 = pi18 ? n47203 : n47204;
  assign n47206 = pi17 ? n47201 : n47205;
  assign n47207 = pi16 ? n47196 : n47206;
  assign n47208 = pi15 ? n47191 : n47207;
  assign n47209 = pi21 ? n32 : n39191;
  assign n47210 = pi20 ? n47209 : n38754;
  assign n47211 = pi20 ? n30868 : n40915;
  assign n47212 = pi19 ? n47210 : n47211;
  assign n47213 = pi18 ? n32 : n47212;
  assign n47214 = pi17 ? n32 : n47213;
  assign n47215 = pi19 ? n46033 : n5760;
  assign n47216 = pi18 ? n37 : n47215;
  assign n47217 = pi17 ? n41644 : n47216;
  assign n47218 = pi16 ? n47214 : n47217;
  assign n47219 = pi21 ? n32 : n42110;
  assign n47220 = pi22 ? n30868 : n33792;
  assign n47221 = pi21 ? n30868 : n47220;
  assign n47222 = pi20 ? n47219 : n47221;
  assign n47223 = pi21 ? n30868 : n40957;
  assign n47224 = pi20 ? n33792 : n47223;
  assign n47225 = pi19 ? n47222 : n47224;
  assign n47226 = pi18 ? n32 : n47225;
  assign n47227 = pi17 ? n32 : n47226;
  assign n47228 = pi20 ? n37 : n25947;
  assign n47229 = pi19 ? n47228 : n5760;
  assign n47230 = pi18 ? n17225 : n47229;
  assign n47231 = pi17 ? n41644 : n47230;
  assign n47232 = pi16 ? n47227 : n47231;
  assign n47233 = pi15 ? n47218 : n47232;
  assign n47234 = pi14 ? n47208 : n47233;
  assign n47235 = pi13 ? n47186 : n47234;
  assign n47236 = pi12 ? n47148 : n47235;
  assign n47237 = pi21 ? n569 : n685;
  assign n47238 = pi20 ? n37 : n47237;
  assign n47239 = pi19 ? n47238 : n7725;
  assign n47240 = pi18 ? n7677 : n47239;
  assign n47241 = pi17 ? n41644 : n47240;
  assign n47242 = pi16 ? n40552 : n47241;
  assign n47243 = pi19 ? n2730 : n3211;
  assign n47244 = pi18 ? n37 : n47243;
  assign n47245 = pi17 ? n41644 : n47244;
  assign n47246 = pi16 ? n40552 : n47245;
  assign n47247 = pi15 ? n47242 : n47246;
  assign n47248 = pi19 ? n37 : n7730;
  assign n47249 = pi22 ? n363 : n18448;
  assign n47250 = pi21 ? n37 : n47249;
  assign n47251 = pi20 ? n37 : n47250;
  assign n47252 = pi19 ? n47251 : n4117;
  assign n47253 = pi18 ? n47248 : n47252;
  assign n47254 = pi17 ? n41633 : n47253;
  assign n47255 = pi16 ? n40552 : n47254;
  assign n47256 = pi20 ? n7730 : n19091;
  assign n47257 = pi19 ? n37 : n47256;
  assign n47258 = pi21 ? n37 : n43595;
  assign n47259 = pi20 ? n9660 : n47258;
  assign n47260 = pi19 ? n47259 : n5831;
  assign n47261 = pi18 ? n47257 : n47260;
  assign n47262 = pi17 ? n41633 : n47261;
  assign n47263 = pi16 ? n40552 : n47262;
  assign n47264 = pi15 ? n47255 : n47263;
  assign n47265 = pi14 ? n47247 : n47264;
  assign n47266 = pi21 ? n46116 : n29133;
  assign n47267 = pi20 ? n20563 : n47266;
  assign n47268 = pi19 ? n47267 : n37;
  assign n47269 = pi18 ? n20563 : n47268;
  assign n47270 = pi19 ? n44060 : n5831;
  assign n47271 = pi18 ? n27500 : n47270;
  assign n47272 = pi17 ? n47269 : n47271;
  assign n47273 = pi16 ? n38959 : n47272;
  assign n47274 = pi20 ? n7730 : n25199;
  assign n47275 = pi19 ? n47274 : n2654;
  assign n47276 = pi18 ? n37 : n47275;
  assign n47277 = pi17 ? n47269 : n47276;
  assign n47278 = pi16 ? n38959 : n47277;
  assign n47279 = pi15 ? n47273 : n47278;
  assign n47280 = pi21 ? n37768 : n20563;
  assign n47281 = pi20 ? n20563 : n47280;
  assign n47282 = pi19 ? n47281 : n37;
  assign n47283 = pi18 ? n20563 : n47282;
  assign n47284 = pi19 ? n37 : n23917;
  assign n47285 = pi18 ? n47284 : n46679;
  assign n47286 = pi17 ? n47283 : n47285;
  assign n47287 = pi16 ? n38950 : n47286;
  assign n47288 = pi20 ? n363 : n18233;
  assign n47289 = pi19 ? n47288 : n32;
  assign n47290 = pi18 ? n47284 : n47289;
  assign n47291 = pi17 ? n47283 : n47290;
  assign n47292 = pi16 ? n38950 : n47291;
  assign n47293 = pi15 ? n47287 : n47292;
  assign n47294 = pi14 ? n47279 : n47293;
  assign n47295 = pi13 ? n47265 : n47294;
  assign n47296 = pi19 ? n38947 : n30868;
  assign n47297 = pi18 ? n32 : n47296;
  assign n47298 = pi17 ? n32 : n47297;
  assign n47299 = pi21 ? n37784 : n30868;
  assign n47300 = pi20 ? n30868 : n47299;
  assign n47301 = pi19 ? n47300 : n5029;
  assign n47302 = pi18 ? n30868 : n47301;
  assign n47303 = pi21 ? n19958 : n685;
  assign n47304 = pi20 ? n363 : n47303;
  assign n47305 = pi19 ? n39861 : n47304;
  assign n47306 = pi20 ? n685 : n18233;
  assign n47307 = pi19 ? n47306 : n32;
  assign n47308 = pi18 ? n47305 : n47307;
  assign n47309 = pi17 ? n47302 : n47308;
  assign n47310 = pi16 ? n47298 : n47309;
  assign n47311 = pi21 ? n46173 : n30868;
  assign n47312 = pi20 ? n30868 : n47311;
  assign n47313 = pi19 ? n47312 : n2242;
  assign n47314 = pi18 ? n30868 : n47313;
  assign n47315 = pi20 ? n9021 : n685;
  assign n47316 = pi19 ? n6524 : n47315;
  assign n47317 = pi18 ? n47316 : n46161;
  assign n47318 = pi17 ? n47314 : n47317;
  assign n47319 = pi16 ? n47196 : n47318;
  assign n47320 = pi15 ? n47310 : n47319;
  assign n47321 = pi22 ? n32 : n46165;
  assign n47322 = pi21 ? n47321 : n30868;
  assign n47323 = pi20 ? n47322 : n30868;
  assign n47324 = pi19 ? n47323 : n30868;
  assign n47325 = pi18 ? n32 : n47324;
  assign n47326 = pi17 ? n32 : n47325;
  assign n47327 = pi21 ? n39926 : n99;
  assign n47328 = pi20 ? n47327 : n99;
  assign n47329 = pi19 ? n43603 : n47328;
  assign n47330 = pi18 ? n30868 : n47329;
  assign n47331 = pi20 ? n7754 : n5085;
  assign n47332 = pi19 ? n99 : n47331;
  assign n47333 = pi21 ? n767 : n99;
  assign n47334 = pi22 ? n316 : n2192;
  assign n47335 = pi21 ? n3445 : n47334;
  assign n47336 = pi20 ? n47333 : n47335;
  assign n47337 = pi19 ? n47336 : n32;
  assign n47338 = pi18 ? n47332 : n47337;
  assign n47339 = pi17 ? n47330 : n47338;
  assign n47340 = pi16 ? n47326 : n47339;
  assign n47341 = pi22 ? n45652 : n36798;
  assign n47342 = pi21 ? n32 : n47341;
  assign n47343 = pi20 ? n47342 : n36798;
  assign n47344 = pi19 ? n47343 : n36798;
  assign n47345 = pi18 ? n32 : n47344;
  assign n47346 = pi17 ? n32 : n47345;
  assign n47347 = pi20 ? n46733 : n139;
  assign n47348 = pi19 ? n33792 : n47347;
  assign n47349 = pi18 ? n33792 : n47348;
  assign n47350 = pi20 ? n347 : n7850;
  assign n47351 = pi19 ? n139 : n47350;
  assign n47352 = pi21 ? n7429 : n5178;
  assign n47353 = pi20 ? n249 : n47352;
  assign n47354 = pi19 ? n47353 : n32;
  assign n47355 = pi18 ? n47351 : n47354;
  assign n47356 = pi17 ? n47349 : n47355;
  assign n47357 = pi16 ? n47346 : n47356;
  assign n47358 = pi15 ? n47340 : n47357;
  assign n47359 = pi14 ? n47320 : n47358;
  assign n47360 = pi22 ? n33792 : n36659;
  assign n47361 = pi21 ? n47360 : n36659;
  assign n47362 = pi20 ? n47361 : n36659;
  assign n47363 = pi19 ? n47362 : n36659;
  assign n47364 = pi22 ? n36659 : n139;
  assign n47365 = pi21 ? n47364 : n139;
  assign n47366 = pi21 ? n139 : n9143;
  assign n47367 = pi20 ? n47365 : n47366;
  assign n47368 = pi19 ? n36659 : n47367;
  assign n47369 = pi18 ? n47363 : n47368;
  assign n47370 = pi21 ? n335 : n316;
  assign n47371 = pi21 ? n248 : n316;
  assign n47372 = pi20 ? n47370 : n47371;
  assign n47373 = pi19 ? n335 : n47372;
  assign n47374 = pi21 ? n8624 : n157;
  assign n47375 = pi20 ? n47374 : n5179;
  assign n47376 = pi19 ? n47375 : n32;
  assign n47377 = pi18 ? n47373 : n47376;
  assign n47378 = pi17 ? n47369 : n47377;
  assign n47379 = pi16 ? n47346 : n47378;
  assign n47380 = pi23 ? n36798 : n36659;
  assign n47381 = pi22 ? n32 : n47380;
  assign n47382 = pi21 ? n32 : n47381;
  assign n47383 = pi20 ? n47382 : n36659;
  assign n47384 = pi19 ? n47383 : n36659;
  assign n47385 = pi18 ? n32 : n47384;
  assign n47386 = pi17 ? n32 : n47385;
  assign n47387 = pi20 ? n46765 : n335;
  assign n47388 = pi19 ? n36659 : n47387;
  assign n47389 = pi18 ? n36659 : n47388;
  assign n47390 = pi20 ? n47370 : n34537;
  assign n47391 = pi19 ? n335 : n47390;
  assign n47392 = pi18 ? n47391 : n31041;
  assign n47393 = pi17 ? n47389 : n47392;
  assign n47394 = pi16 ? n47386 : n47393;
  assign n47395 = pi15 ? n47379 : n47394;
  assign n47396 = pi22 ? n43198 : n36798;
  assign n47397 = pi22 ? n36798 : n43198;
  assign n47398 = pi21 ? n47396 : n47397;
  assign n47399 = pi20 ? n47342 : n47398;
  assign n47400 = pi19 ? n47399 : n43198;
  assign n47401 = pi18 ? n32 : n47400;
  assign n47402 = pi17 ? n32 : n47401;
  assign n47403 = pi21 ? n36798 : n363;
  assign n47404 = pi21 ? n363 : n157;
  assign n47405 = pi20 ? n47403 : n47404;
  assign n47406 = pi19 ? n36781 : n47405;
  assign n47407 = pi18 ? n36781 : n47406;
  assign n47408 = pi17 ? n47407 : n46786;
  assign n47409 = pi16 ? n47402 : n47408;
  assign n47410 = pi22 ? n46275 : n43198;
  assign n47411 = pi21 ? n32 : n47410;
  assign n47412 = pi20 ? n47411 : n43198;
  assign n47413 = pi19 ? n47412 : n43198;
  assign n47414 = pi18 ? n32 : n47413;
  assign n47415 = pi17 ? n32 : n47414;
  assign n47416 = pi20 ? n47403 : n34831;
  assign n47417 = pi19 ? n44208 : n47416;
  assign n47418 = pi18 ? n36781 : n47417;
  assign n47419 = pi17 ? n47418 : n45685;
  assign n47420 = pi16 ? n47415 : n47419;
  assign n47421 = pi15 ? n47409 : n47420;
  assign n47422 = pi14 ? n47395 : n47421;
  assign n47423 = pi13 ? n47359 : n47422;
  assign n47424 = pi12 ? n47295 : n47423;
  assign n47425 = pi11 ? n47236 : n47424;
  assign n47426 = pi10 ? n47075 : n47425;
  assign n47427 = pi09 ? n46850 : n47426;
  assign n47428 = pi21 ? n31924 : n31885;
  assign n47429 = pi20 ? n47428 : n20563;
  assign n47430 = pi19 ? n20563 : n47429;
  assign n47431 = pi18 ? n40497 : n47430;
  assign n47432 = pi21 ? n31294 : n20563;
  assign n47433 = pi21 ? n31924 : n30195;
  assign n47434 = pi20 ? n47432 : n47433;
  assign n47435 = pi20 ? n30195 : n31903;
  assign n47436 = pi19 ? n47434 : n47435;
  assign n47437 = pi20 ? n14844 : n3023;
  assign n47438 = pi19 ? n46822 : n47437;
  assign n47439 = pi18 ? n47436 : n47438;
  assign n47440 = pi17 ? n47431 : n47439;
  assign n47441 = pi16 ? n32 : n47440;
  assign n47442 = pi15 ? n32 : n47441;
  assign n47443 = pi18 ? n40510 : n20563;
  assign n47444 = pi20 ? n30195 : n33964;
  assign n47445 = pi19 ? n32876 : n47444;
  assign n47446 = pi20 ? n3086 : n3067;
  assign n47447 = pi19 ? n37 : n47446;
  assign n47448 = pi18 ? n47445 : n47447;
  assign n47449 = pi17 ? n47443 : n47448;
  assign n47450 = pi16 ? n32 : n47449;
  assign n47451 = pi18 ? n39373 : n20563;
  assign n47452 = pi20 ? n30867 : n31298;
  assign n47453 = pi19 ? n20563 : n47452;
  assign n47454 = pi20 ? n8742 : n3067;
  assign n47455 = pi19 ? n37 : n47454;
  assign n47456 = pi18 ? n47453 : n47455;
  assign n47457 = pi17 ? n47451 : n47456;
  assign n47458 = pi16 ? n32 : n47457;
  assign n47459 = pi15 ? n47450 : n47458;
  assign n47460 = pi14 ? n47442 : n47459;
  assign n47461 = pi13 ? n32 : n47460;
  assign n47462 = pi12 ? n32 : n47461;
  assign n47463 = pi11 ? n32 : n47462;
  assign n47464 = pi10 ? n32 : n47463;
  assign n47465 = pi20 ? n3086 : n17032;
  assign n47466 = pi19 ? n37 : n47465;
  assign n47467 = pi18 ? n33285 : n47466;
  assign n47468 = pi17 ? n46302 : n47467;
  assign n47469 = pi16 ? n32 : n47468;
  assign n47470 = pi17 ? n46832 : n46862;
  assign n47471 = pi16 ? n32 : n47470;
  assign n47472 = pi15 ? n47469 : n47471;
  assign n47473 = pi18 ? n33858 : n46868;
  assign n47474 = pi17 ? n46866 : n47473;
  assign n47475 = pi16 ? n32 : n47474;
  assign n47476 = pi20 ? n3090 : n2566;
  assign n47477 = pi19 ? n37 : n47476;
  assign n47478 = pi18 ? n32288 : n47477;
  assign n47479 = pi17 ? n20563 : n47478;
  assign n47480 = pi16 ? n32 : n47479;
  assign n47481 = pi15 ? n47475 : n47480;
  assign n47482 = pi14 ? n47472 : n47481;
  assign n47483 = pi19 ? n34920 : n33965;
  assign n47484 = pi20 ? n942 : n14835;
  assign n47485 = pi19 ? n9824 : n47484;
  assign n47486 = pi18 ? n47483 : n47485;
  assign n47487 = pi17 ? n20563 : n47486;
  assign n47488 = pi16 ? n46326 : n47487;
  assign n47489 = pi20 ? n577 : n2579;
  assign n47490 = pi19 ? n37 : n47489;
  assign n47491 = pi18 ? n34899 : n47490;
  assign n47492 = pi17 ? n20563 : n47491;
  assign n47493 = pi16 ? n45233 : n47492;
  assign n47494 = pi15 ? n47488 : n47493;
  assign n47495 = pi19 ? n36930 : n37;
  assign n47496 = pi22 ? n43747 : n32;
  assign n47497 = pi21 ? n47496 : n32;
  assign n47498 = pi20 ? n577 : n47497;
  assign n47499 = pi19 ? n37 : n47498;
  assign n47500 = pi18 ? n47495 : n47499;
  assign n47501 = pi17 ? n20563 : n47500;
  assign n47502 = pi16 ? n44635 : n47501;
  assign n47503 = pi22 ? n26981 : n32;
  assign n47504 = pi21 ? n47503 : n32;
  assign n47505 = pi20 ? n649 : n47504;
  assign n47506 = pi19 ? n37 : n47505;
  assign n47507 = pi18 ? n33916 : n47506;
  assign n47508 = pi17 ? n20563 : n47507;
  assign n47509 = pi16 ? n44223 : n47508;
  assign n47510 = pi15 ? n47502 : n47509;
  assign n47511 = pi14 ? n47494 : n47510;
  assign n47512 = pi13 ? n47482 : n47511;
  assign n47513 = pi21 ? n30195 : n30843;
  assign n47514 = pi20 ? n20563 : n47513;
  assign n47515 = pi19 ? n47514 : n37;
  assign n47516 = pi18 ? n47515 : n47506;
  assign n47517 = pi17 ? n20563 : n47516;
  assign n47518 = pi16 ? n45243 : n47517;
  assign n47519 = pi22 ? n20340 : n32;
  assign n47520 = pi21 ? n47519 : n32;
  assign n47521 = pi20 ? n46908 : n47520;
  assign n47522 = pi19 ? n37 : n47521;
  assign n47523 = pi18 ? n37029 : n47522;
  assign n47524 = pi17 ? n20563 : n47523;
  assign n47525 = pi16 ? n46349 : n47524;
  assign n47526 = pi15 ? n47518 : n47525;
  assign n47527 = pi19 ? n47452 : n37;
  assign n47528 = pi20 ? n46915 : n2653;
  assign n47529 = pi19 ? n8802 : n47528;
  assign n47530 = pi18 ? n47527 : n47529;
  assign n47531 = pi17 ? n20563 : n47530;
  assign n47532 = pi16 ? n43664 : n47531;
  assign n47533 = pi20 ? n31770 : n2470;
  assign n47534 = pi19 ? n8802 : n47533;
  assign n47535 = pi18 ? n37 : n47534;
  assign n47536 = pi17 ? n44249 : n47535;
  assign n47537 = pi16 ? n43664 : n47536;
  assign n47538 = pi15 ? n47532 : n47537;
  assign n47539 = pi14 ? n47526 : n47538;
  assign n47540 = pi20 ? n20563 : n30195;
  assign n47541 = pi19 ? n20563 : n47540;
  assign n47542 = pi18 ? n20563 : n47541;
  assign n47543 = pi20 ? n47513 : n37;
  assign n47544 = pi19 ? n47543 : n37;
  assign n47545 = pi20 ? n2094 : n2470;
  assign n47546 = pi19 ? n37 : n47545;
  assign n47547 = pi18 ? n47544 : n47546;
  assign n47548 = pi17 ? n47542 : n47547;
  assign n47549 = pi16 ? n44671 : n47548;
  assign n47550 = pi20 ? n2085 : n2554;
  assign n47551 = pi19 ? n37 : n47550;
  assign n47552 = pi18 ? n42265 : n47551;
  assign n47553 = pi17 ? n20563 : n47552;
  assign n47554 = pi16 ? n43224 : n47553;
  assign n47555 = pi15 ? n47549 : n47554;
  assign n47556 = pi20 ? n2107 : n2679;
  assign n47557 = pi19 ? n37 : n47556;
  assign n47558 = pi18 ? n37 : n47557;
  assign n47559 = pi17 ? n20563 : n47558;
  assign n47560 = pi16 ? n43228 : n47559;
  assign n47561 = pi20 ? n31925 : n30195;
  assign n47562 = pi19 ? n20563 : n47561;
  assign n47563 = pi18 ? n20563 : n47562;
  assign n47564 = pi18 ? n32934 : n46940;
  assign n47565 = pi17 ? n47563 : n47564;
  assign n47566 = pi16 ? n43249 : n47565;
  assign n47567 = pi15 ? n47560 : n47566;
  assign n47568 = pi14 ? n47555 : n47567;
  assign n47569 = pi13 ? n47539 : n47568;
  assign n47570 = pi12 ? n47512 : n47569;
  assign n47571 = pi19 ? n37 : n18182;
  assign n47572 = pi18 ? n32934 : n47571;
  assign n47573 = pi17 ? n47563 : n47572;
  assign n47574 = pi16 ? n44275 : n47573;
  assign n47575 = pi20 ? n20563 : n30867;
  assign n47576 = pi19 ? n20563 : n47575;
  assign n47577 = pi18 ? n20563 : n47576;
  assign n47578 = pi17 ? n47577 : n46954;
  assign n47579 = pi16 ? n42656 : n47578;
  assign n47580 = pi15 ? n47574 : n47579;
  assign n47581 = pi17 ? n47577 : n46963;
  assign n47582 = pi16 ? n42656 : n47581;
  assign n47583 = pi16 ? n42656 : n46970;
  assign n47584 = pi15 ? n47582 : n47583;
  assign n47585 = pi14 ? n47580 : n47584;
  assign n47586 = pi16 ? n42682 : n46974;
  assign n47587 = pi16 ? n42195 : n46976;
  assign n47588 = pi15 ? n47586 : n47587;
  assign n47589 = pi18 ? n20563 : n32872;
  assign n47590 = pi17 ? n47589 : n46982;
  assign n47591 = pi16 ? n43256 : n47590;
  assign n47592 = pi19 ? n38982 : n20563;
  assign n47593 = pi18 ? n32 : n47592;
  assign n47594 = pi17 ? n32 : n47593;
  assign n47595 = pi17 ? n42657 : n46991;
  assign n47596 = pi16 ? n47594 : n47595;
  assign n47597 = pi15 ? n47591 : n47596;
  assign n47598 = pi14 ? n47588 : n47597;
  assign n47599 = pi13 ? n47585 : n47598;
  assign n47600 = pi21 ? n37 : n26687;
  assign n47601 = pi20 ? n47600 : n32;
  assign n47602 = pi19 ? n37 : n47601;
  assign n47603 = pi18 ? n37 : n47602;
  assign n47604 = pi17 ? n42657 : n47603;
  assign n47605 = pi16 ? n42208 : n47604;
  assign n47606 = pi16 ? n42208 : n47008;
  assign n47607 = pi15 ? n47605 : n47606;
  assign n47608 = pi20 ? n2983 : n99;
  assign n47609 = pi19 ? n47608 : n99;
  assign n47610 = pi20 ? n33072 : n32;
  assign n47611 = pi19 ? n99 : n47610;
  assign n47612 = pi18 ? n47609 : n47611;
  assign n47613 = pi17 ? n44732 : n47612;
  assign n47614 = pi16 ? n41632 : n47613;
  assign n47615 = pi20 ? n3032 : n99;
  assign n47616 = pi19 ? n47615 : n99;
  assign n47617 = pi18 ? n47616 : n47611;
  assign n47618 = pi17 ? n47018 : n47617;
  assign n47619 = pi16 ? n41632 : n47618;
  assign n47620 = pi15 ? n47614 : n47619;
  assign n47621 = pi14 ? n47607 : n47620;
  assign n47622 = pi19 ? n47029 : n18701;
  assign n47623 = pi18 ? n99 : n47622;
  assign n47624 = pi17 ? n42647 : n47623;
  assign n47625 = pi16 ? n41643 : n47624;
  assign n47626 = pi19 ? n20563 : n37618;
  assign n47627 = pi18 ? n20563 : n47626;
  assign n47628 = pi19 ? n11445 : n16319;
  assign n47629 = pi18 ? n38578 : n47628;
  assign n47630 = pi17 ? n47627 : n47629;
  assign n47631 = pi16 ? n41643 : n47630;
  assign n47632 = pi15 ? n47625 : n47631;
  assign n47633 = pi21 ? n2957 : n218;
  assign n47634 = pi20 ? n47633 : n99;
  assign n47635 = pi19 ? n47634 : n47046;
  assign n47636 = pi21 ? n5176 : n3523;
  assign n47637 = pi20 ? n47636 : n32;
  assign n47638 = pi19 ? n47049 : n47637;
  assign n47639 = pi18 ? n47635 : n47638;
  assign n47640 = pi17 ? n47044 : n47639;
  assign n47641 = pi16 ? n41643 : n47640;
  assign n47642 = pi19 ? n47064 : n19276;
  assign n47643 = pi18 ? n47063 : n47642;
  assign n47644 = pi17 ? n42663 : n47643;
  assign n47645 = pi16 ? n42701 : n47644;
  assign n47646 = pi15 ? n47641 : n47645;
  assign n47647 = pi14 ? n47632 : n47646;
  assign n47648 = pi13 ? n47621 : n47647;
  assign n47649 = pi12 ? n47599 : n47648;
  assign n47650 = pi11 ? n47570 : n47649;
  assign n47651 = pi19 ? n42915 : n30097;
  assign n47652 = pi18 ? n20563 : n47651;
  assign n47653 = pi21 ? n16438 : n3523;
  assign n47654 = pi20 ? n47653 : n32;
  assign n47655 = pi19 ? n99 : n47654;
  assign n47656 = pi18 ? n34285 : n47655;
  assign n47657 = pi17 ? n47652 : n47656;
  assign n47658 = pi16 ? n42701 : n47657;
  assign n47659 = pi20 ? n41375 : n38969;
  assign n47660 = pi19 ? n32876 : n47659;
  assign n47661 = pi18 ? n20563 : n47660;
  assign n47662 = pi20 ? n3046 : n37;
  assign n47663 = pi19 ? n99 : n47662;
  assign n47664 = pi22 ? n37 : n745;
  assign n47665 = pi21 ? n47664 : n204;
  assign n47666 = pi20 ? n7346 : n47665;
  assign n47667 = pi20 ? n33587 : n32;
  assign n47668 = pi19 ? n47666 : n47667;
  assign n47669 = pi18 ? n47663 : n47668;
  assign n47670 = pi17 ? n47661 : n47669;
  assign n47671 = pi16 ? n42701 : n47670;
  assign n47672 = pi15 ? n47658 : n47671;
  assign n47673 = pi20 ? n47099 : n37;
  assign n47674 = pi19 ? n20563 : n47673;
  assign n47675 = pi18 ? n20563 : n47674;
  assign n47676 = pi19 ? n1017 : n47667;
  assign n47677 = pi18 ? n47103 : n47676;
  assign n47678 = pi17 ? n47675 : n47677;
  assign n47679 = pi16 ? n40025 : n47678;
  assign n47680 = pi20 ? n42433 : n37;
  assign n47681 = pi19 ? n20563 : n47680;
  assign n47682 = pi18 ? n20563 : n47681;
  assign n47683 = pi19 ? n32663 : n20137;
  assign n47684 = pi18 ? n37 : n47683;
  assign n47685 = pi17 ? n47682 : n47684;
  assign n47686 = pi16 ? n41183 : n47685;
  assign n47687 = pi15 ? n47679 : n47686;
  assign n47688 = pi14 ? n47672 : n47687;
  assign n47689 = pi19 ? n34246 : n31299;
  assign n47690 = pi18 ? n20563 : n47689;
  assign n47691 = pi19 ? n12589 : n47093;
  assign n47692 = pi18 ? n17061 : n47691;
  assign n47693 = pi17 ? n47690 : n47692;
  assign n47694 = pi16 ? n41183 : n47693;
  assign n47695 = pi20 ? n37 : n13116;
  assign n47696 = pi19 ? n20563 : n47695;
  assign n47697 = pi18 ? n20563 : n47696;
  assign n47698 = pi20 ? n31614 : n32;
  assign n47699 = pi19 ? n12589 : n47698;
  assign n47700 = pi18 ? n47128 : n47699;
  assign n47701 = pi17 ? n47697 : n47700;
  assign n47702 = pi16 ? n41183 : n47701;
  assign n47703 = pi15 ? n47694 : n47702;
  assign n47704 = pi20 ? n5371 : n32;
  assign n47705 = pi19 ? n12589 : n47704;
  assign n47706 = pi18 ? n47134 : n47705;
  assign n47707 = pi17 ? n42690 : n47706;
  assign n47708 = pi16 ? n41183 : n47707;
  assign n47709 = pi20 ? n23406 : n32;
  assign n47710 = pi19 ? n47140 : n47709;
  assign n47711 = pi18 ? n9770 : n47710;
  assign n47712 = pi17 ? n42196 : n47711;
  assign n47713 = pi16 ? n47058 : n47712;
  assign n47714 = pi15 ? n47708 : n47713;
  assign n47715 = pi14 ? n47703 : n47714;
  assign n47716 = pi13 ? n47688 : n47715;
  assign n47717 = pi19 ? n32876 : n9814;
  assign n47718 = pi18 ? n20563 : n47717;
  assign n47719 = pi19 ? n47153 : n20238;
  assign n47720 = pi18 ? n139 : n47719;
  assign n47721 = pi17 ? n47718 : n47720;
  assign n47722 = pi16 ? n47058 : n47721;
  assign n47723 = pi19 ? n47159 : n32933;
  assign n47724 = pi18 ? n20563 : n47723;
  assign n47725 = pi21 ? n584 : n2007;
  assign n47726 = pi20 ? n47725 : n47163;
  assign n47727 = pi19 ? n47726 : n2004;
  assign n47728 = pi18 ? n47727 : n47167;
  assign n47729 = pi17 ? n47724 : n47728;
  assign n47730 = pi16 ? n47058 : n47729;
  assign n47731 = pi15 ? n47722 : n47730;
  assign n47732 = pi19 ? n47175 : n17906;
  assign n47733 = pi18 ? n47174 : n47732;
  assign n47734 = pi17 ? n43257 : n47733;
  assign n47735 = pi16 ? n47058 : n47734;
  assign n47736 = pi16 ? n47058 : n47183;
  assign n47737 = pi15 ? n47735 : n47736;
  assign n47738 = pi14 ? n47731 : n47737;
  assign n47739 = pi22 ? n233 : n22498;
  assign n47740 = pi21 ? n47739 : n32;
  assign n47741 = pi20 ? n47740 : n32;
  assign n47742 = pi19 ? n19358 : n47741;
  assign n47743 = pi18 ? n45798 : n47742;
  assign n47744 = pi17 ? n42216 : n47743;
  assign n47745 = pi16 ? n40512 : n47744;
  assign n47746 = pi21 ? n32 : n45620;
  assign n47747 = pi20 ? n47746 : n30868;
  assign n47748 = pi19 ? n47747 : n30868;
  assign n47749 = pi18 ? n32 : n47748;
  assign n47750 = pi17 ? n32 : n47749;
  assign n47751 = pi21 ? n30868 : n31294;
  assign n47752 = pi20 ? n30868 : n47751;
  assign n47753 = pi19 ? n47752 : n37;
  assign n47754 = pi18 ? n30868 : n47753;
  assign n47755 = pi19 ? n5024 : n47741;
  assign n47756 = pi18 ? n47203 : n47755;
  assign n47757 = pi17 ? n47754 : n47756;
  assign n47758 = pi16 ? n47750 : n47757;
  assign n47759 = pi15 ? n47745 : n47758;
  assign n47760 = pi20 ? n47746 : n38754;
  assign n47761 = pi19 ? n47760 : n47211;
  assign n47762 = pi18 ? n32 : n47761;
  assign n47763 = pi17 ? n32 : n47762;
  assign n47764 = pi19 ? n46033 : n15882;
  assign n47765 = pi18 ? n37 : n47764;
  assign n47766 = pi17 ? n42203 : n47765;
  assign n47767 = pi16 ? n47763 : n47766;
  assign n47768 = pi22 ? n32 : n37251;
  assign n47769 = pi21 ? n32 : n47768;
  assign n47770 = pi20 ? n47769 : n47221;
  assign n47771 = pi19 ? n47770 : n47224;
  assign n47772 = pi18 ? n32 : n47771;
  assign n47773 = pi17 ? n32 : n47772;
  assign n47774 = pi19 ? n47228 : n15882;
  assign n47775 = pi18 ? n17225 : n47774;
  assign n47776 = pi17 ? n42203 : n47775;
  assign n47777 = pi16 ? n47773 : n47776;
  assign n47778 = pi15 ? n47767 : n47777;
  assign n47779 = pi14 ? n47759 : n47778;
  assign n47780 = pi13 ? n47738 : n47779;
  assign n47781 = pi12 ? n47716 : n47780;
  assign n47782 = pi19 ? n47238 : n9483;
  assign n47783 = pi18 ? n7677 : n47782;
  assign n47784 = pi17 ? n42203 : n47783;
  assign n47785 = pi16 ? n40534 : n47784;
  assign n47786 = pi19 ? n2730 : n4009;
  assign n47787 = pi18 ? n37 : n47786;
  assign n47788 = pi17 ? n42203 : n47787;
  assign n47789 = pi16 ? n40534 : n47788;
  assign n47790 = pi15 ? n47785 : n47789;
  assign n47791 = pi19 ? n5064 : n4117;
  assign n47792 = pi18 ? n47248 : n47791;
  assign n47793 = pi17 ? n42196 : n47792;
  assign n47794 = pi16 ? n40534 : n47793;
  assign n47795 = pi19 ? n47259 : n4117;
  assign n47796 = pi18 ? n47257 : n47795;
  assign n47797 = pi17 ? n42196 : n47796;
  assign n47798 = pi16 ? n40534 : n47797;
  assign n47799 = pi15 ? n47794 : n47798;
  assign n47800 = pi14 ? n47790 : n47799;
  assign n47801 = pi21 ? n46116 : n31924;
  assign n47802 = pi20 ? n20563 : n47801;
  assign n47803 = pi19 ? n47802 : n37;
  assign n47804 = pi18 ? n20563 : n47803;
  assign n47805 = pi17 ? n47804 : n47271;
  assign n47806 = pi16 ? n39375 : n47805;
  assign n47807 = pi19 ? n47274 : n10012;
  assign n47808 = pi18 ? n37 : n47807;
  assign n47809 = pi17 ? n47804 : n47808;
  assign n47810 = pi16 ? n39375 : n47809;
  assign n47811 = pi15 ? n47806 : n47810;
  assign n47812 = pi19 ? n47281 : n32933;
  assign n47813 = pi18 ? n20563 : n47812;
  assign n47814 = pi19 ? n28767 : n7833;
  assign n47815 = pi18 ? n47284 : n47814;
  assign n47816 = pi17 ? n47813 : n47815;
  assign n47817 = pi16 ? n40499 : n47816;
  assign n47818 = pi19 ? n47288 : n1823;
  assign n47819 = pi18 ? n47284 : n47818;
  assign n47820 = pi17 ? n47813 : n47819;
  assign n47821 = pi16 ? n40499 : n47820;
  assign n47822 = pi15 ? n47817 : n47821;
  assign n47823 = pi14 ? n47811 : n47822;
  assign n47824 = pi13 ? n47800 : n47823;
  assign n47825 = pi19 ? n40496 : n30868;
  assign n47826 = pi18 ? n32 : n47825;
  assign n47827 = pi17 ? n32 : n47826;
  assign n47828 = pi20 ? n31903 : n3393;
  assign n47829 = pi19 ? n47300 : n47828;
  assign n47830 = pi18 ? n30868 : n47829;
  assign n47831 = pi19 ? n47306 : n1823;
  assign n47832 = pi18 ? n47305 : n47831;
  assign n47833 = pi17 ? n47830 : n47832;
  assign n47834 = pi16 ? n47827 : n47833;
  assign n47835 = pi21 ? n32 : n47321;
  assign n47836 = pi20 ? n47835 : n30868;
  assign n47837 = pi19 ? n47836 : n30868;
  assign n47838 = pi18 ? n32 : n47837;
  assign n47839 = pi17 ? n32 : n47838;
  assign n47840 = pi21 ? n39315 : n99;
  assign n47841 = pi20 ? n47840 : n2238;
  assign n47842 = pi19 ? n47312 : n47841;
  assign n47843 = pi18 ? n30868 : n47842;
  assign n47844 = pi18 ? n47316 : n46695;
  assign n47845 = pi17 ? n47843 : n47844;
  assign n47846 = pi16 ? n47839 : n47845;
  assign n47847 = pi15 ? n47834 : n47846;
  assign n47848 = pi21 ? n32 : n45598;
  assign n47849 = pi20 ? n47848 : n30868;
  assign n47850 = pi19 ? n47849 : n30868;
  assign n47851 = pi18 ? n32 : n47850;
  assign n47852 = pi17 ? n32 : n47851;
  assign n47853 = pi19 ? n30868 : n47328;
  assign n47854 = pi18 ? n30868 : n47853;
  assign n47855 = pi17 ? n47854 : n47338;
  assign n47856 = pi16 ? n47852 : n47855;
  assign n47857 = pi20 ? n32 : n36798;
  assign n47858 = pi19 ? n47857 : n36798;
  assign n47859 = pi18 ? n32 : n47858;
  assign n47860 = pi17 ? n32 : n47859;
  assign n47861 = pi21 ? n37253 : n139;
  assign n47862 = pi20 ? n47861 : n139;
  assign n47863 = pi19 ? n33792 : n47862;
  assign n47864 = pi18 ? n33792 : n47863;
  assign n47865 = pi17 ? n47864 : n47355;
  assign n47866 = pi16 ? n47860 : n47865;
  assign n47867 = pi15 ? n47856 : n47866;
  assign n47868 = pi14 ? n47847 : n47867;
  assign n47869 = pi22 ? n36659 : n36762;
  assign n47870 = pi21 ? n47869 : n139;
  assign n47871 = pi20 ? n47870 : n47366;
  assign n47872 = pi19 ? n36659 : n47871;
  assign n47873 = pi18 ? n47363 : n47872;
  assign n47874 = pi17 ? n47873 : n47377;
  assign n47875 = pi16 ? n47860 : n47874;
  assign n47876 = pi22 ? n46757 : n36659;
  assign n47877 = pi21 ? n47876 : n36659;
  assign n47878 = pi20 ? n32 : n47877;
  assign n47879 = pi19 ? n47878 : n36659;
  assign n47880 = pi18 ? n32 : n47879;
  assign n47881 = pi17 ? n32 : n47880;
  assign n47882 = pi22 ? n36659 : n36710;
  assign n47883 = pi21 ? n47882 : n335;
  assign n47884 = pi20 ? n47883 : n335;
  assign n47885 = pi19 ? n36659 : n47884;
  assign n47886 = pi18 ? n36659 : n47885;
  assign n47887 = pi18 ? n47391 : n32119;
  assign n47888 = pi17 ? n47886 : n47887;
  assign n47889 = pi16 ? n47881 : n47888;
  assign n47890 = pi15 ? n47875 : n47889;
  assign n47891 = pi20 ? n32 : n47398;
  assign n47892 = pi19 ? n47891 : n43198;
  assign n47893 = pi18 ? n32 : n47892;
  assign n47894 = pi17 ? n32 : n47893;
  assign n47895 = pi22 ? n42171 : n363;
  assign n47896 = pi21 ? n36798 : n47895;
  assign n47897 = pi20 ? n47896 : n47404;
  assign n47898 = pi19 ? n36781 : n47897;
  assign n47899 = pi18 ? n36781 : n47898;
  assign n47900 = pi17 ? n47899 : n46786;
  assign n47901 = pi16 ? n47894 : n47900;
  assign n47902 = pi22 ? n46789 : n43198;
  assign n47903 = pi21 ? n47902 : n43198;
  assign n47904 = pi20 ? n32 : n47903;
  assign n47905 = pi19 ? n47904 : n43198;
  assign n47906 = pi18 ? n32 : n47905;
  assign n47907 = pi17 ? n32 : n47906;
  assign n47908 = pi21 ? n36798 : n42171;
  assign n47909 = pi20 ? n47908 : n34831;
  assign n47910 = pi19 ? n44208 : n47909;
  assign n47911 = pi18 ? n36781 : n47910;
  assign n47912 = pi17 ? n47911 : n45685;
  assign n47913 = pi16 ? n47907 : n47912;
  assign n47914 = pi15 ? n47901 : n47913;
  assign n47915 = pi14 ? n47890 : n47914;
  assign n47916 = pi13 ? n47868 : n47915;
  assign n47917 = pi12 ? n47824 : n47916;
  assign n47918 = pi11 ? n47781 : n47917;
  assign n47919 = pi10 ? n47650 : n47918;
  assign n47920 = pi09 ? n47464 : n47919;
  assign n47921 = pi08 ? n47427 : n47920;
  assign n47922 = pi18 ? n40023 : n20563;
  assign n47923 = pi20 ? n37 : n16991;
  assign n47924 = pi19 ? n37 : n47923;
  assign n47925 = pi18 ? n34258 : n47924;
  assign n47926 = pi17 ? n47922 : n47925;
  assign n47927 = pi16 ? n32 : n47926;
  assign n47928 = pi15 ? n32 : n47927;
  assign n47929 = pi18 ? n41181 : n20563;
  assign n47930 = pi20 ? n3086 : n17001;
  assign n47931 = pi19 ? n33949 : n47930;
  assign n47932 = pi18 ? n20563 : n47931;
  assign n47933 = pi17 ? n47929 : n47932;
  assign n47934 = pi16 ? n32 : n47933;
  assign n47935 = pi18 ? n42239 : n20563;
  assign n47936 = pi20 ? n37 : n17001;
  assign n47937 = pi19 ? n30097 : n47936;
  assign n47938 = pi18 ? n20563 : n47937;
  assign n47939 = pi17 ? n47935 : n47938;
  assign n47940 = pi16 ? n32 : n47939;
  assign n47941 = pi15 ? n47934 : n47940;
  assign n47942 = pi14 ? n47928 : n47941;
  assign n47943 = pi13 ? n32 : n47942;
  assign n47944 = pi12 ? n32 : n47943;
  assign n47945 = pi11 ? n32 : n47944;
  assign n47946 = pi10 ? n32 : n47945;
  assign n47947 = pi18 ? n47056 : n20563;
  assign n47948 = pi21 ? n12003 : n32;
  assign n47949 = pi20 ? n37 : n47948;
  assign n47950 = pi19 ? n37 : n47949;
  assign n47951 = pi18 ? n34869 : n47950;
  assign n47952 = pi17 ? n47947 : n47951;
  assign n47953 = pi16 ? n32 : n47952;
  assign n47954 = pi18 ? n40497 : n20563;
  assign n47955 = pi23 ? n1432 : n5630;
  assign n47956 = pi22 ? n47955 : n32;
  assign n47957 = pi21 ? n47956 : n32;
  assign n47958 = pi20 ? n3625 : n47957;
  assign n47959 = pi19 ? n37 : n47958;
  assign n47960 = pi18 ? n34258 : n47959;
  assign n47961 = pi17 ? n47954 : n47960;
  assign n47962 = pi16 ? n32 : n47961;
  assign n47963 = pi15 ? n47953 : n47962;
  assign n47964 = pi18 ? n45366 : n20563;
  assign n47965 = pi20 ? n3096 : n31331;
  assign n47966 = pi19 ? n37 : n47965;
  assign n47967 = pi18 ? n33245 : n47966;
  assign n47968 = pi17 ? n47964 : n47967;
  assign n47969 = pi16 ? n32 : n47968;
  assign n47970 = pi20 ? n3086 : n16621;
  assign n47971 = pi19 ? n37 : n47970;
  assign n47972 = pi18 ? n34869 : n47971;
  assign n47973 = pi17 ? n45707 : n47972;
  assign n47974 = pi16 ? n32 : n47973;
  assign n47975 = pi15 ? n47969 : n47974;
  assign n47976 = pi14 ? n47963 : n47975;
  assign n47977 = pi21 ? n23334 : n32;
  assign n47978 = pi20 ? n40578 : n47977;
  assign n47979 = pi19 ? n37 : n47978;
  assign n47980 = pi18 ? n34869 : n47979;
  assign n47981 = pi17 ? n46859 : n47980;
  assign n47982 = pi16 ? n32 : n47981;
  assign n47983 = pi20 ? n20157 : n2579;
  assign n47984 = pi19 ? n37 : n47983;
  assign n47985 = pi18 ? n32275 : n47984;
  assign n47986 = pi17 ? n45715 : n47985;
  assign n47987 = pi16 ? n32 : n47986;
  assign n47988 = pi15 ? n47982 : n47987;
  assign n47989 = pi20 ? n649 : n2579;
  assign n47990 = pi19 ? n37 : n47989;
  assign n47991 = pi18 ? n34295 : n47990;
  assign n47992 = pi17 ? n46866 : n47991;
  assign n47993 = pi16 ? n32 : n47992;
  assign n47994 = pi20 ? n649 : n2638;
  assign n47995 = pi19 ? n37 : n47994;
  assign n47996 = pi18 ? n33285 : n47995;
  assign n47997 = pi17 ? n20563 : n47996;
  assign n47998 = pi16 ? n44635 : n47997;
  assign n47999 = pi15 ? n47993 : n47998;
  assign n48000 = pi14 ? n47988 : n47999;
  assign n48001 = pi13 ? n47976 : n48000;
  assign n48002 = pi20 ? n37 : n2638;
  assign n48003 = pi19 ? n37 : n48002;
  assign n48004 = pi18 ? n32275 : n48003;
  assign n48005 = pi17 ? n20563 : n48004;
  assign n48006 = pi16 ? n45740 : n48005;
  assign n48007 = pi20 ? n21635 : n2653;
  assign n48008 = pi19 ? n37 : n48007;
  assign n48009 = pi18 ? n32275 : n48008;
  assign n48010 = pi17 ? n20563 : n48009;
  assign n48011 = pi16 ? n46885 : n48010;
  assign n48012 = pi15 ? n48006 : n48011;
  assign n48013 = pi20 ? n577 : n2653;
  assign n48014 = pi19 ? n37 : n48013;
  assign n48015 = pi18 ? n33299 : n48014;
  assign n48016 = pi17 ? n20563 : n48015;
  assign n48017 = pi16 ? n44653 : n48016;
  assign n48018 = pi18 ? n32295 : n46893;
  assign n48019 = pi17 ? n20563 : n48018;
  assign n48020 = pi16 ? n44223 : n48019;
  assign n48021 = pi15 ? n48017 : n48020;
  assign n48022 = pi14 ? n48012 : n48021;
  assign n48023 = pi20 ? n2094 : n2679;
  assign n48024 = pi19 ? n37 : n48023;
  assign n48025 = pi18 ? n34358 : n48024;
  assign n48026 = pi17 ? n20563 : n48025;
  assign n48027 = pi16 ? n44671 : n48026;
  assign n48028 = pi23 ? n99 : n7420;
  assign n48029 = pi22 ? n37 : n48028;
  assign n48030 = pi21 ? n37 : n48029;
  assign n48031 = pi20 ? n48030 : n2701;
  assign n48032 = pi19 ? n37 : n48031;
  assign n48033 = pi18 ? n32295 : n48032;
  assign n48034 = pi17 ? n20563 : n48033;
  assign n48035 = pi16 ? n43675 : n48034;
  assign n48036 = pi15 ? n48027 : n48035;
  assign n48037 = pi18 ? n34358 : n46940;
  assign n48038 = pi17 ? n20563 : n48037;
  assign n48039 = pi16 ? n43685 : n48038;
  assign n48040 = pi23 ? n1342 : n685;
  assign n48041 = pi22 ? n37 : n48040;
  assign n48042 = pi21 ? n37 : n48041;
  assign n48043 = pi20 ? n48042 : n2638;
  assign n48044 = pi19 ? n37 : n48043;
  assign n48045 = pi18 ? n32899 : n48044;
  assign n48046 = pi17 ? n20563 : n48045;
  assign n48047 = pi16 ? n44688 : n48046;
  assign n48048 = pi15 ? n48039 : n48047;
  assign n48049 = pi14 ? n48036 : n48048;
  assign n48050 = pi13 ? n48022 : n48049;
  assign n48051 = pi12 ? n48001 : n48050;
  assign n48052 = pi23 ? n1432 : n685;
  assign n48053 = pi22 ? n37 : n48052;
  assign n48054 = pi21 ? n37 : n48053;
  assign n48055 = pi20 ? n48054 : n2653;
  assign n48056 = pi19 ? n37 : n48055;
  assign n48057 = pi18 ? n32349 : n48056;
  assign n48058 = pi17 ? n20563 : n48057;
  assign n48059 = pi16 ? n44688 : n48058;
  assign n48060 = pi21 ? n3392 : n14255;
  assign n48061 = pi20 ? n48060 : n1822;
  assign n48062 = pi19 ? n5029 : n48061;
  assign n48063 = pi18 ? n32899 : n48062;
  assign n48064 = pi17 ? n20563 : n48063;
  assign n48065 = pi16 ? n44248 : n48064;
  assign n48066 = pi15 ? n48059 : n48065;
  assign n48067 = pi20 ? n24493 : n1822;
  assign n48068 = pi19 ? n37 : n48067;
  assign n48069 = pi18 ? n34358 : n48068;
  assign n48070 = pi17 ? n20563 : n48069;
  assign n48071 = pi16 ? n44248 : n48070;
  assign n48072 = pi20 ? n2722 : n32;
  assign n48073 = pi19 ? n37 : n48072;
  assign n48074 = pi18 ? n34358 : n48073;
  assign n48075 = pi17 ? n20563 : n48074;
  assign n48076 = pi16 ? n43224 : n48075;
  assign n48077 = pi15 ? n48071 : n48076;
  assign n48078 = pi14 ? n48066 : n48077;
  assign n48079 = pi21 ? n9666 : n2721;
  assign n48080 = pi20 ? n48079 : n32;
  assign n48081 = pi19 ? n37 : n48080;
  assign n48082 = pi18 ? n32349 : n48081;
  assign n48083 = pi17 ? n20563 : n48082;
  assign n48084 = pi16 ? n43228 : n48083;
  assign n48085 = pi18 ? n32377 : n48073;
  assign n48086 = pi17 ? n20563 : n48085;
  assign n48087 = pi16 ? n43249 : n48086;
  assign n48088 = pi15 ? n48084 : n48087;
  assign n48089 = pi21 ? n37 : n3562;
  assign n48090 = pi20 ? n48089 : n32;
  assign n48091 = pi19 ? n37 : n48090;
  assign n48092 = pi18 ? n31939 : n48091;
  assign n48093 = pi17 ? n20563 : n48092;
  assign n48094 = pi16 ? n42646 : n48093;
  assign n48095 = pi21 ? n272 : n6132;
  assign n48096 = pi20 ? n48095 : n32;
  assign n48097 = pi19 ? n37 : n48096;
  assign n48098 = pi18 ? n32377 : n48097;
  assign n48099 = pi17 ? n20563 : n48098;
  assign n48100 = pi16 ? n42646 : n48099;
  assign n48101 = pi15 ? n48094 : n48100;
  assign n48102 = pi14 ? n48088 : n48101;
  assign n48103 = pi13 ? n48078 : n48102;
  assign n48104 = pi18 ? n32377 : n48091;
  assign n48105 = pi17 ? n20563 : n48104;
  assign n48106 = pi16 ? n42656 : n48105;
  assign n48107 = pi20 ? n389 : n32;
  assign n48108 = pi19 ? n37 : n48107;
  assign n48109 = pi18 ? n31939 : n48108;
  assign n48110 = pi17 ? n20563 : n48109;
  assign n48111 = pi16 ? n42682 : n48110;
  assign n48112 = pi15 ? n48106 : n48111;
  assign n48113 = pi19 ? n31280 : n19773;
  assign n48114 = pi21 ? n99 : n7137;
  assign n48115 = pi20 ? n48114 : n32;
  assign n48116 = pi19 ? n99 : n48115;
  assign n48117 = pi18 ? n48113 : n48116;
  assign n48118 = pi17 ? n20563 : n48117;
  assign n48119 = pi16 ? n42195 : n48118;
  assign n48120 = pi19 ? n37927 : n20563;
  assign n48121 = pi18 ? n32 : n48120;
  assign n48122 = pi17 ? n32 : n48121;
  assign n48123 = pi20 ? n30096 : n3039;
  assign n48124 = pi19 ? n48123 : n99;
  assign n48125 = pi18 ? n48124 : n47611;
  assign n48126 = pi17 ? n20563 : n48125;
  assign n48127 = pi16 ? n48122 : n48126;
  assign n48128 = pi15 ? n48119 : n48127;
  assign n48129 = pi14 ? n48112 : n48128;
  assign n48130 = pi20 ? n40755 : n226;
  assign n48131 = pi19 ? n48130 : n99;
  assign n48132 = pi18 ? n48131 : n46450;
  assign n48133 = pi17 ? n20563 : n48132;
  assign n48134 = pi16 ? n48122 : n48133;
  assign n48135 = pi18 ? n20563 : n40793;
  assign n48136 = pi20 ? n40755 : n99;
  assign n48137 = pi19 ? n48136 : n99;
  assign n48138 = pi21 ? n157 : n22911;
  assign n48139 = pi20 ? n48138 : n32;
  assign n48140 = pi19 ? n6542 : n48139;
  assign n48141 = pi18 ? n48137 : n48140;
  assign n48142 = pi17 ? n48135 : n48141;
  assign n48143 = pi16 ? n48122 : n48142;
  assign n48144 = pi15 ? n48134 : n48143;
  assign n48145 = pi19 ? n17013 : n32889;
  assign n48146 = pi21 ? n99 : n1027;
  assign n48147 = pi20 ? n99 : n48146;
  assign n48148 = pi21 ? n1027 : n3523;
  assign n48149 = pi20 ? n48148 : n32;
  assign n48150 = pi19 ? n48147 : n48149;
  assign n48151 = pi18 ? n48145 : n48150;
  assign n48152 = pi17 ? n20563 : n48151;
  assign n48153 = pi16 ? n47594 : n48152;
  assign n48154 = pi19 ? n37 : n33288;
  assign n48155 = pi18 ? n48154 : n48150;
  assign n48156 = pi17 ? n44680 : n48155;
  assign n48157 = pi16 ? n47594 : n48156;
  assign n48158 = pi15 ? n48153 : n48157;
  assign n48159 = pi14 ? n48144 : n48158;
  assign n48160 = pi13 ? n48129 : n48159;
  assign n48161 = pi12 ? n48103 : n48160;
  assign n48162 = pi11 ? n48051 : n48161;
  assign n48163 = pi18 ? n20563 : n38951;
  assign n48164 = pi20 ? n37 : n38343;
  assign n48165 = pi19 ? n48164 : n99;
  assign n48166 = pi20 ? n99 : n22941;
  assign n48167 = pi21 ? n1027 : n13465;
  assign n48168 = pi20 ? n48167 : n32;
  assign n48169 = pi19 ? n48166 : n48168;
  assign n48170 = pi18 ? n48165 : n48169;
  assign n48171 = pi17 ? n48163 : n48170;
  assign n48172 = pi16 ? n41632 : n48171;
  assign n48173 = pi22 ? n39190 : n30868;
  assign n48174 = pi21 ? n20563 : n48173;
  assign n48175 = pi20 ? n20563 : n48174;
  assign n48176 = pi19 ? n20563 : n48175;
  assign n48177 = pi18 ? n20563 : n48176;
  assign n48178 = pi19 ? n37 : n47662;
  assign n48179 = pi19 ? n32636 : n20124;
  assign n48180 = pi18 ? n48178 : n48179;
  assign n48181 = pi17 ? n48177 : n48180;
  assign n48182 = pi16 ? n41632 : n48181;
  assign n48183 = pi15 ? n48172 : n48182;
  assign n48184 = pi21 ? n36489 : n30868;
  assign n48185 = pi20 ? n20563 : n48184;
  assign n48186 = pi19 ? n20563 : n48185;
  assign n48187 = pi18 ? n20563 : n48186;
  assign n48188 = pi19 ? n37 : n28582;
  assign n48189 = pi19 ? n1017 : n20124;
  assign n48190 = pi18 ? n48188 : n48189;
  assign n48191 = pi17 ? n48187 : n48190;
  assign n48192 = pi16 ? n41632 : n48191;
  assign n48193 = pi17 ? n44680 : n47684;
  assign n48194 = pi16 ? n42689 : n48193;
  assign n48195 = pi15 ? n48192 : n48194;
  assign n48196 = pi14 ? n48183 : n48195;
  assign n48197 = pi18 ? n20563 : n40199;
  assign n48198 = pi19 ? n12589 : n47066;
  assign n48199 = pi18 ? n37 : n48198;
  assign n48200 = pi17 ? n48197 : n48199;
  assign n48201 = pi16 ? n42689 : n48200;
  assign n48202 = pi19 ? n9814 : n1806;
  assign n48203 = pi18 ? n48202 : n47699;
  assign n48204 = pi17 ? n43676 : n48203;
  assign n48205 = pi16 ? n42689 : n48204;
  assign n48206 = pi15 ? n48201 : n48205;
  assign n48207 = pi19 ? n12370 : n13192;
  assign n48208 = pi19 ? n12589 : n18375;
  assign n48209 = pi18 ? n48207 : n48208;
  assign n48210 = pi17 ? n43676 : n48209;
  assign n48211 = pi16 ? n41159 : n48210;
  assign n48212 = pi21 ? n28649 : n2678;
  assign n48213 = pi20 ? n48212 : n32;
  assign n48214 = pi19 ? n47140 : n48213;
  assign n48215 = pi18 ? n9815 : n48214;
  assign n48216 = pi17 ? n43676 : n48215;
  assign n48217 = pi16 ? n41159 : n48216;
  assign n48218 = pi15 ? n48211 : n48217;
  assign n48219 = pi14 ? n48206 : n48218;
  assign n48220 = pi13 ? n48196 : n48219;
  assign n48221 = pi22 ? n33792 : n37;
  assign n48222 = pi21 ? n29133 : n48221;
  assign n48223 = pi20 ? n20563 : n48222;
  assign n48224 = pi19 ? n20563 : n48223;
  assign n48225 = pi18 ? n20563 : n48224;
  assign n48226 = pi20 ? n24439 : n32;
  assign n48227 = pi19 ? n47153 : n48226;
  assign n48228 = pi18 ? n9796 : n48227;
  assign n48229 = pi17 ? n48225 : n48228;
  assign n48230 = pi16 ? n41159 : n48229;
  assign n48231 = pi20 ? n638 : n6377;
  assign n48232 = pi19 ? n48231 : n48226;
  assign n48233 = pi18 ? n37 : n48232;
  assign n48234 = pi17 ? n48163 : n48233;
  assign n48235 = pi16 ? n41159 : n48234;
  assign n48236 = pi15 ? n48230 : n48235;
  assign n48237 = pi20 ? n638 : n8927;
  assign n48238 = pi19 ? n48237 : n20585;
  assign n48239 = pi18 ? n7686 : n48238;
  assign n48240 = pi17 ? n42647 : n48239;
  assign n48241 = pi16 ? n41159 : n48240;
  assign n48242 = pi20 ? n37 : n18431;
  assign n48243 = pi19 ? n48242 : n19410;
  assign n48244 = pi18 ? n37 : n48243;
  assign n48245 = pi17 ? n42647 : n48244;
  assign n48246 = pi16 ? n40025 : n48245;
  assign n48247 = pi15 ? n48241 : n48246;
  assign n48248 = pi14 ? n48236 : n48247;
  assign n48249 = pi20 ? n8927 : n18431;
  assign n48250 = pi19 ? n48249 : n19440;
  assign n48251 = pi18 ? n37 : n48250;
  assign n48252 = pi17 ? n42647 : n48251;
  assign n48253 = pi16 ? n40025 : n48252;
  assign n48254 = pi21 ? n46060 : n30868;
  assign n48255 = pi20 ? n32 : n48254;
  assign n48256 = pi19 ? n48255 : n30868;
  assign n48257 = pi18 ? n32 : n48256;
  assign n48258 = pi17 ? n32 : n48257;
  assign n48259 = pi19 ? n30868 : n31267;
  assign n48260 = pi18 ? n30868 : n48259;
  assign n48261 = pi19 ? n19358 : n47180;
  assign n48262 = pi18 ? n6374 : n48261;
  assign n48263 = pi17 ? n48260 : n48262;
  assign n48264 = pi16 ? n48258 : n48263;
  assign n48265 = pi15 ? n48253 : n48264;
  assign n48266 = pi21 ? n28156 : n48173;
  assign n48267 = pi20 ? n32 : n48266;
  assign n48268 = pi19 ? n48267 : n30868;
  assign n48269 = pi18 ? n32 : n48268;
  assign n48270 = pi17 ? n32 : n48269;
  assign n48271 = pi19 ? n13337 : n8918;
  assign n48272 = pi18 ? n37 : n48271;
  assign n48273 = pi17 ? n42657 : n48272;
  assign n48274 = pi16 ? n48270 : n48273;
  assign n48275 = pi22 ? n42109 : n33792;
  assign n48276 = pi21 ? n46060 : n48275;
  assign n48277 = pi20 ? n32 : n48276;
  assign n48278 = pi21 ? n30868 : n33792;
  assign n48279 = pi20 ? n33792 : n48278;
  assign n48280 = pi19 ? n48277 : n48279;
  assign n48281 = pi18 ? n32 : n48280;
  assign n48282 = pi17 ? n32 : n48281;
  assign n48283 = pi19 ? n47228 : n8918;
  assign n48284 = pi18 ? n7677 : n48283;
  assign n48285 = pi17 ? n42657 : n48284;
  assign n48286 = pi16 ? n48282 : n48285;
  assign n48287 = pi15 ? n48274 : n48286;
  assign n48288 = pi14 ? n48265 : n48287;
  assign n48289 = pi13 ? n48248 : n48288;
  assign n48290 = pi12 ? n48220 : n48289;
  assign n48291 = pi19 ? n47238 : n8296;
  assign n48292 = pi18 ? n37 : n48291;
  assign n48293 = pi17 ? n42657 : n48292;
  assign n48294 = pi16 ? n46448 : n48293;
  assign n48295 = pi20 ? n37 : n18212;
  assign n48296 = pi19 ? n48295 : n4009;
  assign n48297 = pi18 ? n37 : n48296;
  assign n48298 = pi17 ? n42647 : n48297;
  assign n48299 = pi16 ? n46448 : n48298;
  assign n48300 = pi15 ? n48294 : n48299;
  assign n48301 = pi19 ? n2723 : n3211;
  assign n48302 = pi18 ? n47248 : n48301;
  assign n48303 = pi17 ? n42647 : n48302;
  assign n48304 = pi16 ? n46448 : n48303;
  assign n48305 = pi20 ? n9660 : n2722;
  assign n48306 = pi19 ? n48305 : n3211;
  assign n48307 = pi18 ? n47257 : n48306;
  assign n48308 = pi17 ? n42647 : n48307;
  assign n48309 = pi16 ? n46448 : n48308;
  assign n48310 = pi15 ? n48304 : n48309;
  assign n48311 = pi14 ? n48300 : n48310;
  assign n48312 = pi20 ? n3393 : n32833;
  assign n48313 = pi19 ? n48312 : n5831;
  assign n48314 = pi18 ? n27500 : n48313;
  assign n48315 = pi17 ? n42647 : n48314;
  assign n48316 = pi16 ? n41183 : n48315;
  assign n48317 = pi20 ? n10503 : n25199;
  assign n48318 = pi22 ? n18256 : n32;
  assign n48319 = pi21 ? n48318 : n32;
  assign n48320 = pi20 ? n48319 : n32;
  assign n48321 = pi19 ? n48317 : n48320;
  assign n48322 = pi18 ? n37 : n48321;
  assign n48323 = pi17 ? n42647 : n48322;
  assign n48324 = pi16 ? n41183 : n48323;
  assign n48325 = pi15 ? n48316 : n48324;
  assign n48326 = pi17 ? n43676 : n47285;
  assign n48327 = pi16 ? n40025 : n48326;
  assign n48328 = pi20 ? n32 : n46699;
  assign n48329 = pi20 ? n40915 : n48184;
  assign n48330 = pi19 ? n48328 : n48329;
  assign n48331 = pi18 ? n32 : n48330;
  assign n48332 = pi17 ? n32 : n48331;
  assign n48333 = pi19 ? n28767 : n1823;
  assign n48334 = pi18 ? n47284 : n48333;
  assign n48335 = pi17 ? n43676 : n48334;
  assign n48336 = pi16 ? n48332 : n48335;
  assign n48337 = pi15 ? n48327 : n48336;
  assign n48338 = pi14 ? n48325 : n48337;
  assign n48339 = pi13 ? n48311 : n48338;
  assign n48340 = pi19 ? n28158 : n30868;
  assign n48341 = pi18 ? n32 : n48340;
  assign n48342 = pi17 ? n32 : n48341;
  assign n48343 = pi20 ? n30868 : n40791;
  assign n48344 = pi19 ? n48343 : n32898;
  assign n48345 = pi18 ? n30868 : n48344;
  assign n48346 = pi21 ? n5015 : n685;
  assign n48347 = pi20 ? n363 : n48346;
  assign n48348 = pi19 ? n7731 : n48347;
  assign n48349 = pi18 ? n48348 : n47831;
  assign n48350 = pi17 ? n48345 : n48349;
  assign n48351 = pi16 ? n48342 : n48350;
  assign n48352 = pi20 ? n30868 : n47327;
  assign n48353 = pi19 ? n30868 : n48352;
  assign n48354 = pi18 ? n30868 : n48353;
  assign n48355 = pi20 ? n157 : n27551;
  assign n48356 = pi19 ? n7845 : n48355;
  assign n48357 = pi18 ? n48356 : n47307;
  assign n48358 = pi17 ? n48354 : n48357;
  assign n48359 = pi16 ? n48258 : n48358;
  assign n48360 = pi15 ? n48351 : n48359;
  assign n48361 = pi19 ? n48328 : n30868;
  assign n48362 = pi18 ? n32 : n48361;
  assign n48363 = pi17 ? n32 : n48362;
  assign n48364 = pi22 ? n158 : n316;
  assign n48365 = pi21 ? n48364 : n316;
  assign n48366 = pi20 ? n99 : n48365;
  assign n48367 = pi19 ? n48366 : n32;
  assign n48368 = pi18 ? n99 : n48367;
  assign n48369 = pi17 ? n48354 : n48368;
  assign n48370 = pi16 ? n48363 : n48369;
  assign n48371 = pi19 ? n45655 : n36798;
  assign n48372 = pi18 ? n32 : n48371;
  assign n48373 = pi17 ? n32 : n48372;
  assign n48374 = pi21 ? n45142 : n33792;
  assign n48375 = pi20 ? n48374 : n33792;
  assign n48376 = pi19 ? n48375 : n33792;
  assign n48377 = pi21 ? n33792 : n139;
  assign n48378 = pi20 ? n33792 : n48377;
  assign n48379 = pi19 ? n33792 : n48378;
  assign n48380 = pi18 ? n48376 : n48379;
  assign n48381 = pi19 ? n139 : n7851;
  assign n48382 = pi21 ? n862 : n157;
  assign n48383 = pi20 ? n48382 : n32082;
  assign n48384 = pi19 ? n48383 : n32;
  assign n48385 = pi18 ? n48381 : n48384;
  assign n48386 = pi17 ? n48380 : n48385;
  assign n48387 = pi16 ? n48373 : n48386;
  assign n48388 = pi15 ? n48370 : n48387;
  assign n48389 = pi14 ? n48360 : n48388;
  assign n48390 = pi21 ? n37899 : n36659;
  assign n48391 = pi20 ? n48390 : n36659;
  assign n48392 = pi19 ? n48391 : n36659;
  assign n48393 = pi21 ? n36659 : n335;
  assign n48394 = pi20 ? n36659 : n48393;
  assign n48395 = pi19 ? n36659 : n48394;
  assign n48396 = pi18 ? n48392 : n48395;
  assign n48397 = pi21 ? n36837 : n316;
  assign n48398 = pi20 ? n47370 : n48397;
  assign n48399 = pi19 ? n335 : n48398;
  assign n48400 = pi20 ? n157 : n47352;
  assign n48401 = pi19 ? n48400 : n32;
  assign n48402 = pi18 ? n48399 : n48401;
  assign n48403 = pi17 ? n48396 : n48402;
  assign n48404 = pi16 ? n48373 : n48403;
  assign n48405 = pi22 ? n47380 : n36659;
  assign n48406 = pi21 ? n32 : n48405;
  assign n48407 = pi20 ? n32 : n48406;
  assign n48408 = pi19 ? n48407 : n36659;
  assign n48409 = pi18 ? n32 : n48408;
  assign n48410 = pi17 ? n32 : n48409;
  assign n48411 = pi18 ? n36659 : n48395;
  assign n48412 = pi17 ? n48411 : n47887;
  assign n48413 = pi16 ? n48410 : n48412;
  assign n48414 = pi15 ? n48404 : n48413;
  assign n48415 = pi21 ? n45653 : n47397;
  assign n48416 = pi20 ? n32 : n48415;
  assign n48417 = pi19 ? n48416 : n43198;
  assign n48418 = pi18 ? n32 : n48417;
  assign n48419 = pi17 ? n32 : n48418;
  assign n48420 = pi21 ? n46280 : n36781;
  assign n48421 = pi20 ? n48420 : n36781;
  assign n48422 = pi19 ? n48421 : n36781;
  assign n48423 = pi21 ? n36781 : n43203;
  assign n48424 = pi20 ? n38923 : n48423;
  assign n48425 = pi19 ? n36781 : n48424;
  assign n48426 = pi18 ? n48422 : n48425;
  assign n48427 = pi22 ? n3944 : n157;
  assign n48428 = pi21 ? n363 : n48427;
  assign n48429 = pi20 ? n48428 : n157;
  assign n48430 = pi19 ? n48429 : n157;
  assign n48431 = pi20 ? n157 : n16339;
  assign n48432 = pi19 ? n48431 : n32;
  assign n48433 = pi18 ? n48430 : n48432;
  assign n48434 = pi17 ? n48426 : n48433;
  assign n48435 = pi16 ? n48419 : n48434;
  assign n48436 = pi21 ? n46276 : n43198;
  assign n48437 = pi20 ? n32 : n48436;
  assign n48438 = pi19 ? n48437 : n43198;
  assign n48439 = pi18 ? n32 : n48438;
  assign n48440 = pi17 ? n32 : n48439;
  assign n48441 = pi21 ? n39972 : n43203;
  assign n48442 = pi20 ? n38923 : n48441;
  assign n48443 = pi19 ? n44208 : n48442;
  assign n48444 = pi18 ? n36781 : n48443;
  assign n48445 = pi20 ? n34831 : n157;
  assign n48446 = pi19 ? n48445 : n157;
  assign n48447 = pi21 ? n10021 : n882;
  assign n48448 = pi20 ? n157 : n48447;
  assign n48449 = pi19 ? n48448 : n32;
  assign n48450 = pi18 ? n48446 : n48449;
  assign n48451 = pi17 ? n48444 : n48450;
  assign n48452 = pi16 ? n48440 : n48451;
  assign n48453 = pi15 ? n48435 : n48452;
  assign n48454 = pi14 ? n48414 : n48453;
  assign n48455 = pi13 ? n48389 : n48454;
  assign n48456 = pi12 ? n48339 : n48455;
  assign n48457 = pi11 ? n48290 : n48456;
  assign n48458 = pi10 ? n48162 : n48457;
  assign n48459 = pi09 ? n47946 : n48458;
  assign n48460 = pi18 ? n41641 : n20563;
  assign n48461 = pi19 ? n31299 : n47923;
  assign n48462 = pi18 ? n34247 : n48461;
  assign n48463 = pi17 ? n48460 : n48462;
  assign n48464 = pi16 ? n32 : n48463;
  assign n48465 = pi15 ? n32 : n48464;
  assign n48466 = pi18 ? n42699 : n20563;
  assign n48467 = pi17 ? n48466 : n47932;
  assign n48468 = pi16 ? n32 : n48467;
  assign n48469 = pi18 ? n46997 : n20563;
  assign n48470 = pi19 ? n33949 : n47936;
  assign n48471 = pi18 ? n20563 : n48470;
  assign n48472 = pi17 ? n48469 : n48471;
  assign n48473 = pi16 ? n32 : n48472;
  assign n48474 = pi15 ? n48468 : n48473;
  assign n48475 = pi14 ? n48465 : n48474;
  assign n48476 = pi13 ? n32 : n48475;
  assign n48477 = pi12 ? n32 : n48476;
  assign n48478 = pi11 ? n32 : n48477;
  assign n48479 = pi10 ? n32 : n48478;
  assign n48480 = pi17 ? n47922 : n47951;
  assign n48481 = pi16 ? n32 : n48480;
  assign n48482 = pi20 ? n3625 : n33398;
  assign n48483 = pi19 ? n37 : n48482;
  assign n48484 = pi18 ? n34258 : n48483;
  assign n48485 = pi17 ? n47954 : n48484;
  assign n48486 = pi16 ? n32 : n48485;
  assign n48487 = pi15 ? n48481 : n48486;
  assign n48488 = pi18 ? n41682 : n20563;
  assign n48489 = pi20 ? n3096 : n3148;
  assign n48490 = pi19 ? n37 : n48489;
  assign n48491 = pi18 ? n33823 : n48490;
  assign n48492 = pi17 ? n48488 : n48491;
  assign n48493 = pi16 ? n32 : n48492;
  assign n48494 = pi20 ? n3086 : n3148;
  assign n48495 = pi19 ? n37 : n48494;
  assign n48496 = pi18 ? n34869 : n48495;
  assign n48497 = pi17 ? n47451 : n48496;
  assign n48498 = pi16 ? n32 : n48497;
  assign n48499 = pi15 ? n48493 : n48498;
  assign n48500 = pi14 ? n48487 : n48499;
  assign n48501 = pi20 ? n40578 : n3023;
  assign n48502 = pi19 ? n37 : n48501;
  assign n48503 = pi18 ? n34869 : n48502;
  assign n48504 = pi17 ? n46302 : n48503;
  assign n48505 = pi16 ? n32 : n48504;
  assign n48506 = pi20 ? n20157 : n33443;
  assign n48507 = pi19 ? n37 : n48506;
  assign n48508 = pi18 ? n32275 : n48507;
  assign n48509 = pi17 ? n46832 : n48508;
  assign n48510 = pi16 ? n32 : n48509;
  assign n48511 = pi15 ? n48505 : n48510;
  assign n48512 = pi20 ? n649 : n17631;
  assign n48513 = pi19 ? n37 : n48512;
  assign n48514 = pi18 ? n33828 : n48513;
  assign n48515 = pi17 ? n47964 : n48514;
  assign n48516 = pi16 ? n32 : n48515;
  assign n48517 = pi21 ? n40091 : n32;
  assign n48518 = pi20 ? n649 : n48517;
  assign n48519 = pi19 ? n37 : n48518;
  assign n48520 = pi18 ? n32288 : n48519;
  assign n48521 = pi17 ? n46866 : n48520;
  assign n48522 = pi16 ? n32 : n48521;
  assign n48523 = pi15 ? n48516 : n48522;
  assign n48524 = pi14 ? n48511 : n48523;
  assign n48525 = pi13 ? n48500 : n48524;
  assign n48526 = pi20 ? n37 : n20890;
  assign n48527 = pi19 ? n37 : n48526;
  assign n48528 = pi18 ? n35812 : n48527;
  assign n48529 = pi17 ? n20563 : n48528;
  assign n48530 = pi16 ? n32 : n48529;
  assign n48531 = pi20 ? n21635 : n3126;
  assign n48532 = pi19 ? n37 : n48531;
  assign n48533 = pi18 ? n32872 : n48532;
  assign n48534 = pi17 ? n20563 : n48533;
  assign n48535 = pi16 ? n46326 : n48534;
  assign n48536 = pi15 ? n48530 : n48535;
  assign n48537 = pi20 ? n577 : n10011;
  assign n48538 = pi19 ? n37 : n48537;
  assign n48539 = pi18 ? n33299 : n48538;
  assign n48540 = pi17 ? n20563 : n48539;
  assign n48541 = pi16 ? n45233 : n48540;
  assign n48542 = pi20 ? n577 : n16621;
  assign n48543 = pi19 ? n37 : n48542;
  assign n48544 = pi18 ? n42358 : n48543;
  assign n48545 = pi17 ? n20563 : n48544;
  assign n48546 = pi16 ? n44635 : n48545;
  assign n48547 = pi15 ? n48541 : n48546;
  assign n48548 = pi14 ? n48536 : n48547;
  assign n48549 = pi20 ? n2094 : n2566;
  assign n48550 = pi19 ? n37 : n48549;
  assign n48551 = pi18 ? n34358 : n48550;
  assign n48552 = pi17 ? n20563 : n48551;
  assign n48553 = pi16 ? n44223 : n48552;
  assign n48554 = pi20 ? n33466 : n2579;
  assign n48555 = pi19 ? n37 : n48554;
  assign n48556 = pi18 ? n32295 : n48555;
  assign n48557 = pi17 ? n20563 : n48556;
  assign n48558 = pi16 ? n45243 : n48557;
  assign n48559 = pi15 ? n48553 : n48558;
  assign n48560 = pi20 ? n2107 : n2579;
  assign n48561 = pi19 ? n37 : n48560;
  assign n48562 = pi18 ? n34358 : n48561;
  assign n48563 = pi17 ? n20563 : n48562;
  assign n48564 = pi16 ? n46349 : n48563;
  assign n48565 = pi20 ? n19934 : n2638;
  assign n48566 = pi19 ? n37 : n48565;
  assign n48567 = pi18 ? n32899 : n48566;
  assign n48568 = pi17 ? n20563 : n48567;
  assign n48569 = pi16 ? n43664 : n48568;
  assign n48570 = pi15 ? n48564 : n48569;
  assign n48571 = pi14 ? n48559 : n48570;
  assign n48572 = pi13 ? n48548 : n48571;
  assign n48573 = pi12 ? n48525 : n48572;
  assign n48574 = pi19 ? n35798 : n37;
  assign n48575 = pi20 ? n19934 : n2653;
  assign n48576 = pi19 ? n37 : n48575;
  assign n48577 = pi18 ? n48574 : n48576;
  assign n48578 = pi17 ? n20563 : n48577;
  assign n48579 = pi16 ? n43664 : n48578;
  assign n48580 = pi18 ? n33916 : n48062;
  assign n48581 = pi17 ? n20563 : n48580;
  assign n48582 = pi16 ? n44671 : n48581;
  assign n48583 = pi15 ? n48579 : n48582;
  assign n48584 = pi18 ? n32315 : n48068;
  assign n48585 = pi17 ? n20563 : n48584;
  assign n48586 = pi16 ? n44671 : n48585;
  assign n48587 = pi18 ? n32315 : n48073;
  assign n48588 = pi17 ? n20563 : n48587;
  assign n48589 = pi16 ? n43675 : n48588;
  assign n48590 = pi15 ? n48586 : n48589;
  assign n48591 = pi14 ? n48583 : n48590;
  assign n48592 = pi18 ? n33924 : n48081;
  assign n48593 = pi17 ? n20563 : n48592;
  assign n48594 = pi16 ? n43685 : n48593;
  assign n48595 = pi16 ? n43685 : n48086;
  assign n48596 = pi15 ? n48594 : n48595;
  assign n48597 = pi18 ? n37649 : n48091;
  assign n48598 = pi17 ? n20563 : n48597;
  assign n48599 = pi16 ? n43219 : n48598;
  assign n48600 = pi18 ? n32369 : n48097;
  assign n48601 = pi17 ? n20563 : n48600;
  assign n48602 = pi16 ? n43219 : n48601;
  assign n48603 = pi15 ? n48599 : n48602;
  assign n48604 = pi14 ? n48596 : n48603;
  assign n48605 = pi13 ? n48591 : n48604;
  assign n48606 = pi20 ? n48089 : n1822;
  assign n48607 = pi19 ? n37 : n48606;
  assign n48608 = pi18 ? n39038 : n48607;
  assign n48609 = pi17 ? n20563 : n48608;
  assign n48610 = pi16 ? n44248 : n48609;
  assign n48611 = pi20 ? n389 : n1822;
  assign n48612 = pi19 ? n37 : n48611;
  assign n48613 = pi18 ? n41334 : n48612;
  assign n48614 = pi17 ? n20563 : n48613;
  assign n48615 = pi16 ? n43224 : n48614;
  assign n48616 = pi15 ? n48610 : n48615;
  assign n48617 = pi19 ? n35317 : n19773;
  assign n48618 = pi20 ? n19208 : n32;
  assign n48619 = pi19 ? n99 : n48618;
  assign n48620 = pi18 ? n48617 : n48619;
  assign n48621 = pi17 ? n20563 : n48620;
  assign n48622 = pi16 ? n43228 : n48621;
  assign n48623 = pi19 ? n32 : n38956;
  assign n48624 = pi18 ? n32 : n48623;
  assign n48625 = pi17 ? n32 : n48624;
  assign n48626 = pi20 ? n33821 : n3039;
  assign n48627 = pi19 ? n48626 : n99;
  assign n48628 = pi18 ? n48627 : n48619;
  assign n48629 = pi17 ? n20563 : n48628;
  assign n48630 = pi16 ? n48625 : n48629;
  assign n48631 = pi15 ? n48622 : n48630;
  assign n48632 = pi14 ? n48616 : n48631;
  assign n48633 = pi16 ? n48625 : n48133;
  assign n48634 = pi20 ? n41913 : n99;
  assign n48635 = pi19 ? n48634 : n99;
  assign n48636 = pi19 ? n6542 : n19182;
  assign n48637 = pi18 ? n48635 : n48636;
  assign n48638 = pi17 ? n48135 : n48637;
  assign n48639 = pi16 ? n48625 : n48638;
  assign n48640 = pi15 ? n48633 : n48639;
  assign n48641 = pi20 ? n33964 : n5077;
  assign n48642 = pi19 ? n48641 : n32889;
  assign n48643 = pi21 ? n1027 : n5178;
  assign n48644 = pi20 ? n48643 : n32;
  assign n48645 = pi19 ? n48147 : n48644;
  assign n48646 = pi18 ? n48642 : n48645;
  assign n48647 = pi17 ? n20563 : n48646;
  assign n48648 = pi16 ? n42646 : n48647;
  assign n48649 = pi19 ? n31299 : n33288;
  assign n48650 = pi18 ? n48649 : n48645;
  assign n48651 = pi17 ? n45246 : n48650;
  assign n48652 = pi16 ? n42656 : n48651;
  assign n48653 = pi15 ? n48648 : n48652;
  assign n48654 = pi14 ? n48640 : n48653;
  assign n48655 = pi13 ? n48632 : n48654;
  assign n48656 = pi12 ? n48605 : n48655;
  assign n48657 = pi11 ? n48573 : n48656;
  assign n48658 = pi18 ? n20563 : n34247;
  assign n48659 = pi19 ? n46822 : n99;
  assign n48660 = pi21 ? n1027 : n26303;
  assign n48661 = pi20 ? n48660 : n32;
  assign n48662 = pi19 ? n48166 : n48661;
  assign n48663 = pi18 ? n48659 : n48662;
  assign n48664 = pi17 ? n48658 : n48663;
  assign n48665 = pi16 ? n42202 : n48664;
  assign n48666 = pi20 ? n9173 : n32;
  assign n48667 = pi19 ? n32636 : n48666;
  assign n48668 = pi18 ? n48178 : n48667;
  assign n48669 = pi17 ? n48177 : n48668;
  assign n48670 = pi16 ? n42202 : n48669;
  assign n48671 = pi15 ? n48665 : n48670;
  assign n48672 = pi21 ? n39164 : n37;
  assign n48673 = pi20 ? n48672 : n37;
  assign n48674 = pi19 ? n48673 : n28582;
  assign n48675 = pi19 ? n1017 : n48666;
  assign n48676 = pi18 ? n48674 : n48675;
  assign n48677 = pi17 ? n48187 : n48676;
  assign n48678 = pi16 ? n42202 : n48677;
  assign n48679 = pi18 ? n20563 : n40191;
  assign n48680 = pi19 ? n32663 : n20532;
  assign n48681 = pi18 ? n32934 : n48680;
  assign n48682 = pi17 ? n48679 : n48681;
  assign n48683 = pi16 ? n43263 : n48682;
  assign n48684 = pi15 ? n48678 : n48683;
  assign n48685 = pi14 ? n48671 : n48684;
  assign n48686 = pi18 ? n20563 : n34865;
  assign n48687 = pi19 ? n12589 : n19276;
  assign n48688 = pi18 ? n32934 : n48687;
  assign n48689 = pi17 ? n48686 : n48688;
  assign n48690 = pi16 ? n43263 : n48689;
  assign n48691 = pi20 ? n32151 : n32;
  assign n48692 = pi19 ? n12589 : n48691;
  assign n48693 = pi18 ? n48202 : n48692;
  assign n48694 = pi17 ? n48197 : n48693;
  assign n48695 = pi16 ? n47594 : n48694;
  assign n48696 = pi15 ? n48690 : n48695;
  assign n48697 = pi18 ? n48207 : n47118;
  assign n48698 = pi17 ? n48197 : n48697;
  assign n48699 = pi16 ? n47594 : n48698;
  assign n48700 = pi21 ? n28649 : n928;
  assign n48701 = pi20 ? n48700 : n32;
  assign n48702 = pi19 ? n47140 : n48701;
  assign n48703 = pi18 ? n9815 : n48702;
  assign n48704 = pi17 ? n48197 : n48703;
  assign n48705 = pi16 ? n47594 : n48704;
  assign n48706 = pi15 ? n48699 : n48705;
  assign n48707 = pi14 ? n48696 : n48706;
  assign n48708 = pi13 ? n48685 : n48707;
  assign n48709 = pi21 ? n31294 : n48221;
  assign n48710 = pi20 ? n20563 : n48709;
  assign n48711 = pi19 ? n20563 : n48710;
  assign n48712 = pi18 ? n20563 : n48711;
  assign n48713 = pi19 ? n47153 : n21212;
  assign n48714 = pi18 ? n9796 : n48713;
  assign n48715 = pi17 ? n48712 : n48714;
  assign n48716 = pi16 ? n47594 : n48715;
  assign n48717 = pi17 ? n48658 : n48233;
  assign n48718 = pi16 ? n47594 : n48717;
  assign n48719 = pi15 ? n48716 : n48718;
  assign n48720 = pi19 ? n20563 : n47514;
  assign n48721 = pi18 ? n20563 : n48720;
  assign n48722 = pi19 ? n48237 : n20208;
  assign n48723 = pi18 ? n7686 : n48722;
  assign n48724 = pi17 ? n48721 : n48723;
  assign n48725 = pi16 ? n47594 : n48724;
  assign n48726 = pi17 ? n48721 : n48244;
  assign n48727 = pi16 ? n42701 : n48726;
  assign n48728 = pi15 ? n48725 : n48727;
  assign n48729 = pi14 ? n48719 : n48728;
  assign n48730 = pi21 ? n19438 : n1009;
  assign n48731 = pi20 ? n48730 : n32;
  assign n48732 = pi19 ? n48249 : n48731;
  assign n48733 = pi18 ? n37 : n48732;
  assign n48734 = pi17 ? n48721 : n48733;
  assign n48735 = pi16 ? n42701 : n48734;
  assign n48736 = pi21 ? n32 : n37805;
  assign n48737 = pi20 ? n32 : n48736;
  assign n48738 = pi19 ? n48737 : n30868;
  assign n48739 = pi18 ? n32 : n48738;
  assign n48740 = pi17 ? n32 : n48739;
  assign n48741 = pi19 ? n30868 : n31914;
  assign n48742 = pi18 ? n30868 : n48741;
  assign n48743 = pi17 ? n48742 : n48262;
  assign n48744 = pi16 ? n48740 : n48743;
  assign n48745 = pi15 ? n48735 : n48744;
  assign n48746 = pi18 ? n20563 : n39626;
  assign n48747 = pi19 ? n13337 : n47187;
  assign n48748 = pi18 ? n37 : n48747;
  assign n48749 = pi17 ? n48746 : n48748;
  assign n48750 = pi16 ? n48740 : n48749;
  assign n48751 = pi21 ? n32 : n37252;
  assign n48752 = pi20 ? n32 : n48751;
  assign n48753 = pi19 ? n48752 : n48279;
  assign n48754 = pi18 ? n32 : n48753;
  assign n48755 = pi17 ? n32 : n48754;
  assign n48756 = pi19 ? n47228 : n47187;
  assign n48757 = pi18 ? n7677 : n48756;
  assign n48758 = pi17 ? n48746 : n48757;
  assign n48759 = pi16 ? n48755 : n48758;
  assign n48760 = pi15 ? n48750 : n48759;
  assign n48761 = pi14 ? n48745 : n48760;
  assign n48762 = pi13 ? n48729 : n48761;
  assign n48763 = pi12 ? n48708 : n48762;
  assign n48764 = pi19 ? n47238 : n9964;
  assign n48765 = pi18 ? n37 : n48764;
  assign n48766 = pi17 ? n48746 : n48765;
  assign n48767 = pi16 ? n40487 : n48766;
  assign n48768 = pi18 ? n20563 : n40067;
  assign n48769 = pi17 ? n48768 : n48297;
  assign n48770 = pi16 ? n40487 : n48769;
  assign n48771 = pi15 ? n48767 : n48770;
  assign n48772 = pi17 ? n48768 : n48302;
  assign n48773 = pi16 ? n40487 : n48772;
  assign n48774 = pi17 ? n48768 : n48307;
  assign n48775 = pi16 ? n40487 : n48774;
  assign n48776 = pi15 ? n48773 : n48775;
  assign n48777 = pi14 ? n48771 : n48776;
  assign n48778 = pi19 ? n48312 : n7050;
  assign n48779 = pi18 ? n27500 : n48778;
  assign n48780 = pi17 ? n48768 : n48779;
  assign n48781 = pi16 ? n46999 : n48780;
  assign n48782 = pi18 ? n20563 : n43367;
  assign n48783 = pi19 ? n48317 : n5831;
  assign n48784 = pi18 ? n37 : n48783;
  assign n48785 = pi17 ? n48782 : n48784;
  assign n48786 = pi16 ? n46999 : n48785;
  assign n48787 = pi15 ? n48781 : n48786;
  assign n48788 = pi17 ? n45775 : n47285;
  assign n48789 = pi16 ? n42689 : n48788;
  assign n48790 = pi20 ? n32 : n47192;
  assign n48791 = pi19 ? n48790 : n48329;
  assign n48792 = pi18 ? n32 : n48791;
  assign n48793 = pi17 ? n32 : n48792;
  assign n48794 = pi16 ? n48793 : n48788;
  assign n48795 = pi15 ? n48789 : n48794;
  assign n48796 = pi14 ? n48787 : n48795;
  assign n48797 = pi13 ? n48777 : n48796;
  assign n48798 = pi19 ? n36868 : n30868;
  assign n48799 = pi18 ? n32 : n48798;
  assign n48800 = pi17 ? n32 : n48799;
  assign n48801 = pi19 ? n48343 : n35776;
  assign n48802 = pi18 ? n30868 : n48801;
  assign n48803 = pi17 ? n48802 : n48349;
  assign n48804 = pi16 ? n48800 : n48803;
  assign n48805 = pi19 ? n46168 : n30868;
  assign n48806 = pi18 ? n32 : n48805;
  assign n48807 = pi17 ? n32 : n48806;
  assign n48808 = pi21 ? n41564 : n99;
  assign n48809 = pi20 ? n30868 : n48808;
  assign n48810 = pi19 ? n30868 : n48809;
  assign n48811 = pi18 ? n30868 : n48810;
  assign n48812 = pi17 ? n48811 : n48357;
  assign n48813 = pi16 ? n48807 : n48812;
  assign n48814 = pi15 ? n48804 : n48813;
  assign n48815 = pi19 ? n46189 : n30868;
  assign n48816 = pi18 ? n32 : n48815;
  assign n48817 = pi17 ? n32 : n48816;
  assign n48818 = pi19 ? n30868 : n38848;
  assign n48819 = pi18 ? n30868 : n48818;
  assign n48820 = pi17 ? n48819 : n48368;
  assign n48821 = pi16 ? n48817 : n48820;
  assign n48822 = pi21 ? n32 : n46727;
  assign n48823 = pi20 ? n32 : n48822;
  assign n48824 = pi19 ? n48823 : n36798;
  assign n48825 = pi18 ? n32 : n48824;
  assign n48826 = pi17 ? n32 : n48825;
  assign n48827 = pi21 ? n33792 : n40429;
  assign n48828 = pi20 ? n33792 : n48827;
  assign n48829 = pi19 ? n33792 : n48828;
  assign n48830 = pi18 ? n48376 : n48829;
  assign n48831 = pi17 ? n48830 : n48385;
  assign n48832 = pi16 ? n48826 : n48831;
  assign n48833 = pi15 ? n48821 : n48832;
  assign n48834 = pi14 ? n48814 : n48833;
  assign n48835 = pi22 ? n38926 : n335;
  assign n48836 = pi21 ? n36659 : n48835;
  assign n48837 = pi20 ? n36659 : n48836;
  assign n48838 = pi19 ? n36659 : n48837;
  assign n48839 = pi18 ? n48392 : n48838;
  assign n48840 = pi21 ? n7429 : n397;
  assign n48841 = pi20 ? n157 : n48840;
  assign n48842 = pi19 ? n48841 : n32;
  assign n48843 = pi18 ? n48399 : n48842;
  assign n48844 = pi17 ? n48839 : n48843;
  assign n48845 = pi16 ? n48826 : n48844;
  assign n48846 = pi21 ? n32 : n46758;
  assign n48847 = pi20 ? n32 : n48846;
  assign n48848 = pi19 ? n48847 : n36659;
  assign n48849 = pi18 ? n32 : n48848;
  assign n48850 = pi17 ? n32 : n48849;
  assign n48851 = pi18 ? n36659 : n48838;
  assign n48852 = pi18 ? n47391 : n32601;
  assign n48853 = pi17 ? n48851 : n48852;
  assign n48854 = pi16 ? n48850 : n48853;
  assign n48855 = pi15 ? n48845 : n48854;
  assign n48856 = pi22 ? n32 : n43198;
  assign n48857 = pi21 ? n32 : n48856;
  assign n48858 = pi20 ? n32 : n48857;
  assign n48859 = pi19 ? n48858 : n43198;
  assign n48860 = pi18 ? n32 : n48859;
  assign n48861 = pi17 ? n32 : n48860;
  assign n48862 = pi21 ? n36781 : n46797;
  assign n48863 = pi20 ? n38923 : n48862;
  assign n48864 = pi19 ? n36781 : n48863;
  assign n48865 = pi18 ? n48422 : n48864;
  assign n48866 = pi20 ? n36813 : n157;
  assign n48867 = pi19 ? n48866 : n157;
  assign n48868 = pi18 ? n48867 : n48432;
  assign n48869 = pi17 ? n48865 : n48868;
  assign n48870 = pi16 ? n48861 : n48869;
  assign n48871 = pi19 ? n46202 : n43198;
  assign n48872 = pi18 ? n32 : n48871;
  assign n48873 = pi17 ? n32 : n48872;
  assign n48874 = pi21 ? n39972 : n46797;
  assign n48875 = pi20 ? n38923 : n48874;
  assign n48876 = pi19 ? n44208 : n48875;
  assign n48877 = pi18 ? n36781 : n48876;
  assign n48878 = pi22 ? n46796 : n157;
  assign n48879 = pi21 ? n48878 : n157;
  assign n48880 = pi20 ? n48879 : n157;
  assign n48881 = pi19 ? n48880 : n157;
  assign n48882 = pi21 ? n10021 : n2320;
  assign n48883 = pi20 ? n157 : n48882;
  assign n48884 = pi19 ? n48883 : n32;
  assign n48885 = pi18 ? n48881 : n48884;
  assign n48886 = pi17 ? n48877 : n48885;
  assign n48887 = pi16 ? n48873 : n48886;
  assign n48888 = pi15 ? n48870 : n48887;
  assign n48889 = pi14 ? n48855 : n48888;
  assign n48890 = pi13 ? n48834 : n48889;
  assign n48891 = pi12 ? n48797 : n48890;
  assign n48892 = pi11 ? n48763 : n48891;
  assign n48893 = pi10 ? n48657 : n48892;
  assign n48894 = pi09 ? n48479 : n48893;
  assign n48895 = pi08 ? n48459 : n48894;
  assign n48896 = pi07 ? n47921 : n48895;
  assign n48897 = pi18 ? n43261 : n20563;
  assign n48898 = pi20 ? n37 : n17948;
  assign n48899 = pi19 ? n37 : n48898;
  assign n48900 = pi18 ? n20563 : n48899;
  assign n48901 = pi17 ? n48897 : n48900;
  assign n48902 = pi16 ? n32 : n48901;
  assign n48903 = pi15 ? n32 : n48902;
  assign n48904 = pi18 ? n48120 : n20563;
  assign n48905 = pi21 ? n37 : n20563;
  assign n48906 = pi20 ? n48905 : n37;
  assign n48907 = pi20 ? n37 : n18573;
  assign n48908 = pi19 ? n48906 : n48907;
  assign n48909 = pi18 ? n20563 : n48908;
  assign n48910 = pi17 ? n48904 : n48909;
  assign n48911 = pi16 ? n32 : n48910;
  assign n48912 = pi18 ? n47592 : n20563;
  assign n48913 = pi17 ? n48912 : n48909;
  assign n48914 = pi16 ? n32 : n48913;
  assign n48915 = pi15 ? n48911 : n48914;
  assign n48916 = pi14 ? n48903 : n48915;
  assign n48917 = pi13 ? n32 : n48916;
  assign n48918 = pi12 ? n32 : n48917;
  assign n48919 = pi11 ? n32 : n48918;
  assign n48920 = pi10 ? n32 : n48919;
  assign n48921 = pi20 ? n37 : n32342;
  assign n48922 = pi19 ? n37 : n48921;
  assign n48923 = pi18 ? n20563 : n48922;
  assign n48924 = pi17 ? n48460 : n48923;
  assign n48925 = pi16 ? n32 : n48924;
  assign n48926 = pi20 ? n3096 : n33325;
  assign n48927 = pi19 ? n37 : n48926;
  assign n48928 = pi18 ? n20563 : n48927;
  assign n48929 = pi17 ? n47922 : n48928;
  assign n48930 = pi16 ? n32 : n48929;
  assign n48931 = pi15 ? n48925 : n48930;
  assign n48932 = pi20 ? n3096 : n18017;
  assign n48933 = pi19 ? n31280 : n48932;
  assign n48934 = pi18 ? n20563 : n48933;
  assign n48935 = pi17 ? n47929 : n48934;
  assign n48936 = pi16 ? n32 : n48935;
  assign n48937 = pi20 ? n3086 : n3849;
  assign n48938 = pi19 ? n31280 : n48937;
  assign n48939 = pi18 ? n20563 : n48938;
  assign n48940 = pi17 ? n47935 : n48939;
  assign n48941 = pi16 ? n32 : n48940;
  assign n48942 = pi15 ? n48936 : n48941;
  assign n48943 = pi14 ? n48931 : n48942;
  assign n48944 = pi20 ? n997 : n3157;
  assign n48945 = pi19 ? n30097 : n48944;
  assign n48946 = pi18 ? n20563 : n48945;
  assign n48947 = pi17 ? n47947 : n48946;
  assign n48948 = pi16 ? n32 : n48947;
  assign n48949 = pi18 ? n46446 : n20563;
  assign n48950 = pi20 ? n37 : n17619;
  assign n48951 = pi19 ? n37 : n48950;
  assign n48952 = pi18 ? n34869 : n48951;
  assign n48953 = pi17 ? n48949 : n48952;
  assign n48954 = pi16 ? n32 : n48953;
  assign n48955 = pi15 ? n48948 : n48954;
  assign n48956 = pi20 ? n37 : n17631;
  assign n48957 = pi19 ? n32933 : n48956;
  assign n48958 = pi18 ? n20563 : n48957;
  assign n48959 = pi17 ? n48488 : n48958;
  assign n48960 = pi16 ? n32 : n48959;
  assign n48961 = pi18 ? n34258 : n48519;
  assign n48962 = pi17 ? n47964 : n48961;
  assign n48963 = pi16 ? n32 : n48962;
  assign n48964 = pi15 ? n48960 : n48963;
  assign n48965 = pi14 ? n48955 : n48964;
  assign n48966 = pi13 ? n48943 : n48965;
  assign n48967 = pi20 ? n649 : n20890;
  assign n48968 = pi19 ? n30097 : n48967;
  assign n48969 = pi18 ? n20563 : n48968;
  assign n48970 = pi17 ? n45707 : n48969;
  assign n48971 = pi16 ? n32 : n48970;
  assign n48972 = pi19 ? n20563 : n37309;
  assign n48973 = pi20 ? n649 : n3126;
  assign n48974 = pi19 ? n37 : n48973;
  assign n48975 = pi18 ? n48972 : n48974;
  assign n48976 = pi17 ? n46859 : n48975;
  assign n48977 = pi16 ? n32 : n48976;
  assign n48978 = pi15 ? n48971 : n48977;
  assign n48979 = pi20 ? n20157 : n23980;
  assign n48980 = pi19 ? n37 : n48979;
  assign n48981 = pi18 ? n34295 : n48980;
  assign n48982 = pi17 ? n45715 : n48981;
  assign n48983 = pi16 ? n32 : n48982;
  assign n48984 = pi20 ? n569 : n16621;
  assign n48985 = pi19 ? n37 : n48984;
  assign n48986 = pi18 ? n33245 : n48985;
  assign n48987 = pi17 ? n46866 : n48986;
  assign n48988 = pi16 ? n32 : n48987;
  assign n48989 = pi15 ? n48983 : n48988;
  assign n48990 = pi14 ? n48978 : n48989;
  assign n48991 = pi20 ? n31220 : n30096;
  assign n48992 = pi19 ? n20563 : n48991;
  assign n48993 = pi20 ? n3393 : n2566;
  assign n48994 = pi19 ? n37 : n48993;
  assign n48995 = pi18 ? n48992 : n48994;
  assign n48996 = pi17 ? n20563 : n48995;
  assign n48997 = pi16 ? n44635 : n48996;
  assign n48998 = pi20 ? n6402 : n2579;
  assign n48999 = pi19 ? n37 : n48998;
  assign n49000 = pi18 ? n38523 : n48999;
  assign n49001 = pi17 ? n20563 : n49000;
  assign n49002 = pi16 ? n45740 : n49001;
  assign n49003 = pi15 ? n48997 : n49002;
  assign n49004 = pi20 ? n6402 : n4116;
  assign n49005 = pi19 ? n37 : n49004;
  assign n49006 = pi18 ? n38523 : n49005;
  assign n49007 = pi17 ? n20563 : n49006;
  assign n49008 = pi16 ? n46885 : n49007;
  assign n49009 = pi18 ? n32275 : n49005;
  assign n49010 = pi17 ? n20563 : n49009;
  assign n49011 = pi16 ? n44653 : n49010;
  assign n49012 = pi15 ? n49008 : n49011;
  assign n49013 = pi14 ? n49003 : n49012;
  assign n49014 = pi13 ? n48990 : n49013;
  assign n49015 = pi12 ? n48966 : n49014;
  assign n49016 = pi20 ? n29133 : n37;
  assign n49017 = pi19 ? n20563 : n49016;
  assign n49018 = pi20 ? n3393 : n5830;
  assign n49019 = pi19 ? n37 : n49018;
  assign n49020 = pi18 ? n49017 : n49019;
  assign n49021 = pi17 ? n20563 : n49020;
  assign n49022 = pi16 ? n44223 : n49021;
  assign n49023 = pi20 ? n363 : n2638;
  assign n49024 = pi19 ? n37 : n49023;
  assign n49025 = pi18 ? n33299 : n49024;
  assign n49026 = pi17 ? n20563 : n49025;
  assign n49027 = pi16 ? n44223 : n49026;
  assign n49028 = pi15 ? n49022 : n49027;
  assign n49029 = pi20 ? n7730 : n2653;
  assign n49030 = pi19 ? n37 : n49029;
  assign n49031 = pi18 ? n33285 : n49030;
  assign n49032 = pi17 ? n20563 : n49031;
  assign n49033 = pi16 ? n44223 : n49032;
  assign n49034 = pi21 ? n5012 : n14255;
  assign n49035 = pi20 ? n49034 : n2653;
  assign n49036 = pi19 ? n37 : n49035;
  assign n49037 = pi18 ? n33285 : n49036;
  assign n49038 = pi17 ? n20563 : n49037;
  assign n49039 = pi16 ? n45243 : n49038;
  assign n49040 = pi15 ? n49033 : n49039;
  assign n49041 = pi14 ? n49028 : n49040;
  assign n49042 = pi21 ? n5012 : n2106;
  assign n49043 = pi20 ? n49042 : n2701;
  assign n49044 = pi19 ? n37 : n49043;
  assign n49045 = pi18 ? n33285 : n49044;
  assign n49046 = pi17 ? n20563 : n49045;
  assign n49047 = pi16 ? n44227 : n49046;
  assign n49048 = pi20 ? n48089 : n2679;
  assign n49049 = pi19 ? n37 : n49048;
  assign n49050 = pi18 ? n32295 : n49049;
  assign n49051 = pi17 ? n20563 : n49050;
  assign n49052 = pi16 ? n44227 : n49051;
  assign n49053 = pi15 ? n49047 : n49052;
  assign n49054 = pi18 ? n32295 : n48607;
  assign n49055 = pi17 ? n20563 : n49054;
  assign n49056 = pi16 ? n43664 : n49055;
  assign n49057 = pi21 ? n37 : n6132;
  assign n49058 = pi20 ? n49057 : n2701;
  assign n49059 = pi19 ? n37 : n49058;
  assign n49060 = pi18 ? n33299 : n49059;
  assign n49061 = pi17 ? n20563 : n49060;
  assign n49062 = pi16 ? n43664 : n49061;
  assign n49063 = pi15 ? n49056 : n49062;
  assign n49064 = pi14 ? n49053 : n49063;
  assign n49065 = pi13 ? n49041 : n49064;
  assign n49066 = pi21 ? n37 : n4015;
  assign n49067 = pi20 ? n49066 : n1822;
  assign n49068 = pi19 ? n37 : n49067;
  assign n49069 = pi18 ? n33299 : n49068;
  assign n49070 = pi17 ? n20563 : n49069;
  assign n49071 = pi16 ? n44671 : n49070;
  assign n49072 = pi19 ? n20563 : n35209;
  assign n49073 = pi20 ? n19208 : n1822;
  assign n49074 = pi19 ? n99 : n49073;
  assign n49075 = pi18 ? n49072 : n49074;
  assign n49076 = pi17 ? n20563 : n49075;
  assign n49077 = pi16 ? n43675 : n49076;
  assign n49078 = pi15 ? n49071 : n49077;
  assign n49079 = pi19 ? n37309 : n17013;
  assign n49080 = pi19 ? n3050 : n20979;
  assign n49081 = pi18 ? n49079 : n49080;
  assign n49082 = pi17 ? n20563 : n49081;
  assign n49083 = pi16 ? n43675 : n49082;
  assign n49084 = pi19 ? n37309 : n34261;
  assign n49085 = pi19 ? n99 : n19172;
  assign n49086 = pi18 ? n49084 : n49085;
  assign n49087 = pi17 ? n20563 : n49086;
  assign n49088 = pi16 ? n44688 : n49087;
  assign n49089 = pi15 ? n49083 : n49088;
  assign n49090 = pi14 ? n49078 : n49089;
  assign n49091 = pi19 ? n38333 : n26407;
  assign n49092 = pi21 ? n775 : n5145;
  assign n49093 = pi20 ? n49092 : n32;
  assign n49094 = pi19 ? n2242 : n49093;
  assign n49095 = pi18 ? n49091 : n49094;
  assign n49096 = pi17 ? n20563 : n49095;
  assign n49097 = pi16 ? n44688 : n49096;
  assign n49098 = pi20 ? n20563 : n42418;
  assign n49099 = pi19 ? n49098 : n26407;
  assign n49100 = pi21 ? n7815 : n5178;
  assign n49101 = pi20 ? n49100 : n32;
  assign n49102 = pi19 ? n1666 : n49101;
  assign n49103 = pi18 ? n49099 : n49102;
  assign n49104 = pi17 ? n20563 : n49103;
  assign n49105 = pi16 ? n44688 : n49104;
  assign n49106 = pi15 ? n49097 : n49105;
  assign n49107 = pi19 ? n31221 : n17013;
  assign n49108 = pi20 ? n99 : n42885;
  assign n49109 = pi19 ? n49108 : n22006;
  assign n49110 = pi18 ? n49107 : n49109;
  assign n49111 = pi17 ? n20563 : n49110;
  assign n49112 = pi16 ? n43219 : n49111;
  assign n49113 = pi21 ? n99 : n15439;
  assign n49114 = pi20 ? n49113 : n32;
  assign n49115 = pi19 ? n26407 : n49114;
  assign n49116 = pi18 ? n32899 : n49115;
  assign n49117 = pi17 ? n20563 : n49116;
  assign n49118 = pi16 ? n44248 : n49117;
  assign n49119 = pi15 ? n49112 : n49118;
  assign n49120 = pi14 ? n49106 : n49119;
  assign n49121 = pi13 ? n49090 : n49120;
  assign n49122 = pi12 ? n49065 : n49121;
  assign n49123 = pi11 ? n49015 : n49122;
  assign n49124 = pi20 ? n37 : n14524;
  assign n49125 = pi19 ? n32348 : n49124;
  assign n49126 = pi20 ? n22666 : n1912;
  assign n49127 = pi21 ? n204 : n14168;
  assign n49128 = pi20 ? n49127 : n32;
  assign n49129 = pi19 ? n49126 : n49128;
  assign n49130 = pi18 ? n49125 : n49129;
  assign n49131 = pi17 ? n20563 : n49130;
  assign n49132 = pi16 ? n43249 : n49131;
  assign n49133 = pi19 ? n38333 : n37;
  assign n49134 = pi21 ? n204 : n2230;
  assign n49135 = pi20 ? n49134 : n32;
  assign n49136 = pi19 ? n20743 : n49135;
  assign n49137 = pi18 ? n49133 : n49136;
  assign n49138 = pi17 ? n20563 : n49137;
  assign n49139 = pi16 ? n43249 : n49138;
  assign n49140 = pi15 ? n49132 : n49139;
  assign n49141 = pi20 ? n40791 : n42418;
  assign n49142 = pi19 ? n49141 : n37;
  assign n49143 = pi18 ? n49142 : n49136;
  assign n49144 = pi17 ? n20563 : n49143;
  assign n49145 = pi16 ? n43249 : n49144;
  assign n49146 = pi20 ? n942 : n3096;
  assign n49147 = pi19 ? n49146 : n19276;
  assign n49148 = pi18 ? n32899 : n49147;
  assign n49149 = pi17 ? n20563 : n49148;
  assign n49150 = pi16 ? n44275 : n49149;
  assign n49151 = pi15 ? n49145 : n49150;
  assign n49152 = pi14 ? n49140 : n49151;
  assign n49153 = pi20 ? n8742 : n139;
  assign n49154 = pi19 ? n49153 : n19276;
  assign n49155 = pi18 ? n35300 : n49154;
  assign n49156 = pi17 ? n20563 : n49155;
  assign n49157 = pi16 ? n48625 : n49156;
  assign n49158 = pi19 ? n14962 : n46508;
  assign n49159 = pi18 ? n32377 : n49158;
  assign n49160 = pi17 ? n20563 : n49159;
  assign n49161 = pi16 ? n42195 : n49160;
  assign n49162 = pi15 ? n49157 : n49161;
  assign n49163 = pi21 ? n28649 : n3339;
  assign n49164 = pi20 ? n49163 : n32;
  assign n49165 = pi19 ? n8765 : n49164;
  assign n49166 = pi18 ? n32349 : n49165;
  assign n49167 = pi17 ? n20563 : n49166;
  assign n49168 = pi16 ? n42195 : n49167;
  assign n49169 = pi21 ? n28649 : n2637;
  assign n49170 = pi20 ? n49169 : n32;
  assign n49171 = pi19 ? n8765 : n49170;
  assign n49172 = pi18 ? n32349 : n49171;
  assign n49173 = pi17 ? n20563 : n49172;
  assign n49174 = pi16 ? n42195 : n49173;
  assign n49175 = pi15 ? n49168 : n49174;
  assign n49176 = pi14 ? n49162 : n49175;
  assign n49177 = pi13 ? n49152 : n49176;
  assign n49178 = pi21 ? n48221 : n37;
  assign n49179 = pi20 ? n20563 : n49178;
  assign n49180 = pi19 ? n49179 : n37;
  assign n49181 = pi19 ? n24788 : n39518;
  assign n49182 = pi18 ? n49180 : n49181;
  assign n49183 = pi17 ? n20563 : n49182;
  assign n49184 = pi16 ? n42195 : n49183;
  assign n49185 = pi20 ? n24379 : n32;
  assign n49186 = pi19 ? n7685 : n49185;
  assign n49187 = pi18 ? n32349 : n49186;
  assign n49188 = pi17 ? n20563 : n49187;
  assign n49189 = pi16 ? n42195 : n49188;
  assign n49190 = pi15 ? n49184 : n49189;
  assign n49191 = pi20 ? n37 : n31770;
  assign n49192 = pi21 ? n12635 : n928;
  assign n49193 = pi20 ? n49192 : n32;
  assign n49194 = pi19 ? n49191 : n49193;
  assign n49195 = pi18 ? n31939 : n49194;
  assign n49196 = pi17 ? n20563 : n49195;
  assign n49197 = pi16 ? n42202 : n49196;
  assign n49198 = pi21 ? n37 : n4902;
  assign n49199 = pi20 ? n37 : n49198;
  assign n49200 = pi19 ? n49199 : n20238;
  assign n49201 = pi18 ? n32377 : n49200;
  assign n49202 = pi17 ? n20563 : n49201;
  assign n49203 = pi16 ? n42202 : n49202;
  assign n49204 = pi15 ? n49197 : n49203;
  assign n49205 = pi14 ? n49190 : n49204;
  assign n49206 = pi22 ? n30865 : n39190;
  assign n49207 = pi21 ? n49206 : n30868;
  assign n49208 = pi20 ? n49207 : n30868;
  assign n49209 = pi19 ? n32 : n49208;
  assign n49210 = pi18 ? n32 : n49209;
  assign n49211 = pi17 ? n32 : n49210;
  assign n49212 = pi18 ? n30868 : n42015;
  assign n49213 = pi20 ? n31104 : n32;
  assign n49214 = pi19 ? n7685 : n49213;
  assign n49215 = pi18 ? n32377 : n49214;
  assign n49216 = pi17 ? n49212 : n49215;
  assign n49217 = pi16 ? n49211 : n49216;
  assign n49218 = pi20 ? n37806 : n30868;
  assign n49219 = pi19 ? n32 : n49218;
  assign n49220 = pi18 ? n32 : n49219;
  assign n49221 = pi17 ? n32 : n49220;
  assign n49222 = pi20 ? n37 : n31760;
  assign n49223 = pi19 ? n49222 : n47180;
  assign n49224 = pi18 ? n31939 : n49223;
  assign n49225 = pi17 ? n49212 : n49224;
  assign n49226 = pi16 ? n49221 : n49225;
  assign n49227 = pi15 ? n49217 : n49226;
  assign n49228 = pi22 ? n37804 : n42109;
  assign n49229 = pi21 ? n49228 : n33792;
  assign n49230 = pi20 ? n49229 : n40958;
  assign n49231 = pi19 ? n32 : n49230;
  assign n49232 = pi18 ? n32 : n49231;
  assign n49233 = pi17 ? n32 : n49232;
  assign n49234 = pi20 ? n40958 : n20563;
  assign n49235 = pi19 ? n49234 : n20563;
  assign n49236 = pi18 ? n49235 : n20563;
  assign n49237 = pi19 ? n8928 : n9432;
  assign n49238 = pi18 ? n31939 : n49237;
  assign n49239 = pi17 ? n49236 : n49238;
  assign n49240 = pi16 ? n49233 : n49239;
  assign n49241 = pi21 ? n40917 : n20563;
  assign n49242 = pi20 ? n37806 : n49241;
  assign n49243 = pi19 ? n32 : n49242;
  assign n49244 = pi18 ? n32 : n49243;
  assign n49245 = pi17 ? n32 : n49244;
  assign n49246 = pi21 ? n48173 : n20563;
  assign n49247 = pi20 ? n49246 : n20563;
  assign n49248 = pi19 ? n49247 : n20563;
  assign n49249 = pi18 ? n49248 : n20563;
  assign n49250 = pi19 ? n2095 : n16945;
  assign n49251 = pi18 ? n31939 : n49250;
  assign n49252 = pi17 ? n49249 : n49251;
  assign n49253 = pi16 ? n49245 : n49252;
  assign n49254 = pi15 ? n49240 : n49253;
  assign n49255 = pi14 ? n49227 : n49254;
  assign n49256 = pi13 ? n49205 : n49255;
  assign n49257 = pi12 ? n49177 : n49256;
  assign n49258 = pi19 ? n2108 : n9457;
  assign n49259 = pi18 ? n32377 : n49258;
  assign n49260 = pi17 ? n20563 : n49259;
  assign n49261 = pi16 ? n41632 : n49260;
  assign n49262 = pi21 ? n37 : n28506;
  assign n49263 = pi20 ? n37 : n49262;
  assign n49264 = pi19 ? n49263 : n9964;
  assign n49265 = pi18 ? n31939 : n49264;
  assign n49266 = pi17 ? n20563 : n49265;
  assign n49267 = pi16 ? n41632 : n49266;
  assign n49268 = pi15 ? n49261 : n49267;
  assign n49269 = pi19 ? n2723 : n9483;
  assign n49270 = pi18 ? n31939 : n49269;
  assign n49271 = pi17 ? n20563 : n49270;
  assign n49272 = pi16 ? n41632 : n49271;
  assign n49273 = pi20 ? n31266 : n181;
  assign n49274 = pi20 ? n2973 : n3393;
  assign n49275 = pi19 ? n49273 : n49274;
  assign n49276 = pi20 ? n22881 : n19084;
  assign n49277 = pi19 ? n49276 : n7050;
  assign n49278 = pi18 ? n49275 : n49277;
  assign n49279 = pi17 ? n20563 : n49278;
  assign n49280 = pi16 ? n41632 : n49279;
  assign n49281 = pi15 ? n49272 : n49280;
  assign n49282 = pi14 ? n49268 : n49281;
  assign n49283 = pi19 ? n31267 : n35667;
  assign n49284 = pi19 ? n32794 : n7050;
  assign n49285 = pi18 ? n49283 : n49284;
  assign n49286 = pi17 ? n20563 : n49285;
  assign n49287 = pi16 ? n43263 : n49286;
  assign n49288 = pi20 ? n20563 : n297;
  assign n49289 = pi20 ? n1003 : n27484;
  assign n49290 = pi19 ? n49288 : n49289;
  assign n49291 = pi19 ? n32794 : n5831;
  assign n49292 = pi18 ? n49290 : n49291;
  assign n49293 = pi17 ? n20563 : n49292;
  assign n49294 = pi16 ? n43263 : n49293;
  assign n49295 = pi15 ? n49287 : n49294;
  assign n49296 = pi20 ? n24865 : n24220;
  assign n49297 = pi19 ? n49296 : n2654;
  assign n49298 = pi18 ? n32377 : n49297;
  assign n49299 = pi17 ? n20563 : n49298;
  assign n49300 = pi16 ? n43263 : n49299;
  assign n49301 = pi20 ? n24865 : n25199;
  assign n49302 = pi19 ? n49301 : n2654;
  assign n49303 = pi18 ? n32377 : n49302;
  assign n49304 = pi17 ? n20563 : n49303;
  assign n49305 = pi16 ? n43263 : n49304;
  assign n49306 = pi15 ? n49300 : n49305;
  assign n49307 = pi14 ? n49295 : n49306;
  assign n49308 = pi13 ? n49282 : n49307;
  assign n49309 = pi20 ? n43010 : n30868;
  assign n49310 = pi19 ? n49309 : n30868;
  assign n49311 = pi18 ? n49310 : n30868;
  assign n49312 = pi21 ? n30868 : n29133;
  assign n49313 = pi20 ? n49312 : n37;
  assign n49314 = pi19 ? n49313 : n21611;
  assign n49315 = pi22 ? n685 : n4537;
  assign n49316 = pi21 ? n49315 : n316;
  assign n49317 = pi20 ? n2729 : n49316;
  assign n49318 = pi19 ? n49317 : n2702;
  assign n49319 = pi18 ? n49314 : n49318;
  assign n49320 = pi17 ? n49311 : n49319;
  assign n49321 = pi16 ? n43263 : n49320;
  assign n49322 = pi19 ? n32 : n30868;
  assign n49323 = pi18 ? n32 : n49322;
  assign n49324 = pi17 ? n32 : n49323;
  assign n49325 = pi20 ? n787 : n34537;
  assign n49326 = pi19 ? n49325 : n1823;
  assign n49327 = pi18 ? n46193 : n49326;
  assign n49328 = pi17 ? n30868 : n49327;
  assign n49329 = pi16 ? n49324 : n49328;
  assign n49330 = pi15 ? n49321 : n49329;
  assign n49331 = pi20 ? n32 : n47835;
  assign n49332 = pi19 ? n49331 : n30868;
  assign n49333 = pi18 ? n32 : n49332;
  assign n49334 = pi17 ? n32 : n49333;
  assign n49335 = pi22 ? n37809 : n30868;
  assign n49336 = pi21 ? n30868 : n49335;
  assign n49337 = pi21 ? n37240 : n745;
  assign n49338 = pi20 ? n49336 : n49337;
  assign n49339 = pi22 ? n37809 : n812;
  assign n49340 = pi21 ? n49339 : n825;
  assign n49341 = pi22 ? n745 : n37809;
  assign n49342 = pi21 ? n49341 : n3520;
  assign n49343 = pi20 ? n49340 : n49342;
  assign n49344 = pi19 ? n49338 : n49343;
  assign n49345 = pi22 ? n745 : n158;
  assign n49346 = pi21 ? n49345 : n157;
  assign n49347 = pi21 ? n819 : n8643;
  assign n49348 = pi20 ? n49346 : n49347;
  assign n49349 = pi19 ? n49348 : n1823;
  assign n49350 = pi18 ? n49344 : n49349;
  assign n49351 = pi17 ? n30868 : n49350;
  assign n49352 = pi16 ? n49334 : n49351;
  assign n49353 = pi19 ? n32 : n46729;
  assign n49354 = pi18 ? n32 : n49353;
  assign n49355 = pi17 ? n32 : n49354;
  assign n49356 = pi20 ? n36798 : n48374;
  assign n49357 = pi19 ? n49356 : n33792;
  assign n49358 = pi18 ? n49357 : n33792;
  assign n49359 = pi20 ? n33792 : n139;
  assign n49360 = pi19 ? n49359 : n139;
  assign n49361 = pi21 ? n248 : n13408;
  assign n49362 = pi20 ? n875 : n49361;
  assign n49363 = pi19 ? n49362 : n32;
  assign n49364 = pi18 ? n49360 : n49363;
  assign n49365 = pi17 ? n49358 : n49364;
  assign n49366 = pi16 ? n49355 : n49365;
  assign n49367 = pi15 ? n49352 : n49366;
  assign n49368 = pi14 ? n49330 : n49367;
  assign n49369 = pi21 ? n36798 : n36659;
  assign n49370 = pi20 ? n46728 : n49369;
  assign n49371 = pi19 ? n32 : n49370;
  assign n49372 = pi18 ? n32 : n49371;
  assign n49373 = pi17 ? n32 : n49372;
  assign n49374 = pi21 ? n46260 : n48405;
  assign n49375 = pi20 ? n49374 : n36659;
  assign n49376 = pi19 ? n49375 : n36659;
  assign n49377 = pi18 ? n49376 : n36659;
  assign n49378 = pi20 ? n36659 : n335;
  assign n49379 = pi19 ? n49378 : n335;
  assign n49380 = pi21 ? n316 : n13408;
  assign n49381 = pi20 ? n36837 : n49380;
  assign n49382 = pi19 ? n49381 : n32;
  assign n49383 = pi18 ? n49379 : n49382;
  assign n49384 = pi17 ? n49377 : n49383;
  assign n49385 = pi16 ? n49373 : n49384;
  assign n49386 = pi21 ? n48856 : n43198;
  assign n49387 = pi20 ? n49386 : n43198;
  assign n49388 = pi19 ? n32 : n49387;
  assign n49389 = pi18 ? n32 : n49388;
  assign n49390 = pi17 ? n32 : n49389;
  assign n49391 = pi20 ? n43198 : n36659;
  assign n49392 = pi19 ? n49391 : n36659;
  assign n49393 = pi18 ? n49392 : n36659;
  assign n49394 = pi21 ? n36837 : n1091;
  assign n49395 = pi20 ? n49394 : n5205;
  assign n49396 = pi19 ? n49395 : n32;
  assign n49397 = pi18 ? n49379 : n49396;
  assign n49398 = pi17 ? n49393 : n49397;
  assign n49399 = pi16 ? n49390 : n49398;
  assign n49400 = pi15 ? n49385 : n49399;
  assign n49401 = pi21 ? n43198 : n36798;
  assign n49402 = pi20 ? n49386 : n49401;
  assign n49403 = pi19 ? n32 : n49402;
  assign n49404 = pi18 ? n32 : n49403;
  assign n49405 = pi17 ? n32 : n49404;
  assign n49406 = pi23 ? n43198 : n36781;
  assign n49407 = pi22 ? n49406 : n36798;
  assign n49408 = pi21 ? n47397 : n49407;
  assign n49409 = pi20 ? n49408 : n38923;
  assign n49410 = pi19 ? n49409 : n36781;
  assign n49411 = pi18 ? n49410 : n36781;
  assign n49412 = pi23 ? n36781 : n36798;
  assign n49413 = pi22 ? n49412 : n36781;
  assign n49414 = pi21 ? n36781 : n49413;
  assign n49415 = pi21 ? n43203 : n363;
  assign n49416 = pi20 ? n49414 : n49415;
  assign n49417 = pi20 ? n36813 : n34831;
  assign n49418 = pi19 ? n49416 : n49417;
  assign n49419 = pi20 ? n157 : n18285;
  assign n49420 = pi19 ? n49419 : n32;
  assign n49421 = pi18 ? n49418 : n49420;
  assign n49422 = pi17 ? n49411 : n49421;
  assign n49423 = pi16 ? n49405 : n49422;
  assign n49424 = pi21 ? n43198 : n36781;
  assign n49425 = pi20 ? n43198 : n49424;
  assign n49426 = pi19 ? n49425 : n36781;
  assign n49427 = pi18 ? n49426 : n36781;
  assign n49428 = pi20 ? n42170 : n49415;
  assign n49429 = pi19 ? n49428 : n157;
  assign n49430 = pi18 ? n49429 : n46785;
  assign n49431 = pi17 ? n49427 : n49430;
  assign n49432 = pi16 ? n49390 : n49431;
  assign n49433 = pi15 ? n49423 : n49432;
  assign n49434 = pi14 ? n49400 : n49433;
  assign n49435 = pi13 ? n49368 : n49434;
  assign n49436 = pi12 ? n49308 : n49435;
  assign n49437 = pi11 ? n49257 : n49436;
  assign n49438 = pi10 ? n49123 : n49437;
  assign n49439 = pi09 ? n48920 : n49438;
  assign n49440 = pi18 ? n42644 : n20563;
  assign n49441 = pi21 ? n37 : n31890;
  assign n49442 = pi20 ? n49441 : n37;
  assign n49443 = pi19 ? n49442 : n48898;
  assign n49444 = pi18 ? n20563 : n49443;
  assign n49445 = pi17 ? n49440 : n49444;
  assign n49446 = pi16 ? n32 : n49445;
  assign n49447 = pi15 ? n32 : n49446;
  assign n49448 = pi18 ? n42654 : n20563;
  assign n49449 = pi17 ? n49448 : n48909;
  assign n49450 = pi16 ? n32 : n49449;
  assign n49451 = pi18 ? n42680 : n20563;
  assign n49452 = pi23 ? n139 : n8184;
  assign n49453 = pi22 ? n49452 : n32;
  assign n49454 = pi21 ? n49453 : n32;
  assign n49455 = pi20 ? n37 : n49454;
  assign n49456 = pi19 ? n48906 : n49455;
  assign n49457 = pi18 ? n20563 : n49456;
  assign n49458 = pi17 ? n49451 : n49457;
  assign n49459 = pi16 ? n32 : n49458;
  assign n49460 = pi15 ? n49450 : n49459;
  assign n49461 = pi14 ? n49447 : n49460;
  assign n49462 = pi13 ? n32 : n49461;
  assign n49463 = pi12 ? n32 : n49462;
  assign n49464 = pi11 ? n32 : n49463;
  assign n49465 = pi10 ? n32 : n49464;
  assign n49466 = pi22 ? n27388 : n32;
  assign n49467 = pi21 ? n49466 : n32;
  assign n49468 = pi20 ? n37 : n49467;
  assign n49469 = pi19 ? n37 : n49468;
  assign n49470 = pi18 ? n20563 : n49469;
  assign n49471 = pi17 ? n48897 : n49470;
  assign n49472 = pi16 ? n32 : n49471;
  assign n49473 = pi17 ? n48460 : n48928;
  assign n49474 = pi16 ? n32 : n49473;
  assign n49475 = pi15 ? n49472 : n49474;
  assign n49476 = pi17 ? n48466 : n48934;
  assign n49477 = pi16 ? n32 : n49476;
  assign n49478 = pi20 ? n3086 : n16991;
  assign n49479 = pi19 ? n32871 : n49478;
  assign n49480 = pi18 ? n20563 : n49479;
  assign n49481 = pi17 ? n48469 : n49480;
  assign n49482 = pi16 ? n32 : n49481;
  assign n49483 = pi15 ? n49477 : n49482;
  assign n49484 = pi14 ? n49475 : n49483;
  assign n49485 = pi18 ? n40485 : n20563;
  assign n49486 = pi20 ? n997 : n18040;
  assign n49487 = pi19 ? n32287 : n49486;
  assign n49488 = pi18 ? n20563 : n49487;
  assign n49489 = pi17 ? n49485 : n49488;
  assign n49490 = pi16 ? n32 : n49489;
  assign n49491 = pi20 ? n20563 : n36977;
  assign n49492 = pi19 ? n20563 : n49491;
  assign n49493 = pi20 ? n37 : n32927;
  assign n49494 = pi19 ? n37 : n49493;
  assign n49495 = pi18 ? n49492 : n49494;
  assign n49496 = pi17 ? n47929 : n49495;
  assign n49497 = pi16 ? n32 : n49496;
  assign n49498 = pi15 ? n49490 : n49497;
  assign n49499 = pi20 ? n37 : n5772;
  assign n49500 = pi19 ? n32933 : n49499;
  assign n49501 = pi18 ? n20563 : n49500;
  assign n49502 = pi17 ? n48488 : n49501;
  assign n49503 = pi16 ? n32 : n49502;
  assign n49504 = pi20 ? n649 : n5784;
  assign n49505 = pi19 ? n37 : n49504;
  assign n49506 = pi18 ? n34865 : n49505;
  assign n49507 = pi17 ? n48488 : n49506;
  assign n49508 = pi16 ? n32 : n49507;
  assign n49509 = pi15 ? n49503 : n49508;
  assign n49510 = pi14 ? n49498 : n49509;
  assign n49511 = pi13 ? n49484 : n49510;
  assign n49512 = pi20 ? n649 : n21388;
  assign n49513 = pi19 ? n30097 : n49512;
  assign n49514 = pi18 ? n20563 : n49513;
  assign n49515 = pi17 ? n47451 : n49514;
  assign n49516 = pi16 ? n32 : n49515;
  assign n49517 = pi20 ? n649 : n32960;
  assign n49518 = pi19 ? n37 : n49517;
  assign n49519 = pi18 ? n38963 : n49518;
  assign n49520 = pi17 ? n46302 : n49519;
  assign n49521 = pi16 ? n32 : n49520;
  assign n49522 = pi15 ? n49516 : n49521;
  assign n49523 = pi20 ? n20157 : n7733;
  assign n49524 = pi19 ? n37 : n49523;
  assign n49525 = pi18 ? n34295 : n49524;
  assign n49526 = pi17 ? n46832 : n49525;
  assign n49527 = pi16 ? n32 : n49526;
  assign n49528 = pi20 ? n569 : n17591;
  assign n49529 = pi19 ? n37 : n49528;
  assign n49530 = pi18 ? n33823 : n49529;
  assign n49531 = pi17 ? n47964 : n49530;
  assign n49532 = pi16 ? n32 : n49531;
  assign n49533 = pi15 ? n49527 : n49532;
  assign n49534 = pi14 ? n49522 : n49533;
  assign n49535 = pi20 ? n36929 : n30096;
  assign n49536 = pi19 ? n20563 : n49535;
  assign n49537 = pi20 ? n3393 : n3176;
  assign n49538 = pi19 ? n37 : n49537;
  assign n49539 = pi18 ? n49536 : n49538;
  assign n49540 = pi17 ? n46866 : n49539;
  assign n49541 = pi16 ? n32 : n49540;
  assign n49542 = pi19 ? n20563 : n40123;
  assign n49543 = pi20 ? n6402 : n6417;
  assign n49544 = pi19 ? n37 : n49543;
  assign n49545 = pi18 ? n49542 : n49544;
  assign n49546 = pi17 ? n20563 : n49545;
  assign n49547 = pi16 ? n32 : n49546;
  assign n49548 = pi15 ? n49541 : n49547;
  assign n49549 = pi18 ? n39585 : n49005;
  assign n49550 = pi17 ? n20563 : n49549;
  assign n49551 = pi16 ? n46326 : n49550;
  assign n49552 = pi18 ? n32872 : n49005;
  assign n49553 = pi17 ? n20563 : n49552;
  assign n49554 = pi16 ? n45233 : n49553;
  assign n49555 = pi15 ? n49551 : n49554;
  assign n49556 = pi14 ? n49548 : n49555;
  assign n49557 = pi13 ? n49534 : n49556;
  assign n49558 = pi12 ? n49511 : n49557;
  assign n49559 = pi21 ? n31294 : n29133;
  assign n49560 = pi20 ? n49559 : n37;
  assign n49561 = pi19 ? n20563 : n49560;
  assign n49562 = pi18 ? n49561 : n49019;
  assign n49563 = pi17 ? n20563 : n49562;
  assign n49564 = pi16 ? n44635 : n49563;
  assign n49565 = pi18 ? n33858 : n49024;
  assign n49566 = pi17 ? n20563 : n49565;
  assign n49567 = pi16 ? n44635 : n49566;
  assign n49568 = pi15 ? n49564 : n49567;
  assign n49569 = pi18 ? n32288 : n49030;
  assign n49570 = pi17 ? n20563 : n49569;
  assign n49571 = pi16 ? n44635 : n49570;
  assign n49572 = pi18 ? n34891 : n49036;
  assign n49573 = pi17 ? n20563 : n49572;
  assign n49574 = pi16 ? n45740 : n49573;
  assign n49575 = pi15 ? n49571 : n49574;
  assign n49576 = pi14 ? n49568 : n49575;
  assign n49577 = pi16 ? n44644 : n49046;
  assign n49578 = pi20 ? n48089 : n2701;
  assign n49579 = pi19 ? n37 : n49578;
  assign n49580 = pi18 ? n42358 : n49579;
  assign n49581 = pi17 ? n20563 : n49580;
  assign n49582 = pi16 ? n44653 : n49581;
  assign n49583 = pi15 ? n49577 : n49582;
  assign n49584 = pi16 ? n44653 : n49055;
  assign n49585 = pi16 ? n44653 : n49061;
  assign n49586 = pi15 ? n49584 : n49585;
  assign n49587 = pi14 ? n49583 : n49586;
  assign n49588 = pi13 ? n49576 : n49587;
  assign n49589 = pi20 ? n49066 : n2653;
  assign n49590 = pi19 ? n37 : n49589;
  assign n49591 = pi18 ? n33299 : n49590;
  assign n49592 = pi17 ? n20563 : n49591;
  assign n49593 = pi16 ? n44223 : n49592;
  assign n49594 = pi18 ? n32 : n28159;
  assign n49595 = pi17 ? n32 : n49594;
  assign n49596 = pi20 ? n19208 : n2653;
  assign n49597 = pi19 ? n99 : n49596;
  assign n49598 = pi18 ? n49072 : n49597;
  assign n49599 = pi17 ? n20563 : n49598;
  assign n49600 = pi16 ? n49595 : n49599;
  assign n49601 = pi15 ? n49593 : n49600;
  assign n49602 = pi19 ? n38962 : n17013;
  assign n49603 = pi20 ? n20978 : n1822;
  assign n49604 = pi19 ? n3050 : n49603;
  assign n49605 = pi18 ? n49602 : n49604;
  assign n49606 = pi17 ? n20563 : n49605;
  assign n49607 = pi16 ? n49595 : n49606;
  assign n49608 = pi19 ? n38962 : n34261;
  assign n49609 = pi20 ? n19171 : n1822;
  assign n49610 = pi19 ? n99 : n49609;
  assign n49611 = pi18 ? n49608 : n49610;
  assign n49612 = pi17 ? n20563 : n49611;
  assign n49613 = pi16 ? n44227 : n49612;
  assign n49614 = pi15 ? n49607 : n49613;
  assign n49615 = pi14 ? n49601 : n49614;
  assign n49616 = pi21 ? n36489 : n39164;
  assign n49617 = pi20 ? n20563 : n49616;
  assign n49618 = pi19 ? n49617 : n26407;
  assign n49619 = pi21 ? n775 : n6535;
  assign n49620 = pi20 ? n49619 : n32;
  assign n49621 = pi19 ? n2242 : n49620;
  assign n49622 = pi18 ? n49618 : n49621;
  assign n49623 = pi17 ? n20563 : n49622;
  assign n49624 = pi16 ? n44227 : n49623;
  assign n49625 = pi21 ? n30868 : n39164;
  assign n49626 = pi20 ? n20563 : n49625;
  assign n49627 = pi19 ? n49626 : n26407;
  assign n49628 = pi21 ? n775 : n397;
  assign n49629 = pi20 ? n49628 : n32;
  assign n49630 = pi19 ? n99 : n49629;
  assign n49631 = pi18 ? n49627 : n49630;
  assign n49632 = pi17 ? n20563 : n49631;
  assign n49633 = pi16 ? n44227 : n49632;
  assign n49634 = pi15 ? n49624 : n49633;
  assign n49635 = pi19 ? n35854 : n17013;
  assign n49636 = pi19 ? n49108 : n21475;
  assign n49637 = pi18 ? n49635 : n49636;
  assign n49638 = pi17 ? n20563 : n49637;
  assign n49639 = pi16 ? n43664 : n49638;
  assign n49640 = pi21 ? n99 : n9584;
  assign n49641 = pi20 ? n49640 : n32;
  assign n49642 = pi19 ? n26407 : n49641;
  assign n49643 = pi18 ? n33916 : n49642;
  assign n49644 = pi17 ? n20563 : n49643;
  assign n49645 = pi16 ? n43664 : n49644;
  assign n49646 = pi15 ? n49639 : n49645;
  assign n49647 = pi14 ? n49634 : n49646;
  assign n49648 = pi13 ? n49615 : n49647;
  assign n49649 = pi12 ? n49588 : n49648;
  assign n49650 = pi11 ? n49558 : n49649;
  assign n49651 = pi19 ? n35798 : n49124;
  assign n49652 = pi19 ? n20743 : n49128;
  assign n49653 = pi18 ? n49651 : n49652;
  assign n49654 = pi17 ? n20563 : n49653;
  assign n49655 = pi16 ? n43675 : n49654;
  assign n49656 = pi16 ? n43675 : n49138;
  assign n49657 = pi15 ? n49655 : n49656;
  assign n49658 = pi21 ? n30868 : n39182;
  assign n49659 = pi20 ? n40791 : n49658;
  assign n49660 = pi19 ? n49659 : n37;
  assign n49661 = pi18 ? n49660 : n49136;
  assign n49662 = pi17 ? n20563 : n49661;
  assign n49663 = pi16 ? n43675 : n49662;
  assign n49664 = pi19 ? n49146 : n20107;
  assign n49665 = pi18 ? n37029 : n49664;
  assign n49666 = pi17 ? n20563 : n49665;
  assign n49667 = pi16 ? n43685 : n49666;
  assign n49668 = pi15 ? n49663 : n49667;
  assign n49669 = pi14 ? n49657 : n49668;
  assign n49670 = pi18 ? n37029 : n49154;
  assign n49671 = pi17 ? n20563 : n49670;
  assign n49672 = pi16 ? n44688 : n49671;
  assign n49673 = pi21 ? n204 : n7041;
  assign n49674 = pi20 ? n49673 : n32;
  assign n49675 = pi19 ? n14962 : n49674;
  assign n49676 = pi18 ? n39038 : n49675;
  assign n49677 = pi17 ? n20563 : n49676;
  assign n49678 = pi16 ? n43228 : n49677;
  assign n49679 = pi15 ? n49672 : n49678;
  assign n49680 = pi21 ? n28649 : n4101;
  assign n49681 = pi20 ? n49680 : n32;
  assign n49682 = pi19 ? n8765 : n49681;
  assign n49683 = pi18 ? n35300 : n49682;
  assign n49684 = pi17 ? n20563 : n49683;
  assign n49685 = pi16 ? n43224 : n49684;
  assign n49686 = pi21 ? n28649 : n5829;
  assign n49687 = pi20 ? n49686 : n32;
  assign n49688 = pi19 ? n8765 : n49687;
  assign n49689 = pi18 ? n35300 : n49688;
  assign n49690 = pi17 ? n20563 : n49689;
  assign n49691 = pi16 ? n43224 : n49690;
  assign n49692 = pi15 ? n49685 : n49691;
  assign n49693 = pi14 ? n49679 : n49692;
  assign n49694 = pi13 ? n49669 : n49693;
  assign n49695 = pi16 ? n43224 : n49183;
  assign n49696 = pi18 ? n48574 : n49186;
  assign n49697 = pi17 ? n20563 : n49696;
  assign n49698 = pi16 ? n43228 : n49697;
  assign n49699 = pi15 ? n49695 : n49698;
  assign n49700 = pi18 ? n41334 : n49194;
  assign n49701 = pi17 ? n20563 : n49700;
  assign n49702 = pi16 ? n42646 : n49701;
  assign n49703 = pi19 ? n49199 : n21212;
  assign n49704 = pi18 ? n34949 : n49703;
  assign n49705 = pi17 ? n20563 : n49704;
  assign n49706 = pi16 ? n42646 : n49705;
  assign n49707 = pi15 ? n49702 : n49706;
  assign n49708 = pi14 ? n49699 : n49707;
  assign n49709 = pi20 ? n45599 : n30868;
  assign n49710 = pi19 ? n32 : n49709;
  assign n49711 = pi18 ? n32 : n49710;
  assign n49712 = pi17 ? n32 : n49711;
  assign n49713 = pi18 ? n34949 : n49214;
  assign n49714 = pi17 ? n49212 : n49713;
  assign n49715 = pi16 ? n49712 : n49714;
  assign n49716 = pi18 ? n35318 : n49223;
  assign n49717 = pi17 ? n49212 : n49716;
  assign n49718 = pi16 ? n49712 : n49717;
  assign n49719 = pi15 ? n49715 : n49718;
  assign n49720 = pi23 ? n32 : n33792;
  assign n49721 = pi22 ? n32 : n49720;
  assign n49722 = pi21 ? n49721 : n33792;
  assign n49723 = pi20 ? n49722 : n40958;
  assign n49724 = pi19 ? n32 : n49723;
  assign n49725 = pi18 ? n32 : n49724;
  assign n49726 = pi17 ? n32 : n49725;
  assign n49727 = pi19 ? n8928 : n17906;
  assign n49728 = pi18 ? n37649 : n49727;
  assign n49729 = pi17 ? n49236 : n49728;
  assign n49730 = pi16 ? n49726 : n49729;
  assign n49731 = pi19 ? n2095 : n9432;
  assign n49732 = pi18 ? n37649 : n49731;
  assign n49733 = pi17 ? n20563 : n49732;
  assign n49734 = pi16 ? n42682 : n49733;
  assign n49735 = pi15 ? n49730 : n49734;
  assign n49736 = pi14 ? n49719 : n49735;
  assign n49737 = pi13 ? n49708 : n49736;
  assign n49738 = pi12 ? n49694 : n49737;
  assign n49739 = pi18 ? n32369 : n49258;
  assign n49740 = pi17 ? n20563 : n49739;
  assign n49741 = pi16 ? n42682 : n49740;
  assign n49742 = pi19 ? n49263 : n10352;
  assign n49743 = pi18 ? n37649 : n49742;
  assign n49744 = pi17 ? n20563 : n49743;
  assign n49745 = pi16 ? n42682 : n49744;
  assign n49746 = pi15 ? n49741 : n49745;
  assign n49747 = pi19 ? n2723 : n8296;
  assign n49748 = pi18 ? n37649 : n49747;
  assign n49749 = pi17 ? n20563 : n49748;
  assign n49750 = pi16 ? n42682 : n49749;
  assign n49751 = pi20 ? n31925 : n181;
  assign n49752 = pi19 ? n49751 : n49274;
  assign n49753 = pi19 ? n49276 : n36391;
  assign n49754 = pi18 ? n49752 : n49753;
  assign n49755 = pi17 ? n20563 : n49754;
  assign n49756 = pi16 ? n42682 : n49755;
  assign n49757 = pi15 ? n49750 : n49756;
  assign n49758 = pi14 ? n49746 : n49757;
  assign n49759 = pi19 ? n31926 : n35667;
  assign n49760 = pi19 ? n32794 : n36391;
  assign n49761 = pi18 ? n49759 : n49760;
  assign n49762 = pi17 ? n20563 : n49761;
  assign n49763 = pi16 ? n42656 : n49762;
  assign n49764 = pi22 ? n30195 : n139;
  assign n49765 = pi21 ? n49764 : n297;
  assign n49766 = pi20 ? n20563 : n49765;
  assign n49767 = pi20 ? n1003 : n27962;
  assign n49768 = pi19 ? n49766 : n49767;
  assign n49769 = pi18 ? n49768 : n49291;
  assign n49770 = pi17 ? n20563 : n49769;
  assign n49771 = pi16 ? n44275 : n49770;
  assign n49772 = pi15 ? n49763 : n49771;
  assign n49773 = pi19 ? n49296 : n48320;
  assign n49774 = pi18 ? n32369 : n49773;
  assign n49775 = pi17 ? n20563 : n49774;
  assign n49776 = pi16 ? n44275 : n49775;
  assign n49777 = pi18 ? n32369 : n49302;
  assign n49778 = pi17 ? n20563 : n49777;
  assign n49779 = pi16 ? n44275 : n49778;
  assign n49780 = pi15 ? n49776 : n49779;
  assign n49781 = pi14 ? n49772 : n49780;
  assign n49782 = pi13 ? n49758 : n49781;
  assign n49783 = pi21 ? n30868 : n31924;
  assign n49784 = pi20 ? n49783 : n37;
  assign n49785 = pi19 ? n49784 : n21611;
  assign n49786 = pi18 ? n49785 : n49318;
  assign n49787 = pi17 ? n49311 : n49786;
  assign n49788 = pi16 ? n44275 : n49787;
  assign n49789 = pi19 ? n32 : n47193;
  assign n49790 = pi18 ? n32 : n49789;
  assign n49791 = pi17 ? n32 : n49790;
  assign n49792 = pi19 ? n40417 : n99;
  assign n49793 = pi18 ? n49792 : n49326;
  assign n49794 = pi17 ? n30868 : n49793;
  assign n49795 = pi16 ? n49791 : n49794;
  assign n49796 = pi15 ? n49788 : n49795;
  assign n49797 = pi19 ? n32 : n47323;
  assign n49798 = pi18 ? n32 : n49797;
  assign n49799 = pi17 ? n32 : n49798;
  assign n49800 = pi23 ? n30868 : n139;
  assign n49801 = pi21 ? n30868 : n49800;
  assign n49802 = pi20 ? n30868 : n49801;
  assign n49803 = pi22 ? n49800 : n139;
  assign n49804 = pi21 ? n49803 : n139;
  assign n49805 = pi22 ? n139 : n49800;
  assign n49806 = pi21 ? n49805 : n248;
  assign n49807 = pi20 ? n49804 : n49806;
  assign n49808 = pi19 ? n49802 : n49807;
  assign n49809 = pi21 ? n248 : n8643;
  assign n49810 = pi20 ? n249 : n49809;
  assign n49811 = pi19 ? n49810 : n1823;
  assign n49812 = pi18 ? n49808 : n49811;
  assign n49813 = pi17 ? n30868 : n49812;
  assign n49814 = pi16 ? n49799 : n49813;
  assign n49815 = pi21 ? n32 : n41600;
  assign n49816 = pi20 ? n49815 : n36798;
  assign n49817 = pi19 ? n32 : n49816;
  assign n49818 = pi18 ? n32 : n49817;
  assign n49819 = pi17 ? n32 : n49818;
  assign n49820 = pi22 ? n1484 : n2834;
  assign n49821 = pi21 ? n248 : n49820;
  assign n49822 = pi20 ? n875 : n49821;
  assign n49823 = pi19 ? n49822 : n32;
  assign n49824 = pi18 ? n46208 : n49823;
  assign n49825 = pi17 ? n49358 : n49824;
  assign n49826 = pi16 ? n49819 : n49825;
  assign n49827 = pi15 ? n49814 : n49826;
  assign n49828 = pi14 ? n49796 : n49827;
  assign n49829 = pi20 ? n48822 : n49369;
  assign n49830 = pi19 ? n32 : n49829;
  assign n49831 = pi18 ? n32 : n49830;
  assign n49832 = pi17 ? n32 : n49831;
  assign n49833 = pi22 ? n36659 : n37276;
  assign n49834 = pi21 ? n49833 : n36659;
  assign n49835 = pi20 ? n49834 : n36659;
  assign n49836 = pi19 ? n49835 : n36659;
  assign n49837 = pi18 ? n49836 : n36659;
  assign n49838 = pi20 ? n36659 : n46244;
  assign n49839 = pi19 ? n49838 : n335;
  assign n49840 = pi18 ? n49839 : n49382;
  assign n49841 = pi17 ? n49837 : n49840;
  assign n49842 = pi16 ? n49832 : n49841;
  assign n49843 = pi23 ? n46274 : n43198;
  assign n49844 = pi22 ? n49843 : n43198;
  assign n49845 = pi21 ? n32 : n49844;
  assign n49846 = pi20 ? n49845 : n43198;
  assign n49847 = pi19 ? n32 : n49846;
  assign n49848 = pi18 ? n32 : n49847;
  assign n49849 = pi17 ? n32 : n49848;
  assign n49850 = pi18 ? n49839 : n49396;
  assign n49851 = pi17 ? n49393 : n49850;
  assign n49852 = pi16 ? n49849 : n49851;
  assign n49853 = pi15 ? n49842 : n49852;
  assign n49854 = pi20 ? n48857 : n49401;
  assign n49855 = pi19 ? n32 : n49854;
  assign n49856 = pi18 ? n32 : n49855;
  assign n49857 = pi17 ? n32 : n49856;
  assign n49858 = pi22 ? n36798 : n43199;
  assign n49859 = pi21 ? n49858 : n39972;
  assign n49860 = pi20 ? n49859 : n38923;
  assign n49861 = pi19 ? n49860 : n36781;
  assign n49862 = pi18 ? n49861 : n36781;
  assign n49863 = pi20 ? n36781 : n49415;
  assign n49864 = pi19 ? n49863 : n49417;
  assign n49865 = pi18 ? n49864 : n49420;
  assign n49866 = pi17 ? n49862 : n49865;
  assign n49867 = pi16 ? n49857 : n49866;
  assign n49868 = pi19 ? n32 : n47412;
  assign n49869 = pi18 ? n32 : n49868;
  assign n49870 = pi17 ? n32 : n49869;
  assign n49871 = pi21 ? n43644 : n47895;
  assign n49872 = pi20 ? n42170 : n49871;
  assign n49873 = pi19 ? n49872 : n157;
  assign n49874 = pi21 ? n46267 : n3523;
  assign n49875 = pi20 ? n157 : n49874;
  assign n49876 = pi19 ? n49875 : n32;
  assign n49877 = pi18 ? n49873 : n49876;
  assign n49878 = pi17 ? n49427 : n49877;
  assign n49879 = pi16 ? n49870 : n49878;
  assign n49880 = pi15 ? n49867 : n49879;
  assign n49881 = pi14 ? n49853 : n49880;
  assign n49882 = pi13 ? n49828 : n49881;
  assign n49883 = pi12 ? n49782 : n49882;
  assign n49884 = pi11 ? n49738 : n49883;
  assign n49885 = pi10 ? n49650 : n49884;
  assign n49886 = pi09 ? n49465 : n49885;
  assign n49887 = pi08 ? n49439 : n49886;
  assign n49888 = pi18 ? n44246 : n20563;
  assign n49889 = pi19 ? n37 : n18847;
  assign n49890 = pi18 ? n20563 : n49889;
  assign n49891 = pi17 ? n49888 : n49890;
  assign n49892 = pi16 ? n32 : n49891;
  assign n49893 = pi15 ? n32 : n49892;
  assign n49894 = pi18 ? n43222 : n20563;
  assign n49895 = pi20 ? n37 : n5624;
  assign n49896 = pi19 ? n48906 : n49895;
  assign n49897 = pi18 ? n20563 : n49896;
  assign n49898 = pi17 ? n49894 : n49897;
  assign n49899 = pi16 ? n32 : n49898;
  assign n49900 = pi18 ? n48623 : n20563;
  assign n49901 = pi17 ? n49900 : n49897;
  assign n49902 = pi16 ? n32 : n49901;
  assign n49903 = pi15 ? n49899 : n49902;
  assign n49904 = pi14 ? n49893 : n49903;
  assign n49905 = pi13 ? n32 : n49904;
  assign n49906 = pi12 ? n32 : n49905;
  assign n49907 = pi11 ? n32 : n49906;
  assign n49908 = pi10 ? n32 : n49907;
  assign n49909 = pi22 ? n5011 : n5631;
  assign n49910 = pi21 ? n49909 : n32;
  assign n49911 = pi20 ? n37 : n49910;
  assign n49912 = pi19 ? n37 : n49911;
  assign n49913 = pi18 ? n20563 : n49912;
  assign n49914 = pi17 ? n49440 : n49913;
  assign n49915 = pi16 ? n32 : n49914;
  assign n49916 = pi21 ? n37 : n36249;
  assign n49917 = pi20 ? n49916 : n37;
  assign n49918 = pi22 ? n364 : n2468;
  assign n49919 = pi21 ? n49918 : n32;
  assign n49920 = pi20 ? n3096 : n49919;
  assign n49921 = pi19 ? n49917 : n49920;
  assign n49922 = pi18 ? n20563 : n49921;
  assign n49923 = pi17 ? n48897 : n49922;
  assign n49924 = pi16 ? n32 : n49923;
  assign n49925 = pi15 ? n49915 : n49924;
  assign n49926 = pi20 ? n3086 : n33325;
  assign n49927 = pi19 ? n32898 : n49926;
  assign n49928 = pi18 ? n20563 : n49927;
  assign n49929 = pi17 ? n48904 : n49928;
  assign n49930 = pi16 ? n32 : n49929;
  assign n49931 = pi20 ? n37 : n3953;
  assign n49932 = pi19 ? n32898 : n49931;
  assign n49933 = pi18 ? n20563 : n49932;
  assign n49934 = pi17 ? n48912 : n49933;
  assign n49935 = pi16 ? n32 : n49934;
  assign n49936 = pi15 ? n49930 : n49935;
  assign n49937 = pi14 ? n49925 : n49936;
  assign n49938 = pi18 ? n42206 : n20563;
  assign n49939 = pi19 ? n31267 : n49931;
  assign n49940 = pi18 ? n20563 : n49939;
  assign n49941 = pi17 ? n49938 : n49940;
  assign n49942 = pi16 ? n32 : n49941;
  assign n49943 = pi22 ? n6961 : n32;
  assign n49944 = pi21 ? n49943 : n32;
  assign n49945 = pi20 ? n37 : n49944;
  assign n49946 = pi19 ? n30097 : n49945;
  assign n49947 = pi18 ? n48972 : n49946;
  assign n49948 = pi17 ? n48466 : n49947;
  assign n49949 = pi16 ? n32 : n49948;
  assign n49950 = pi15 ? n49942 : n49949;
  assign n49951 = pi20 ? n37439 : n37;
  assign n49952 = pi19 ? n49951 : n49945;
  assign n49953 = pi18 ? n20563 : n49952;
  assign n49954 = pi17 ? n47929 : n49953;
  assign n49955 = pi16 ? n32 : n49954;
  assign n49956 = pi21 ? n41221 : n32;
  assign n49957 = pi20 ? n649 : n49956;
  assign n49958 = pi19 ? n31280 : n49957;
  assign n49959 = pi18 ? n20563 : n49958;
  assign n49960 = pi17 ? n47929 : n49959;
  assign n49961 = pi16 ? n32 : n49960;
  assign n49962 = pi15 ? n49955 : n49961;
  assign n49963 = pi14 ? n49950 : n49962;
  assign n49964 = pi13 ? n49937 : n49963;
  assign n49965 = pi20 ? n577 : n5784;
  assign n49966 = pi19 ? n31267 : n49965;
  assign n49967 = pi18 ? n20563 : n49966;
  assign n49968 = pi17 ? n47935 : n49967;
  assign n49969 = pi16 ? n32 : n49968;
  assign n49970 = pi20 ? n649 : n33391;
  assign n49971 = pi19 ? n30097 : n49970;
  assign n49972 = pi18 ? n48972 : n49971;
  assign n49973 = pi17 ? n47947 : n49972;
  assign n49974 = pi16 ? n32 : n49973;
  assign n49975 = pi15 ? n49969 : n49974;
  assign n49976 = pi20 ? n649 : n47948;
  assign n49977 = pi19 ? n37 : n49976;
  assign n49978 = pi18 ? n34869 : n49977;
  assign n49979 = pi17 ? n48949 : n49978;
  assign n49980 = pi16 ? n32 : n49979;
  assign n49981 = pi22 ? n1150 : n32;
  assign n49982 = pi21 ? n49981 : n32;
  assign n49983 = pi20 ? n649 : n49982;
  assign n49984 = pi19 ? n30097 : n49983;
  assign n49985 = pi18 ? n20563 : n49984;
  assign n49986 = pi17 ? n48488 : n49985;
  assign n49987 = pi16 ? n32 : n49986;
  assign n49988 = pi15 ? n49980 : n49987;
  assign n49989 = pi14 ? n49975 : n49988;
  assign n49990 = pi20 ? n3393 : n31964;
  assign n49991 = pi19 ? n37 : n49990;
  assign n49992 = pi18 ? n20563 : n49991;
  assign n49993 = pi17 ? n47964 : n49992;
  assign n49994 = pi16 ? n32 : n49993;
  assign n49995 = pi20 ? n6402 : n7724;
  assign n49996 = pi19 ? n37 : n49995;
  assign n49997 = pi18 ? n34258 : n49996;
  assign n49998 = pi17 ? n45707 : n49997;
  assign n49999 = pi16 ? n32 : n49998;
  assign n50000 = pi15 ? n49994 : n49999;
  assign n50001 = pi17 ? n46859 : n49997;
  assign n50002 = pi16 ? n32 : n50001;
  assign n50003 = pi20 ? n3393 : n7724;
  assign n50004 = pi19 ? n37 : n50003;
  assign n50005 = pi18 ? n33260 : n50004;
  assign n50006 = pi17 ? n45715 : n50005;
  assign n50007 = pi16 ? n32 : n50006;
  assign n50008 = pi15 ? n50002 : n50007;
  assign n50009 = pi14 ? n50000 : n50008;
  assign n50010 = pi13 ? n49989 : n50009;
  assign n50011 = pi12 ? n49964 : n50010;
  assign n50012 = pi22 ? n363 : n583;
  assign n50013 = pi21 ? n37 : n50012;
  assign n50014 = pi20 ? n50013 : n3210;
  assign n50015 = pi19 ? n37 : n50014;
  assign n50016 = pi18 ? n34258 : n50015;
  assign n50017 = pi17 ? n46866 : n50016;
  assign n50018 = pi16 ? n32 : n50017;
  assign n50019 = pi19 ? n37 : n20896;
  assign n50020 = pi18 ? n34295 : n50019;
  assign n50021 = pi17 ? n46866 : n50020;
  assign n50022 = pi16 ? n32 : n50021;
  assign n50023 = pi15 ? n50018 : n50022;
  assign n50024 = pi20 ? n20563 : n30120;
  assign n50025 = pi19 ? n20563 : n50024;
  assign n50026 = pi20 ? n363 : n5830;
  assign n50027 = pi19 ? n37 : n50026;
  assign n50028 = pi18 ? n50025 : n50027;
  assign n50029 = pi17 ? n46312 : n50028;
  assign n50030 = pi16 ? n32 : n50029;
  assign n50031 = pi18 ? n34869 : n49019;
  assign n50032 = pi17 ? n20563 : n50031;
  assign n50033 = pi16 ? n32 : n50032;
  assign n50034 = pi15 ? n50030 : n50033;
  assign n50035 = pi14 ? n50023 : n50034;
  assign n50036 = pi19 ? n37 : n19607;
  assign n50037 = pi18 ? n34295 : n50036;
  assign n50038 = pi17 ? n20563 : n50037;
  assign n50039 = pi16 ? n46326 : n50038;
  assign n50040 = pi20 ? n382 : n2653;
  assign n50041 = pi19 ? n37 : n50040;
  assign n50042 = pi18 ? n33245 : n50041;
  assign n50043 = pi17 ? n20563 : n50042;
  assign n50044 = pi16 ? n45233 : n50043;
  assign n50045 = pi15 ? n50039 : n50044;
  assign n50046 = pi20 ? n24493 : n2653;
  assign n50047 = pi19 ? n37 : n50046;
  assign n50048 = pi18 ? n33260 : n50047;
  assign n50049 = pi17 ? n20563 : n50048;
  assign n50050 = pi16 ? n45233 : n50049;
  assign n50051 = pi20 ? n24493 : n2638;
  assign n50052 = pi19 ? n37 : n50051;
  assign n50053 = pi18 ? n34295 : n50052;
  assign n50054 = pi17 ? n20563 : n50053;
  assign n50055 = pi16 ? n45233 : n50054;
  assign n50056 = pi15 ? n50050 : n50055;
  assign n50057 = pi14 ? n50045 : n50056;
  assign n50058 = pi13 ? n50035 : n50057;
  assign n50059 = pi22 ? n112 : n316;
  assign n50060 = pi21 ? n37 : n50059;
  assign n50061 = pi20 ? n50060 : n2653;
  assign n50062 = pi19 ? n37 : n50061;
  assign n50063 = pi18 ? n34295 : n50062;
  assign n50064 = pi17 ? n20563 : n50063;
  assign n50065 = pi16 ? n44635 : n50064;
  assign n50066 = pi18 ? n32 : n37957;
  assign n50067 = pi17 ? n32 : n50066;
  assign n50068 = pi20 ? n31266 : n5077;
  assign n50069 = pi19 ? n20563 : n50068;
  assign n50070 = pi21 ? n99 : n25813;
  assign n50071 = pi20 ? n50070 : n2653;
  assign n50072 = pi19 ? n18853 : n50071;
  assign n50073 = pi18 ? n50069 : n50072;
  assign n50074 = pi17 ? n20563 : n50073;
  assign n50075 = pi16 ? n50067 : n50074;
  assign n50076 = pi15 ? n50065 : n50075;
  assign n50077 = pi20 ? n50070 : n1822;
  assign n50078 = pi19 ? n21611 : n50077;
  assign n50079 = pi18 ? n33260 : n50078;
  assign n50080 = pi17 ? n20563 : n50079;
  assign n50081 = pi16 ? n44644 : n50080;
  assign n50082 = pi22 ? n1656 : n316;
  assign n50083 = pi21 ? n99 : n50082;
  assign n50084 = pi20 ? n50083 : n1822;
  assign n50085 = pi19 ? n99 : n50084;
  assign n50086 = pi18 ? n32275 : n50085;
  assign n50087 = pi17 ? n20563 : n50086;
  assign n50088 = pi16 ? n44644 : n50087;
  assign n50089 = pi15 ? n50081 : n50088;
  assign n50090 = pi14 ? n50076 : n50089;
  assign n50091 = pi20 ? n20563 : n42006;
  assign n50092 = pi20 ? n31220 : n3039;
  assign n50093 = pi19 ? n50091 : n50092;
  assign n50094 = pi22 ? n1656 : n396;
  assign n50095 = pi21 ? n99 : n50094;
  assign n50096 = pi20 ? n50095 : n32;
  assign n50097 = pi19 ? n99 : n50096;
  assign n50098 = pi18 ? n50093 : n50097;
  assign n50099 = pi17 ? n20563 : n50098;
  assign n50100 = pi16 ? n44644 : n50099;
  assign n50101 = pi20 ? n20563 : n43010;
  assign n50102 = pi20 ? n31220 : n220;
  assign n50103 = pi19 ? n50101 : n50102;
  assign n50104 = pi18 ? n50103 : n47611;
  assign n50105 = pi17 ? n20563 : n50104;
  assign n50106 = pi16 ? n44644 : n50105;
  assign n50107 = pi15 ? n50100 : n50106;
  assign n50108 = pi21 ? n3759 : n397;
  assign n50109 = pi20 ? n50108 : n32;
  assign n50110 = pi19 ? n99 : n50109;
  assign n50111 = pi18 ? n33285 : n50110;
  assign n50112 = pi17 ? n20563 : n50111;
  assign n50113 = pi16 ? n45243 : n50112;
  assign n50114 = pi21 ? n99 : n21980;
  assign n50115 = pi20 ? n50114 : n32;
  assign n50116 = pi19 ? n26407 : n50115;
  assign n50117 = pi18 ? n33285 : n50116;
  assign n50118 = pi17 ? n20563 : n50117;
  assign n50119 = pi16 ? n45243 : n50118;
  assign n50120 = pi15 ? n50113 : n50119;
  assign n50121 = pi14 ? n50107 : n50120;
  assign n50122 = pi13 ? n50090 : n50121;
  assign n50123 = pi12 ? n50058 : n50122;
  assign n50124 = pi11 ? n50011 : n50123;
  assign n50125 = pi21 ? n204 : n10099;
  assign n50126 = pi20 ? n50125 : n32;
  assign n50127 = pi19 ? n20743 : n50126;
  assign n50128 = pi18 ? n33285 : n50127;
  assign n50129 = pi17 ? n20563 : n50128;
  assign n50130 = pi16 ? n46349 : n50129;
  assign n50131 = pi19 ? n20743 : n21990;
  assign n50132 = pi18 ? n32275 : n50131;
  assign n50133 = pi17 ? n20563 : n50132;
  assign n50134 = pi16 ? n46349 : n50133;
  assign n50135 = pi15 ? n50130 : n50134;
  assign n50136 = pi20 ? n40791 : n43010;
  assign n50137 = pi19 ? n50136 : n31280;
  assign n50138 = pi19 ? n20743 : n22516;
  assign n50139 = pi18 ? n50137 : n50138;
  assign n50140 = pi17 ? n20563 : n50139;
  assign n50141 = pi16 ? n46349 : n50140;
  assign n50142 = pi19 ? n3096 : n22006;
  assign n50143 = pi18 ? n32275 : n50142;
  assign n50144 = pi17 ? n20563 : n50143;
  assign n50145 = pi16 ? n49595 : n50144;
  assign n50146 = pi15 ? n50141 : n50145;
  assign n50147 = pi14 ? n50135 : n50146;
  assign n50148 = pi21 ? n204 : n5758;
  assign n50149 = pi20 ? n50148 : n32;
  assign n50150 = pi19 ? n9795 : n50149;
  assign n50151 = pi18 ? n33299 : n50150;
  assign n50152 = pi17 ? n20563 : n50151;
  assign n50153 = pi16 ? n49595 : n50152;
  assign n50154 = pi19 ? n8765 : n47667;
  assign n50155 = pi18 ? n33299 : n50154;
  assign n50156 = pi17 ? n20563 : n50155;
  assign n50157 = pi16 ? n43664 : n50156;
  assign n50158 = pi15 ? n50153 : n50157;
  assign n50159 = pi21 ? n28649 : n13315;
  assign n50160 = pi20 ? n50159 : n32;
  assign n50161 = pi19 ? n8765 : n50160;
  assign n50162 = pi18 ? n33285 : n50161;
  assign n50163 = pi17 ? n20563 : n50162;
  assign n50164 = pi16 ? n43664 : n50163;
  assign n50165 = pi22 ? n6833 : n233;
  assign n50166 = pi21 ? n50165 : n6416;
  assign n50167 = pi20 ? n50166 : n32;
  assign n50168 = pi19 ? n42722 : n50167;
  assign n50169 = pi18 ? n33285 : n50168;
  assign n50170 = pi17 ? n20563 : n50169;
  assign n50171 = pi16 ? n43664 : n50170;
  assign n50172 = pi15 ? n50164 : n50171;
  assign n50173 = pi14 ? n50158 : n50172;
  assign n50174 = pi13 ? n50147 : n50173;
  assign n50175 = pi21 ? n19386 : n5829;
  assign n50176 = pi20 ? n50175 : n32;
  assign n50177 = pi19 ? n24788 : n50176;
  assign n50178 = pi18 ? n33285 : n50177;
  assign n50179 = pi17 ? n20563 : n50178;
  assign n50180 = pi16 ? n43664 : n50179;
  assign n50181 = pi21 ? n6376 : n5829;
  assign n50182 = pi20 ? n50181 : n32;
  assign n50183 = pi19 ? n7685 : n50182;
  assign n50184 = pi18 ? n33285 : n50183;
  assign n50185 = pi17 ? n20563 : n50184;
  assign n50186 = pi16 ? n44671 : n50185;
  assign n50187 = pi15 ? n50180 : n50186;
  assign n50188 = pi19 ? n24788 : n49185;
  assign n50189 = pi18 ? n33299 : n50188;
  assign n50190 = pi17 ? n20563 : n50189;
  assign n50191 = pi16 ? n43219 : n50190;
  assign n50192 = pi21 ? n11336 : n928;
  assign n50193 = pi20 ? n50192 : n32;
  assign n50194 = pi19 ? n7685 : n50193;
  assign n50195 = pi18 ? n33285 : n50194;
  assign n50196 = pi17 ? n20563 : n50195;
  assign n50197 = pi16 ? n43219 : n50196;
  assign n50198 = pi15 ? n50191 : n50197;
  assign n50199 = pi14 ? n50187 : n50198;
  assign n50200 = pi19 ? n32 : n47747;
  assign n50201 = pi18 ? n32 : n50200;
  assign n50202 = pi17 ? n32 : n50201;
  assign n50203 = pi19 ? n7685 : n12493;
  assign n50204 = pi18 ? n33285 : n50203;
  assign n50205 = pi17 ? n49212 : n50204;
  assign n50206 = pi16 ? n50202 : n50205;
  assign n50207 = pi20 ? n38981 : n40791;
  assign n50208 = pi19 ? n32 : n50207;
  assign n50209 = pi18 ? n32 : n50208;
  assign n50210 = pi17 ? n32 : n50209;
  assign n50211 = pi19 ? n7685 : n18413;
  assign n50212 = pi18 ? n33299 : n50211;
  assign n50213 = pi17 ? n49212 : n50212;
  assign n50214 = pi16 ? n50210 : n50213;
  assign n50215 = pi15 ? n50206 : n50214;
  assign n50216 = pi19 ? n8928 : n47180;
  assign n50217 = pi18 ? n32295 : n50216;
  assign n50218 = pi17 ? n20563 : n50217;
  assign n50219 = pi16 ? n43219 : n50218;
  assign n50220 = pi19 ? n7676 : n12129;
  assign n50221 = pi18 ? n32295 : n50220;
  assign n50222 = pi17 ? n20563 : n50221;
  assign n50223 = pi16 ? n43249 : n50222;
  assign n50224 = pi15 ? n50219 : n50223;
  assign n50225 = pi14 ? n50215 : n50224;
  assign n50226 = pi13 ? n50199 : n50225;
  assign n50227 = pi12 ? n50174 : n50226;
  assign n50228 = pi19 ? n2108 : n11244;
  assign n50229 = pi18 ? n33299 : n50228;
  assign n50230 = pi17 ? n20563 : n50229;
  assign n50231 = pi16 ? n43249 : n50230;
  assign n50232 = pi19 ? n2108 : n10327;
  assign n50233 = pi18 ? n32295 : n50232;
  assign n50234 = pi17 ? n20563 : n50233;
  assign n50235 = pi16 ? n43249 : n50234;
  assign n50236 = pi15 ? n50231 : n50235;
  assign n50237 = pi22 ? n112 : n3944;
  assign n50238 = pi21 ? n37 : n50237;
  assign n50239 = pi20 ? n37 : n50238;
  assign n50240 = pi19 ? n50239 : n8296;
  assign n50241 = pi18 ? n32295 : n50240;
  assign n50242 = pi17 ? n20563 : n50241;
  assign n50243 = pi16 ? n43249 : n50242;
  assign n50244 = pi20 ? n20563 : n36489;
  assign n50245 = pi21 ? n7327 : n10488;
  assign n50246 = pi20 ? n2973 : n50245;
  assign n50247 = pi19 ? n50244 : n50246;
  assign n50248 = pi21 ? n5015 : n767;
  assign n50249 = pi20 ? n22881 : n50248;
  assign n50250 = pi19 ? n50249 : n9483;
  assign n50251 = pi18 ? n50247 : n50250;
  assign n50252 = pi17 ? n20563 : n50251;
  assign n50253 = pi16 ? n44248 : n50252;
  assign n50254 = pi15 ? n50243 : n50253;
  assign n50255 = pi14 ? n50236 : n50254;
  assign n50256 = pi21 ? n3392 : n10488;
  assign n50257 = pi20 ? n37 : n50256;
  assign n50258 = pi19 ? n20563 : n50257;
  assign n50259 = pi21 ? n1476 : n32;
  assign n50260 = pi20 ? n50259 : n32;
  assign n50261 = pi19 ? n32794 : n50260;
  assign n50262 = pi18 ? n50258 : n50261;
  assign n50263 = pi17 ? n20563 : n50262;
  assign n50264 = pi16 ? n44248 : n50263;
  assign n50265 = pi20 ? n20563 : n45016;
  assign n50266 = pi22 ? n20563 : n139;
  assign n50267 = pi21 ? n50266 : n37;
  assign n50268 = pi20 ? n50267 : n37;
  assign n50269 = pi19 ? n50265 : n50268;
  assign n50270 = pi19 ? n32794 : n3211;
  assign n50271 = pi18 ? n50269 : n50270;
  assign n50272 = pi17 ? n20563 : n50271;
  assign n50273 = pi16 ? n43219 : n50272;
  assign n50274 = pi15 ? n50264 : n50273;
  assign n50275 = pi19 ? n47274 : n5831;
  assign n50276 = pi18 ? n33299 : n50275;
  assign n50277 = pi17 ? n20563 : n50276;
  assign n50278 = pi16 ? n43219 : n50277;
  assign n50279 = pi14 ? n50274 : n50278;
  assign n50280 = pi13 ? n50255 : n50279;
  assign n50281 = pi19 ? n43011 : n21611;
  assign n50282 = pi21 ? n685 : n316;
  assign n50283 = pi20 ? n2729 : n50282;
  assign n50284 = pi19 ? n50283 : n2654;
  assign n50285 = pi18 ? n50281 : n50284;
  assign n50286 = pi17 ? n49311 : n50285;
  assign n50287 = pi16 ? n44248 : n50286;
  assign n50288 = pi19 ? n30868 : n99;
  assign n50289 = pi20 ? n2243 : n34537;
  assign n50290 = pi19 ? n50289 : n2654;
  assign n50291 = pi18 ? n50288 : n50290;
  assign n50292 = pi17 ? n30868 : n50291;
  assign n50293 = pi16 ? n50202 : n50292;
  assign n50294 = pi15 ? n50287 : n50293;
  assign n50295 = pi19 ? n32 : n47857;
  assign n50296 = pi18 ? n32 : n50295;
  assign n50297 = pi17 ? n32 : n50296;
  assign n50298 = pi21 ? n45142 : n36798;
  assign n50299 = pi20 ? n50298 : n36798;
  assign n50300 = pi21 ? n36798 : n33792;
  assign n50301 = pi20 ? n50298 : n50300;
  assign n50302 = pi19 ? n50299 : n50301;
  assign n50303 = pi18 ? n36798 : n50302;
  assign n50304 = pi20 ? n46733 : n4665;
  assign n50305 = pi19 ? n33792 : n50304;
  assign n50306 = pi20 ? n282 : n34537;
  assign n50307 = pi19 ? n50306 : n1823;
  assign n50308 = pi18 ? n50305 : n50307;
  assign n50309 = pi17 ? n50303 : n50308;
  assign n50310 = pi16 ? n50297 : n50309;
  assign n50311 = pi20 ? n36798 : n45143;
  assign n50312 = pi19 ? n50311 : n33792;
  assign n50313 = pi18 ? n50312 : n33792;
  assign n50314 = pi21 ? n248 : n397;
  assign n50315 = pi20 ? n139 : n50314;
  assign n50316 = pi19 ? n50315 : n32;
  assign n50317 = pi18 ? n47348 : n50316;
  assign n50318 = pi17 ? n50313 : n50317;
  assign n50319 = pi16 ? n50297 : n50318;
  assign n50320 = pi15 ? n50310 : n50319;
  assign n50321 = pi14 ? n50294 : n50320;
  assign n50322 = pi22 ? n36783 : n36659;
  assign n50323 = pi21 ? n50322 : n36659;
  assign n50324 = pi20 ? n32 : n50323;
  assign n50325 = pi19 ? n32 : n50324;
  assign n50326 = pi18 ? n32 : n50325;
  assign n50327 = pi17 ? n32 : n50326;
  assign n50328 = pi21 ? n335 : n36837;
  assign n50329 = pi20 ? n50328 : n48840;
  assign n50330 = pi19 ? n50329 : n32;
  assign n50331 = pi18 ? n47388 : n50330;
  assign n50332 = pi17 ? n36659 : n50331;
  assign n50333 = pi16 ? n50327 : n50332;
  assign n50334 = pi20 ? n32 : n43198;
  assign n50335 = pi19 ? n32 : n50334;
  assign n50336 = pi18 ? n32 : n50335;
  assign n50337 = pi17 ? n32 : n50336;
  assign n50338 = pi22 ? n43198 : n36659;
  assign n50339 = pi23 ? n36659 : n43198;
  assign n50340 = pi22 ? n36659 : n50339;
  assign n50341 = pi21 ? n50338 : n50340;
  assign n50342 = pi21 ? n50338 : n36659;
  assign n50343 = pi20 ? n50341 : n50342;
  assign n50344 = pi19 ? n50343 : n36659;
  assign n50345 = pi18 ? n50344 : n36659;
  assign n50346 = pi22 ? n316 : n19696;
  assign n50347 = pi21 ? n316 : n50346;
  assign n50348 = pi20 ? n335 : n50347;
  assign n50349 = pi19 ? n50348 : n32;
  assign n50350 = pi18 ? n47388 : n50349;
  assign n50351 = pi17 ? n50345 : n50350;
  assign n50352 = pi16 ? n50337 : n50351;
  assign n50353 = pi15 ? n50333 : n50352;
  assign n50354 = pi21 ? n36798 : n38901;
  assign n50355 = pi20 ? n39973 : n50354;
  assign n50356 = pi19 ? n50355 : n36781;
  assign n50357 = pi18 ? n50356 : n36781;
  assign n50358 = pi23 ? n157 : n363;
  assign n50359 = pi22 ? n157 : n50358;
  assign n50360 = pi21 ? n363 : n50359;
  assign n50361 = pi20 ? n40442 : n50360;
  assign n50362 = pi19 ? n36781 : n50361;
  assign n50363 = pi21 ? n6132 : n3523;
  assign n50364 = pi20 ? n157 : n50363;
  assign n50365 = pi19 ? n50364 : n32;
  assign n50366 = pi18 ? n50362 : n50365;
  assign n50367 = pi17 ? n50357 : n50366;
  assign n50368 = pi16 ? n50297 : n50367;
  assign n50369 = pi19 ? n46282 : n36781;
  assign n50370 = pi18 ? n50369 : n36781;
  assign n50371 = pi20 ? n42170 : n38902;
  assign n50372 = pi19 ? n50371 : n45691;
  assign n50373 = pi21 ? n10021 : n3523;
  assign n50374 = pi20 ? n157 : n50373;
  assign n50375 = pi19 ? n50374 : n32;
  assign n50376 = pi18 ? n50372 : n50375;
  assign n50377 = pi17 ? n50370 : n50376;
  assign n50378 = pi16 ? n50337 : n50377;
  assign n50379 = pi15 ? n50368 : n50378;
  assign n50380 = pi14 ? n50353 : n50379;
  assign n50381 = pi13 ? n50321 : n50380;
  assign n50382 = pi12 ? n50280 : n50381;
  assign n50383 = pi11 ? n50227 : n50382;
  assign n50384 = pi10 ? n50124 : n50383;
  assign n50385 = pi09 ? n49908 : n50384;
  assign n50386 = pi18 ? n43683 : n20563;
  assign n50387 = pi17 ? n50386 : n49890;
  assign n50388 = pi16 ? n32 : n50387;
  assign n50389 = pi15 ? n32 : n50388;
  assign n50390 = pi18 ? n44686 : n20563;
  assign n50391 = pi17 ? n50390 : n49897;
  assign n50392 = pi16 ? n32 : n50391;
  assign n50393 = pi18 ? n43217 : n20563;
  assign n50394 = pi17 ? n50393 : n49897;
  assign n50395 = pi16 ? n32 : n50394;
  assign n50396 = pi15 ? n50392 : n50395;
  assign n50397 = pi14 ? n50389 : n50396;
  assign n50398 = pi13 ? n32 : n50397;
  assign n50399 = pi12 ? n32 : n50398;
  assign n50400 = pi11 ? n32 : n50399;
  assign n50401 = pi10 ? n32 : n50400;
  assign n50402 = pi22 ? n7024 : n5631;
  assign n50403 = pi21 ? n50402 : n32;
  assign n50404 = pi20 ? n37 : n50403;
  assign n50405 = pi19 ? n37 : n50404;
  assign n50406 = pi18 ? n20563 : n50405;
  assign n50407 = pi17 ? n49888 : n50406;
  assign n50408 = pi16 ? n32 : n50407;
  assign n50409 = pi17 ? n49440 : n49922;
  assign n50410 = pi16 ? n32 : n50409;
  assign n50411 = pi15 ? n50408 : n50410;
  assign n50412 = pi20 ? n3086 : n33886;
  assign n50413 = pi19 ? n32898 : n50412;
  assign n50414 = pi18 ? n20563 : n50413;
  assign n50415 = pi17 ? n49448 : n50414;
  assign n50416 = pi16 ? n32 : n50415;
  assign n50417 = pi22 ? n295 : n32;
  assign n50418 = pi21 ? n50417 : n32;
  assign n50419 = pi20 ? n37 : n50418;
  assign n50420 = pi19 ? n32898 : n50419;
  assign n50421 = pi18 ? n20563 : n50420;
  assign n50422 = pi17 ? n49451 : n50421;
  assign n50423 = pi16 ? n32 : n50422;
  assign n50424 = pi15 ? n50416 : n50423;
  assign n50425 = pi14 ? n50411 : n50424;
  assign n50426 = pi18 ? n42193 : n20563;
  assign n50427 = pi22 ? n583 : n625;
  assign n50428 = pi21 ? n50427 : n32;
  assign n50429 = pi20 ? n37 : n50428;
  assign n50430 = pi19 ? n31267 : n50429;
  assign n50431 = pi18 ? n20563 : n50430;
  assign n50432 = pi17 ? n50426 : n50431;
  assign n50433 = pi16 ? n32 : n50432;
  assign n50434 = pi21 ? n626 : n32;
  assign n50435 = pi20 ? n37 : n50434;
  assign n50436 = pi19 ? n30097 : n50435;
  assign n50437 = pi18 ? n48972 : n50436;
  assign n50438 = pi17 ? n48904 : n50437;
  assign n50439 = pi16 ? n32 : n50438;
  assign n50440 = pi15 ? n50433 : n50439;
  assign n50441 = pi19 ? n49951 : n50435;
  assign n50442 = pi18 ? n20563 : n50441;
  assign n50443 = pi17 ? n48466 : n50442;
  assign n50444 = pi16 ? n32 : n50443;
  assign n50445 = pi20 ? n649 : n50434;
  assign n50446 = pi19 ? n32871 : n50445;
  assign n50447 = pi18 ? n20563 : n50446;
  assign n50448 = pi17 ? n48466 : n50447;
  assign n50449 = pi16 ? n32 : n50448;
  assign n50450 = pi15 ? n50444 : n50449;
  assign n50451 = pi14 ? n50440 : n50450;
  assign n50452 = pi13 ? n50425 : n50451;
  assign n50453 = pi20 ? n577 : n18928;
  assign n50454 = pi19 ? n31267 : n50453;
  assign n50455 = pi18 ? n20563 : n50454;
  assign n50456 = pi17 ? n48469 : n50455;
  assign n50457 = pi16 ? n32 : n50456;
  assign n50458 = pi22 ? n10400 : n688;
  assign n50459 = pi21 ? n50458 : n32;
  assign n50460 = pi20 ? n649 : n50459;
  assign n50461 = pi19 ? n30097 : n50460;
  assign n50462 = pi18 ? n48972 : n50461;
  assign n50463 = pi17 ? n49485 : n50462;
  assign n50464 = pi16 ? n32 : n50463;
  assign n50465 = pi15 ? n50457 : n50464;
  assign n50466 = pi22 ? n10400 : n706;
  assign n50467 = pi21 ? n50466 : n32;
  assign n50468 = pi20 ? n649 : n50467;
  assign n50469 = pi19 ? n37 : n50468;
  assign n50470 = pi18 ? n34869 : n50469;
  assign n50471 = pi17 ? n47929 : n50470;
  assign n50472 = pi16 ? n32 : n50471;
  assign n50473 = pi20 ? n649 : n3937;
  assign n50474 = pi19 ? n33949 : n50473;
  assign n50475 = pi18 ? n20563 : n50474;
  assign n50476 = pi17 ? n48488 : n50475;
  assign n50477 = pi16 ? n32 : n50476;
  assign n50478 = pi15 ? n50472 : n50477;
  assign n50479 = pi14 ? n50465 : n50478;
  assign n50480 = pi22 ? n18448 : n32;
  assign n50481 = pi21 ? n50480 : n32;
  assign n50482 = pi20 ? n3393 : n50481;
  assign n50483 = pi19 ? n37 : n50482;
  assign n50484 = pi18 ? n20563 : n50483;
  assign n50485 = pi17 ? n48488 : n50484;
  assign n50486 = pi16 ? n32 : n50485;
  assign n50487 = pi17 ? n47451 : n49997;
  assign n50488 = pi16 ? n32 : n50487;
  assign n50489 = pi15 ? n50486 : n50488;
  assign n50490 = pi17 ? n46302 : n49997;
  assign n50491 = pi16 ? n32 : n50490;
  assign n50492 = pi17 ? n46832 : n50005;
  assign n50493 = pi16 ? n32 : n50492;
  assign n50494 = pi15 ? n50491 : n50493;
  assign n50495 = pi14 ? n50489 : n50494;
  assign n50496 = pi13 ? n50479 : n50495;
  assign n50497 = pi12 ? n50452 : n50496;
  assign n50498 = pi20 ? n19091 : n3210;
  assign n50499 = pi19 ? n32933 : n50498;
  assign n50500 = pi18 ? n34865 : n50499;
  assign n50501 = pi17 ? n47964 : n50500;
  assign n50502 = pi16 ? n32 : n50501;
  assign n50503 = pi21 ? n37 : n30195;
  assign n50504 = pi20 ? n20563 : n50503;
  assign n50505 = pi19 ? n20563 : n50504;
  assign n50506 = pi18 ? n50505 : n50019;
  assign n50507 = pi17 ? n47964 : n50506;
  assign n50508 = pi16 ? n32 : n50507;
  assign n50509 = pi15 ? n50502 : n50508;
  assign n50510 = pi21 ? n37 : n31924;
  assign n50511 = pi20 ? n20563 : n50510;
  assign n50512 = pi19 ? n20563 : n50511;
  assign n50513 = pi18 ? n50512 : n50027;
  assign n50514 = pi17 ? n46839 : n50513;
  assign n50515 = pi16 ? n32 : n50514;
  assign n50516 = pi20 ? n3393 : n2638;
  assign n50517 = pi19 ? n37 : n50516;
  assign n50518 = pi18 ? n39073 : n50517;
  assign n50519 = pi17 ? n45707 : n50518;
  assign n50520 = pi16 ? n32 : n50519;
  assign n50521 = pi15 ? n50515 : n50520;
  assign n50522 = pi14 ? n50509 : n50521;
  assign n50523 = pi17 ? n46859 : n50037;
  assign n50524 = pi16 ? n32 : n50523;
  assign n50525 = pi18 ? n33823 : n50041;
  assign n50526 = pi17 ? n45715 : n50525;
  assign n50527 = pi16 ? n32 : n50526;
  assign n50528 = pi15 ? n50524 : n50527;
  assign n50529 = pi18 ? n40228 : n50047;
  assign n50530 = pi17 ? n45715 : n50529;
  assign n50531 = pi16 ? n32 : n50530;
  assign n50532 = pi18 ? n45413 : n20563;
  assign n50533 = pi18 ? n33828 : n50052;
  assign n50534 = pi17 ? n50532 : n50533;
  assign n50535 = pi16 ? n32 : n50534;
  assign n50536 = pi15 ? n50531 : n50535;
  assign n50537 = pi14 ? n50528 : n50536;
  assign n50538 = pi13 ? n50522 : n50537;
  assign n50539 = pi20 ? n382 : n10011;
  assign n50540 = pi19 ? n37 : n50539;
  assign n50541 = pi18 ? n40067 : n50540;
  assign n50542 = pi17 ? n46312 : n50541;
  assign n50543 = pi16 ? n32 : n50542;
  assign n50544 = pi20 ? n31913 : n5077;
  assign n50545 = pi19 ? n20563 : n50544;
  assign n50546 = pi20 ? n24957 : n2653;
  assign n50547 = pi19 ? n18853 : n50546;
  assign n50548 = pi18 ? n50545 : n50547;
  assign n50549 = pi17 ? n20563 : n50548;
  assign n50550 = pi16 ? n32 : n50549;
  assign n50551 = pi15 ? n50543 : n50550;
  assign n50552 = pi19 ? n21611 : n50546;
  assign n50553 = pi18 ? n33260 : n50552;
  assign n50554 = pi17 ? n20563 : n50553;
  assign n50555 = pi16 ? n46326 : n50554;
  assign n50556 = pi19 ? n99 : n50077;
  assign n50557 = pi18 ? n32275 : n50556;
  assign n50558 = pi17 ? n20563 : n50557;
  assign n50559 = pi16 ? n46326 : n50558;
  assign n50560 = pi15 ? n50555 : n50559;
  assign n50561 = pi14 ? n50551 : n50560;
  assign n50562 = pi20 ? n32313 : n3039;
  assign n50563 = pi19 ? n50091 : n50562;
  assign n50564 = pi20 ? n50083 : n32;
  assign n50565 = pi19 ? n99 : n50564;
  assign n50566 = pi18 ? n50563 : n50565;
  assign n50567 = pi17 ? n20563 : n50566;
  assign n50568 = pi16 ? n46326 : n50567;
  assign n50569 = pi20 ? n32313 : n220;
  assign n50570 = pi19 ? n50101 : n50569;
  assign n50571 = pi18 ? n50570 : n48619;
  assign n50572 = pi17 ? n20563 : n50571;
  assign n50573 = pi16 ? n46326 : n50572;
  assign n50574 = pi15 ? n50568 : n50573;
  assign n50575 = pi20 ? n41893 : n32;
  assign n50576 = pi19 ? n99 : n50575;
  assign n50577 = pi18 ? n32288 : n50576;
  assign n50578 = pi17 ? n20563 : n50577;
  assign n50579 = pi16 ? n45740 : n50578;
  assign n50580 = pi21 ? n99 : n7637;
  assign n50581 = pi20 ? n50580 : n32;
  assign n50582 = pi19 ? n26407 : n50581;
  assign n50583 = pi18 ? n32288 : n50582;
  assign n50584 = pi17 ? n20563 : n50583;
  assign n50585 = pi16 ? n46885 : n50584;
  assign n50586 = pi15 ? n50579 : n50585;
  assign n50587 = pi14 ? n50574 : n50586;
  assign n50588 = pi13 ? n50561 : n50587;
  assign n50589 = pi12 ? n50538 : n50588;
  assign n50590 = pi11 ? n50497 : n50589;
  assign n50591 = pi20 ? n36572 : n32;
  assign n50592 = pi19 ? n20743 : n50591;
  assign n50593 = pi18 ? n33285 : n50592;
  assign n50594 = pi17 ? n20563 : n50593;
  assign n50595 = pi16 ? n46885 : n50594;
  assign n50596 = pi22 ? n37 : n30869;
  assign n50597 = pi21 ? n20563 : n50596;
  assign n50598 = pi20 ? n50597 : n37;
  assign n50599 = pi19 ? n20563 : n50598;
  assign n50600 = pi21 ? n204 : n11235;
  assign n50601 = pi20 ? n50600 : n32;
  assign n50602 = pi19 ? n20743 : n50601;
  assign n50603 = pi18 ? n50599 : n50602;
  assign n50604 = pi17 ? n20563 : n50603;
  assign n50605 = pi16 ? n46885 : n50604;
  assign n50606 = pi15 ? n50595 : n50605;
  assign n50607 = pi18 ? n50137 : n50131;
  assign n50608 = pi17 ? n20563 : n50607;
  assign n50609 = pi16 ? n46885 : n50608;
  assign n50610 = pi16 ? n44653 : n50144;
  assign n50611 = pi15 ? n50609 : n50610;
  assign n50612 = pi14 ? n50606 : n50611;
  assign n50613 = pi21 ? n204 : n13280;
  assign n50614 = pi20 ? n50613 : n32;
  assign n50615 = pi19 ? n9795 : n50614;
  assign n50616 = pi18 ? n33858 : n50615;
  assign n50617 = pi17 ? n20563 : n50616;
  assign n50618 = pi16 ? n44653 : n50617;
  assign n50619 = pi19 ? n8765 : n20124;
  assign n50620 = pi18 ? n33858 : n50619;
  assign n50621 = pi17 ? n20563 : n50620;
  assign n50622 = pi16 ? n44223 : n50621;
  assign n50623 = pi15 ? n50618 : n50622;
  assign n50624 = pi18 ? n32288 : n49682;
  assign n50625 = pi17 ? n20563 : n50624;
  assign n50626 = pi16 ? n44223 : n50625;
  assign n50627 = pi21 ? n50165 : n4109;
  assign n50628 = pi20 ? n50627 : n32;
  assign n50629 = pi19 ? n42722 : n50628;
  assign n50630 = pi18 ? n32288 : n50629;
  assign n50631 = pi17 ? n20563 : n50630;
  assign n50632 = pi16 ? n44223 : n50631;
  assign n50633 = pi15 ? n50626 : n50632;
  assign n50634 = pi14 ? n50623 : n50633;
  assign n50635 = pi13 ? n50612 : n50634;
  assign n50636 = pi21 ? n31294 : n36618;
  assign n50637 = pi20 ? n50636 : n37;
  assign n50638 = pi19 ? n20563 : n50637;
  assign n50639 = pi21 ? n19386 : n33622;
  assign n50640 = pi20 ? n50639 : n32;
  assign n50641 = pi19 ? n24788 : n50640;
  assign n50642 = pi18 ? n50638 : n50641;
  assign n50643 = pi17 ? n20563 : n50642;
  assign n50644 = pi16 ? n44223 : n50643;
  assign n50645 = pi21 ? n6376 : n760;
  assign n50646 = pi20 ? n50645 : n32;
  assign n50647 = pi19 ? n7685 : n50646;
  assign n50648 = pi18 ? n33285 : n50647;
  assign n50649 = pi17 ? n20563 : n50648;
  assign n50650 = pi16 ? n44223 : n50649;
  assign n50651 = pi15 ? n50644 : n50650;
  assign n50652 = pi21 ? n6376 : n2835;
  assign n50653 = pi20 ? n50652 : n32;
  assign n50654 = pi19 ? n24788 : n50653;
  assign n50655 = pi18 ? n38549 : n50654;
  assign n50656 = pi17 ? n20563 : n50655;
  assign n50657 = pi16 ? n43664 : n50656;
  assign n50658 = pi21 ? n11336 : n882;
  assign n50659 = pi20 ? n50658 : n32;
  assign n50660 = pi19 ? n7685 : n50659;
  assign n50661 = pi18 ? n33285 : n50660;
  assign n50662 = pi17 ? n20563 : n50661;
  assign n50663 = pi16 ? n46349 : n50662;
  assign n50664 = pi15 ? n50657 : n50663;
  assign n50665 = pi14 ? n50651 : n50664;
  assign n50666 = pi22 ? n32 : n40342;
  assign n50667 = pi21 ? n50666 : n30868;
  assign n50668 = pi20 ? n32 : n50667;
  assign n50669 = pi19 ? n32 : n50668;
  assign n50670 = pi18 ? n32 : n50669;
  assign n50671 = pi17 ? n32 : n50670;
  assign n50672 = pi19 ? n7685 : n12102;
  assign n50673 = pi18 ? n33285 : n50672;
  assign n50674 = pi17 ? n49212 : n50673;
  assign n50675 = pi16 ? n50671 : n50674;
  assign n50676 = pi21 ? n39394 : n30868;
  assign n50677 = pi20 ? n32 : n50676;
  assign n50678 = pi19 ? n32 : n50677;
  assign n50679 = pi18 ? n32 : n50678;
  assign n50680 = pi17 ? n32 : n50679;
  assign n50681 = pi19 ? n7685 : n20238;
  assign n50682 = pi18 ? n38549 : n50681;
  assign n50683 = pi17 ? n49212 : n50682;
  assign n50684 = pi16 ? n50680 : n50683;
  assign n50685 = pi15 ? n50675 : n50684;
  assign n50686 = pi18 ? n42358 : n50216;
  assign n50687 = pi17 ? n20563 : n50686;
  assign n50688 = pi16 ? n49595 : n50687;
  assign n50689 = pi19 ? n7676 : n11696;
  assign n50690 = pi18 ? n42358 : n50689;
  assign n50691 = pi17 ? n20563 : n50690;
  assign n50692 = pi16 ? n43219 : n50691;
  assign n50693 = pi15 ? n50688 : n50692;
  assign n50694 = pi14 ? n50685 : n50693;
  assign n50695 = pi13 ? n50665 : n50694;
  assign n50696 = pi12 ? n50635 : n50695;
  assign n50697 = pi19 ? n2108 : n11696;
  assign n50698 = pi18 ? n33299 : n50697;
  assign n50699 = pi17 ? n20563 : n50698;
  assign n50700 = pi16 ? n43675 : n50699;
  assign n50701 = pi18 ? n42358 : n50232;
  assign n50702 = pi17 ? n20563 : n50701;
  assign n50703 = pi16 ? n43675 : n50702;
  assign n50704 = pi15 ? n50700 : n50703;
  assign n50705 = pi18 ? n47689 : n50240;
  assign n50706 = pi17 ? n20563 : n50705;
  assign n50707 = pi16 ? n43675 : n50706;
  assign n50708 = pi22 ? n30867 : n99;
  assign n50709 = pi21 ? n50708 : n37;
  assign n50710 = pi21 ? n2175 : n10488;
  assign n50711 = pi20 ? n50709 : n50710;
  assign n50712 = pi19 ? n50244 : n50711;
  assign n50713 = pi18 ? n50712 : n50250;
  assign n50714 = pi17 ? n20563 : n50713;
  assign n50715 = pi16 ? n44671 : n50714;
  assign n50716 = pi15 ? n50707 : n50715;
  assign n50717 = pi14 ? n50704 : n50716;
  assign n50718 = pi20 ? n31298 : n50256;
  assign n50719 = pi19 ? n20563 : n50718;
  assign n50720 = pi19 ? n32794 : n9483;
  assign n50721 = pi18 ? n50719 : n50720;
  assign n50722 = pi17 ? n20563 : n50721;
  assign n50723 = pi16 ? n44671 : n50722;
  assign n50724 = pi20 ? n50267 : n13147;
  assign n50725 = pi19 ? n50265 : n50724;
  assign n50726 = pi18 ? n50725 : n50270;
  assign n50727 = pi17 ? n20563 : n50726;
  assign n50728 = pi16 ? n44671 : n50727;
  assign n50729 = pi15 ? n50723 : n50728;
  assign n50730 = pi21 ? n37805 : n40913;
  assign n50731 = pi20 ? n32 : n50730;
  assign n50732 = pi19 ? n32 : n50731;
  assign n50733 = pi18 ? n32 : n50732;
  assign n50734 = pi17 ? n32 : n50733;
  assign n50735 = pi21 ? n46116 : n20563;
  assign n50736 = pi21 ? n40913 : n20563;
  assign n50737 = pi20 ? n50735 : n50736;
  assign n50738 = pi19 ? n50737 : n20563;
  assign n50739 = pi18 ? n50738 : n20563;
  assign n50740 = pi19 ? n47274 : n7050;
  assign n50741 = pi18 ? n33858 : n50740;
  assign n50742 = pi17 ? n50739 : n50741;
  assign n50743 = pi16 ? n50734 : n50742;
  assign n50744 = pi17 ? n20563 : n50741;
  assign n50745 = pi16 ? n49595 : n50744;
  assign n50746 = pi15 ? n50743 : n50745;
  assign n50747 = pi14 ? n50729 : n50746;
  assign n50748 = pi13 ? n50717 : n50747;
  assign n50749 = pi21 ? n31200 : n99;
  assign n50750 = pi20 ? n50749 : n99;
  assign n50751 = pi19 ? n43011 : n50750;
  assign n50752 = pi19 ? n50283 : n48320;
  assign n50753 = pi18 ? n50751 : n50752;
  assign n50754 = pi17 ? n49311 : n50753;
  assign n50755 = pi16 ? n49595 : n50754;
  assign n50756 = pi19 ? n32 : n48255;
  assign n50757 = pi18 ? n32 : n50756;
  assign n50758 = pi17 ? n32 : n50757;
  assign n50759 = pi22 ? n37240 : n99;
  assign n50760 = pi21 ? n50759 : n99;
  assign n50761 = pi20 ? n50760 : n99;
  assign n50762 = pi19 ? n30868 : n50761;
  assign n50763 = pi18 ? n50762 : n50290;
  assign n50764 = pi17 ? n30868 : n50763;
  assign n50765 = pi16 ? n50758 : n50764;
  assign n50766 = pi15 ? n50755 : n50765;
  assign n50767 = pi22 ? n32 : n36831;
  assign n50768 = pi21 ? n50767 : n36798;
  assign n50769 = pi20 ? n32 : n50768;
  assign n50770 = pi19 ? n32 : n50769;
  assign n50771 = pi18 ? n32 : n50770;
  assign n50772 = pi17 ? n32 : n50771;
  assign n50773 = pi21 ? n44143 : n139;
  assign n50774 = pi20 ? n50773 : n248;
  assign n50775 = pi19 ? n33792 : n50774;
  assign n50776 = pi18 ? n50775 : n50307;
  assign n50777 = pi17 ? n50303 : n50776;
  assign n50778 = pi16 ? n50772 : n50777;
  assign n50779 = pi20 ? n139 : n47371;
  assign n50780 = pi19 ? n50779 : n32;
  assign n50781 = pi18 ? n47348 : n50780;
  assign n50782 = pi17 ? n50313 : n50781;
  assign n50783 = pi16 ? n50772 : n50782;
  assign n50784 = pi15 ? n50778 : n50783;
  assign n50785 = pi14 ? n50766 : n50784;
  assign n50786 = pi22 ? n32 : n49843;
  assign n50787 = pi21 ? n50786 : n43198;
  assign n50788 = pi20 ? n32 : n50787;
  assign n50789 = pi19 ? n32 : n50788;
  assign n50790 = pi18 ? n32 : n50789;
  assign n50791 = pi17 ? n32 : n50790;
  assign n50792 = pi23 ? n43198 : n36659;
  assign n50793 = pi22 ? n50792 : n50339;
  assign n50794 = pi21 ? n50793 : n36659;
  assign n50795 = pi22 ? n36659 : n43198;
  assign n50796 = pi22 ? n50792 : n36659;
  assign n50797 = pi21 ? n50795 : n50796;
  assign n50798 = pi20 ? n50794 : n50797;
  assign n50799 = pi19 ? n50798 : n36659;
  assign n50800 = pi18 ? n50799 : n36659;
  assign n50801 = pi22 ? n36659 : n38926;
  assign n50802 = pi21 ? n50801 : n335;
  assign n50803 = pi20 ? n50802 : n335;
  assign n50804 = pi19 ? n36659 : n50803;
  assign n50805 = pi20 ? n50328 : n9752;
  assign n50806 = pi19 ? n50805 : n32;
  assign n50807 = pi18 ? n50804 : n50806;
  assign n50808 = pi17 ? n50800 : n50807;
  assign n50809 = pi16 ? n50791 : n50808;
  assign n50810 = pi21 ? n32 : n43198;
  assign n50811 = pi20 ? n32 : n50810;
  assign n50812 = pi19 ? n32 : n50811;
  assign n50813 = pi18 ? n32 : n50812;
  assign n50814 = pi17 ? n32 : n50813;
  assign n50815 = pi21 ? n50796 : n36659;
  assign n50816 = pi20 ? n50342 : n50815;
  assign n50817 = pi19 ? n50816 : n36659;
  assign n50818 = pi18 ? n50817 : n36659;
  assign n50819 = pi18 ? n50804 : n50349;
  assign n50820 = pi17 ? n50818 : n50819;
  assign n50821 = pi16 ? n50814 : n50820;
  assign n50822 = pi15 ? n50809 : n50821;
  assign n50823 = pi18 ? n32 : n45656;
  assign n50824 = pi17 ? n32 : n50823;
  assign n50825 = pi22 ? n36781 : n40004;
  assign n50826 = pi21 ? n50825 : n363;
  assign n50827 = pi20 ? n50826 : n34841;
  assign n50828 = pi19 ? n36781 : n50827;
  assign n50829 = pi21 ? n6132 : n5178;
  assign n50830 = pi20 ? n157 : n50829;
  assign n50831 = pi19 ? n50830 : n32;
  assign n50832 = pi18 ? n50828 : n50831;
  assign n50833 = pi17 ? n50357 : n50832;
  assign n50834 = pi16 ? n50824 : n50833;
  assign n50835 = pi19 ? n32 : n48437;
  assign n50836 = pi18 ? n32 : n50835;
  assign n50837 = pi17 ? n32 : n50836;
  assign n50838 = pi21 ? n36798 : n48878;
  assign n50839 = pi20 ? n50838 : n157;
  assign n50840 = pi19 ? n50371 : n50839;
  assign n50841 = pi18 ? n50840 : n50375;
  assign n50842 = pi17 ? n50370 : n50841;
  assign n50843 = pi16 ? n50837 : n50842;
  assign n50844 = pi15 ? n50834 : n50843;
  assign n50845 = pi14 ? n50822 : n50844;
  assign n50846 = pi13 ? n50785 : n50845;
  assign n50847 = pi12 ? n50748 : n50846;
  assign n50848 = pi11 ? n50696 : n50847;
  assign n50849 = pi10 ? n50590 : n50848;
  assign n50850 = pi09 ? n50401 : n50849;
  assign n50851 = pi08 ? n50385 : n50850;
  assign n50852 = pi07 ? n49887 : n50851;
  assign n50853 = pi06 ? n48896 : n50852;
  assign n50854 = pi20 ? n31220 : n48905;
  assign n50855 = pi19 ? n50854 : n31221;
  assign n50856 = pi21 ? n12243 : n32;
  assign n50857 = pi20 ? n37 : n50856;
  assign n50858 = pi19 ? n37 : n50857;
  assign n50859 = pi18 ? n50855 : n50858;
  assign n50860 = pi17 ? n39456 : n50859;
  assign n50861 = pi16 ? n32 : n50860;
  assign n50862 = pi15 ? n32 : n50861;
  assign n50863 = pi20 ? n31266 : n20563;
  assign n50864 = pi19 ? n50863 : n32898;
  assign n50865 = pi20 ? n3086 : n50856;
  assign n50866 = pi19 ? n37 : n50865;
  assign n50867 = pi18 ? n50864 : n50866;
  assign n50868 = pi17 ? n34859 : n50867;
  assign n50869 = pi16 ? n32 : n50868;
  assign n50870 = pi22 ? n139 : n23268;
  assign n50871 = pi21 ? n50870 : n32;
  assign n50872 = pi20 ? n37 : n50871;
  assign n50873 = pi19 ? n37 : n50872;
  assign n50874 = pi18 ? n34295 : n50873;
  assign n50875 = pi17 ? n35764 : n50874;
  assign n50876 = pi16 ? n32 : n50875;
  assign n50877 = pi15 ? n50869 : n50876;
  assign n50878 = pi14 ? n50862 : n50877;
  assign n50879 = pi13 ? n32 : n50878;
  assign n50880 = pi12 ? n32 : n50879;
  assign n50881 = pi11 ? n32 : n50880;
  assign n50882 = pi10 ? n32 : n50881;
  assign n50883 = pi20 ? n37 : n31266;
  assign n50884 = pi22 ? n37 : n46851;
  assign n50885 = pi21 ? n50884 : n32;
  assign n50886 = pi20 ? n3086 : n50885;
  assign n50887 = pi19 ? n50883 : n50886;
  assign n50888 = pi18 ? n34258 : n50887;
  assign n50889 = pi17 ? n49888 : n50888;
  assign n50890 = pi16 ? n32 : n50889;
  assign n50891 = pi21 ? n42702 : n32;
  assign n50892 = pi20 ? n13121 : n50891;
  assign n50893 = pi19 ? n50883 : n50892;
  assign n50894 = pi18 ? n34869 : n50893;
  assign n50895 = pi17 ? n49888 : n50894;
  assign n50896 = pi16 ? n32 : n50895;
  assign n50897 = pi15 ? n50890 : n50896;
  assign n50898 = pi22 ? n37 : n2468;
  assign n50899 = pi21 ? n50898 : n32;
  assign n50900 = pi20 ? n8742 : n50899;
  assign n50901 = pi19 ? n37 : n50900;
  assign n50902 = pi18 ? n34295 : n50901;
  assign n50903 = pi17 ? n49894 : n50902;
  assign n50904 = pi16 ? n32 : n50903;
  assign n50905 = pi18 ? n43226 : n20563;
  assign n50906 = pi20 ? n31220 : n20563;
  assign n50907 = pi19 ? n50906 : n32348;
  assign n50908 = pi22 ? n112 : n2468;
  assign n50909 = pi21 ? n50908 : n32;
  assign n50910 = pi20 ? n37 : n50909;
  assign n50911 = pi19 ? n37 : n50910;
  assign n50912 = pi18 ? n50907 : n50911;
  assign n50913 = pi17 ? n50905 : n50912;
  assign n50914 = pi16 ? n32 : n50913;
  assign n50915 = pi15 ? n50904 : n50914;
  assign n50916 = pi14 ? n50897 : n50915;
  assign n50917 = pi20 ? n37 : n18895;
  assign n50918 = pi19 ? n37 : n50917;
  assign n50919 = pi18 ? n34295 : n50918;
  assign n50920 = pi17 ? n49440 : n50919;
  assign n50921 = pi16 ? n32 : n50920;
  assign n50922 = pi19 ? n37 : n50435;
  assign n50923 = pi18 ? n34869 : n50922;
  assign n50924 = pi17 ? n49448 : n50923;
  assign n50925 = pi16 ? n32 : n50924;
  assign n50926 = pi15 ? n50921 : n50925;
  assign n50927 = pi20 ? n48905 : n30096;
  assign n50928 = pi19 ? n50927 : n50435;
  assign n50929 = pi18 ? n20563 : n50928;
  assign n50930 = pi17 ? n48904 : n50929;
  assign n50931 = pi16 ? n32 : n50930;
  assign n50932 = pi20 ? n48905 : n31220;
  assign n50933 = pi19 ? n50932 : n50445;
  assign n50934 = pi18 ? n20563 : n50933;
  assign n50935 = pi17 ? n48904 : n50934;
  assign n50936 = pi16 ? n32 : n50935;
  assign n50937 = pi15 ? n50931 : n50936;
  assign n50938 = pi14 ? n50926 : n50937;
  assign n50939 = pi13 ? n50916 : n50938;
  assign n50940 = pi20 ? n3299 : n18928;
  assign n50941 = pi19 ? n32898 : n50940;
  assign n50942 = pi18 ? n20563 : n50941;
  assign n50943 = pi17 ? n48912 : n50942;
  assign n50944 = pi16 ? n32 : n50943;
  assign n50945 = pi20 ? n649 : n22333;
  assign n50946 = pi19 ? n32348 : n50945;
  assign n50947 = pi18 ? n20563 : n50946;
  assign n50948 = pi17 ? n49938 : n50947;
  assign n50949 = pi16 ? n32 : n50948;
  assign n50950 = pi15 ? n50944 : n50949;
  assign n50951 = pi20 ? n649 : n25406;
  assign n50952 = pi19 ? n31280 : n50951;
  assign n50953 = pi18 ? n20563 : n50952;
  assign n50954 = pi17 ? n48466 : n50953;
  assign n50955 = pi16 ? n32 : n50954;
  assign n50956 = pi21 ? n37 : n7986;
  assign n50957 = pi20 ? n50956 : n34390;
  assign n50958 = pi19 ? n31267 : n50957;
  assign n50959 = pi18 ? n20563 : n50958;
  assign n50960 = pi17 ? n47929 : n50959;
  assign n50961 = pi16 ? n32 : n50960;
  assign n50962 = pi15 ? n50955 : n50961;
  assign n50963 = pi14 ? n50950 : n50962;
  assign n50964 = pi20 ? n37 : n18971;
  assign n50965 = pi19 ? n32348 : n50964;
  assign n50966 = pi18 ? n20563 : n50965;
  assign n50967 = pi17 ? n47929 : n50966;
  assign n50968 = pi16 ? n32 : n50967;
  assign n50969 = pi21 ? n43816 : n32;
  assign n50970 = pi20 ? n37 : n50969;
  assign n50971 = pi19 ? n32348 : n50970;
  assign n50972 = pi18 ? n20563 : n50971;
  assign n50973 = pi17 ? n47935 : n50972;
  assign n50974 = pi16 ? n32 : n50973;
  assign n50975 = pi15 ? n50968 : n50974;
  assign n50976 = pi20 ? n37 : n8295;
  assign n50977 = pi19 ? n31267 : n50976;
  assign n50978 = pi18 ? n20563 : n50977;
  assign n50979 = pi17 ? n47947 : n50978;
  assign n50980 = pi16 ? n32 : n50979;
  assign n50981 = pi20 ? n3393 : n8295;
  assign n50982 = pi19 ? n31280 : n50981;
  assign n50983 = pi18 ? n20563 : n50982;
  assign n50984 = pi17 ? n48949 : n50983;
  assign n50985 = pi16 ? n32 : n50984;
  assign n50986 = pi15 ? n50980 : n50985;
  assign n50987 = pi14 ? n50975 : n50986;
  assign n50988 = pi13 ? n50963 : n50987;
  assign n50989 = pi12 ? n50939 : n50988;
  assign n50990 = pi20 ? n37 : n9482;
  assign n50991 = pi19 ? n31280 : n50990;
  assign n50992 = pi18 ? n20563 : n50991;
  assign n50993 = pi17 ? n48488 : n50992;
  assign n50994 = pi16 ? n32 : n50993;
  assign n50995 = pi20 ? n7730 : n32960;
  assign n50996 = pi19 ? n31280 : n50995;
  assign n50997 = pi18 ? n20563 : n50996;
  assign n50998 = pi17 ? n48488 : n50997;
  assign n50999 = pi16 ? n32 : n50998;
  assign n51000 = pi15 ? n50994 : n50999;
  assign n51001 = pi20 ? n7730 : n7733;
  assign n51002 = pi19 ? n31267 : n51001;
  assign n51003 = pi18 ? n20563 : n51002;
  assign n51004 = pi17 ? n47443 : n51003;
  assign n51005 = pi16 ? n32 : n51004;
  assign n51006 = pi23 ? n8310 : n531;
  assign n51007 = pi22 ? n51006 : n32;
  assign n51008 = pi21 ? n51007 : n32;
  assign n51009 = pi20 ? n24865 : n51008;
  assign n51010 = pi19 ? n31280 : n51009;
  assign n51011 = pi18 ? n20563 : n51010;
  assign n51012 = pi17 ? n47451 : n51011;
  assign n51013 = pi16 ? n32 : n51012;
  assign n51014 = pi15 ? n51005 : n51013;
  assign n51015 = pi14 ? n51000 : n51014;
  assign n51016 = pi20 ? n5077 : n3303;
  assign n51017 = pi19 ? n37 : n51016;
  assign n51018 = pi18 ? n20563 : n51017;
  assign n51019 = pi17 ? n46302 : n51018;
  assign n51020 = pi16 ? n32 : n51019;
  assign n51021 = pi22 ? n41366 : n32;
  assign n51022 = pi21 ? n51021 : n32;
  assign n51023 = pi20 ? n25804 : n51022;
  assign n51024 = pi19 ? n30097 : n51023;
  assign n51025 = pi18 ? n20563 : n51024;
  assign n51026 = pi17 ? n46832 : n51025;
  assign n51027 = pi16 ? n32 : n51026;
  assign n51028 = pi15 ? n51020 : n51027;
  assign n51029 = pi23 ? n35938 : n687;
  assign n51030 = pi22 ? n51029 : n32;
  assign n51031 = pi21 ? n51030 : n32;
  assign n51032 = pi20 ? n24493 : n51031;
  assign n51033 = pi19 ? n30097 : n51032;
  assign n51034 = pi18 ? n20563 : n51033;
  assign n51035 = pi17 ? n46832 : n51034;
  assign n51036 = pi16 ? n32 : n51035;
  assign n51037 = pi18 ? n38948 : n20563;
  assign n51038 = pi20 ? n24493 : n12192;
  assign n51039 = pi19 ? n31280 : n51038;
  assign n51040 = pi18 ? n20563 : n51039;
  assign n51041 = pi17 ? n51037 : n51040;
  assign n51042 = pi16 ? n32 : n51041;
  assign n51043 = pi15 ? n51036 : n51042;
  assign n51044 = pi14 ? n51028 : n51043;
  assign n51045 = pi13 ? n51015 : n51044;
  assign n51046 = pi21 ? n181 : n381;
  assign n51047 = pi20 ? n51046 : n10011;
  assign n51048 = pi19 ? n30097 : n51047;
  assign n51049 = pi18 ? n20563 : n51048;
  assign n51050 = pi17 ? n46839 : n51049;
  assign n51051 = pi16 ? n32 : n51050;
  assign n51052 = pi19 ? n34261 : n50546;
  assign n51053 = pi18 ? n20563 : n51052;
  assign n51054 = pi17 ? n45707 : n51053;
  assign n51055 = pi16 ? n32 : n51054;
  assign n51056 = pi15 ? n51051 : n51055;
  assign n51057 = pi20 ? n30096 : n99;
  assign n51058 = pi19 ? n51057 : n50546;
  assign n51059 = pi18 ? n20563 : n51058;
  assign n51060 = pi17 ? n46859 : n51059;
  assign n51061 = pi16 ? n32 : n51060;
  assign n51062 = pi20 ? n24957 : n1822;
  assign n51063 = pi19 ? n34261 : n51062;
  assign n51064 = pi18 ? n34869 : n51063;
  assign n51065 = pi17 ? n46859 : n51064;
  assign n51066 = pi16 ? n32 : n51065;
  assign n51067 = pi15 ? n51061 : n51066;
  assign n51068 = pi14 ? n51056 : n51067;
  assign n51069 = pi20 ? n20563 : n38381;
  assign n51070 = pi19 ? n20563 : n51069;
  assign n51071 = pi20 ? n14524 : n219;
  assign n51072 = pi20 ? n24957 : n32;
  assign n51073 = pi19 ? n51071 : n51072;
  assign n51074 = pi18 ? n51070 : n51073;
  assign n51075 = pi17 ? n46866 : n51074;
  assign n51076 = pi16 ? n32 : n51075;
  assign n51077 = pi20 ? n20563 : n39805;
  assign n51078 = pi19 ? n20563 : n51077;
  assign n51079 = pi19 ? n27249 : n51072;
  assign n51080 = pi18 ? n51078 : n51079;
  assign n51081 = pi17 ? n46866 : n51080;
  assign n51082 = pi16 ? n32 : n51081;
  assign n51083 = pi15 ? n51076 : n51082;
  assign n51084 = pi21 ? n99 : n5235;
  assign n51085 = pi20 ? n51084 : n32;
  assign n51086 = pi19 ? n45708 : n51085;
  assign n51087 = pi18 ? n34258 : n51086;
  assign n51088 = pi17 ? n50532 : n51087;
  assign n51089 = pi16 ? n32 : n51088;
  assign n51090 = pi21 ? n916 : n22491;
  assign n51091 = pi20 ? n51090 : n32;
  assign n51092 = pi19 ? n17013 : n51091;
  assign n51093 = pi18 ? n34258 : n51092;
  assign n51094 = pi17 ? n46312 : n51093;
  assign n51095 = pi16 ? n32 : n51094;
  assign n51096 = pi15 ? n51089 : n51095;
  assign n51097 = pi14 ? n51083 : n51096;
  assign n51098 = pi13 ? n51068 : n51097;
  assign n51099 = pi12 ? n51045 : n51098;
  assign n51100 = pi11 ? n50989 : n51099;
  assign n51101 = pi21 ? n916 : n1071;
  assign n51102 = pi20 ? n51101 : n32;
  assign n51103 = pi19 ? n37 : n51102;
  assign n51104 = pi18 ? n33245 : n51103;
  assign n51105 = pi17 ? n46312 : n51104;
  assign n51106 = pi16 ? n32 : n51105;
  assign n51107 = pi21 ? n139 : n11235;
  assign n51108 = pi20 ? n51107 : n32;
  assign n51109 = pi19 ? n9814 : n51108;
  assign n51110 = pi18 ? n33245 : n51109;
  assign n51111 = pi17 ? n46312 : n51110;
  assign n51112 = pi16 ? n32 : n51111;
  assign n51113 = pi15 ? n51106 : n51112;
  assign n51114 = pi19 ? n20563 : n49098;
  assign n51115 = pi20 ? n40755 : n3096;
  assign n51116 = pi21 ? n916 : n10417;
  assign n51117 = pi20 ? n51116 : n32;
  assign n51118 = pi19 ? n51115 : n51117;
  assign n51119 = pi18 ? n51114 : n51118;
  assign n51120 = pi17 ? n46312 : n51119;
  assign n51121 = pi16 ? n32 : n51120;
  assign n51122 = pi21 ? n916 : n12381;
  assign n51123 = pi20 ? n51122 : n32;
  assign n51124 = pi19 ? n9824 : n51123;
  assign n51125 = pi18 ? n33245 : n51124;
  assign n51126 = pi17 ? n20563 : n51125;
  assign n51127 = pi16 ? n45233 : n51126;
  assign n51128 = pi15 ? n51121 : n51127;
  assign n51129 = pi14 ? n51113 : n51128;
  assign n51130 = pi22 ? n4883 : n625;
  assign n51131 = pi21 ? n916 : n51130;
  assign n51132 = pi20 ? n51131 : n32;
  assign n51133 = pi19 ? n9814 : n51132;
  assign n51134 = pi18 ? n34258 : n51133;
  assign n51135 = pi17 ? n20563 : n51134;
  assign n51136 = pi16 ? n44635 : n51135;
  assign n51137 = pi21 ? n14952 : n13280;
  assign n51138 = pi20 ? n51137 : n32;
  assign n51139 = pi19 ? n9765 : n51138;
  assign n51140 = pi18 ? n34869 : n51139;
  assign n51141 = pi17 ? n20563 : n51140;
  assign n51142 = pi16 ? n44635 : n51141;
  assign n51143 = pi15 ? n51136 : n51142;
  assign n51144 = pi21 ? n297 : n335;
  assign n51145 = pi20 ? n37 : n51144;
  assign n51146 = pi21 ? n14952 : n4926;
  assign n51147 = pi20 ? n51146 : n32;
  assign n51148 = pi19 ? n51145 : n51147;
  assign n51149 = pi18 ? n34869 : n51148;
  assign n51150 = pi17 ? n20563 : n51149;
  assign n51151 = pi16 ? n44635 : n51150;
  assign n51152 = pi21 ? n6376 : n7723;
  assign n51153 = pi20 ? n51152 : n32;
  assign n51154 = pi19 ? n7685 : n51153;
  assign n51155 = pi18 ? n34869 : n51154;
  assign n51156 = pi17 ? n20563 : n51155;
  assign n51157 = pi16 ? n44635 : n51156;
  assign n51158 = pi15 ? n51151 : n51157;
  assign n51159 = pi14 ? n51143 : n51158;
  assign n51160 = pi13 ? n51129 : n51159;
  assign n51161 = pi21 ? n45016 : n37;
  assign n51162 = pi20 ? n20563 : n51161;
  assign n51163 = pi19 ? n20563 : n51162;
  assign n51164 = pi21 ? n19386 : n12825;
  assign n51165 = pi20 ? n51164 : n32;
  assign n51166 = pi19 ? n37 : n51165;
  assign n51167 = pi18 ? n51163 : n51166;
  assign n51168 = pi17 ? n20563 : n51167;
  assign n51169 = pi16 ? n46885 : n51168;
  assign n51170 = pi21 ? n19386 : n6416;
  assign n51171 = pi20 ? n51170 : n32;
  assign n51172 = pi19 ? n37 : n51171;
  assign n51173 = pi18 ? n39432 : n51172;
  assign n51174 = pi17 ? n20563 : n51173;
  assign n51175 = pi16 ? n46885 : n51174;
  assign n51176 = pi15 ? n51169 : n51175;
  assign n51177 = pi20 ? n33635 : n32;
  assign n51178 = pi19 ? n7676 : n51177;
  assign n51179 = pi18 ? n33245 : n51178;
  assign n51180 = pi17 ? n20563 : n51179;
  assign n51181 = pi16 ? n50067 : n51180;
  assign n51182 = pi21 ? n20563 : n46116;
  assign n51183 = pi21 ? n45049 : n40917;
  assign n51184 = pi20 ? n51182 : n51183;
  assign n51185 = pi21 ? n46116 : n40917;
  assign n51186 = pi19 ? n51184 : n51185;
  assign n51187 = pi21 ? n39191 : n20563;
  assign n51188 = pi21 ? n20563 : n40917;
  assign n51189 = pi20 ? n51187 : n51188;
  assign n51190 = pi20 ? n51185 : n51182;
  assign n51191 = pi19 ? n51189 : n51190;
  assign n51192 = pi18 ? n51186 : n51191;
  assign n51193 = pi22 ? n10098 : n32;
  assign n51194 = pi21 ? n233 : n51193;
  assign n51195 = pi20 ? n51194 : n32;
  assign n51196 = pi19 ? n7676 : n51195;
  assign n51197 = pi18 ? n33245 : n51196;
  assign n51198 = pi17 ? n51192 : n51197;
  assign n51199 = pi16 ? n50067 : n51198;
  assign n51200 = pi15 ? n51181 : n51199;
  assign n51201 = pi14 ? n51176 : n51200;
  assign n51202 = pi21 ? n39801 : n20563;
  assign n51203 = pi20 ? n51202 : n20563;
  assign n51204 = pi19 ? n48343 : n51203;
  assign n51205 = pi18 ? n51204 : n20563;
  assign n51206 = pi19 ? n7685 : n19353;
  assign n51207 = pi18 ? n34295 : n51206;
  assign n51208 = pi17 ? n51205 : n51207;
  assign n51209 = pi16 ? n50067 : n51208;
  assign n51210 = pi18 ? n32 : n46190;
  assign n51211 = pi17 ? n32 : n51210;
  assign n51212 = pi22 ? n42109 : n20563;
  assign n51213 = pi21 ? n40913 : n51212;
  assign n51214 = pi22 ? n36615 : n39190;
  assign n51215 = pi22 ? n30868 : n36615;
  assign n51216 = pi21 ? n51214 : n51215;
  assign n51217 = pi20 ? n51213 : n51216;
  assign n51218 = pi21 ? n37768 : n40960;
  assign n51219 = pi19 ? n51217 : n51218;
  assign n51220 = pi21 ? n41489 : n20563;
  assign n51221 = pi21 ? n20563 : n40960;
  assign n51222 = pi20 ? n51220 : n51221;
  assign n51223 = pi21 ? n20563 : n37768;
  assign n51224 = pi20 ? n51218 : n51223;
  assign n51225 = pi19 ? n51222 : n51224;
  assign n51226 = pi18 ? n51219 : n51225;
  assign n51227 = pi19 ? n7676 : n20208;
  assign n51228 = pi18 ? n34295 : n51227;
  assign n51229 = pi17 ? n51226 : n51228;
  assign n51230 = pi16 ? n51211 : n51229;
  assign n51231 = pi15 ? n51209 : n51230;
  assign n51232 = pi22 ? n45597 : n20563;
  assign n51233 = pi21 ? n32 : n51232;
  assign n51234 = pi20 ? n32 : n51233;
  assign n51235 = pi19 ? n32 : n51234;
  assign n51236 = pi18 ? n32 : n51235;
  assign n51237 = pi17 ? n32 : n51236;
  assign n51238 = pi19 ? n7676 : n13794;
  assign n51239 = pi18 ? n33245 : n51238;
  assign n51240 = pi17 ? n20563 : n51239;
  assign n51241 = pi16 ? n51237 : n51240;
  assign n51242 = pi19 ? n5029 : n12129;
  assign n51243 = pi18 ? n33245 : n51242;
  assign n51244 = pi17 ? n20563 : n51243;
  assign n51245 = pi16 ? n46349 : n51244;
  assign n51246 = pi15 ? n51241 : n51245;
  assign n51247 = pi14 ? n51231 : n51246;
  assign n51248 = pi13 ? n51201 : n51247;
  assign n51249 = pi12 ? n51160 : n51248;
  assign n51250 = pi19 ? n5029 : n10327;
  assign n51251 = pi18 ? n34295 : n51250;
  assign n51252 = pi17 ? n20563 : n51251;
  assign n51253 = pi16 ? n46349 : n51252;
  assign n51254 = pi15 ? n51245 : n51253;
  assign n51255 = pi19 ? n23917 : n8296;
  assign n51256 = pi18 ? n33245 : n51255;
  assign n51257 = pi17 ? n20563 : n51256;
  assign n51258 = pi16 ? n44653 : n51257;
  assign n51259 = pi20 ? n43010 : n3812;
  assign n51260 = pi19 ? n20563 : n51259;
  assign n51261 = pi22 ? n11911 : n157;
  assign n51262 = pi21 ? n363 : n51261;
  assign n51263 = pi20 ? n37 : n51262;
  assign n51264 = pi19 ? n51263 : n8296;
  assign n51265 = pi18 ? n51260 : n51264;
  assign n51266 = pi17 ? n20563 : n51265;
  assign n51267 = pi16 ? n44653 : n51266;
  assign n51268 = pi15 ? n51258 : n51267;
  assign n51269 = pi14 ? n51254 : n51268;
  assign n51270 = pi22 ? n20563 : n36781;
  assign n51271 = pi21 ? n51270 : n37;
  assign n51272 = pi20 ? n20563 : n51271;
  assign n51273 = pi19 ? n20563 : n51272;
  assign n51274 = pi21 ? n37 : n44124;
  assign n51275 = pi20 ? n37 : n51274;
  assign n51276 = pi19 ? n51275 : n9483;
  assign n51277 = pi18 ? n51273 : n51276;
  assign n51278 = pi17 ? n20563 : n51277;
  assign n51279 = pi16 ? n44653 : n51278;
  assign n51280 = pi21 ? n33792 : n20563;
  assign n51281 = pi21 ? n29133 : n297;
  assign n51282 = pi20 ? n51280 : n51281;
  assign n51283 = pi19 ? n20563 : n51282;
  assign n51284 = pi19 ? n31455 : n7725;
  assign n51285 = pi18 ? n51283 : n51284;
  assign n51286 = pi17 ? n20563 : n51285;
  assign n51287 = pi16 ? n44653 : n51286;
  assign n51288 = pi15 ? n51279 : n51287;
  assign n51289 = pi19 ? n32 : n48790;
  assign n51290 = pi18 ? n32 : n51289;
  assign n51291 = pi17 ? n32 : n51290;
  assign n51292 = pi20 ? n39805 : n30868;
  assign n51293 = pi19 ? n51292 : n20563;
  assign n51294 = pi18 ? n51293 : n20563;
  assign n51295 = pi21 ? n99 : n2721;
  assign n51296 = pi20 ? n37 : n51295;
  assign n51297 = pi19 ? n51296 : n7050;
  assign n51298 = pi18 ? n33245 : n51297;
  assign n51299 = pi17 ? n51294 : n51298;
  assign n51300 = pi16 ? n51291 : n51299;
  assign n51301 = pi20 ? n20563 : n30868;
  assign n51302 = pi19 ? n51301 : n20563;
  assign n51303 = pi18 ? n51302 : n20563;
  assign n51304 = pi21 ? n3392 : n2721;
  assign n51305 = pi20 ? n37 : n51304;
  assign n51306 = pi19 ? n51305 : n5831;
  assign n51307 = pi18 ? n33245 : n51306;
  assign n51308 = pi17 ? n51303 : n51307;
  assign n51309 = pi16 ? n44644 : n51308;
  assign n51310 = pi15 ? n51300 : n51309;
  assign n51311 = pi14 ? n51288 : n51310;
  assign n51312 = pi13 ? n51269 : n51311;
  assign n51313 = pi22 ? n30868 : n36781;
  assign n51314 = pi21 ? n51313 : n99;
  assign n51315 = pi20 ? n30868 : n51314;
  assign n51316 = pi19 ? n30868 : n51315;
  assign n51317 = pi21 ? n139 : n3562;
  assign n51318 = pi20 ? n99 : n51317;
  assign n51319 = pi19 ? n51318 : n2654;
  assign n51320 = pi18 ? n51316 : n51319;
  assign n51321 = pi17 ? n30868 : n51320;
  assign n51322 = pi16 ? n44644 : n51321;
  assign n51323 = pi19 ? n32 : n48737;
  assign n51324 = pi18 ? n32 : n51323;
  assign n51325 = pi17 ? n32 : n51324;
  assign n51326 = pi20 ? n99 : n34069;
  assign n51327 = pi19 ? n51326 : n2654;
  assign n51328 = pi18 ? n51316 : n51327;
  assign n51329 = pi17 ? n30868 : n51328;
  assign n51330 = pi16 ? n51325 : n51329;
  assign n51331 = pi15 ? n51322 : n51330;
  assign n51332 = pi19 ? n32 : n48823;
  assign n51333 = pi18 ? n32 : n51332;
  assign n51334 = pi17 ? n32 : n51333;
  assign n51335 = pi21 ? n36798 : n139;
  assign n51336 = pi20 ? n33792 : n51335;
  assign n51337 = pi19 ? n46204 : n51336;
  assign n51338 = pi19 ? n50779 : n35482;
  assign n51339 = pi18 ? n51337 : n51338;
  assign n51340 = pi17 ? n36798 : n51339;
  assign n51341 = pi16 ? n51334 : n51340;
  assign n51342 = pi20 ? n45143 : n50298;
  assign n51343 = pi19 ? n51342 : n48375;
  assign n51344 = pi18 ? n51343 : n33792;
  assign n51345 = pi19 ? n33792 : n49359;
  assign n51346 = pi18 ? n51345 : n50780;
  assign n51347 = pi17 ? n51344 : n51346;
  assign n51348 = pi16 ? n51334 : n51347;
  assign n51349 = pi15 ? n51341 : n51348;
  assign n51350 = pi14 ? n51331 : n51349;
  assign n51351 = pi19 ? n32 : n48858;
  assign n51352 = pi18 ? n32 : n51351;
  assign n51353 = pi17 ? n32 : n51352;
  assign n51354 = pi21 ? n43198 : n50338;
  assign n51355 = pi20 ? n51354 : n43198;
  assign n51356 = pi21 ? n43198 : n36659;
  assign n51357 = pi20 ? n51356 : n36659;
  assign n51358 = pi19 ? n51355 : n51357;
  assign n51359 = pi18 ? n51358 : n36659;
  assign n51360 = pi21 ? n36837 : n10417;
  assign n51361 = pi20 ? n335 : n51360;
  assign n51362 = pi19 ? n51361 : n32;
  assign n51363 = pi18 ? n48395 : n51362;
  assign n51364 = pi17 ? n51359 : n51363;
  assign n51365 = pi16 ? n51353 : n51364;
  assign n51366 = pi23 ? n36830 : n36781;
  assign n51367 = pi22 ? n32 : n51366;
  assign n51368 = pi21 ? n32 : n51367;
  assign n51369 = pi20 ? n32 : n51368;
  assign n51370 = pi19 ? n32 : n51369;
  assign n51371 = pi18 ? n32 : n51370;
  assign n51372 = pi17 ? n32 : n51371;
  assign n51373 = pi21 ? n36837 : n39815;
  assign n51374 = pi20 ? n335 : n51373;
  assign n51375 = pi19 ? n51374 : n32;
  assign n51376 = pi18 ? n48395 : n51375;
  assign n51377 = pi17 ? n36659 : n51376;
  assign n51378 = pi16 ? n51372 : n51377;
  assign n51379 = pi15 ? n51365 : n51378;
  assign n51380 = pi20 ? n50354 : n42170;
  assign n51381 = pi19 ? n51380 : n36781;
  assign n51382 = pi18 ? n51381 : n36781;
  assign n51383 = pi20 ? n36781 : n48423;
  assign n51384 = pi19 ? n36781 : n51383;
  assign n51385 = pi20 ? n363 : n5179;
  assign n51386 = pi19 ? n51385 : n32;
  assign n51387 = pi18 ? n51384 : n51386;
  assign n51388 = pi17 ? n51382 : n51387;
  assign n51389 = pi16 ? n51334 : n51388;
  assign n51390 = pi20 ? n46281 : n43198;
  assign n51391 = pi20 ? n49424 : n36781;
  assign n51392 = pi19 ? n51390 : n51391;
  assign n51393 = pi18 ? n51392 : n36781;
  assign n51394 = pi20 ? n36781 : n36798;
  assign n51395 = pi19 ? n36781 : n51394;
  assign n51396 = pi21 ? n48427 : n157;
  assign n51397 = pi20 ? n51396 : n19275;
  assign n51398 = pi19 ? n51397 : n32;
  assign n51399 = pi18 ? n51395 : n51398;
  assign n51400 = pi17 ? n51393 : n51399;
  assign n51401 = pi16 ? n51353 : n51400;
  assign n51402 = pi15 ? n51389 : n51401;
  assign n51403 = pi14 ? n51379 : n51402;
  assign n51404 = pi13 ? n51350 : n51403;
  assign n51405 = pi12 ? n51312 : n51404;
  assign n51406 = pi11 ? n51249 : n51405;
  assign n51407 = pi10 ? n51100 : n51406;
  assign n51408 = pi09 ? n50882 : n51407;
  assign n51409 = pi17 ? n37958 : n50859;
  assign n51410 = pi16 ? n32 : n51409;
  assign n51411 = pi15 ? n32 : n51410;
  assign n51412 = pi17 ? n37323 : n50867;
  assign n51413 = pi16 ? n32 : n51412;
  assign n51414 = pi20 ? n37 : n19778;
  assign n51415 = pi19 ? n37 : n51414;
  assign n51416 = pi18 ? n34295 : n51415;
  assign n51417 = pi17 ? n37323 : n51416;
  assign n51418 = pi16 ? n32 : n51417;
  assign n51419 = pi15 ? n51413 : n51418;
  assign n51420 = pi14 ? n51411 : n51419;
  assign n51421 = pi13 ? n32 : n51420;
  assign n51422 = pi12 ? n32 : n51421;
  assign n51423 = pi11 ? n32 : n51422;
  assign n51424 = pi10 ? n32 : n51423;
  assign n51425 = pi20 ? n3086 : n19794;
  assign n51426 = pi19 ? n50883 : n51425;
  assign n51427 = pi18 ? n34258 : n51426;
  assign n51428 = pi17 ? n35764 : n51427;
  assign n51429 = pi16 ? n32 : n51428;
  assign n51430 = pi20 ? n3086 : n50891;
  assign n51431 = pi19 ? n50883 : n51430;
  assign n51432 = pi18 ? n34869 : n51431;
  assign n51433 = pi17 ? n35764 : n51432;
  assign n51434 = pi16 ? n32 : n51433;
  assign n51435 = pi15 ? n51429 : n51434;
  assign n51436 = pi22 ? n37 : n261;
  assign n51437 = pi21 ? n51436 : n32;
  assign n51438 = pi20 ? n8742 : n51437;
  assign n51439 = pi19 ? n37 : n51438;
  assign n51440 = pi18 ? n34295 : n51439;
  assign n51441 = pi17 ? n50390 : n51440;
  assign n51442 = pi16 ? n32 : n51441;
  assign n51443 = pi22 ? n295 : n261;
  assign n51444 = pi21 ? n51443 : n32;
  assign n51445 = pi20 ? n37 : n51444;
  assign n51446 = pi19 ? n37 : n51445;
  assign n51447 = pi18 ? n50907 : n51446;
  assign n51448 = pi17 ? n50393 : n51447;
  assign n51449 = pi16 ? n32 : n51448;
  assign n51450 = pi15 ? n51442 : n51449;
  assign n51451 = pi14 ? n51435 : n51450;
  assign n51452 = pi20 ? n37 : n19505;
  assign n51453 = pi19 ? n37 : n51452;
  assign n51454 = pi18 ? n34295 : n51453;
  assign n51455 = pi17 ? n49888 : n51454;
  assign n51456 = pi16 ? n32 : n51455;
  assign n51457 = pi20 ? n37 : n35231;
  assign n51458 = pi21 ? n43748 : n32;
  assign n51459 = pi20 ? n37 : n51458;
  assign n51460 = pi19 ? n51457 : n51459;
  assign n51461 = pi18 ? n34869 : n51460;
  assign n51462 = pi17 ? n49894 : n51461;
  assign n51463 = pi16 ? n32 : n51462;
  assign n51464 = pi15 ? n51456 : n51463;
  assign n51465 = pi20 ? n48905 : n33821;
  assign n51466 = pi19 ? n51465 : n51459;
  assign n51467 = pi18 ? n20563 : n51466;
  assign n51468 = pi17 ? n49448 : n51467;
  assign n51469 = pi16 ? n32 : n51468;
  assign n51470 = pi20 ? n649 : n20801;
  assign n51471 = pi19 ? n50932 : n51470;
  assign n51472 = pi18 ? n20563 : n51471;
  assign n51473 = pi17 ? n49448 : n51472;
  assign n51474 = pi16 ? n32 : n51473;
  assign n51475 = pi15 ? n51469 : n51474;
  assign n51476 = pi14 ? n51464 : n51475;
  assign n51477 = pi13 ? n51451 : n51476;
  assign n51478 = pi21 ? n26982 : n32;
  assign n51479 = pi20 ? n3299 : n51478;
  assign n51480 = pi19 ? n32898 : n51479;
  assign n51481 = pi18 ? n20563 : n51480;
  assign n51482 = pi17 ? n49451 : n51481;
  assign n51483 = pi16 ? n32 : n51482;
  assign n51484 = pi22 ? n363 : n20340;
  assign n51485 = pi21 ? n51484 : n32;
  assign n51486 = pi20 ? n649 : n51485;
  assign n51487 = pi19 ? n32348 : n51486;
  assign n51488 = pi18 ? n20563 : n51487;
  assign n51489 = pi17 ? n50426 : n51488;
  assign n51490 = pi16 ? n32 : n51489;
  assign n51491 = pi15 ? n51483 : n51490;
  assign n51492 = pi20 ? n649 : n25399;
  assign n51493 = pi19 ? n31280 : n51492;
  assign n51494 = pi18 ? n20563 : n51493;
  assign n51495 = pi17 ? n48904 : n51494;
  assign n51496 = pi16 ? n32 : n51495;
  assign n51497 = pi20 ? n50956 : n34952;
  assign n51498 = pi19 ? n31267 : n51497;
  assign n51499 = pi18 ? n20563 : n51498;
  assign n51500 = pi17 ? n48466 : n51499;
  assign n51501 = pi16 ? n32 : n51500;
  assign n51502 = pi15 ? n51496 : n51501;
  assign n51503 = pi14 ? n51491 : n51502;
  assign n51504 = pi20 ? n37 : n4749;
  assign n51505 = pi19 ? n32348 : n51504;
  assign n51506 = pi18 ? n20563 : n51505;
  assign n51507 = pi17 ? n48466 : n51506;
  assign n51508 = pi16 ? n32 : n51507;
  assign n51509 = pi23 ? n5612 : n204;
  assign n51510 = pi22 ? n51509 : n532;
  assign n51511 = pi21 ? n51510 : n32;
  assign n51512 = pi20 ? n37 : n51511;
  assign n51513 = pi19 ? n32348 : n51512;
  assign n51514 = pi18 ? n20563 : n51513;
  assign n51515 = pi17 ? n48469 : n51514;
  assign n51516 = pi16 ? n32 : n51515;
  assign n51517 = pi15 ? n51508 : n51516;
  assign n51518 = pi20 ? n37 : n22920;
  assign n51519 = pi19 ? n31267 : n51518;
  assign n51520 = pi18 ? n20563 : n51519;
  assign n51521 = pi17 ? n49485 : n51520;
  assign n51522 = pi16 ? n32 : n51521;
  assign n51523 = pi17 ? n47929 : n50983;
  assign n51524 = pi16 ? n32 : n51523;
  assign n51525 = pi15 ? n51522 : n51524;
  assign n51526 = pi14 ? n51517 : n51525;
  assign n51527 = pi13 ? n51503 : n51526;
  assign n51528 = pi12 ? n51477 : n51527;
  assign n51529 = pi19 ? n32871 : n50990;
  assign n51530 = pi18 ? n20563 : n51529;
  assign n51531 = pi17 ? n47929 : n51530;
  assign n51532 = pi16 ? n32 : n51531;
  assign n51533 = pi17 ? n47929 : n50997;
  assign n51534 = pi16 ? n32 : n51533;
  assign n51535 = pi15 ? n51532 : n51534;
  assign n51536 = pi17 ? n47929 : n51003;
  assign n51537 = pi16 ? n32 : n51536;
  assign n51538 = pi20 ? n24865 : n31964;
  assign n51539 = pi19 ? n31280 : n51538;
  assign n51540 = pi18 ? n20563 : n51539;
  assign n51541 = pi17 ? n47935 : n51540;
  assign n51542 = pi16 ? n32 : n51541;
  assign n51543 = pi15 ? n51537 : n51542;
  assign n51544 = pi14 ? n51535 : n51543;
  assign n51545 = pi23 ? n31328 : n99;
  assign n51546 = pi22 ? n37 : n51545;
  assign n51547 = pi21 ? n37 : n51546;
  assign n51548 = pi20 ? n51547 : n3303;
  assign n51549 = pi19 ? n31299 : n51548;
  assign n51550 = pi18 ? n20563 : n51549;
  assign n51551 = pi17 ? n47947 : n51550;
  assign n51552 = pi16 ? n32 : n51551;
  assign n51553 = pi20 ? n25804 : n3303;
  assign n51554 = pi19 ? n32287 : n51553;
  assign n51555 = pi18 ? n20563 : n51554;
  assign n51556 = pi17 ? n47954 : n51555;
  assign n51557 = pi16 ? n32 : n51556;
  assign n51558 = pi15 ? n51552 : n51557;
  assign n51559 = pi20 ? n24493 : n6417;
  assign n51560 = pi19 ? n30097 : n51559;
  assign n51561 = pi18 ? n20563 : n51560;
  assign n51562 = pi17 ? n47954 : n51561;
  assign n51563 = pi16 ? n32 : n51562;
  assign n51564 = pi25 ? n684 : n32;
  assign n51565 = pi24 ? n51564 : n32;
  assign n51566 = pi23 ? n316 : n51565;
  assign n51567 = pi22 ? n51566 : n32;
  assign n51568 = pi21 ? n51567 : n32;
  assign n51569 = pi20 ? n24493 : n51568;
  assign n51570 = pi19 ? n31280 : n51569;
  assign n51571 = pi18 ? n20563 : n51570;
  assign n51572 = pi17 ? n48488 : n51571;
  assign n51573 = pi16 ? n32 : n51572;
  assign n51574 = pi15 ? n51563 : n51573;
  assign n51575 = pi14 ? n51558 : n51574;
  assign n51576 = pi13 ? n51544 : n51575;
  assign n51577 = pi20 ? n51046 : n3210;
  assign n51578 = pi19 ? n33949 : n51577;
  assign n51579 = pi18 ? n20563 : n51578;
  assign n51580 = pi17 ? n47443 : n51579;
  assign n51581 = pi16 ? n32 : n51580;
  assign n51582 = pi20 ? n31298 : n14844;
  assign n51583 = pi20 ? n24957 : n10011;
  assign n51584 = pi19 ? n51582 : n51583;
  assign n51585 = pi18 ? n20563 : n51584;
  assign n51586 = pi17 ? n47451 : n51585;
  assign n51587 = pi16 ? n32 : n51586;
  assign n51588 = pi15 ? n51581 : n51587;
  assign n51589 = pi19 ? n51057 : n51583;
  assign n51590 = pi18 ? n20563 : n51589;
  assign n51591 = pi17 ? n46302 : n51590;
  assign n51592 = pi16 ? n32 : n51591;
  assign n51593 = pi18 ? n36931 : n51052;
  assign n51594 = pi17 ? n46302 : n51593;
  assign n51595 = pi16 ? n32 : n51594;
  assign n51596 = pi15 ? n51592 : n51595;
  assign n51597 = pi14 ? n51588 : n51596;
  assign n51598 = pi21 ? n20563 : n37124;
  assign n51599 = pi20 ? n20563 : n51598;
  assign n51600 = pi19 ? n20563 : n51599;
  assign n51601 = pi20 ? n37 : n219;
  assign n51602 = pi19 ? n51601 : n51062;
  assign n51603 = pi18 ? n51600 : n51602;
  assign n51604 = pi17 ? n47964 : n51603;
  assign n51605 = pi16 ? n32 : n51604;
  assign n51606 = pi22 ? n30869 : n99;
  assign n51607 = pi21 ? n51606 : n181;
  assign n51608 = pi20 ? n51607 : n99;
  assign n51609 = pi19 ? n51608 : n51062;
  assign n51610 = pi18 ? n51078 : n51609;
  assign n51611 = pi17 ? n47964 : n51610;
  assign n51612 = pi16 ? n32 : n51611;
  assign n51613 = pi15 ? n51605 : n51612;
  assign n51614 = pi21 ? n99 : n916;
  assign n51615 = pi20 ? n51614 : n32;
  assign n51616 = pi19 ? n45708 : n51615;
  assign n51617 = pi18 ? n34865 : n51616;
  assign n51618 = pi17 ? n51037 : n51617;
  assign n51619 = pi16 ? n32 : n51618;
  assign n51620 = pi20 ? n30593 : n32;
  assign n51621 = pi19 ? n17013 : n51620;
  assign n51622 = pi18 ? n34865 : n51621;
  assign n51623 = pi17 ? n46839 : n51622;
  assign n51624 = pi16 ? n32 : n51623;
  assign n51625 = pi15 ? n51619 : n51624;
  assign n51626 = pi14 ? n51613 : n51625;
  assign n51627 = pi13 ? n51597 : n51626;
  assign n51628 = pi12 ? n51576 : n51627;
  assign n51629 = pi11 ? n51528 : n51628;
  assign n51630 = pi19 ? n37 : n51620;
  assign n51631 = pi18 ? n35777 : n51630;
  assign n51632 = pi17 ? n46839 : n51631;
  assign n51633 = pi16 ? n32 : n51632;
  assign n51634 = pi21 ? n139 : n29992;
  assign n51635 = pi20 ? n51634 : n32;
  assign n51636 = pi19 ? n9814 : n51635;
  assign n51637 = pi18 ? n35777 : n51636;
  assign n51638 = pi17 ? n46859 : n51637;
  assign n51639 = pi16 ? n32 : n51638;
  assign n51640 = pi15 ? n51633 : n51639;
  assign n51641 = pi21 ? n30868 : n31200;
  assign n51642 = pi20 ? n20563 : n51641;
  assign n51643 = pi19 ? n20563 : n51642;
  assign n51644 = pi21 ? n916 : n29992;
  assign n51645 = pi20 ? n51644 : n32;
  assign n51646 = pi19 ? n51115 : n51645;
  assign n51647 = pi18 ? n51643 : n51646;
  assign n51648 = pi17 ? n46859 : n51647;
  assign n51649 = pi16 ? n32 : n51648;
  assign n51650 = pi21 ? n916 : n1027;
  assign n51651 = pi20 ? n51650 : n32;
  assign n51652 = pi19 ? n9824 : n51651;
  assign n51653 = pi18 ? n40199 : n51652;
  assign n51654 = pi17 ? n45715 : n51653;
  assign n51655 = pi16 ? n32 : n51654;
  assign n51656 = pi15 ? n51649 : n51655;
  assign n51657 = pi14 ? n51640 : n51656;
  assign n51658 = pi21 ? n916 : n10106;
  assign n51659 = pi20 ? n51658 : n32;
  assign n51660 = pi19 ? n9814 : n51659;
  assign n51661 = pi18 ? n34258 : n51660;
  assign n51662 = pi17 ? n46866 : n51661;
  assign n51663 = pi16 ? n32 : n51662;
  assign n51664 = pi21 ? n14952 : n8916;
  assign n51665 = pi20 ? n51664 : n32;
  assign n51666 = pi19 ? n9765 : n51665;
  assign n51667 = pi18 ? n34869 : n51666;
  assign n51668 = pi17 ? n46866 : n51667;
  assign n51669 = pi16 ? n32 : n51668;
  assign n51670 = pi15 ? n51663 : n51669;
  assign n51671 = pi21 ? n14952 : n5758;
  assign n51672 = pi20 ? n51671 : n32;
  assign n51673 = pi19 ? n51145 : n51672;
  assign n51674 = pi18 ? n34869 : n51673;
  assign n51675 = pi17 ? n46866 : n51674;
  assign n51676 = pi16 ? n32 : n51675;
  assign n51677 = pi18 ? n38951 : n51154;
  assign n51678 = pi17 ? n46866 : n51677;
  assign n51679 = pi16 ? n32 : n51678;
  assign n51680 = pi15 ? n51676 : n51679;
  assign n51681 = pi14 ? n51670 : n51680;
  assign n51682 = pi13 ? n51657 : n51681;
  assign n51683 = pi21 ? n45016 : n30843;
  assign n51684 = pi20 ? n20563 : n51683;
  assign n51685 = pi19 ? n20563 : n51684;
  assign n51686 = pi21 ? n19386 : n7041;
  assign n51687 = pi20 ? n51686 : n32;
  assign n51688 = pi19 ? n37 : n51687;
  assign n51689 = pi18 ? n51685 : n51688;
  assign n51690 = pi17 ? n46312 : n51689;
  assign n51691 = pi16 ? n32 : n51690;
  assign n51692 = pi21 ? n19386 : n4101;
  assign n51693 = pi20 ? n51692 : n32;
  assign n51694 = pi19 ? n37 : n51693;
  assign n51695 = pi18 ? n40191 : n51694;
  assign n51696 = pi17 ? n20563 : n51695;
  assign n51697 = pi16 ? n45233 : n51696;
  assign n51698 = pi15 ? n51691 : n51697;
  assign n51699 = pi18 ? n35777 : n51178;
  assign n51700 = pi17 ? n20563 : n51699;
  assign n51701 = pi16 ? n32 : n51700;
  assign n51702 = pi20 ? n32 : n47848;
  assign n51703 = pi19 ? n32 : n51702;
  assign n51704 = pi18 ? n32 : n51703;
  assign n51705 = pi17 ? n32 : n51704;
  assign n51706 = pi21 ? n40249 : n30868;
  assign n51707 = pi20 ? n30868 : n51706;
  assign n51708 = pi21 ? n40913 : n36489;
  assign n51709 = pi21 ? n46116 : n40912;
  assign n51710 = pi20 ? n51708 : n51709;
  assign n51711 = pi19 ? n51707 : n51710;
  assign n51712 = pi21 ? n45049 : n36489;
  assign n51713 = pi20 ? n51187 : n51712;
  assign n51714 = pi22 ? n39190 : n40386;
  assign n51715 = pi21 ? n51714 : n40917;
  assign n51716 = pi20 ? n51715 : n46116;
  assign n51717 = pi19 ? n51713 : n51716;
  assign n51718 = pi18 ? n51711 : n51717;
  assign n51719 = pi19 ? n7676 : n20549;
  assign n51720 = pi18 ? n35777 : n51719;
  assign n51721 = pi17 ? n51718 : n51720;
  assign n51722 = pi16 ? n51705 : n51721;
  assign n51723 = pi15 ? n51701 : n51722;
  assign n51724 = pi14 ? n51698 : n51723;
  assign n51725 = pi21 ? n233 : n19697;
  assign n51726 = pi20 ? n51725 : n32;
  assign n51727 = pi19 ? n7685 : n51726;
  assign n51728 = pi18 ? n43367 : n51727;
  assign n51729 = pi17 ? n51205 : n51728;
  assign n51730 = pi16 ? n32 : n51729;
  assign n51731 = pi21 ? n32 : n49721;
  assign n51732 = pi20 ? n32 : n51731;
  assign n51733 = pi19 ? n32 : n51732;
  assign n51734 = pi18 ? n32 : n51733;
  assign n51735 = pi17 ? n32 : n51734;
  assign n51736 = pi21 ? n45526 : n33792;
  assign n51737 = pi20 ? n33792 : n51736;
  assign n51738 = pi21 ? n40955 : n45016;
  assign n51739 = pi21 ? n37768 : n45008;
  assign n51740 = pi20 ? n51738 : n51739;
  assign n51741 = pi19 ? n51737 : n51740;
  assign n51742 = pi21 ? n40954 : n45016;
  assign n51743 = pi20 ? n51220 : n51742;
  assign n51744 = pi22 ? n37173 : n36615;
  assign n51745 = pi21 ? n51744 : n40960;
  assign n51746 = pi20 ? n51745 : n37768;
  assign n51747 = pi19 ? n51743 : n51746;
  assign n51748 = pi18 ? n51741 : n51747;
  assign n51749 = pi19 ? n7676 : n22583;
  assign n51750 = pi18 ? n43367 : n51749;
  assign n51751 = pi17 ? n51748 : n51750;
  assign n51752 = pi16 ? n51735 : n51751;
  assign n51753 = pi15 ? n51730 : n51752;
  assign n51754 = pi23 ? n32 : n36659;
  assign n51755 = pi22 ? n32 : n51754;
  assign n51756 = pi21 ? n32 : n51755;
  assign n51757 = pi20 ? n32 : n51756;
  assign n51758 = pi19 ? n32 : n51757;
  assign n51759 = pi18 ? n32 : n51758;
  assign n51760 = pi17 ? n32 : n51759;
  assign n51761 = pi21 ? n36659 : n43571;
  assign n51762 = pi22 ? n37783 : n36659;
  assign n51763 = pi21 ? n20563 : n51762;
  assign n51764 = pi20 ? n51761 : n51763;
  assign n51765 = pi19 ? n51764 : n20563;
  assign n51766 = pi18 ? n51765 : n20563;
  assign n51767 = pi19 ? n7676 : n14724;
  assign n51768 = pi18 ? n33823 : n51767;
  assign n51769 = pi17 ? n51766 : n51768;
  assign n51770 = pi16 ? n51760 : n51769;
  assign n51771 = pi20 ? n39328 : n32;
  assign n51772 = pi19 ? n5029 : n51771;
  assign n51773 = pi18 ? n33823 : n51772;
  assign n51774 = pi17 ? n20563 : n51773;
  assign n51775 = pi16 ? n46885 : n51774;
  assign n51776 = pi15 ? n51770 : n51775;
  assign n51777 = pi14 ? n51753 : n51776;
  assign n51778 = pi13 ? n51724 : n51777;
  assign n51779 = pi12 ? n51682 : n51778;
  assign n51780 = pi18 ? n33823 : n51242;
  assign n51781 = pi17 ? n20563 : n51780;
  assign n51782 = pi16 ? n45740 : n51781;
  assign n51783 = pi18 ? n35799 : n51250;
  assign n51784 = pi17 ? n20563 : n51783;
  assign n51785 = pi16 ? n45740 : n51784;
  assign n51786 = pi15 ? n51782 : n51785;
  assign n51787 = pi19 ? n23917 : n9457;
  assign n51788 = pi18 ? n39432 : n51787;
  assign n51789 = pi17 ? n20563 : n51788;
  assign n51790 = pi16 ? n44635 : n51789;
  assign n51791 = pi20 ? n43010 : n40263;
  assign n51792 = pi19 ? n20563 : n51791;
  assign n51793 = pi21 ? n363 : n244;
  assign n51794 = pi20 ? n37 : n51793;
  assign n51795 = pi19 ? n51794 : n9964;
  assign n51796 = pi18 ? n51792 : n51795;
  assign n51797 = pi17 ? n20563 : n51796;
  assign n51798 = pi16 ? n44635 : n51797;
  assign n51799 = pi15 ? n51790 : n51798;
  assign n51800 = pi14 ? n51786 : n51799;
  assign n51801 = pi21 ? n51270 : n30843;
  assign n51802 = pi20 ? n20563 : n51801;
  assign n51803 = pi19 ? n20563 : n51802;
  assign n51804 = pi18 ? n51803 : n51276;
  assign n51805 = pi17 ? n20563 : n51804;
  assign n51806 = pi16 ? n44635 : n51805;
  assign n51807 = pi21 ? n39292 : n49764;
  assign n51808 = pi20 ? n51280 : n51807;
  assign n51809 = pi19 ? n20563 : n51808;
  assign n51810 = pi19 ? n31455 : n37549;
  assign n51811 = pi18 ? n51809 : n51810;
  assign n51812 = pi17 ? n20563 : n51811;
  assign n51813 = pi16 ? n46326 : n51812;
  assign n51814 = pi15 ? n51806 : n51813;
  assign n51815 = pi20 ? n32 : n47746;
  assign n51816 = pi19 ? n32 : n51815;
  assign n51817 = pi18 ? n32 : n51816;
  assign n51818 = pi17 ? n32 : n51817;
  assign n51819 = pi19 ? n51296 : n8991;
  assign n51820 = pi18 ? n39432 : n51819;
  assign n51821 = pi17 ? n51294 : n51820;
  assign n51822 = pi16 ? n51818 : n51821;
  assign n51823 = pi19 ? n32 : n49331;
  assign n51824 = pi18 ? n32 : n51823;
  assign n51825 = pi17 ? n32 : n51824;
  assign n51826 = pi22 ? n50358 : n685;
  assign n51827 = pi21 ? n3392 : n51826;
  assign n51828 = pi20 ? n37 : n51827;
  assign n51829 = pi19 ? n51828 : n7050;
  assign n51830 = pi18 ? n39432 : n51829;
  assign n51831 = pi17 ? n51303 : n51830;
  assign n51832 = pi16 ? n51825 : n51831;
  assign n51833 = pi15 ? n51822 : n51832;
  assign n51834 = pi14 ? n51814 : n51833;
  assign n51835 = pi13 ? n51800 : n51834;
  assign n51836 = pi21 ? n51313 : n39315;
  assign n51837 = pi20 ? n30868 : n51836;
  assign n51838 = pi19 ? n30868 : n51837;
  assign n51839 = pi19 ? n51318 : n10012;
  assign n51840 = pi18 ? n51838 : n51839;
  assign n51841 = pi17 ? n30868 : n51840;
  assign n51842 = pi16 ? n32 : n51841;
  assign n51843 = pi19 ? n51326 : n10012;
  assign n51844 = pi18 ? n51838 : n51843;
  assign n51845 = pi17 ? n30868 : n51844;
  assign n51846 = pi16 ? n32 : n51845;
  assign n51847 = pi15 ? n51842 : n51846;
  assign n51848 = pi20 ? n41601 : n36798;
  assign n51849 = pi19 ? n51848 : n36798;
  assign n51850 = pi18 ? n51849 : n36798;
  assign n51851 = pi21 ? n36798 : n36762;
  assign n51852 = pi20 ? n33792 : n51851;
  assign n51853 = pi19 ? n46204 : n51852;
  assign n51854 = pi19 ? n50779 : n2654;
  assign n51855 = pi18 ? n51853 : n51854;
  assign n51856 = pi17 ? n51850 : n51855;
  assign n51857 = pi16 ? n32 : n51856;
  assign n51858 = pi21 ? n41600 : n45142;
  assign n51859 = pi20 ? n51858 : n50298;
  assign n51860 = pi19 ? n51859 : n48375;
  assign n51861 = pi18 ? n51860 : n33792;
  assign n51862 = pi21 ? n40428 : n139;
  assign n51863 = pi20 ? n33792 : n51862;
  assign n51864 = pi19 ? n33792 : n51863;
  assign n51865 = pi18 ? n51864 : n51854;
  assign n51866 = pi17 ? n51861 : n51865;
  assign n51867 = pi16 ? n32 : n51866;
  assign n51868 = pi15 ? n51857 : n51867;
  assign n51869 = pi14 ? n51847 : n51868;
  assign n51870 = pi21 ? n49844 : n50338;
  assign n51871 = pi20 ? n51870 : n43198;
  assign n51872 = pi19 ? n51871 : n51357;
  assign n51873 = pi18 ? n51872 : n36659;
  assign n51874 = pi20 ? n36659 : n37903;
  assign n51875 = pi19 ? n36659 : n51874;
  assign n51876 = pi21 ? n36837 : n10410;
  assign n51877 = pi20 ? n335 : n51876;
  assign n51878 = pi19 ? n51877 : n32;
  assign n51879 = pi18 ? n51875 : n51878;
  assign n51880 = pi17 ? n51873 : n51879;
  assign n51881 = pi16 ? n32 : n51880;
  assign n51882 = pi22 ? n46275 : n36659;
  assign n51883 = pi21 ? n51882 : n36659;
  assign n51884 = pi20 ? n51883 : n36659;
  assign n51885 = pi19 ? n51884 : n36659;
  assign n51886 = pi18 ? n51885 : n36659;
  assign n51887 = pi18 ? n51875 : n51375;
  assign n51888 = pi17 ? n51886 : n51887;
  assign n51889 = pi16 ? n32 : n51888;
  assign n51890 = pi15 ? n51881 : n51889;
  assign n51891 = pi21 ? n46727 : n38901;
  assign n51892 = pi20 ? n51891 : n42170;
  assign n51893 = pi19 ? n51892 : n36781;
  assign n51894 = pi18 ? n51893 : n36781;
  assign n51895 = pi23 ? n36781 : n363;
  assign n51896 = pi22 ? n36798 : n51895;
  assign n51897 = pi21 ? n36781 : n51896;
  assign n51898 = pi20 ? n36781 : n51897;
  assign n51899 = pi19 ? n36781 : n51898;
  assign n51900 = pi18 ? n51899 : n51386;
  assign n51901 = pi17 ? n51894 : n51900;
  assign n51902 = pi16 ? n32 : n51901;
  assign n51903 = pi21 ? n48856 : n46280;
  assign n51904 = pi20 ? n51903 : n43198;
  assign n51905 = pi19 ? n51904 : n51391;
  assign n51906 = pi18 ? n51905 : n36781;
  assign n51907 = pi23 ? n36798 : n157;
  assign n51908 = pi22 ? n51907 : n157;
  assign n51909 = pi21 ? n51908 : n157;
  assign n51910 = pi21 ? n204 : n3494;
  assign n51911 = pi20 ? n51909 : n51910;
  assign n51912 = pi19 ? n51911 : n32;
  assign n51913 = pi18 ? n51395 : n51912;
  assign n51914 = pi17 ? n51906 : n51913;
  assign n51915 = pi16 ? n32 : n51914;
  assign n51916 = pi15 ? n51902 : n51915;
  assign n51917 = pi14 ? n51890 : n51916;
  assign n51918 = pi13 ? n51869 : n51917;
  assign n51919 = pi12 ? n51835 : n51918;
  assign n51920 = pi11 ? n51779 : n51919;
  assign n51921 = pi10 ? n51629 : n51920;
  assign n51922 = pi09 ? n51424 : n51921;
  assign n51923 = pi08 ? n51408 : n51922;
  assign n51924 = pi22 ? n139 : n18038;
  assign n51925 = pi21 ? n51924 : n32;
  assign n51926 = pi20 ? n37 : n51925;
  assign n51927 = pi19 ? n37 : n51926;
  assign n51928 = pi18 ? n50855 : n51927;
  assign n51929 = pi17 ? n38984 : n51928;
  assign n51930 = pi16 ? n32 : n51929;
  assign n51931 = pi15 ? n32 : n51930;
  assign n51932 = pi20 ? n31925 : n20563;
  assign n51933 = pi19 ? n51932 : n32898;
  assign n51934 = pi20 ? n8742 : n51925;
  assign n51935 = pi19 ? n37 : n51934;
  assign n51936 = pi18 ? n51933 : n51935;
  assign n51937 = pi17 ? n40057 : n51936;
  assign n51938 = pi16 ? n32 : n51937;
  assign n51939 = pi23 ? n8184 : n586;
  assign n51940 = pi22 ? n139 : n51939;
  assign n51941 = pi21 ? n51940 : n32;
  assign n51942 = pi20 ? n37 : n51941;
  assign n51943 = pi19 ? n37 : n51942;
  assign n51944 = pi18 ? n34295 : n51943;
  assign n51945 = pi17 ? n36870 : n51944;
  assign n51946 = pi16 ? n32 : n51945;
  assign n51947 = pi15 ? n51938 : n51946;
  assign n51948 = pi14 ? n51931 : n51947;
  assign n51949 = pi13 ? n32 : n51948;
  assign n51950 = pi12 ? n32 : n51949;
  assign n51951 = pi11 ? n32 : n51950;
  assign n51952 = pi10 ? n32 : n51951;
  assign n51953 = pi20 ? n37 : n20563;
  assign n51954 = pi21 ? n27288 : n32;
  assign n51955 = pi20 ? n8742 : n51954;
  assign n51956 = pi19 ? n51953 : n51955;
  assign n51957 = pi18 ? n34258 : n51956;
  assign n51958 = pi17 ? n39456 : n51957;
  assign n51959 = pi16 ? n32 : n51958;
  assign n51960 = pi23 ? n1432 : n1149;
  assign n51961 = pi22 ? n139 : n51960;
  assign n51962 = pi21 ? n51961 : n32;
  assign n51963 = pi20 ? n3086 : n51962;
  assign n51964 = pi19 ? n50883 : n51963;
  assign n51965 = pi18 ? n34869 : n51964;
  assign n51966 = pi17 ? n39456 : n51965;
  assign n51967 = pi16 ? n32 : n51966;
  assign n51968 = pi15 ? n51959 : n51967;
  assign n51969 = pi23 ? n31328 : n531;
  assign n51970 = pi22 ? n37 : n51969;
  assign n51971 = pi21 ? n51970 : n32;
  assign n51972 = pi20 ? n37 : n51971;
  assign n51973 = pi19 ? n37 : n51972;
  assign n51974 = pi18 ? n34295 : n51973;
  assign n51975 = pi17 ? n36162 : n51974;
  assign n51976 = pi16 ? n32 : n51975;
  assign n51977 = pi22 ? n37 : n171;
  assign n51978 = pi21 ? n51977 : n32;
  assign n51979 = pi20 ? n37 : n51978;
  assign n51980 = pi19 ? n37 : n51979;
  assign n51981 = pi18 ? n50907 : n51980;
  assign n51982 = pi17 ? n35764 : n51981;
  assign n51983 = pi16 ? n32 : n51982;
  assign n51984 = pi15 ? n51976 : n51983;
  assign n51985 = pi14 ? n51968 : n51984;
  assign n51986 = pi17 ? n36215 : n51454;
  assign n51987 = pi16 ? n32 : n51986;
  assign n51988 = pi21 ? n36249 : n30843;
  assign n51989 = pi20 ? n37 : n51988;
  assign n51990 = pi20 ? n37 : n20794;
  assign n51991 = pi19 ? n51989 : n51990;
  assign n51992 = pi18 ? n34869 : n51991;
  assign n51993 = pi17 ? n49894 : n51992;
  assign n51994 = pi16 ? n32 : n51993;
  assign n51995 = pi15 ? n51987 : n51994;
  assign n51996 = pi20 ? n48905 : n31266;
  assign n51997 = pi20 ? n37 : n20801;
  assign n51998 = pi19 ? n51996 : n51997;
  assign n51999 = pi18 ? n20563 : n51998;
  assign n52000 = pi17 ? n49894 : n51999;
  assign n52001 = pi16 ? n32 : n52000;
  assign n52002 = pi17 ? n49894 : n51472;
  assign n52003 = pi16 ? n32 : n52002;
  assign n52004 = pi15 ? n52001 : n52003;
  assign n52005 = pi14 ? n51995 : n52004;
  assign n52006 = pi13 ? n51985 : n52005;
  assign n52007 = pi20 ? n37 : n8261;
  assign n52008 = pi19 ? n32898 : n52007;
  assign n52009 = pi18 ? n20563 : n52008;
  assign n52010 = pi17 ? n50905 : n52009;
  assign n52011 = pi16 ? n32 : n52010;
  assign n52012 = pi20 ? n649 : n34943;
  assign n52013 = pi19 ? n32348 : n52012;
  assign n52014 = pi18 ? n20563 : n52013;
  assign n52015 = pi17 ? n49440 : n52014;
  assign n52016 = pi16 ? n32 : n52015;
  assign n52017 = pi15 ? n52011 : n52016;
  assign n52018 = pi20 ? n31220 : n36250;
  assign n52019 = pi20 ? n649 : n6214;
  assign n52020 = pi19 ? n52018 : n52019;
  assign n52021 = pi18 ? n20563 : n52020;
  assign n52022 = pi17 ? n49448 : n52021;
  assign n52023 = pi16 ? n32 : n52022;
  assign n52024 = pi20 ? n3393 : n34952;
  assign n52025 = pi19 ? n31221 : n52024;
  assign n52026 = pi18 ? n20563 : n52025;
  assign n52027 = pi17 ? n48904 : n52026;
  assign n52028 = pi16 ? n32 : n52027;
  assign n52029 = pi15 ? n52023 : n52028;
  assign n52030 = pi14 ? n52017 : n52029;
  assign n52031 = pi22 ? n3944 : n532;
  assign n52032 = pi21 ? n52031 : n32;
  assign n52033 = pi20 ? n37 : n52032;
  assign n52034 = pi19 ? n32898 : n52033;
  assign n52035 = pi18 ? n20563 : n52034;
  assign n52036 = pi17 ? n48904 : n52035;
  assign n52037 = pi16 ? n32 : n52036;
  assign n52038 = pi22 ? n3472 : n1407;
  assign n52039 = pi21 ? n52038 : n32;
  assign n52040 = pi20 ? n37 : n52039;
  assign n52041 = pi19 ? n32898 : n52040;
  assign n52042 = pi18 ? n20563 : n52041;
  assign n52043 = pi17 ? n48912 : n52042;
  assign n52044 = pi16 ? n32 : n52043;
  assign n52045 = pi15 ? n52037 : n52044;
  assign n52046 = pi20 ? n37 : n9456;
  assign n52047 = pi19 ? n31267 : n52046;
  assign n52048 = pi18 ? n20563 : n52047;
  assign n52049 = pi17 ? n49938 : n52048;
  assign n52050 = pi16 ? n32 : n52049;
  assign n52051 = pi19 ? n31280 : n52046;
  assign n52052 = pi18 ? n20563 : n52051;
  assign n52053 = pi17 ? n48466 : n52052;
  assign n52054 = pi16 ? n32 : n52053;
  assign n52055 = pi15 ? n52050 : n52054;
  assign n52056 = pi14 ? n52045 : n52055;
  assign n52057 = pi13 ? n52030 : n52056;
  assign n52058 = pi12 ? n52006 : n52057;
  assign n52059 = pi19 ? n32348 : n22873;
  assign n52060 = pi18 ? n20563 : n52059;
  assign n52061 = pi17 ? n48466 : n52060;
  assign n52062 = pi16 ? n32 : n52061;
  assign n52063 = pi22 ? n3944 : n706;
  assign n52064 = pi21 ? n52063 : n32;
  assign n52065 = pi20 ? n7730 : n52064;
  assign n52066 = pi19 ? n32898 : n52065;
  assign n52067 = pi18 ? n20563 : n52066;
  assign n52068 = pi17 ? n48466 : n52067;
  assign n52069 = pi16 ? n32 : n52068;
  assign n52070 = pi15 ? n52062 : n52069;
  assign n52071 = pi20 ? n7730 : n14352;
  assign n52072 = pi19 ? n32898 : n52071;
  assign n52073 = pi18 ? n20563 : n52072;
  assign n52074 = pi17 ? n48466 : n52073;
  assign n52075 = pi16 ? n32 : n52074;
  assign n52076 = pi22 ? n5061 : n32;
  assign n52077 = pi21 ? n52076 : n32;
  assign n52078 = pi20 ? n5013 : n52077;
  assign n52079 = pi19 ? n32348 : n52078;
  assign n52080 = pi18 ? n20563 : n52079;
  assign n52081 = pi17 ? n48469 : n52080;
  assign n52082 = pi16 ? n32 : n52081;
  assign n52083 = pi15 ? n52075 : n52082;
  assign n52084 = pi14 ? n52070 : n52083;
  assign n52085 = pi20 ? n5077 : n7035;
  assign n52086 = pi19 ? n31267 : n52085;
  assign n52087 = pi18 ? n20563 : n52086;
  assign n52088 = pi17 ? n47922 : n52087;
  assign n52089 = pi16 ? n32 : n52088;
  assign n52090 = pi20 ? n25804 : n3210;
  assign n52091 = pi19 ? n31267 : n52090;
  assign n52092 = pi18 ? n20563 : n52091;
  assign n52093 = pi17 ? n47922 : n52092;
  assign n52094 = pi16 ? n32 : n52093;
  assign n52095 = pi15 ? n52089 : n52094;
  assign n52096 = pi20 ? n24493 : n3210;
  assign n52097 = pi19 ? n31267 : n52096;
  assign n52098 = pi18 ? n20563 : n52097;
  assign n52099 = pi17 ? n47922 : n52098;
  assign n52100 = pi16 ? n32 : n52099;
  assign n52101 = pi14 ? n52095 : n52100;
  assign n52102 = pi13 ? n52084 : n52101;
  assign n52103 = pi21 ? n181 : n20977;
  assign n52104 = pi20 ? n52103 : n3210;
  assign n52105 = pi19 ? n32348 : n52104;
  assign n52106 = pi18 ? n20563 : n52105;
  assign n52107 = pi17 ? n47929 : n52106;
  assign n52108 = pi16 ? n32 : n52107;
  assign n52109 = pi21 ? n99 : n48364;
  assign n52110 = pi20 ? n52109 : n10011;
  assign n52111 = pi19 ? n45406 : n52110;
  assign n52112 = pi18 ? n20563 : n52111;
  assign n52113 = pi17 ? n47935 : n52112;
  assign n52114 = pi16 ? n32 : n52113;
  assign n52115 = pi15 ? n52108 : n52114;
  assign n52116 = pi19 ? n37618 : n52110;
  assign n52117 = pi18 ? n20563 : n52116;
  assign n52118 = pi17 ? n48949 : n52117;
  assign n52119 = pi16 ? n32 : n52118;
  assign n52120 = pi19 ? n45406 : n50546;
  assign n52121 = pi18 ? n20563 : n52120;
  assign n52122 = pi17 ? n48949 : n52121;
  assign n52123 = pi16 ? n32 : n52122;
  assign n52124 = pi15 ? n52119 : n52123;
  assign n52125 = pi14 ? n52115 : n52124;
  assign n52126 = pi20 ? n24957 : n2679;
  assign n52127 = pi19 ? n45406 : n52126;
  assign n52128 = pi18 ? n20563 : n52127;
  assign n52129 = pi17 ? n47954 : n52128;
  assign n52130 = pi16 ? n32 : n52129;
  assign n52131 = pi21 ? n36489 : n29133;
  assign n52132 = pi20 ? n52131 : n99;
  assign n52133 = pi19 ? n52132 : n52126;
  assign n52134 = pi18 ? n51078 : n52133;
  assign n52135 = pi17 ? n47954 : n52134;
  assign n52136 = pi16 ? n32 : n52135;
  assign n52137 = pi15 ? n52130 : n52136;
  assign n52138 = pi20 ? n51614 : n2701;
  assign n52139 = pi19 ? n39128 : n52138;
  assign n52140 = pi18 ? n20563 : n52139;
  assign n52141 = pi17 ? n48488 : n52140;
  assign n52142 = pi16 ? n32 : n52141;
  assign n52143 = pi21 ? n916 : n8842;
  assign n52144 = pi20 ? n52143 : n1822;
  assign n52145 = pi19 ? n31267 : n52144;
  assign n52146 = pi18 ? n20563 : n52145;
  assign n52147 = pi17 ? n47443 : n52146;
  assign n52148 = pi16 ? n32 : n52147;
  assign n52149 = pi15 ? n52142 : n52148;
  assign n52150 = pi14 ? n52137 : n52149;
  assign n52151 = pi13 ? n52125 : n52150;
  assign n52152 = pi12 ? n52102 : n52151;
  assign n52153 = pi11 ? n52058 : n52152;
  assign n52154 = pi21 ? n1056 : n11808;
  assign n52155 = pi20 ? n52154 : n1822;
  assign n52156 = pi19 ? n31280 : n52155;
  assign n52157 = pi18 ? n20563 : n52156;
  assign n52158 = pi17 ? n47443 : n52157;
  assign n52159 = pi16 ? n32 : n52158;
  assign n52160 = pi20 ? n31220 : n3096;
  assign n52161 = pi21 ? n919 : n3763;
  assign n52162 = pi20 ? n52161 : n32;
  assign n52163 = pi19 ? n52160 : n52162;
  assign n52164 = pi18 ? n20563 : n52163;
  assign n52165 = pi17 ? n46302 : n52164;
  assign n52166 = pi16 ? n32 : n52165;
  assign n52167 = pi15 ? n52159 : n52166;
  assign n52168 = pi19 ? n20563 : n50101;
  assign n52169 = pi21 ? n39801 : n37;
  assign n52170 = pi20 ? n52169 : n3096;
  assign n52171 = pi21 ? n919 : n16438;
  assign n52172 = pi20 ? n52171 : n32;
  assign n52173 = pi19 ? n52170 : n52172;
  assign n52174 = pi18 ? n52168 : n52173;
  assign n52175 = pi17 ? n46302 : n52174;
  assign n52176 = pi16 ? n32 : n52175;
  assign n52177 = pi20 ? n31220 : n3086;
  assign n52178 = pi19 ? n52177 : n52172;
  assign n52179 = pi18 ? n20563 : n52178;
  assign n52180 = pi17 ? n46832 : n52179;
  assign n52181 = pi16 ? n32 : n52180;
  assign n52182 = pi15 ? n52176 : n52181;
  assign n52183 = pi14 ? n52167 : n52182;
  assign n52184 = pi21 ? n1793 : n36058;
  assign n52185 = pi20 ? n52184 : n32;
  assign n52186 = pi19 ? n52177 : n52185;
  assign n52187 = pi18 ? n20563 : n52186;
  assign n52188 = pi17 ? n47964 : n52187;
  assign n52189 = pi16 ? n32 : n52188;
  assign n52190 = pi21 ? n9828 : n14168;
  assign n52191 = pi20 ? n52190 : n32;
  assign n52192 = pi19 ? n52160 : n52191;
  assign n52193 = pi18 ? n20563 : n52192;
  assign n52194 = pi17 ? n47964 : n52193;
  assign n52195 = pi16 ? n32 : n52194;
  assign n52196 = pi15 ? n52189 : n52195;
  assign n52197 = pi20 ? n31220 : n577;
  assign n52198 = pi19 ? n52197 : n51665;
  assign n52199 = pi18 ? n20563 : n52198;
  assign n52200 = pi17 ? n46839 : n52199;
  assign n52201 = pi16 ? n32 : n52200;
  assign n52202 = pi21 ? n2061 : n6366;
  assign n52203 = pi20 ? n52202 : n32;
  assign n52204 = pi19 ? n52197 : n52203;
  assign n52205 = pi18 ? n20563 : n52204;
  assign n52206 = pi17 ? n46839 : n52205;
  assign n52207 = pi16 ? n32 : n52206;
  assign n52208 = pi15 ? n52201 : n52207;
  assign n52209 = pi14 ? n52196 : n52208;
  assign n52210 = pi13 ? n52183 : n52209;
  assign n52211 = pi21 ? n2061 : n29061;
  assign n52212 = pi20 ? n52211 : n32;
  assign n52213 = pi19 ? n31280 : n52212;
  assign n52214 = pi18 ? n20563 : n52213;
  assign n52215 = pi17 ? n46839 : n52214;
  assign n52216 = pi16 ? n32 : n52215;
  assign n52217 = pi22 ? n99 : n2060;
  assign n52218 = pi21 ? n52217 : n4101;
  assign n52219 = pi20 ? n52218 : n32;
  assign n52220 = pi19 ? n31267 : n52219;
  assign n52221 = pi18 ? n20563 : n52220;
  assign n52222 = pi17 ? n45715 : n52221;
  assign n52223 = pi16 ? n32 : n52222;
  assign n52224 = pi15 ? n52216 : n52223;
  assign n52225 = pi20 ? n30096 : n649;
  assign n52226 = pi19 ? n52225 : n20549;
  assign n52227 = pi18 ? n20563 : n52226;
  assign n52228 = pi17 ? n45707 : n52227;
  assign n52229 = pi16 ? n32 : n52228;
  assign n52230 = pi20 ? n48254 : n30868;
  assign n52231 = pi21 ? n40912 : n36489;
  assign n52232 = pi20 ? n40915 : n52231;
  assign n52233 = pi19 ? n52230 : n52232;
  assign n52234 = pi21 ? n40912 : n39801;
  assign n52235 = pi20 ? n52234 : n51187;
  assign n52236 = pi21 ? n45049 : n40912;
  assign n52237 = pi20 ? n52234 : n52236;
  assign n52238 = pi19 ? n52235 : n52237;
  assign n52239 = pi18 ? n52233 : n52238;
  assign n52240 = pi17 ? n52239 : n52227;
  assign n52241 = pi16 ? n32 : n52240;
  assign n52242 = pi15 ? n52229 : n52241;
  assign n52243 = pi14 ? n52224 : n52242;
  assign n52244 = pi21 ? n40960 : n30868;
  assign n52245 = pi20 ? n38376 : n52244;
  assign n52246 = pi22 ? n30868 : n37173;
  assign n52247 = pi21 ? n52246 : n20563;
  assign n52248 = pi20 ? n52247 : n20563;
  assign n52249 = pi19 ? n52245 : n52248;
  assign n52250 = pi18 ? n52249 : n20563;
  assign n52251 = pi23 ? n685 : n14362;
  assign n52252 = pi22 ? n52251 : n32;
  assign n52253 = pi21 ? n233 : n52252;
  assign n52254 = pi20 ? n52253 : n32;
  assign n52255 = pi19 ? n7676 : n52254;
  assign n52256 = pi18 ? n20563 : n52255;
  assign n52257 = pi17 ? n52250 : n52256;
  assign n52258 = pi16 ? n32 : n52257;
  assign n52259 = pi22 ? n32 : n33792;
  assign n52260 = pi21 ? n52259 : n33792;
  assign n52261 = pi20 ? n52260 : n33792;
  assign n52262 = pi19 ? n52261 : n33792;
  assign n52263 = pi19 ? n40958 : n33792;
  assign n52264 = pi18 ? n52262 : n52263;
  assign n52265 = pi20 ? n45016 : n20563;
  assign n52266 = pi19 ? n52265 : n34246;
  assign n52267 = pi19 ? n8802 : n19353;
  assign n52268 = pi18 ? n52266 : n52267;
  assign n52269 = pi17 ? n52264 : n52268;
  assign n52270 = pi16 ? n32 : n52269;
  assign n52271 = pi15 ? n52258 : n52270;
  assign n52272 = pi21 ? n29133 : n584;
  assign n52273 = pi20 ? n37308 : n52272;
  assign n52274 = pi19 ? n52273 : n14724;
  assign n52275 = pi18 ? n20563 : n52274;
  assign n52276 = pi17 ? n46312 : n52275;
  assign n52277 = pi16 ? n32 : n52276;
  assign n52278 = pi19 ? n6403 : n51771;
  assign n52279 = pi18 ? n20563 : n52278;
  assign n52280 = pi17 ? n46312 : n52279;
  assign n52281 = pi16 ? n32 : n52280;
  assign n52282 = pi15 ? n52277 : n52281;
  assign n52283 = pi14 ? n52271 : n52282;
  assign n52284 = pi13 ? n52243 : n52283;
  assign n52285 = pi12 ? n52210 : n52284;
  assign n52286 = pi19 ? n6403 : n12515;
  assign n52287 = pi18 ? n20563 : n52286;
  assign n52288 = pi17 ? n46312 : n52287;
  assign n52289 = pi16 ? n32 : n52288;
  assign n52290 = pi23 ? n20627 : n335;
  assign n52291 = pi22 ? n37 : n52290;
  assign n52292 = pi21 ? n37 : n52291;
  assign n52293 = pi20 ? n30096 : n52292;
  assign n52294 = pi20 ? n38879 : n32;
  assign n52295 = pi19 ? n52293 : n52294;
  assign n52296 = pi18 ? n20563 : n52295;
  assign n52297 = pi17 ? n46312 : n52296;
  assign n52298 = pi16 ? n32 : n52297;
  assign n52299 = pi15 ? n52289 : n52298;
  assign n52300 = pi20 ? n30096 : n363;
  assign n52301 = pi19 ? n52300 : n9464;
  assign n52302 = pi18 ? n20563 : n52301;
  assign n52303 = pi17 ? n46866 : n52302;
  assign n52304 = pi16 ? n32 : n52303;
  assign n52305 = pi20 ? n43010 : n38754;
  assign n52306 = pi19 ? n20563 : n52305;
  assign n52307 = pi23 ? n3491 : n363;
  assign n52308 = pi22 ? n37 : n52307;
  assign n52309 = pi21 ? n363 : n52308;
  assign n52310 = pi20 ? n30096 : n52309;
  assign n52311 = pi22 ? n1457 : n317;
  assign n52312 = pi21 ? n52311 : n32;
  assign n52313 = pi20 ? n52312 : n32;
  assign n52314 = pi19 ? n52310 : n52313;
  assign n52315 = pi18 ? n52306 : n52314;
  assign n52316 = pi17 ? n46859 : n52315;
  assign n52317 = pi16 ? n32 : n52316;
  assign n52318 = pi15 ? n52304 : n52317;
  assign n52319 = pi14 ? n52299 : n52318;
  assign n52320 = pi22 ? n363 : n861;
  assign n52321 = pi21 ? n37 : n52320;
  assign n52322 = pi20 ? n30096 : n52321;
  assign n52323 = pi21 ? n4296 : n32;
  assign n52324 = pi20 ? n52323 : n32;
  assign n52325 = pi19 ? n52322 : n52324;
  assign n52326 = pi18 ? n20563 : n52325;
  assign n52327 = pi17 ? n46859 : n52326;
  assign n52328 = pi16 ? n32 : n52327;
  assign n52329 = pi20 ? n51280 : n47158;
  assign n52330 = pi19 ? n20563 : n52329;
  assign n52331 = pi20 ? n30096 : n51274;
  assign n52332 = pi19 ? n52331 : n40815;
  assign n52333 = pi18 ? n52330 : n52332;
  assign n52334 = pi17 ? n46859 : n52333;
  assign n52335 = pi16 ? n32 : n52334;
  assign n52336 = pi15 ? n52328 : n52335;
  assign n52337 = pi21 ? n39394 : n48173;
  assign n52338 = pi20 ? n52337 : n30868;
  assign n52339 = pi21 ? n36489 : n39801;
  assign n52340 = pi20 ? n52339 : n20563;
  assign n52341 = pi19 ? n52338 : n52340;
  assign n52342 = pi18 ? n52341 : n20563;
  assign n52343 = pi22 ? n363 : n448;
  assign n52344 = pi21 ? n99 : n52343;
  assign n52345 = pi20 ? n31220 : n52344;
  assign n52346 = pi19 ? n52345 : n9483;
  assign n52347 = pi18 ? n20563 : n52346;
  assign n52348 = pi17 ? n52342 : n52347;
  assign n52349 = pi16 ? n32 : n52348;
  assign n52350 = pi20 ? n39395 : n30868;
  assign n52351 = pi19 ? n52350 : n20563;
  assign n52352 = pi18 ? n52351 : n20563;
  assign n52353 = pi22 ? n335 : n18448;
  assign n52354 = pi21 ? n3392 : n52353;
  assign n52355 = pi20 ? n31220 : n52354;
  assign n52356 = pi19 ? n52355 : n3211;
  assign n52357 = pi18 ? n20563 : n52356;
  assign n52358 = pi17 ? n52352 : n52357;
  assign n52359 = pi16 ? n32 : n52358;
  assign n52360 = pi15 ? n52349 : n52359;
  assign n52361 = pi14 ? n52336 : n52360;
  assign n52362 = pi13 ? n52319 : n52361;
  assign n52363 = pi20 ? n45621 : n30868;
  assign n52364 = pi19 ? n52363 : n30868;
  assign n52365 = pi18 ? n52364 : n30868;
  assign n52366 = pi21 ? n139 : n45681;
  assign n52367 = pi20 ? n38250 : n52366;
  assign n52368 = pi19 ? n52367 : n3211;
  assign n52369 = pi18 ? n30868 : n52368;
  assign n52370 = pi17 ? n52365 : n52369;
  assign n52371 = pi16 ? n32 : n52370;
  assign n52372 = pi21 ? n30868 : n746;
  assign n52373 = pi22 ? n157 : n233;
  assign n52374 = pi21 ? n777 : n52373;
  assign n52375 = pi20 ? n52372 : n52374;
  assign n52376 = pi19 ? n52375 : n10012;
  assign n52377 = pi18 ? n30868 : n52376;
  assign n52378 = pi17 ? n52365 : n52377;
  assign n52379 = pi16 ? n32 : n52378;
  assign n52380 = pi15 ? n52371 : n52379;
  assign n52381 = pi20 ? n45654 : n36798;
  assign n52382 = pi19 ? n52381 : n36798;
  assign n52383 = pi18 ? n52382 : n36798;
  assign n52384 = pi20 ? n33792 : n50300;
  assign n52385 = pi19 ? n46204 : n52384;
  assign n52386 = pi20 ? n48377 : n47371;
  assign n52387 = pi19 ? n52386 : n2654;
  assign n52388 = pi18 ? n52385 : n52387;
  assign n52389 = pi17 ? n52383 : n52388;
  assign n52390 = pi16 ? n32 : n52389;
  assign n52391 = pi23 ? n36782 : n33792;
  assign n52392 = pi22 ? n52391 : n33792;
  assign n52393 = pi21 ? n32 : n52392;
  assign n52394 = pi20 ? n52393 : n33792;
  assign n52395 = pi23 ? n33792 : n36781;
  assign n52396 = pi22 ? n33792 : n52395;
  assign n52397 = pi21 ? n52396 : n33792;
  assign n52398 = pi20 ? n52397 : n33792;
  assign n52399 = pi19 ? n52394 : n52398;
  assign n52400 = pi18 ? n52399 : n33792;
  assign n52401 = pi18 ? n33792 : n52387;
  assign n52402 = pi17 ? n52400 : n52401;
  assign n52403 = pi16 ? n32 : n52402;
  assign n52404 = pi15 ? n52390 : n52403;
  assign n52405 = pi14 ? n52380 : n52404;
  assign n52406 = pi20 ? n48436 : n43198;
  assign n52407 = pi19 ? n52406 : n49391;
  assign n52408 = pi18 ? n52407 : n36659;
  assign n52409 = pi21 ? n335 : n1027;
  assign n52410 = pi20 ? n48393 : n52409;
  assign n52411 = pi19 ? n52410 : n1823;
  assign n52412 = pi18 ? n36659 : n52411;
  assign n52413 = pi17 ? n52408 : n52412;
  assign n52414 = pi16 ? n32 : n52413;
  assign n52415 = pi23 ? n36830 : n36659;
  assign n52416 = pi22 ? n52415 : n36659;
  assign n52417 = pi21 ? n32 : n52416;
  assign n52418 = pi20 ? n52417 : n36659;
  assign n52419 = pi19 ? n52418 : n49835;
  assign n52420 = pi18 ? n52419 : n36659;
  assign n52421 = pi23 ? n363 : n36659;
  assign n52422 = pi22 ? n52421 : n18461;
  assign n52423 = pi21 ? n36659 : n52422;
  assign n52424 = pi21 ? n7986 : n25977;
  assign n52425 = pi20 ? n52423 : n52424;
  assign n52426 = pi19 ? n52425 : n32;
  assign n52427 = pi18 ? n36659 : n52426;
  assign n52428 = pi17 ? n52420 : n52427;
  assign n52429 = pi16 ? n32 : n52428;
  assign n52430 = pi15 ? n52414 : n52429;
  assign n52431 = pi23 ? n46274 : n36781;
  assign n52432 = pi22 ? n52431 : n36781;
  assign n52433 = pi21 ? n32 : n52432;
  assign n52434 = pi20 ? n52433 : n42170;
  assign n52435 = pi21 ? n43200 : n36781;
  assign n52436 = pi20 ? n52435 : n36781;
  assign n52437 = pi19 ? n52434 : n52436;
  assign n52438 = pi18 ? n52437 : n36781;
  assign n52439 = pi21 ? n36781 : n40441;
  assign n52440 = pi21 ? n5054 : n397;
  assign n52441 = pi20 ? n52439 : n52440;
  assign n52442 = pi19 ? n52441 : n32;
  assign n52443 = pi18 ? n36781 : n52442;
  assign n52444 = pi17 ? n52438 : n52443;
  assign n52445 = pi16 ? n32 : n52444;
  assign n52446 = pi20 ? n50810 : n43198;
  assign n52447 = pi21 ? n43198 : n46283;
  assign n52448 = pi20 ? n52447 : n36781;
  assign n52449 = pi19 ? n52446 : n52448;
  assign n52450 = pi18 ? n52449 : n36781;
  assign n52451 = pi23 ? n157 : n36798;
  assign n52452 = pi22 ? n36798 : n52451;
  assign n52453 = pi21 ? n36781 : n52452;
  assign n52454 = pi20 ? n52453 : n20106;
  assign n52455 = pi19 ? n52454 : n32;
  assign n52456 = pi18 ? n51395 : n52455;
  assign n52457 = pi17 ? n52450 : n52456;
  assign n52458 = pi16 ? n32 : n52457;
  assign n52459 = pi15 ? n52445 : n52458;
  assign n52460 = pi14 ? n52430 : n52459;
  assign n52461 = pi13 ? n52405 : n52460;
  assign n52462 = pi12 ? n52362 : n52461;
  assign n52463 = pi11 ? n52285 : n52462;
  assign n52464 = pi10 ? n52153 : n52463;
  assign n52465 = pi09 ? n51952 : n52464;
  assign n52466 = pi17 ? n39398 : n51928;
  assign n52467 = pi16 ? n32 : n52466;
  assign n52468 = pi15 ? n32 : n52467;
  assign n52469 = pi18 ? n51933 : n51927;
  assign n52470 = pi17 ? n40551 : n52469;
  assign n52471 = pi16 ? n32 : n52470;
  assign n52472 = pi22 ? n139 : n2026;
  assign n52473 = pi21 ? n52472 : n32;
  assign n52474 = pi20 ? n37 : n52473;
  assign n52475 = pi19 ? n37 : n52474;
  assign n52476 = pi18 ? n34295 : n52475;
  assign n52477 = pi17 ? n38330 : n52476;
  assign n52478 = pi16 ? n32 : n52477;
  assign n52479 = pi15 ? n52471 : n52478;
  assign n52480 = pi14 ? n52468 : n52479;
  assign n52481 = pi13 ? n32 : n52480;
  assign n52482 = pi12 ? n32 : n52481;
  assign n52483 = pi11 ? n32 : n52482;
  assign n52484 = pi10 ? n32 : n52483;
  assign n52485 = pi22 ? n37 : n10164;
  assign n52486 = pi21 ? n52485 : n32;
  assign n52487 = pi20 ? n8742 : n52486;
  assign n52488 = pi19 ? n51953 : n52487;
  assign n52489 = pi18 ? n34258 : n52488;
  assign n52490 = pi17 ? n36870 : n52489;
  assign n52491 = pi16 ? n32 : n52490;
  assign n52492 = pi21 ? n43713 : n32;
  assign n52493 = pi20 ? n3086 : n52492;
  assign n52494 = pi19 ? n50883 : n52493;
  assign n52495 = pi18 ? n34869 : n52494;
  assign n52496 = pi17 ? n36870 : n52495;
  assign n52497 = pi16 ? n32 : n52496;
  assign n52498 = pi15 ? n52491 : n52497;
  assign n52499 = pi22 ? n37 : n1217;
  assign n52500 = pi21 ? n52499 : n32;
  assign n52501 = pi20 ? n37 : n52500;
  assign n52502 = pi19 ? n37 : n52501;
  assign n52503 = pi18 ? n34295 : n52502;
  assign n52504 = pi17 ? n39000 : n52503;
  assign n52505 = pi16 ? n32 : n52504;
  assign n52506 = pi20 ? n37 : n35792;
  assign n52507 = pi19 ? n37 : n52506;
  assign n52508 = pi18 ? n50907 : n52507;
  assign n52509 = pi17 ? n37336 : n52508;
  assign n52510 = pi16 ? n32 : n52509;
  assign n52511 = pi15 ? n52505 : n52510;
  assign n52512 = pi14 ? n52498 : n52511;
  assign n52513 = pi20 ? n37 : n6079;
  assign n52514 = pi19 ? n37 : n52513;
  assign n52515 = pi18 ? n34295 : n52514;
  assign n52516 = pi17 ? n37336 : n52515;
  assign n52517 = pi16 ? n32 : n52516;
  assign n52518 = pi20 ? n37 : n37439;
  assign n52519 = pi20 ? n37 : n22279;
  assign n52520 = pi19 ? n52518 : n52519;
  assign n52521 = pi18 ? n34869 : n52520;
  assign n52522 = pi17 ? n36215 : n52521;
  assign n52523 = pi16 ? n32 : n52522;
  assign n52524 = pi15 ? n52517 : n52523;
  assign n52525 = pi20 ? n37 : n21760;
  assign n52526 = pi19 ? n51996 : n52525;
  assign n52527 = pi18 ? n20563 : n52526;
  assign n52528 = pi17 ? n36215 : n52527;
  assign n52529 = pi16 ? n32 : n52528;
  assign n52530 = pi20 ? n649 : n21760;
  assign n52531 = pi19 ? n50932 : n52530;
  assign n52532 = pi18 ? n20563 : n52531;
  assign n52533 = pi17 ? n50390 : n52532;
  assign n52534 = pi16 ? n32 : n52533;
  assign n52535 = pi15 ? n52529 : n52534;
  assign n52536 = pi14 ? n52524 : n52535;
  assign n52537 = pi13 ? n52512 : n52536;
  assign n52538 = pi20 ? n37 : n9414;
  assign n52539 = pi19 ? n32898 : n52538;
  assign n52540 = pi18 ? n20563 : n52539;
  assign n52541 = pi17 ? n50393 : n52540;
  assign n52542 = pi16 ? n32 : n52541;
  assign n52543 = pi20 ? n649 : n9926;
  assign n52544 = pi19 ? n32348 : n52543;
  assign n52545 = pi18 ? n20563 : n52544;
  assign n52546 = pi17 ? n49888 : n52545;
  assign n52547 = pi16 ? n32 : n52546;
  assign n52548 = pi15 ? n52542 : n52547;
  assign n52549 = pi20 ? n649 : n35840;
  assign n52550 = pi19 ? n52018 : n52549;
  assign n52551 = pi18 ? n20563 : n52550;
  assign n52552 = pi17 ? n49894 : n52551;
  assign n52553 = pi16 ? n32 : n52552;
  assign n52554 = pi21 ? n12731 : n32;
  assign n52555 = pi20 ? n3393 : n52554;
  assign n52556 = pi19 ? n31221 : n52555;
  assign n52557 = pi18 ? n20563 : n52556;
  assign n52558 = pi17 ? n49448 : n52557;
  assign n52559 = pi16 ? n32 : n52558;
  assign n52560 = pi15 ? n52553 : n52559;
  assign n52561 = pi14 ? n52548 : n52560;
  assign n52562 = pi22 ? n3944 : n2564;
  assign n52563 = pi21 ? n52562 : n32;
  assign n52564 = pi20 ? n37 : n52563;
  assign n52565 = pi19 ? n32898 : n52564;
  assign n52566 = pi18 ? n20563 : n52565;
  assign n52567 = pi17 ? n49448 : n52566;
  assign n52568 = pi16 ? n32 : n52567;
  assign n52569 = pi21 ? n16230 : n32;
  assign n52570 = pi20 ? n37 : n52569;
  assign n52571 = pi19 ? n32898 : n52570;
  assign n52572 = pi18 ? n20563 : n52571;
  assign n52573 = pi17 ? n49451 : n52572;
  assign n52574 = pi16 ? n32 : n52573;
  assign n52575 = pi15 ? n52568 : n52574;
  assign n52576 = pi17 ? n50426 : n52048;
  assign n52577 = pi16 ? n32 : n52576;
  assign n52578 = pi17 ? n48904 : n52052;
  assign n52579 = pi16 ? n32 : n52578;
  assign n52580 = pi15 ? n52577 : n52579;
  assign n52581 = pi14 ? n52575 : n52580;
  assign n52582 = pi13 ? n52561 : n52581;
  assign n52583 = pi12 ? n52537 : n52582;
  assign n52584 = pi19 ? n31904 : n22873;
  assign n52585 = pi18 ? n20563 : n52584;
  assign n52586 = pi17 ? n48904 : n52585;
  assign n52587 = pi16 ? n32 : n52586;
  assign n52588 = pi17 ? n48904 : n52067;
  assign n52589 = pi16 ? n32 : n52588;
  assign n52590 = pi15 ? n52587 : n52589;
  assign n52591 = pi17 ? n48904 : n52073;
  assign n52592 = pi16 ? n32 : n52591;
  assign n52593 = pi17 ? n48912 : n52080;
  assign n52594 = pi16 ? n32 : n52593;
  assign n52595 = pi15 ? n52592 : n52594;
  assign n52596 = pi14 ? n52590 : n52595;
  assign n52597 = pi17 ? n48460 : n52087;
  assign n52598 = pi16 ? n32 : n52597;
  assign n52599 = pi17 ? n48460 : n52092;
  assign n52600 = pi16 ? n32 : n52599;
  assign n52601 = pi15 ? n52598 : n52600;
  assign n52602 = pi17 ? n48460 : n52098;
  assign n52603 = pi16 ? n32 : n52602;
  assign n52604 = pi14 ? n52601 : n52603;
  assign n52605 = pi13 ? n52596 : n52604;
  assign n52606 = pi20 ? n52103 : n4008;
  assign n52607 = pi19 ? n31904 : n52606;
  assign n52608 = pi18 ? n20563 : n52607;
  assign n52609 = pi17 ? n48466 : n52608;
  assign n52610 = pi16 ? n32 : n52609;
  assign n52611 = pi18 ? n41168 : n20563;
  assign n52612 = pi20 ? n52109 : n3210;
  assign n52613 = pi19 ? n39670 : n52612;
  assign n52614 = pi18 ? n20563 : n52613;
  assign n52615 = pi17 ? n52611 : n52614;
  assign n52616 = pi16 ? n32 : n52615;
  assign n52617 = pi15 ? n52610 : n52616;
  assign n52618 = pi19 ? n37618 : n52612;
  assign n52619 = pi18 ? n20563 : n52618;
  assign n52620 = pi17 ? n52611 : n52619;
  assign n52621 = pi16 ? n32 : n52620;
  assign n52622 = pi19 ? n45406 : n24958;
  assign n52623 = pi18 ? n20563 : n52622;
  assign n52624 = pi17 ? n52611 : n52623;
  assign n52625 = pi16 ? n32 : n52624;
  assign n52626 = pi15 ? n52621 : n52625;
  assign n52627 = pi14 ? n52617 : n52626;
  assign n52628 = pi19 ? n39670 : n50546;
  assign n52629 = pi18 ? n20563 : n52628;
  assign n52630 = pi17 ? n52611 : n52629;
  assign n52631 = pi16 ? n32 : n52630;
  assign n52632 = pi22 ? n20563 : n30869;
  assign n52633 = pi21 ? n36489 : n52632;
  assign n52634 = pi20 ? n52633 : n99;
  assign n52635 = pi19 ? n52634 : n50546;
  assign n52636 = pi18 ? n51078 : n52635;
  assign n52637 = pi17 ? n52611 : n52636;
  assign n52638 = pi16 ? n32 : n52637;
  assign n52639 = pi15 ? n52631 : n52638;
  assign n52640 = pi20 ? n32313 : n5077;
  assign n52641 = pi20 ? n51614 : n2679;
  assign n52642 = pi19 ? n52640 : n52641;
  assign n52643 = pi18 ? n20563 : n52642;
  assign n52644 = pi17 ? n47922 : n52643;
  assign n52645 = pi16 ? n32 : n52644;
  assign n52646 = pi21 ? n916 : n46526;
  assign n52647 = pi20 ? n52646 : n2701;
  assign n52648 = pi19 ? n31267 : n52647;
  assign n52649 = pi18 ? n20563 : n52648;
  assign n52650 = pi17 ? n47935 : n52649;
  assign n52651 = pi16 ? n32 : n52650;
  assign n52652 = pi15 ? n52645 : n52651;
  assign n52653 = pi14 ? n52639 : n52652;
  assign n52654 = pi13 ? n52627 : n52653;
  assign n52655 = pi12 ? n52605 : n52654;
  assign n52656 = pi11 ? n52583 : n52655;
  assign n52657 = pi19 ? n32871 : n52155;
  assign n52658 = pi18 ? n20563 : n52657;
  assign n52659 = pi17 ? n47935 : n52658;
  assign n52660 = pi16 ? n32 : n52659;
  assign n52661 = pi20 ? n34919 : n3096;
  assign n52662 = pi22 ? n204 : n27667;
  assign n52663 = pi21 ? n139 : n52662;
  assign n52664 = pi20 ? n52663 : n1822;
  assign n52665 = pi19 ? n52661 : n52664;
  assign n52666 = pi18 ? n20563 : n52665;
  assign n52667 = pi17 ? n47947 : n52666;
  assign n52668 = pi16 ? n32 : n52667;
  assign n52669 = pi15 ? n52660 : n52668;
  assign n52670 = pi21 ? n39801 : n30195;
  assign n52671 = pi20 ? n52670 : n3096;
  assign n52672 = pi24 ? n685 : n51564;
  assign n52673 = pi23 ? n204 : n52672;
  assign n52674 = pi22 ? n204 : n52673;
  assign n52675 = pi21 ? n139 : n52674;
  assign n52676 = pi20 ? n52675 : n32;
  assign n52677 = pi19 ? n52671 : n52676;
  assign n52678 = pi18 ? n52168 : n52677;
  assign n52679 = pi17 ? n47947 : n52678;
  assign n52680 = pi16 ? n32 : n52679;
  assign n52681 = pi21 ? n1531 : n16438;
  assign n52682 = pi20 ? n52681 : n32;
  assign n52683 = pi19 ? n52177 : n52682;
  assign n52684 = pi18 ? n20563 : n52683;
  assign n52685 = pi17 ? n48949 : n52684;
  assign n52686 = pi16 ? n32 : n52685;
  assign n52687 = pi15 ? n52680 : n52686;
  assign n52688 = pi14 ? n52669 : n52687;
  assign n52689 = pi22 ? n204 : n44992;
  assign n52690 = pi21 ? n1793 : n52689;
  assign n52691 = pi20 ? n52690 : n32;
  assign n52692 = pi19 ? n52177 : n52691;
  assign n52693 = pi18 ? n20563 : n52692;
  assign n52694 = pi17 ? n47954 : n52693;
  assign n52695 = pi16 ? n32 : n52694;
  assign n52696 = pi21 ? n9828 : n19726;
  assign n52697 = pi20 ? n52696 : n32;
  assign n52698 = pi19 ? n52160 : n52697;
  assign n52699 = pi18 ? n20563 : n52698;
  assign n52700 = pi17 ? n47954 : n52699;
  assign n52701 = pi16 ? n32 : n52700;
  assign n52702 = pi15 ? n52695 : n52701;
  assign n52703 = pi21 ? n14952 : n23543;
  assign n52704 = pi20 ? n52703 : n32;
  assign n52705 = pi19 ? n52197 : n52704;
  assign n52706 = pi18 ? n20563 : n52705;
  assign n52707 = pi17 ? n47443 : n52706;
  assign n52708 = pi16 ? n32 : n52707;
  assign n52709 = pi21 ? n2061 : n15889;
  assign n52710 = pi20 ? n52709 : n32;
  assign n52711 = pi19 ? n52197 : n52710;
  assign n52712 = pi18 ? n20563 : n52711;
  assign n52713 = pi17 ? n47443 : n52712;
  assign n52714 = pi16 ? n32 : n52713;
  assign n52715 = pi15 ? n52708 : n52714;
  assign n52716 = pi14 ? n52702 : n52715;
  assign n52717 = pi13 ? n52688 : n52716;
  assign n52718 = pi21 ? n2061 : n5758;
  assign n52719 = pi20 ? n52718 : n32;
  assign n52720 = pi19 ? n31280 : n52719;
  assign n52721 = pi18 ? n20563 : n52720;
  assign n52722 = pi17 ? n47443 : n52721;
  assign n52723 = pi16 ? n32 : n52722;
  assign n52724 = pi17 ? n46832 : n52221;
  assign n52725 = pi16 ? n32 : n52724;
  assign n52726 = pi15 ? n52723 : n52725;
  assign n52727 = pi20 ? n33821 : n649;
  assign n52728 = pi20 ? n38214 : n32;
  assign n52729 = pi19 ? n52727 : n52728;
  assign n52730 = pi18 ? n20563 : n52729;
  assign n52731 = pi17 ? n47451 : n52730;
  assign n52732 = pi16 ? n32 : n52731;
  assign n52733 = pi20 ? n46188 : n30868;
  assign n52734 = pi19 ? n52733 : n52232;
  assign n52735 = pi20 ? n52339 : n51187;
  assign n52736 = pi19 ? n52735 : n52237;
  assign n52737 = pi18 ? n52734 : n52736;
  assign n52738 = pi17 ? n52737 : n52730;
  assign n52739 = pi16 ? n32 : n52738;
  assign n52740 = pi15 ? n52732 : n52739;
  assign n52741 = pi14 ? n52726 : n52740;
  assign n52742 = pi22 ? n49720 : n33792;
  assign n52743 = pi21 ? n32 : n52742;
  assign n52744 = pi21 ? n36615 : n30868;
  assign n52745 = pi20 ? n52743 : n52744;
  assign n52746 = pi21 ? n52246 : n40954;
  assign n52747 = pi20 ? n52746 : n20563;
  assign n52748 = pi19 ? n52745 : n52747;
  assign n52749 = pi18 ? n52748 : n20563;
  assign n52750 = pi20 ? n31298 : n649;
  assign n52751 = pi19 ? n52750 : n52254;
  assign n52752 = pi18 ? n20563 : n52751;
  assign n52753 = pi17 ? n52749 : n52752;
  assign n52754 = pi16 ? n32 : n52753;
  assign n52755 = pi20 ? n52743 : n33792;
  assign n52756 = pi19 ? n52755 : n33792;
  assign n52757 = pi18 ? n52756 : n52263;
  assign n52758 = pi22 ? n20563 : n36617;
  assign n52759 = pi21 ? n20563 : n52758;
  assign n52760 = pi20 ? n20563 : n52759;
  assign n52761 = pi19 ? n52265 : n52760;
  assign n52762 = pi20 ? n31298 : n3299;
  assign n52763 = pi19 ? n52762 : n19353;
  assign n52764 = pi18 ? n52761 : n52763;
  assign n52765 = pi17 ? n52757 : n52764;
  assign n52766 = pi16 ? n32 : n52765;
  assign n52767 = pi15 ? n52754 : n52766;
  assign n52768 = pi17 ? n46859 : n52275;
  assign n52769 = pi16 ? n32 : n52768;
  assign n52770 = pi20 ? n31298 : n6402;
  assign n52771 = pi21 ? n5113 : n33225;
  assign n52772 = pi20 ? n52771 : n32;
  assign n52773 = pi19 ? n52770 : n52772;
  assign n52774 = pi18 ? n20563 : n52773;
  assign n52775 = pi17 ? n46839 : n52774;
  assign n52776 = pi16 ? n32 : n52775;
  assign n52777 = pi15 ? n52769 : n52776;
  assign n52778 = pi14 ? n52767 : n52777;
  assign n52779 = pi13 ? n52741 : n52778;
  assign n52780 = pi12 ? n52717 : n52779;
  assign n52781 = pi21 ? n3445 : n2700;
  assign n52782 = pi20 ? n52781 : n32;
  assign n52783 = pi19 ? n52770 : n52782;
  assign n52784 = pi18 ? n20563 : n52783;
  assign n52785 = pi17 ? n46839 : n52784;
  assign n52786 = pi16 ? n32 : n52785;
  assign n52787 = pi21 ? n37 : n21622;
  assign n52788 = pi20 ? n32286 : n52787;
  assign n52789 = pi19 ? n52788 : n13794;
  assign n52790 = pi18 ? n20563 : n52789;
  assign n52791 = pi17 ? n46839 : n52790;
  assign n52792 = pi16 ? n32 : n52791;
  assign n52793 = pi15 ? n52786 : n52792;
  assign n52794 = pi20 ? n32286 : n363;
  assign n52795 = pi22 ? n686 : n316;
  assign n52796 = pi21 ? n52795 : n32;
  assign n52797 = pi20 ? n52796 : n32;
  assign n52798 = pi19 ? n52794 : n52797;
  assign n52799 = pi18 ? n20563 : n52798;
  assign n52800 = pi17 ? n47964 : n52799;
  assign n52801 = pi16 ? n32 : n52800;
  assign n52802 = pi22 ? n37 : n364;
  assign n52803 = pi21 ? n363 : n52802;
  assign n52804 = pi20 ? n32286 : n52803;
  assign n52805 = pi22 ? n1457 : n316;
  assign n52806 = pi21 ? n52805 : n32;
  assign n52807 = pi20 ? n52806 : n32;
  assign n52808 = pi19 ? n52804 : n52807;
  assign n52809 = pi18 ? n52306 : n52808;
  assign n52810 = pi17 ? n47964 : n52809;
  assign n52811 = pi16 ? n32 : n52810;
  assign n52812 = pi15 ? n52801 : n52811;
  assign n52813 = pi14 ? n52793 : n52812;
  assign n52814 = pi20 ? n32286 : n52321;
  assign n52815 = pi22 ? n2244 : n21502;
  assign n52816 = pi21 ? n52815 : n32;
  assign n52817 = pi20 ? n52816 : n32;
  assign n52818 = pi19 ? n52814 : n52817;
  assign n52819 = pi18 ? n20563 : n52818;
  assign n52820 = pi17 ? n47964 : n52819;
  assign n52821 = pi16 ? n32 : n52820;
  assign n52822 = pi22 ? n40386 : n39190;
  assign n52823 = pi21 ? n52822 : n20563;
  assign n52824 = pi20 ? n48736 : n52823;
  assign n52825 = pi21 ? n39191 : n45049;
  assign n52826 = pi20 ? n52825 : n20563;
  assign n52827 = pi19 ? n52824 : n52826;
  assign n52828 = pi18 ? n52827 : n20563;
  assign n52829 = pi20 ? n32286 : n51274;
  assign n52830 = pi19 ? n52829 : n40815;
  assign n52831 = pi18 ? n52330 : n52830;
  assign n52832 = pi17 ? n52828 : n52831;
  assign n52833 = pi16 ? n32 : n52832;
  assign n52834 = pi15 ? n52821 : n52833;
  assign n52835 = pi20 ? n48736 : n30868;
  assign n52836 = pi19 ? n52835 : n52340;
  assign n52837 = pi18 ? n52836 : n20563;
  assign n52838 = pi17 ? n52837 : n52347;
  assign n52839 = pi16 ? n32 : n52838;
  assign n52840 = pi20 ? n36867 : n30868;
  assign n52841 = pi19 ? n52840 : n20563;
  assign n52842 = pi18 ? n52841 : n20563;
  assign n52843 = pi20 ? n35316 : n52354;
  assign n52844 = pi19 ? n52843 : n3211;
  assign n52845 = pi18 ? n20563 : n52844;
  assign n52846 = pi17 ? n52842 : n52845;
  assign n52847 = pi16 ? n32 : n52846;
  assign n52848 = pi15 ? n52839 : n52847;
  assign n52849 = pi14 ? n52834 : n52848;
  assign n52850 = pi13 ? n52813 : n52849;
  assign n52851 = pi20 ? n46167 : n30868;
  assign n52852 = pi19 ? n52851 : n30868;
  assign n52853 = pi18 ? n52852 : n30868;
  assign n52854 = pi17 ? n52853 : n52369;
  assign n52855 = pi16 ? n32 : n52854;
  assign n52856 = pi21 ? n30868 : n50759;
  assign n52857 = pi20 ? n52856 : n52374;
  assign n52858 = pi19 ? n52857 : n10012;
  assign n52859 = pi18 ? n30868 : n52858;
  assign n52860 = pi17 ? n52853 : n52859;
  assign n52861 = pi16 ? n32 : n52860;
  assign n52862 = pi15 ? n52855 : n52861;
  assign n52863 = pi21 ? n32 : n50767;
  assign n52864 = pi20 ? n52863 : n36798;
  assign n52865 = pi19 ? n52864 : n36798;
  assign n52866 = pi18 ? n52865 : n36798;
  assign n52867 = pi20 ? n32257 : n32;
  assign n52868 = pi19 ? n52386 : n52867;
  assign n52869 = pi18 ? n52385 : n52868;
  assign n52870 = pi17 ? n52866 : n52869;
  assign n52871 = pi16 ? n32 : n52870;
  assign n52872 = pi21 ? n32 : n50786;
  assign n52873 = pi23 ? n43198 : n33792;
  assign n52874 = pi22 ? n43198 : n52873;
  assign n52875 = pi23 ? n33792 : n43198;
  assign n52876 = pi22 ? n52875 : n33792;
  assign n52877 = pi21 ? n52874 : n52876;
  assign n52878 = pi20 ? n52872 : n52877;
  assign n52879 = pi22 ? n52875 : n52873;
  assign n52880 = pi21 ? n33792 : n52879;
  assign n52881 = pi20 ? n52880 : n33792;
  assign n52882 = pi19 ? n52878 : n52881;
  assign n52883 = pi18 ? n52882 : n33792;
  assign n52884 = pi20 ? n37842 : n47371;
  assign n52885 = pi19 ? n52884 : n2654;
  assign n52886 = pi18 ? n33792 : n52885;
  assign n52887 = pi17 ? n52883 : n52886;
  assign n52888 = pi16 ? n32 : n52887;
  assign n52889 = pi15 ? n52871 : n52888;
  assign n52890 = pi14 ? n52862 : n52889;
  assign n52891 = pi20 ? n52872 : n43198;
  assign n52892 = pi19 ? n52891 : n49391;
  assign n52893 = pi18 ? n52892 : n36659;
  assign n52894 = pi21 ? n36659 : n46243;
  assign n52895 = pi20 ? n52894 : n52409;
  assign n52896 = pi21 ? n39932 : n32;
  assign n52897 = pi20 ? n52896 : n32;
  assign n52898 = pi19 ? n52895 : n52897;
  assign n52899 = pi18 ? n36659 : n52898;
  assign n52900 = pi17 ? n52893 : n52899;
  assign n52901 = pi16 ? n32 : n52900;
  assign n52902 = pi20 ? n46225 : n36659;
  assign n52903 = pi19 ? n52902 : n36659;
  assign n52904 = pi18 ? n52903 : n36659;
  assign n52905 = pi22 ? n36659 : n18461;
  assign n52906 = pi21 ? n36659 : n52905;
  assign n52907 = pi20 ? n52906 : n52424;
  assign n52908 = pi19 ? n52907 : n32;
  assign n52909 = pi18 ? n36659 : n52908;
  assign n52910 = pi17 ? n52904 : n52909;
  assign n52911 = pi16 ? n32 : n52910;
  assign n52912 = pi15 ? n52901 : n52911;
  assign n52913 = pi20 ? n46277 : n42170;
  assign n52914 = pi19 ? n52913 : n36781;
  assign n52915 = pi18 ? n52914 : n36781;
  assign n52916 = pi17 ? n52915 : n52443;
  assign n52917 = pi16 ? n32 : n52916;
  assign n52918 = pi21 ? n32 : n46790;
  assign n52919 = pi20 ? n52918 : n43198;
  assign n52920 = pi19 ? n52919 : n52448;
  assign n52921 = pi18 ? n52920 : n36781;
  assign n52922 = pi20 ? n42170 : n20106;
  assign n52923 = pi19 ? n52922 : n32;
  assign n52924 = pi18 ? n51395 : n52923;
  assign n52925 = pi17 ? n52921 : n52924;
  assign n52926 = pi16 ? n32 : n52925;
  assign n52927 = pi15 ? n52917 : n52926;
  assign n52928 = pi14 ? n52912 : n52927;
  assign n52929 = pi13 ? n52890 : n52928;
  assign n52930 = pi12 ? n52850 : n52929;
  assign n52931 = pi11 ? n52780 : n52930;
  assign n52932 = pi10 ? n52656 : n52931;
  assign n52933 = pi09 ? n52484 : n52932;
  assign n52934 = pi08 ? n52465 : n52933;
  assign n52935 = pi07 ? n51923 : n52934;
  assign n52936 = pi21 ? n297 : n32;
  assign n52937 = pi20 ? n37 : n52936;
  assign n52938 = pi19 ? n37 : n52937;
  assign n52939 = pi18 ? n38951 : n52938;
  assign n52940 = pi17 ? n45367 : n52939;
  assign n52941 = pi16 ? n32 : n52940;
  assign n52942 = pi15 ? n32 : n52941;
  assign n52943 = pi20 ? n37 : n7308;
  assign n52944 = pi19 ? n37 : n52943;
  assign n52945 = pi18 ? n35777 : n52944;
  assign n52946 = pi17 ? n38958 : n52945;
  assign n52947 = pi16 ? n32 : n52946;
  assign n52948 = pi20 ? n38477 : n20563;
  assign n52949 = pi19 ? n20563 : n52948;
  assign n52950 = pi21 ? n9143 : n32;
  assign n52951 = pi20 ? n37 : n52950;
  assign n52952 = pi19 ? n32898 : n52951;
  assign n52953 = pi18 ? n52949 : n52952;
  assign n52954 = pi17 ? n38958 : n52953;
  assign n52955 = pi16 ? n32 : n52954;
  assign n52956 = pi15 ? n52947 : n52955;
  assign n52957 = pi14 ? n52942 : n52956;
  assign n52958 = pi13 ? n32 : n52957;
  assign n52959 = pi12 ? n32 : n52958;
  assign n52960 = pi11 ? n32 : n52959;
  assign n52961 = pi10 ? n32 : n52960;
  assign n52962 = pi21 ? n36249 : n20563;
  assign n52963 = pi20 ? n52962 : n20563;
  assign n52964 = pi19 ? n32294 : n52963;
  assign n52965 = pi21 ? n44672 : n32;
  assign n52966 = pi20 ? n3086 : n52965;
  assign n52967 = pi19 ? n37 : n52966;
  assign n52968 = pi18 ? n52964 : n52967;
  assign n52969 = pi17 ? n38330 : n52968;
  assign n52970 = pi16 ? n32 : n52969;
  assign n52971 = pi21 ? n894 : n32;
  assign n52972 = pi20 ? n3086 : n52971;
  assign n52973 = pi19 ? n37 : n52972;
  assign n52974 = pi18 ? n32294 : n52973;
  assign n52975 = pi17 ? n37929 : n52974;
  assign n52976 = pi16 ? n32 : n52975;
  assign n52977 = pi15 ? n52970 : n52976;
  assign n52978 = pi20 ? n31266 : n38477;
  assign n52979 = pi19 ? n52978 : n32898;
  assign n52980 = pi21 ? n7195 : n32;
  assign n52981 = pi20 ? n37 : n52980;
  assign n52982 = pi19 ? n37 : n52981;
  assign n52983 = pi18 ? n52979 : n52982;
  assign n52984 = pi17 ? n40057 : n52983;
  assign n52985 = pi16 ? n32 : n52984;
  assign n52986 = pi19 ? n50863 : n32348;
  assign n52987 = pi22 ? n37 : n1167;
  assign n52988 = pi21 ? n52987 : n32;
  assign n52989 = pi20 ? n37 : n52988;
  assign n52990 = pi19 ? n37 : n52989;
  assign n52991 = pi18 ? n52986 : n52990;
  assign n52992 = pi17 ? n37936 : n52991;
  assign n52993 = pi16 ? n32 : n52992;
  assign n52994 = pi15 ? n52985 : n52993;
  assign n52995 = pi14 ? n52977 : n52994;
  assign n52996 = pi22 ? n37 : n7513;
  assign n52997 = pi21 ? n52996 : n32;
  assign n52998 = pi20 ? n37 : n52997;
  assign n52999 = pi19 ? n37 : n52998;
  assign n53000 = pi18 ? n34258 : n52999;
  assign n53001 = pi17 ? n37958 : n53000;
  assign n53002 = pi16 ? n32 : n53001;
  assign n53003 = pi20 ? n36250 : n48905;
  assign n53004 = pi22 ? n335 : n7513;
  assign n53005 = pi21 ? n53004 : n32;
  assign n53006 = pi20 ? n52272 : n53005;
  assign n53007 = pi19 ? n53003 : n53006;
  assign n53008 = pi18 ? n34258 : n53007;
  assign n53009 = pi17 ? n36162 : n53008;
  assign n53010 = pi16 ? n32 : n53009;
  assign n53011 = pi15 ? n53002 : n53010;
  assign n53012 = pi20 ? n20563 : n48905;
  assign n53013 = pi19 ? n53012 : n32898;
  assign n53014 = pi20 ? n3299 : n22279;
  assign n53015 = pi19 ? n37 : n53014;
  assign n53016 = pi18 ? n53013 : n53015;
  assign n53017 = pi17 ? n36162 : n53016;
  assign n53018 = pi16 ? n32 : n53017;
  assign n53019 = pi18 ? n28159 : n52949;
  assign n53020 = pi19 ? n50854 : n31267;
  assign n53021 = pi20 ? n37 : n20319;
  assign n53022 = pi19 ? n37 : n53021;
  assign n53023 = pi18 ? n53020 : n53022;
  assign n53024 = pi17 ? n53019 : n53023;
  assign n53025 = pi16 ? n32 : n53024;
  assign n53026 = pi15 ? n53018 : n53025;
  assign n53027 = pi14 ? n53011 : n53026;
  assign n53028 = pi13 ? n52995 : n53027;
  assign n53029 = pi20 ? n30096 : n20563;
  assign n53030 = pi19 ? n53029 : n49016;
  assign n53031 = pi22 ? n37 : n16771;
  assign n53032 = pi21 ? n53031 : n32;
  assign n53033 = pi20 ? n37 : n53032;
  assign n53034 = pi19 ? n37 : n53033;
  assign n53035 = pi18 ? n53030 : n53034;
  assign n53036 = pi17 ? n35764 : n53035;
  assign n53037 = pi16 ? n32 : n53036;
  assign n53038 = pi20 ? n37 : n36285;
  assign n53039 = pi19 ? n37 : n53038;
  assign n53040 = pi18 ? n34295 : n53039;
  assign n53041 = pi17 ? n36215 : n53040;
  assign n53042 = pi16 ? n32 : n53041;
  assign n53043 = pi15 ? n53037 : n53042;
  assign n53044 = pi22 ? n335 : n6146;
  assign n53045 = pi21 ? n53044 : n32;
  assign n53046 = pi20 ? n37 : n53045;
  assign n53047 = pi19 ? n50883 : n53046;
  assign n53048 = pi18 ? n34258 : n53047;
  assign n53049 = pi17 ? n49894 : n53048;
  assign n53050 = pi16 ? n32 : n53049;
  assign n53051 = pi20 ? n37 : n52962;
  assign n53052 = pi22 ? n295 : n1378;
  assign n53053 = pi21 ? n53052 : n32;
  assign n53054 = pi20 ? n37 : n53053;
  assign n53055 = pi19 ? n53051 : n53054;
  assign n53056 = pi18 ? n20563 : n53055;
  assign n53057 = pi17 ? n49894 : n53056;
  assign n53058 = pi16 ? n32 : n53057;
  assign n53059 = pi15 ? n53050 : n53058;
  assign n53060 = pi14 ? n53043 : n53059;
  assign n53061 = pi20 ? n37308 : n20563;
  assign n53062 = pi19 ? n53061 : n31267;
  assign n53063 = pi22 ? n363 : n2564;
  assign n53064 = pi21 ? n53063 : n32;
  assign n53065 = pi20 ? n37 : n53064;
  assign n53066 = pi19 ? n37 : n53065;
  assign n53067 = pi18 ? n53062 : n53066;
  assign n53068 = pi17 ? n49894 : n53067;
  assign n53069 = pi16 ? n32 : n53068;
  assign n53070 = pi19 ? n51953 : n30097;
  assign n53071 = pi21 ? n16779 : n32;
  assign n53072 = pi20 ? n37 : n53071;
  assign n53073 = pi19 ? n37 : n53072;
  assign n53074 = pi18 ? n53070 : n53073;
  assign n53075 = pi17 ? n50905 : n53074;
  assign n53076 = pi16 ? n32 : n53075;
  assign n53077 = pi15 ? n53069 : n53076;
  assign n53078 = pi18 ? n34295 : n53073;
  assign n53079 = pi17 ? n49440 : n53078;
  assign n53080 = pi16 ? n32 : n53079;
  assign n53081 = pi20 ? n37 : n32313;
  assign n53082 = pi20 ? n37 : n10311;
  assign n53083 = pi19 ? n53081 : n53082;
  assign n53084 = pi18 ? n34258 : n53083;
  assign n53085 = pi17 ? n49448 : n53084;
  assign n53086 = pi16 ? n32 : n53085;
  assign n53087 = pi15 ? n53080 : n53086;
  assign n53088 = pi14 ? n53077 : n53087;
  assign n53089 = pi13 ? n53060 : n53088;
  assign n53090 = pi12 ? n53028 : n53089;
  assign n53091 = pi21 ? n2193 : n32;
  assign n53092 = pi20 ? n37 : n53091;
  assign n53093 = pi19 ? n51996 : n53092;
  assign n53094 = pi18 ? n20563 : n53093;
  assign n53095 = pi17 ? n49448 : n53094;
  assign n53096 = pi16 ? n32 : n53095;
  assign n53097 = pi20 ? n49916 : n31266;
  assign n53098 = pi20 ? n37 : n34943;
  assign n53099 = pi19 ? n53097 : n53098;
  assign n53100 = pi18 ? n34869 : n53099;
  assign n53101 = pi17 ? n49448 : n53100;
  assign n53102 = pi16 ? n32 : n53101;
  assign n53103 = pi15 ? n53096 : n53102;
  assign n53104 = pi20 ? n48905 : n20563;
  assign n53105 = pi19 ? n53104 : n31280;
  assign n53106 = pi20 ? n49916 : n30096;
  assign n53107 = pi19 ? n53106 : n53098;
  assign n53108 = pi18 ? n53105 : n53107;
  assign n53109 = pi17 ? n49448 : n53108;
  assign n53110 = pi16 ? n32 : n53109;
  assign n53111 = pi22 ? n27994 : n532;
  assign n53112 = pi21 ? n53111 : n32;
  assign n53113 = pi20 ? n37 : n53112;
  assign n53114 = pi19 ? n49917 : n53113;
  assign n53115 = pi18 ? n53105 : n53114;
  assign n53116 = pi17 ? n49451 : n53115;
  assign n53117 = pi16 ? n32 : n53116;
  assign n53118 = pi15 ? n53110 : n53117;
  assign n53119 = pi14 ? n53103 : n53118;
  assign n53120 = pi22 ? n157 : n625;
  assign n53121 = pi21 ? n53120 : n32;
  assign n53122 = pi20 ? n24493 : n53121;
  assign n53123 = pi19 ? n50932 : n53122;
  assign n53124 = pi18 ? n34869 : n53123;
  assign n53125 = pi17 ? n48897 : n53124;
  assign n53126 = pi16 ? n32 : n53125;
  assign n53127 = pi20 ? n21635 : n4008;
  assign n53128 = pi19 ? n50932 : n53127;
  assign n53129 = pi18 ? n34869 : n53128;
  assign n53130 = pi17 ? n48897 : n53129;
  assign n53131 = pi16 ? n32 : n53130;
  assign n53132 = pi15 ? n53126 : n53131;
  assign n53133 = pi20 ? n24493 : n12149;
  assign n53134 = pi19 ? n51996 : n53133;
  assign n53135 = pi18 ? n20563 : n53134;
  assign n53136 = pi17 ? n48897 : n53135;
  assign n53137 = pi16 ? n32 : n53136;
  assign n53138 = pi21 ? n37 : n777;
  assign n53139 = pi20 ? n53138 : n4008;
  assign n53140 = pi19 ? n51996 : n53139;
  assign n53141 = pi18 ? n20563 : n53140;
  assign n53142 = pi17 ? n48897 : n53141;
  assign n53143 = pi16 ? n32 : n53142;
  assign n53144 = pi15 ? n53137 : n53143;
  assign n53145 = pi14 ? n53132 : n53144;
  assign n53146 = pi13 ? n53119 : n53145;
  assign n53147 = pi19 ? n50927 : n53139;
  assign n53148 = pi18 ? n20563 : n53147;
  assign n53149 = pi17 ? n48904 : n53148;
  assign n53150 = pi16 ? n32 : n53149;
  assign n53151 = pi18 ? n42687 : n20563;
  assign n53152 = pi20 ? n2238 : n7733;
  assign n53153 = pi19 ? n31221 : n53152;
  assign n53154 = pi18 ? n34869 : n53153;
  assign n53155 = pi17 ? n53151 : n53154;
  assign n53156 = pi16 ? n32 : n53155;
  assign n53157 = pi15 ? n53150 : n53156;
  assign n53158 = pi20 ? n20563 : n5077;
  assign n53159 = pi20 ? n1665 : n3977;
  assign n53160 = pi19 ? n53158 : n53159;
  assign n53161 = pi18 ? n20563 : n53160;
  assign n53162 = pi17 ? n53151 : n53161;
  assign n53163 = pi16 ? n32 : n53162;
  assign n53164 = pi23 ? n3491 : n316;
  assign n53165 = pi22 ? n99 : n53164;
  assign n53166 = pi21 ? n99 : n53165;
  assign n53167 = pi20 ? n53166 : n3210;
  assign n53168 = pi19 ? n31221 : n53167;
  assign n53169 = pi18 ? n20563 : n53168;
  assign n53170 = pi17 ? n53151 : n53169;
  assign n53171 = pi16 ? n32 : n53170;
  assign n53172 = pi15 ? n53163 : n53171;
  assign n53173 = pi14 ? n53157 : n53172;
  assign n53174 = pi24 ? n99 : n316;
  assign n53175 = pi23 ? n53174 : n316;
  assign n53176 = pi22 ? n99 : n53175;
  assign n53177 = pi21 ? n99 : n53176;
  assign n53178 = pi20 ? n53177 : n10011;
  assign n53179 = pi19 ? n32898 : n53178;
  assign n53180 = pi18 ? n20563 : n53179;
  assign n53181 = pi17 ? n53151 : n53180;
  assign n53182 = pi16 ? n32 : n53181;
  assign n53183 = pi20 ? n20563 : n36516;
  assign n53184 = pi23 ? n11962 : n204;
  assign n53185 = pi22 ? n99 : n53184;
  assign n53186 = pi21 ? n99 : n53185;
  assign n53187 = pi20 ? n53186 : n2638;
  assign n53188 = pi19 ? n53183 : n53187;
  assign n53189 = pi18 ? n20563 : n53188;
  assign n53190 = pi17 ? n53151 : n53189;
  assign n53191 = pi16 ? n32 : n53190;
  assign n53192 = pi15 ? n53182 : n53191;
  assign n53193 = pi21 ? n181 : n204;
  assign n53194 = pi20 ? n53193 : n2638;
  assign n53195 = pi19 ? n32348 : n53194;
  assign n53196 = pi18 ? n20563 : n53195;
  assign n53197 = pi17 ? n49485 : n53196;
  assign n53198 = pi16 ? n32 : n53197;
  assign n53199 = pi21 ? n297 : n8842;
  assign n53200 = pi20 ? n53199 : n2653;
  assign n53201 = pi19 ? n32898 : n53200;
  assign n53202 = pi18 ? n20563 : n53201;
  assign n53203 = pi17 ? n49485 : n53202;
  assign n53204 = pi16 ? n32 : n53203;
  assign n53205 = pi15 ? n53198 : n53204;
  assign n53206 = pi14 ? n53192 : n53205;
  assign n53207 = pi13 ? n53173 : n53206;
  assign n53208 = pi12 ? n53146 : n53207;
  assign n53209 = pi11 ? n53090 : n53208;
  assign n53210 = pi21 ? n3073 : n8842;
  assign n53211 = pi20 ? n53210 : n2653;
  assign n53212 = pi19 ? n32898 : n53211;
  assign n53213 = pi18 ? n20563 : n53212;
  assign n53214 = pi17 ? n49485 : n53213;
  assign n53215 = pi16 ? n32 : n53214;
  assign n53216 = pi21 ? n139 : n3763;
  assign n53217 = pi20 ? n53216 : n1822;
  assign n53218 = pi19 ? n32898 : n53217;
  assign n53219 = pi18 ? n20563 : n53218;
  assign n53220 = pi17 ? n49485 : n53219;
  assign n53221 = pi16 ? n32 : n53220;
  assign n53222 = pi15 ? n53215 : n53221;
  assign n53223 = pi21 ? n139 : n16438;
  assign n53224 = pi20 ? n53223 : n32;
  assign n53225 = pi19 ? n32898 : n53224;
  assign n53226 = pi18 ? n20563 : n53225;
  assign n53227 = pi17 ? n49485 : n53226;
  assign n53228 = pi16 ? n32 : n53227;
  assign n53229 = pi18 ? n41157 : n20563;
  assign n53230 = pi21 ? n297 : n16438;
  assign n53231 = pi20 ? n53230 : n32;
  assign n53232 = pi19 ? n32348 : n53231;
  assign n53233 = pi18 ? n20563 : n53232;
  assign n53234 = pi17 ? n53229 : n53233;
  assign n53235 = pi16 ? n32 : n53234;
  assign n53236 = pi15 ? n53228 : n53235;
  assign n53237 = pi14 ? n53222 : n53236;
  assign n53238 = pi21 ? n29133 : n99;
  assign n53239 = pi20 ? n20563 : n53238;
  assign n53240 = pi21 ? n297 : n1389;
  assign n53241 = pi20 ? n53240 : n32;
  assign n53242 = pi19 ? n53239 : n53241;
  assign n53243 = pi18 ? n20563 : n53242;
  assign n53244 = pi17 ? n47922 : n53243;
  assign n53245 = pi16 ? n32 : n53244;
  assign n53246 = pi22 ? n673 : n759;
  assign n53247 = pi21 ? n139 : n53246;
  assign n53248 = pi20 ? n53247 : n32;
  assign n53249 = pi19 ? n32898 : n53248;
  assign n53250 = pi18 ? n20563 : n53249;
  assign n53251 = pi17 ? n47922 : n53250;
  assign n53252 = pi16 ? n32 : n53251;
  assign n53253 = pi15 ? n53245 : n53252;
  assign n53254 = pi22 ? n1457 : n396;
  assign n53255 = pi21 ? n9143 : n53254;
  assign n53256 = pi20 ? n53255 : n32;
  assign n53257 = pi19 ? n32898 : n53256;
  assign n53258 = pi18 ? n20563 : n53257;
  assign n53259 = pi17 ? n47929 : n53258;
  assign n53260 = pi16 ? n32 : n53259;
  assign n53261 = pi21 ? n335 : n52311;
  assign n53262 = pi20 ? n53261 : n32;
  assign n53263 = pi19 ? n32898 : n53262;
  assign n53264 = pi18 ? n20563 : n53263;
  assign n53265 = pi17 ? n47929 : n53264;
  assign n53266 = pi16 ? n32 : n53265;
  assign n53267 = pi15 ? n53260 : n53266;
  assign n53268 = pi14 ? n53253 : n53267;
  assign n53269 = pi13 ? n53237 : n53268;
  assign n53270 = pi21 ? n335 : n9186;
  assign n53271 = pi20 ? n53270 : n32;
  assign n53272 = pi19 ? n51162 : n53271;
  assign n53273 = pi18 ? n20563 : n53272;
  assign n53274 = pi17 ? n47929 : n53273;
  assign n53275 = pi16 ? n32 : n53274;
  assign n53276 = pi22 ? n27667 : n32;
  assign n53277 = pi21 ? n363 : n53276;
  assign n53278 = pi20 ? n53277 : n32;
  assign n53279 = pi19 ? n31221 : n53278;
  assign n53280 = pi18 ? n20563 : n53279;
  assign n53281 = pi17 ? n48949 : n53280;
  assign n53282 = pi16 ? n32 : n53281;
  assign n53283 = pi15 ? n53275 : n53282;
  assign n53284 = pi21 ? n38041 : n12825;
  assign n53285 = pi20 ? n53284 : n32;
  assign n53286 = pi19 ? n31221 : n53285;
  assign n53287 = pi18 ? n20563 : n53286;
  assign n53288 = pi17 ? n47935 : n53287;
  assign n53289 = pi16 ? n32 : n53288;
  assign n53290 = pi20 ? n32 : n30868;
  assign n53291 = pi20 ? n42005 : n51708;
  assign n53292 = pi19 ? n53290 : n53291;
  assign n53293 = pi20 ? n43935 : n42006;
  assign n53294 = pi19 ? n53293 : n50244;
  assign n53295 = pi18 ? n53292 : n53294;
  assign n53296 = pi20 ? n43935 : n20563;
  assign n53297 = pi19 ? n53296 : n20563;
  assign n53298 = pi21 ? n157 : n4101;
  assign n53299 = pi20 ? n53298 : n32;
  assign n53300 = pi19 ? n31221 : n53299;
  assign n53301 = pi18 ? n53297 : n53300;
  assign n53302 = pi17 ? n53295 : n53301;
  assign n53303 = pi16 ? n32 : n53302;
  assign n53304 = pi15 ? n53289 : n53303;
  assign n53305 = pi14 ? n53283 : n53304;
  assign n53306 = pi20 ? n32 : n33792;
  assign n53307 = pi21 ? n40957 : n33792;
  assign n53308 = pi21 ? n40955 : n20563;
  assign n53309 = pi20 ? n53307 : n53308;
  assign n53310 = pi19 ? n53306 : n53309;
  assign n53311 = pi18 ? n53310 : n20563;
  assign n53312 = pi20 ? n40791 : n31220;
  assign n53313 = pi23 ? n233 : n157;
  assign n53314 = pi22 ? n335 : n53313;
  assign n53315 = pi21 ? n53314 : n6416;
  assign n53316 = pi20 ? n53315 : n32;
  assign n53317 = pi19 ? n53312 : n53316;
  assign n53318 = pi18 ? n20563 : n53317;
  assign n53319 = pi17 ? n53311 : n53318;
  assign n53320 = pi16 ? n32 : n53319;
  assign n53321 = pi19 ? n53306 : n33792;
  assign n53322 = pi20 ? n53307 : n33792;
  assign n53323 = pi19 ? n33792 : n53322;
  assign n53324 = pi18 ? n53321 : n53323;
  assign n53325 = pi19 ? n53307 : n20563;
  assign n53326 = pi21 ? n20563 : n33792;
  assign n53327 = pi20 ? n53326 : n31220;
  assign n53328 = pi21 ? n6376 : n3339;
  assign n53329 = pi20 ? n53328 : n32;
  assign n53330 = pi19 ? n53327 : n53329;
  assign n53331 = pi18 ? n53325 : n53330;
  assign n53332 = pi17 ? n53324 : n53331;
  assign n53333 = pi16 ? n32 : n53332;
  assign n53334 = pi15 ? n53320 : n53333;
  assign n53335 = pi22 ? n363 : n1449;
  assign n53336 = pi21 ? n53335 : n5829;
  assign n53337 = pi20 ? n53336 : n32;
  assign n53338 = pi19 ? n31221 : n53337;
  assign n53339 = pi18 ? n20563 : n53338;
  assign n53340 = pi17 ? n47451 : n53339;
  assign n53341 = pi16 ? n32 : n53340;
  assign n53342 = pi22 ? n20563 : n99;
  assign n53343 = pi21 ? n20563 : n53342;
  assign n53344 = pi20 ? n20563 : n53343;
  assign n53345 = pi22 ? n52307 : n29708;
  assign n53346 = pi21 ? n53345 : n5370;
  assign n53347 = pi20 ? n53346 : n32;
  assign n53348 = pi19 ? n53344 : n53347;
  assign n53349 = pi18 ? n20563 : n53348;
  assign n53350 = pi17 ? n47443 : n53349;
  assign n53351 = pi16 ? n32 : n53350;
  assign n53352 = pi15 ? n53341 : n53351;
  assign n53353 = pi14 ? n53334 : n53352;
  assign n53354 = pi13 ? n53305 : n53353;
  assign n53355 = pi12 ? n53269 : n53354;
  assign n53356 = pi21 ? n20563 : n50266;
  assign n53357 = pi20 ? n20563 : n53356;
  assign n53358 = pi23 ? n8184 : n157;
  assign n53359 = pi22 ? n53358 : n685;
  assign n53360 = pi21 ? n53359 : n928;
  assign n53361 = pi20 ? n53360 : n32;
  assign n53362 = pi19 ? n53357 : n53361;
  assign n53363 = pi18 ? n20563 : n53362;
  assign n53364 = pi17 ? n47443 : n53363;
  assign n53365 = pi16 ? n32 : n53364;
  assign n53366 = pi22 ? n20563 : n335;
  assign n53367 = pi21 ? n20563 : n53366;
  assign n53368 = pi20 ? n20563 : n53367;
  assign n53369 = pi23 ? n3134 : n157;
  assign n53370 = pi22 ? n53369 : n685;
  assign n53371 = pi21 ? n53370 : n1009;
  assign n53372 = pi20 ? n53371 : n32;
  assign n53373 = pi19 ? n53368 : n53372;
  assign n53374 = pi18 ? n20563 : n53373;
  assign n53375 = pi17 ? n47443 : n53374;
  assign n53376 = pi16 ? n32 : n53375;
  assign n53377 = pi15 ? n53365 : n53376;
  assign n53378 = pi22 ? n5061 : n316;
  assign n53379 = pi21 ? n53378 : n32;
  assign n53380 = pi20 ? n53379 : n32;
  assign n53381 = pi19 ? n53368 : n53380;
  assign n53382 = pi18 ? n20563 : n53381;
  assign n53383 = pi17 ? n47954 : n53382;
  assign n53384 = pi16 ? n32 : n53383;
  assign n53385 = pi22 ? n20563 : n363;
  assign n53386 = pi21 ? n20563 : n53385;
  assign n53387 = pi20 ? n20563 : n53386;
  assign n53388 = pi20 ? n42628 : n32;
  assign n53389 = pi19 ? n53387 : n53388;
  assign n53390 = pi18 ? n20563 : n53389;
  assign n53391 = pi17 ? n47954 : n53390;
  assign n53392 = pi16 ? n32 : n53391;
  assign n53393 = pi15 ? n53384 : n53392;
  assign n53394 = pi14 ? n53377 : n53393;
  assign n53395 = pi22 ? n30868 : n363;
  assign n53396 = pi21 ? n20563 : n53395;
  assign n53397 = pi20 ? n20563 : n53396;
  assign n53398 = pi22 ? n1457 : n2192;
  assign n53399 = pi21 ? n53398 : n32;
  assign n53400 = pi20 ? n53399 : n32;
  assign n53401 = pi19 ? n53397 : n53400;
  assign n53402 = pi18 ? n20563 : n53401;
  assign n53403 = pi17 ? n47954 : n53402;
  assign n53404 = pi16 ? n32 : n53403;
  assign n53405 = pi20 ? n47835 : n40915;
  assign n53406 = pi19 ? n53405 : n30868;
  assign n53407 = pi18 ? n53406 : n43012;
  assign n53408 = pi22 ? n30868 : n157;
  assign n53409 = pi21 ? n20563 : n53408;
  assign n53410 = pi20 ? n20563 : n53409;
  assign n53411 = pi21 ? n9584 : n32;
  assign n53412 = pi20 ? n53411 : n32;
  assign n53413 = pi19 ? n53410 : n53412;
  assign n53414 = pi18 ? n20563 : n53413;
  assign n53415 = pi17 ? n53407 : n53414;
  assign n53416 = pi16 ? n32 : n53415;
  assign n53417 = pi15 ? n53404 : n53416;
  assign n53418 = pi20 ? n42005 : n50736;
  assign n53419 = pi19 ? n53405 : n53418;
  assign n53420 = pi18 ? n53419 : n20563;
  assign n53421 = pi22 ? n33792 : n157;
  assign n53422 = pi21 ? n20563 : n53421;
  assign n53423 = pi20 ? n20563 : n53422;
  assign n53424 = pi19 ? n53423 : n9964;
  assign n53425 = pi18 ? n20563 : n53424;
  assign n53426 = pi17 ? n53420 : n53425;
  assign n53427 = pi16 ? n32 : n53426;
  assign n53428 = pi21 ? n49206 : n20563;
  assign n53429 = pi20 ? n32 : n53428;
  assign n53430 = pi19 ? n53429 : n20563;
  assign n53431 = pi18 ? n53430 : n20563;
  assign n53432 = pi22 ? n36659 : n204;
  assign n53433 = pi21 ? n36489 : n53432;
  assign n53434 = pi20 ? n20563 : n53433;
  assign n53435 = pi19 ? n53434 : n4009;
  assign n53436 = pi18 ? n20563 : n53435;
  assign n53437 = pi17 ? n53431 : n53436;
  assign n53438 = pi16 ? n32 : n53437;
  assign n53439 = pi15 ? n53427 : n53438;
  assign n53440 = pi14 ? n53417 : n53439;
  assign n53441 = pi13 ? n53394 : n53440;
  assign n53442 = pi19 ? n37807 : n30868;
  assign n53443 = pi18 ? n53442 : n30868;
  assign n53444 = pi21 ? n30868 : n51564;
  assign n53445 = pi20 ? n30868 : n53444;
  assign n53446 = pi19 ? n53445 : n4009;
  assign n53447 = pi18 ? n30868 : n53446;
  assign n53448 = pi17 ? n53443 : n53447;
  assign n53449 = pi16 ? n32 : n53448;
  assign n53450 = pi23 ? n99 : n33792;
  assign n53451 = pi22 ? n30868 : n53450;
  assign n53452 = pi21 ? n30868 : n53451;
  assign n53453 = pi21 ? n47220 : n51564;
  assign n53454 = pi20 ? n53452 : n53453;
  assign n53455 = pi19 ? n53454 : n5831;
  assign n53456 = pi18 ? n30868 : n53455;
  assign n53457 = pi17 ? n53443 : n53456;
  assign n53458 = pi16 ? n32 : n53457;
  assign n53459 = pi15 ? n53449 : n53458;
  assign n53460 = pi21 ? n47341 : n36798;
  assign n53461 = pi20 ? n32 : n53460;
  assign n53462 = pi19 ? n53461 : n36798;
  assign n53463 = pi22 ? n33792 : n36798;
  assign n53464 = pi21 ? n53463 : n36798;
  assign n53465 = pi20 ? n33792 : n53464;
  assign n53466 = pi19 ? n36798 : n53465;
  assign n53467 = pi18 ? n53462 : n53466;
  assign n53468 = pi21 ? n36798 : n53463;
  assign n53469 = pi20 ? n53468 : n33792;
  assign n53470 = pi19 ? n53469 : n33792;
  assign n53471 = pi22 ? n33792 : n43198;
  assign n53472 = pi21 ? n53471 : n13481;
  assign n53473 = pi20 ? n33792 : n53472;
  assign n53474 = pi19 ? n53473 : n2654;
  assign n53475 = pi18 ? n53470 : n53474;
  assign n53476 = pi17 ? n53467 : n53475;
  assign n53477 = pi16 ? n32 : n53476;
  assign n53478 = pi21 ? n47410 : n43198;
  assign n53479 = pi20 ? n32 : n53478;
  assign n53480 = pi22 ? n52873 : n33792;
  assign n53481 = pi21 ? n43198 : n53480;
  assign n53482 = pi20 ? n53471 : n53481;
  assign n53483 = pi19 ? n53479 : n53482;
  assign n53484 = pi22 ? n43198 : n33792;
  assign n53485 = pi21 ? n33792 : n53484;
  assign n53486 = pi20 ? n33792 : n53485;
  assign n53487 = pi19 ? n53486 : n33792;
  assign n53488 = pi18 ? n53483 : n53487;
  assign n53489 = pi21 ? n47360 : n13481;
  assign n53490 = pi20 ? n33792 : n53489;
  assign n53491 = pi19 ? n53490 : n2654;
  assign n53492 = pi18 ? n33792 : n53491;
  assign n53493 = pi17 ? n53488 : n53492;
  assign n53494 = pi16 ? n32 : n53493;
  assign n53495 = pi15 ? n53477 : n53494;
  assign n53496 = pi14 ? n53459 : n53495;
  assign n53497 = pi21 ? n50338 : n50796;
  assign n53498 = pi20 ? n36659 : n53497;
  assign n53499 = pi19 ? n53479 : n53498;
  assign n53500 = pi18 ? n53499 : n36659;
  assign n53501 = pi21 ? n36659 : n13481;
  assign n53502 = pi20 ? n36659 : n53501;
  assign n53503 = pi19 ? n53502 : n1823;
  assign n53504 = pi18 ? n36659 : n53503;
  assign n53505 = pi17 ? n53500 : n53504;
  assign n53506 = pi16 ? n32 : n53505;
  assign n53507 = pi22 ? n32 : n52415;
  assign n53508 = pi22 ? n50339 : n36659;
  assign n53509 = pi21 ? n53507 : n53508;
  assign n53510 = pi20 ? n32 : n53509;
  assign n53511 = pi21 ? n37277 : n36659;
  assign n53512 = pi20 ? n37878 : n53511;
  assign n53513 = pi19 ? n53510 : n53512;
  assign n53514 = pi21 ? n37878 : n42146;
  assign n53515 = pi20 ? n42147 : n53514;
  assign n53516 = pi21 ? n36781 : n37878;
  assign n53517 = pi20 ? n53516 : n42147;
  assign n53518 = pi19 ? n53515 : n53517;
  assign n53519 = pi18 ? n53513 : n53518;
  assign n53520 = pi22 ? n36781 : n37288;
  assign n53521 = pi21 ? n37878 : n53520;
  assign n53522 = pi20 ? n40002 : n53521;
  assign n53523 = pi22 ? n37288 : n36659;
  assign n53524 = pi21 ? n37288 : n53523;
  assign n53525 = pi20 ? n37288 : n53524;
  assign n53526 = pi19 ? n53522 : n53525;
  assign n53527 = pi21 ? n42146 : n53520;
  assign n53528 = pi21 ? n37878 : n13481;
  assign n53529 = pi20 ? n53527 : n53528;
  assign n53530 = pi19 ? n53529 : n35482;
  assign n53531 = pi18 ? n53526 : n53530;
  assign n53532 = pi17 ? n53519 : n53531;
  assign n53533 = pi16 ? n32 : n53532;
  assign n53534 = pi15 ? n53506 : n53533;
  assign n53535 = pi21 ? n51367 : n36781;
  assign n53536 = pi20 ? n32 : n53535;
  assign n53537 = pi22 ? n43199 : n36781;
  assign n53538 = pi21 ? n53537 : n36781;
  assign n53539 = pi20 ? n36781 : n53538;
  assign n53540 = pi19 ? n53536 : n53539;
  assign n53541 = pi18 ? n53540 : n36781;
  assign n53542 = pi22 ? n13481 : n2192;
  assign n53543 = pi21 ? n39972 : n53542;
  assign n53544 = pi20 ? n36781 : n53543;
  assign n53545 = pi19 ? n53544 : n32;
  assign n53546 = pi18 ? n36781 : n53545;
  assign n53547 = pi17 ? n53541 : n53546;
  assign n53548 = pi16 ? n32 : n53547;
  assign n53549 = pi20 ? n32 : n49386;
  assign n53550 = pi23 ? n36798 : n43198;
  assign n53551 = pi22 ? n36798 : n53550;
  assign n53552 = pi21 ? n53551 : n43198;
  assign n53553 = pi20 ? n53552 : n47396;
  assign n53554 = pi19 ? n53549 : n53553;
  assign n53555 = pi21 ? n47397 : n36798;
  assign n53556 = pi20 ? n53555 : n36798;
  assign n53557 = pi19 ? n53556 : n36798;
  assign n53558 = pi18 ? n53554 : n53557;
  assign n53559 = pi22 ? n51564 : n317;
  assign n53560 = pi21 ? n43198 : n53559;
  assign n53561 = pi20 ? n36798 : n53560;
  assign n53562 = pi19 ? n53561 : n32;
  assign n53563 = pi18 ? n36798 : n53562;
  assign n53564 = pi17 ? n53558 : n53563;
  assign n53565 = pi16 ? n32 : n53564;
  assign n53566 = pi15 ? n53548 : n53565;
  assign n53567 = pi14 ? n53534 : n53566;
  assign n53568 = pi13 ? n53496 : n53567;
  assign n53569 = pi12 ? n53441 : n53568;
  assign n53570 = pi11 ? n53355 : n53569;
  assign n53571 = pi10 ? n53209 : n53570;
  assign n53572 = pi09 ? n52961 : n53571;
  assign n53573 = pi18 ? n34258 : n52938;
  assign n53574 = pi17 ? n40511 : n53573;
  assign n53575 = pi16 ? n32 : n53574;
  assign n53576 = pi15 ? n32 : n53575;
  assign n53577 = pi21 ? n35230 : n29133;
  assign n53578 = pi20 ? n53577 : n37;
  assign n53579 = pi19 ? n53578 : n52943;
  assign n53580 = pi18 ? n34869 : n53579;
  assign n53581 = pi17 ? n39374 : n53580;
  assign n53582 = pi16 ? n32 : n53581;
  assign n53583 = pi15 ? n53582 : n52955;
  assign n53584 = pi14 ? n53576 : n53583;
  assign n53585 = pi13 ? n32 : n53584;
  assign n53586 = pi12 ? n32 : n53585;
  assign n53587 = pi11 ? n32 : n53586;
  assign n53588 = pi10 ? n32 : n53587;
  assign n53589 = pi17 ? n38958 : n52968;
  assign n53590 = pi16 ? n32 : n53589;
  assign n53591 = pi17 ? n40046 : n52974;
  assign n53592 = pi16 ? n32 : n53591;
  assign n53593 = pi15 ? n53590 : n53592;
  assign n53594 = pi22 ? n295 : n25629;
  assign n53595 = pi21 ? n53594 : n32;
  assign n53596 = pi20 ? n37 : n53595;
  assign n53597 = pi19 ? n37 : n53596;
  assign n53598 = pi18 ? n52979 : n53597;
  assign n53599 = pi17 ? n40551 : n53598;
  assign n53600 = pi16 ? n32 : n53599;
  assign n53601 = pi20 ? n31913 : n20563;
  assign n53602 = pi19 ? n53601 : n31904;
  assign n53603 = pi18 ? n53602 : n52990;
  assign n53604 = pi17 ? n45393 : n53603;
  assign n53605 = pi16 ? n32 : n53604;
  assign n53606 = pi15 ? n53600 : n53605;
  assign n53607 = pi14 ? n53593 : n53606;
  assign n53608 = pi21 ? n11616 : n32;
  assign n53609 = pi20 ? n37 : n53608;
  assign n53610 = pi19 ? n37 : n53609;
  assign n53611 = pi18 ? n34258 : n53610;
  assign n53612 = pi17 ? n37929 : n53611;
  assign n53613 = pi16 ? n32 : n53612;
  assign n53614 = pi20 ? n52272 : n22814;
  assign n53615 = pi19 ? n53003 : n53614;
  assign n53616 = pi18 ? n34247 : n53615;
  assign n53617 = pi17 ? n37958 : n53616;
  assign n53618 = pi16 ? n32 : n53617;
  assign n53619 = pi15 ? n53613 : n53618;
  assign n53620 = pi20 ? n3299 : n22814;
  assign n53621 = pi19 ? n37 : n53620;
  assign n53622 = pi18 ? n53013 : n53621;
  assign n53623 = pi17 ? n37958 : n53622;
  assign n53624 = pi16 ? n32 : n53623;
  assign n53625 = pi18 ? n38999 : n52949;
  assign n53626 = pi20 ? n4971 : n10262;
  assign n53627 = pi19 ? n37 : n53626;
  assign n53628 = pi18 ? n53020 : n53627;
  assign n53629 = pi17 ? n53625 : n53628;
  assign n53630 = pi16 ? n32 : n53629;
  assign n53631 = pi15 ? n53624 : n53630;
  assign n53632 = pi14 ? n53619 : n53631;
  assign n53633 = pi13 ? n53607 : n53632;
  assign n53634 = pi19 ? n37 : n25331;
  assign n53635 = pi18 ? n53030 : n53634;
  assign n53636 = pi17 ? n37336 : n53635;
  assign n53637 = pi16 ? n32 : n53636;
  assign n53638 = pi20 ? n37 : n36983;
  assign n53639 = pi19 ? n37 : n53638;
  assign n53640 = pi18 ? n34295 : n53639;
  assign n53641 = pi17 ? n37336 : n53640;
  assign n53642 = pi16 ? n32 : n53641;
  assign n53643 = pi15 ? n53637 : n53642;
  assign n53644 = pi22 ? n335 : n1484;
  assign n53645 = pi21 ? n53644 : n32;
  assign n53646 = pi20 ? n37 : n53645;
  assign n53647 = pi19 ? n50883 : n53646;
  assign n53648 = pi18 ? n34258 : n53647;
  assign n53649 = pi17 ? n36215 : n53648;
  assign n53650 = pi16 ? n32 : n53649;
  assign n53651 = pi22 ? n295 : n6114;
  assign n53652 = pi21 ? n53651 : n32;
  assign n53653 = pi20 ? n37 : n53652;
  assign n53654 = pi19 ? n53051 : n53653;
  assign n53655 = pi18 ? n20563 : n53654;
  assign n53656 = pi17 ? n36215 : n53655;
  assign n53657 = pi16 ? n32 : n53656;
  assign n53658 = pi15 ? n53650 : n53657;
  assign n53659 = pi14 ? n53643 : n53658;
  assign n53660 = pi22 ? n363 : n3174;
  assign n53661 = pi21 ? n53660 : n32;
  assign n53662 = pi20 ? n37 : n53661;
  assign n53663 = pi19 ? n37 : n53662;
  assign n53664 = pi18 ? n53062 : n53663;
  assign n53665 = pi17 ? n50390 : n53664;
  assign n53666 = pi16 ? n32 : n53665;
  assign n53667 = pi22 ? n14245 : n730;
  assign n53668 = pi21 ? n53667 : n32;
  assign n53669 = pi20 ? n37 : n53668;
  assign n53670 = pi19 ? n37 : n53669;
  assign n53671 = pi18 ? n53070 : n53670;
  assign n53672 = pi17 ? n50393 : n53671;
  assign n53673 = pi16 ? n32 : n53672;
  assign n53674 = pi15 ? n53666 : n53673;
  assign n53675 = pi22 ? n14245 : n10784;
  assign n53676 = pi21 ? n53675 : n32;
  assign n53677 = pi20 ? n37 : n53676;
  assign n53678 = pi19 ? n37 : n53677;
  assign n53679 = pi18 ? n34295 : n53678;
  assign n53680 = pi17 ? n49888 : n53679;
  assign n53681 = pi16 ? n32 : n53680;
  assign n53682 = pi17 ? n49894 : n53084;
  assign n53683 = pi16 ? n32 : n53682;
  assign n53684 = pi15 ? n53681 : n53683;
  assign n53685 = pi14 ? n53674 : n53684;
  assign n53686 = pi13 ? n53659 : n53685;
  assign n53687 = pi12 ? n53633 : n53686;
  assign n53688 = pi17 ? n49894 : n53094;
  assign n53689 = pi16 ? n32 : n53688;
  assign n53690 = pi17 ? n49894 : n53100;
  assign n53691 = pi16 ? n32 : n53690;
  assign n53692 = pi15 ? n53689 : n53691;
  assign n53693 = pi17 ? n49894 : n53108;
  assign n53694 = pi16 ? n32 : n53693;
  assign n53695 = pi22 ? n158 : n532;
  assign n53696 = pi21 ? n53695 : n32;
  assign n53697 = pi20 ? n37 : n53696;
  assign n53698 = pi19 ? n49917 : n53697;
  assign n53699 = pi18 ? n53105 : n53698;
  assign n53700 = pi17 ? n49900 : n53699;
  assign n53701 = pi16 ? n32 : n53700;
  assign n53702 = pi15 ? n53694 : n53701;
  assign n53703 = pi14 ? n53692 : n53702;
  assign n53704 = pi17 ? n49440 : n53124;
  assign n53705 = pi16 ? n32 : n53704;
  assign n53706 = pi20 ? n21635 : n12149;
  assign n53707 = pi19 ? n50932 : n53706;
  assign n53708 = pi18 ? n34869 : n53707;
  assign n53709 = pi17 ? n49440 : n53708;
  assign n53710 = pi16 ? n32 : n53709;
  assign n53711 = pi15 ? n53705 : n53710;
  assign n53712 = pi20 ? n24493 : n4008;
  assign n53713 = pi19 ? n51996 : n53712;
  assign n53714 = pi18 ? n20563 : n53713;
  assign n53715 = pi17 ? n49440 : n53714;
  assign n53716 = pi16 ? n32 : n53715;
  assign n53717 = pi17 ? n49440 : n53141;
  assign n53718 = pi16 ? n32 : n53717;
  assign n53719 = pi15 ? n53716 : n53718;
  assign n53720 = pi14 ? n53711 : n53719;
  assign n53721 = pi13 ? n53703 : n53720;
  assign n53722 = pi20 ? n53138 : n5667;
  assign n53723 = pi19 ? n50927 : n53722;
  assign n53724 = pi18 ? n20563 : n53723;
  assign n53725 = pi17 ? n49448 : n53724;
  assign n53726 = pi16 ? n32 : n53725;
  assign n53727 = pi18 ? n42200 : n20563;
  assign n53728 = pi19 ? n31221 : n24938;
  assign n53729 = pi18 ? n34869 : n53728;
  assign n53730 = pi17 ? n53727 : n53729;
  assign n53731 = pi16 ? n32 : n53730;
  assign n53732 = pi15 ? n53726 : n53731;
  assign n53733 = pi21 ? n31200 : n181;
  assign n53734 = pi20 ? n20563 : n53733;
  assign n53735 = pi23 ? n15293 : n316;
  assign n53736 = pi22 ? n53735 : n32;
  assign n53737 = pi21 ? n53736 : n32;
  assign n53738 = pi20 ? n1665 : n53737;
  assign n53739 = pi19 ? n53734 : n53738;
  assign n53740 = pi18 ? n20563 : n53739;
  assign n53741 = pi17 ? n53727 : n53740;
  assign n53742 = pi16 ? n32 : n53741;
  assign n53743 = pi22 ? n99 : n1784;
  assign n53744 = pi21 ? n99 : n53743;
  assign n53745 = pi20 ? n53744 : n3210;
  assign n53746 = pi19 ? n31221 : n53745;
  assign n53747 = pi18 ? n20563 : n53746;
  assign n53748 = pi17 ? n53727 : n53747;
  assign n53749 = pi16 ? n32 : n53748;
  assign n53750 = pi15 ? n53742 : n53749;
  assign n53751 = pi14 ? n53732 : n53750;
  assign n53752 = pi20 ? n53744 : n10011;
  assign n53753 = pi19 ? n32898 : n53752;
  assign n53754 = pi18 ? n20563 : n53753;
  assign n53755 = pi17 ? n53727 : n53754;
  assign n53756 = pi16 ? n32 : n53755;
  assign n53757 = pi22 ? n99 : n448;
  assign n53758 = pi21 ? n99 : n53757;
  assign n53759 = pi23 ? n1598 : n687;
  assign n53760 = pi22 ? n53759 : n32;
  assign n53761 = pi21 ? n53760 : n32;
  assign n53762 = pi20 ? n53758 : n53761;
  assign n53763 = pi19 ? n53183 : n53762;
  assign n53764 = pi18 ? n20563 : n53763;
  assign n53765 = pi17 ? n53727 : n53764;
  assign n53766 = pi16 ? n32 : n53765;
  assign n53767 = pi15 ? n53756 : n53766;
  assign n53768 = pi21 ? n7263 : n32;
  assign n53769 = pi20 ? n53193 : n53768;
  assign n53770 = pi19 ? n35798 : n53769;
  assign n53771 = pi18 ? n20563 : n53770;
  assign n53772 = pi17 ? n49938 : n53771;
  assign n53773 = pi16 ? n32 : n53772;
  assign n53774 = pi21 ? n297 : n46526;
  assign n53775 = pi20 ? n53774 : n18612;
  assign n53776 = pi19 ? n32898 : n53775;
  assign n53777 = pi18 ? n20563 : n53776;
  assign n53778 = pi17 ? n49938 : n53777;
  assign n53779 = pi16 ? n32 : n53778;
  assign n53780 = pi15 ? n53773 : n53779;
  assign n53781 = pi14 ? n53767 : n53780;
  assign n53782 = pi13 ? n53751 : n53781;
  assign n53783 = pi12 ? n53721 : n53782;
  assign n53784 = pi11 ? n53687 : n53783;
  assign n53785 = pi21 ? n37 : n25463;
  assign n53786 = pi20 ? n53785 : n2653;
  assign n53787 = pi19 ? n33822 : n53786;
  assign n53788 = pi18 ? n20563 : n53787;
  assign n53789 = pi17 ? n49938 : n53788;
  assign n53790 = pi16 ? n32 : n53789;
  assign n53791 = pi21 ? n139 : n25463;
  assign n53792 = pi20 ? n53791 : n2701;
  assign n53793 = pi19 ? n33822 : n53792;
  assign n53794 = pi18 ? n20563 : n53793;
  assign n53795 = pi17 ? n49938 : n53794;
  assign n53796 = pi16 ? n32 : n53795;
  assign n53797 = pi15 ? n53790 : n53796;
  assign n53798 = pi21 ? n139 : n17463;
  assign n53799 = pi20 ? n53798 : n1822;
  assign n53800 = pi19 ? n33822 : n53799;
  assign n53801 = pi18 ? n20563 : n53800;
  assign n53802 = pi17 ? n49938 : n53801;
  assign n53803 = pi16 ? n32 : n53802;
  assign n53804 = pi21 ? n297 : n17463;
  assign n53805 = pi20 ? n53804 : n1822;
  assign n53806 = pi19 ? n32348 : n53805;
  assign n53807 = pi18 ? n20563 : n53806;
  assign n53808 = pi17 ? n48466 : n53807;
  assign n53809 = pi16 ? n32 : n53808;
  assign n53810 = pi15 ? n53803 : n53809;
  assign n53811 = pi14 ? n53797 : n53810;
  assign n53812 = pi17 ? n48466 : n53243;
  assign n53813 = pi16 ? n32 : n53812;
  assign n53814 = pi23 ? n8184 : n233;
  assign n53815 = pi22 ? n53814 : n6415;
  assign n53816 = pi21 ? n139 : n53815;
  assign n53817 = pi20 ? n53816 : n32;
  assign n53818 = pi19 ? n32898 : n53817;
  assign n53819 = pi18 ? n20563 : n53818;
  assign n53820 = pi17 ? n48466 : n53819;
  assign n53821 = pi16 ? n32 : n53820;
  assign n53822 = pi15 ? n53813 : n53821;
  assign n53823 = pi22 ? n16717 : n3338;
  assign n53824 = pi21 ? n9143 : n53823;
  assign n53825 = pi20 ? n53824 : n32;
  assign n53826 = pi19 ? n32898 : n53825;
  assign n53827 = pi18 ? n20563 : n53826;
  assign n53828 = pi17 ? n48466 : n53827;
  assign n53829 = pi16 ? n32 : n53828;
  assign n53830 = pi21 ? n335 : n1397;
  assign n53831 = pi20 ? n53830 : n32;
  assign n53832 = pi19 ? n32898 : n53831;
  assign n53833 = pi18 ? n20563 : n53832;
  assign n53834 = pi17 ? n48466 : n53833;
  assign n53835 = pi16 ? n32 : n53834;
  assign n53836 = pi15 ? n53829 : n53835;
  assign n53837 = pi14 ? n53822 : n53836;
  assign n53838 = pi13 ? n53811 : n53837;
  assign n53839 = pi23 ? n27397 : n685;
  assign n53840 = pi22 ? n53839 : n1407;
  assign n53841 = pi21 ? n335 : n53840;
  assign n53842 = pi20 ? n53841 : n32;
  assign n53843 = pi19 ? n51162 : n53842;
  assign n53844 = pi18 ? n20563 : n53843;
  assign n53845 = pi17 ? n48466 : n53844;
  assign n53846 = pi16 ? n32 : n53845;
  assign n53847 = pi21 ? n363 : n16822;
  assign n53848 = pi20 ? n53847 : n32;
  assign n53849 = pi19 ? n31221 : n53848;
  assign n53850 = pi18 ? n20563 : n53849;
  assign n53851 = pi17 ? n53229 : n53850;
  assign n53852 = pi16 ? n32 : n53851;
  assign n53853 = pi15 ? n53846 : n53852;
  assign n53854 = pi22 ? n1070 : n317;
  assign n53855 = pi21 ? n14865 : n53854;
  assign n53856 = pi20 ? n53855 : n32;
  assign n53857 = pi19 ? n31221 : n53856;
  assign n53858 = pi18 ? n20563 : n53857;
  assign n53859 = pi17 ? n49485 : n53858;
  assign n53860 = pi16 ? n32 : n53859;
  assign n53861 = pi19 ? n45600 : n53291;
  assign n53862 = pi18 ? n53861 : n53294;
  assign n53863 = pi21 ? n157 : n53854;
  assign n53864 = pi20 ? n53863 : n32;
  assign n53865 = pi19 ? n31221 : n53864;
  assign n53866 = pi18 ? n53297 : n53865;
  assign n53867 = pi17 ? n53862 : n53866;
  assign n53868 = pi16 ? n32 : n53867;
  assign n53869 = pi15 ? n53860 : n53868;
  assign n53870 = pi14 ? n53853 : n53869;
  assign n53871 = pi20 ? n32 : n49722;
  assign n53872 = pi19 ? n53871 : n53309;
  assign n53873 = pi18 ? n53872 : n20563;
  assign n53874 = pi22 ? n335 : n23156;
  assign n53875 = pi21 ? n53874 : n6416;
  assign n53876 = pi20 ? n53875 : n32;
  assign n53877 = pi19 ? n53312 : n53876;
  assign n53878 = pi18 ? n20563 : n53877;
  assign n53879 = pi17 ? n53873 : n53878;
  assign n53880 = pi16 ? n32 : n53879;
  assign n53881 = pi19 ? n53871 : n33792;
  assign n53882 = pi18 ? n53881 : n53323;
  assign n53883 = pi19 ? n53327 : n50182;
  assign n53884 = pi18 ? n53325 : n53883;
  assign n53885 = pi17 ? n53882 : n53884;
  assign n53886 = pi16 ? n32 : n53885;
  assign n53887 = pi15 ? n53880 : n53886;
  assign n53888 = pi22 ? n363 : n7780;
  assign n53889 = pi21 ? n53888 : n5829;
  assign n53890 = pi20 ? n53889 : n32;
  assign n53891 = pi19 ? n31221 : n53890;
  assign n53892 = pi18 ? n20563 : n53891;
  assign n53893 = pi17 ? n47935 : n53892;
  assign n53894 = pi16 ? n32 : n53893;
  assign n53895 = pi22 ? n52307 : n1449;
  assign n53896 = pi21 ? n53895 : n928;
  assign n53897 = pi20 ? n53896 : n32;
  assign n53898 = pi19 ? n53344 : n53897;
  assign n53899 = pi18 ? n20563 : n53898;
  assign n53900 = pi17 ? n47935 : n53899;
  assign n53901 = pi16 ? n32 : n53900;
  assign n53902 = pi15 ? n53894 : n53901;
  assign n53903 = pi14 ? n53887 : n53902;
  assign n53904 = pi13 ? n53870 : n53903;
  assign n53905 = pi12 ? n53838 : n53904;
  assign n53906 = pi17 ? n47929 : n53363;
  assign n53907 = pi16 ? n32 : n53906;
  assign n53908 = pi24 ? n139 : n36659;
  assign n53909 = pi23 ? n53908 : n157;
  assign n53910 = pi22 ? n53909 : n685;
  assign n53911 = pi21 ? n53910 : n1009;
  assign n53912 = pi20 ? n53911 : n32;
  assign n53913 = pi19 ? n53368 : n53912;
  assign n53914 = pi18 ? n20563 : n53913;
  assign n53915 = pi17 ? n47929 : n53914;
  assign n53916 = pi16 ? n32 : n53915;
  assign n53917 = pi15 ? n53907 : n53916;
  assign n53918 = pi17 ? n52611 : n53382;
  assign n53919 = pi16 ? n32 : n53918;
  assign n53920 = pi17 ? n52611 : n53390;
  assign n53921 = pi16 ? n32 : n53920;
  assign n53922 = pi15 ? n53919 : n53921;
  assign n53923 = pi14 ? n53917 : n53922;
  assign n53924 = pi17 ? n52611 : n53402;
  assign n53925 = pi16 ? n32 : n53924;
  assign n53926 = pi21 ? n45620 : n39801;
  assign n53927 = pi20 ? n32 : n53926;
  assign n53928 = pi19 ? n53927 : n30868;
  assign n53929 = pi18 ? n53928 : n43012;
  assign n53930 = pi23 ? n204 : n14626;
  assign n53931 = pi22 ? n53930 : n396;
  assign n53932 = pi21 ? n53931 : n32;
  assign n53933 = pi20 ? n53932 : n32;
  assign n53934 = pi19 ? n53410 : n53933;
  assign n53935 = pi18 ? n20563 : n53934;
  assign n53936 = pi17 ? n53929 : n53935;
  assign n53937 = pi16 ? n32 : n53936;
  assign n53938 = pi15 ? n53925 : n53937;
  assign n53939 = pi19 ? n53927 : n53418;
  assign n53940 = pi18 ? n53939 : n20563;
  assign n53941 = pi17 ? n53940 : n53425;
  assign n53942 = pi16 ? n32 : n53941;
  assign n53943 = pi21 ? n45598 : n20563;
  assign n53944 = pi20 ? n32 : n53943;
  assign n53945 = pi19 ? n53944 : n20563;
  assign n53946 = pi18 ? n53945 : n20563;
  assign n53947 = pi17 ? n53946 : n53436;
  assign n53948 = pi16 ? n32 : n53947;
  assign n53949 = pi15 ? n53942 : n53948;
  assign n53950 = pi14 ? n53938 : n53949;
  assign n53951 = pi13 ? n53923 : n53950;
  assign n53952 = pi20 ? n32 : n47322;
  assign n53953 = pi19 ? n53952 : n30868;
  assign n53954 = pi18 ? n53953 : n30868;
  assign n53955 = pi17 ? n53954 : n53447;
  assign n53956 = pi16 ? n32 : n53955;
  assign n53957 = pi20 ? n41565 : n53453;
  assign n53958 = pi19 ? n53957 : n5831;
  assign n53959 = pi18 ? n30868 : n53958;
  assign n53960 = pi17 ? n53954 : n53959;
  assign n53961 = pi16 ? n32 : n53960;
  assign n53962 = pi15 ? n53956 : n53961;
  assign n53963 = pi20 ? n32 : n49815;
  assign n53964 = pi19 ? n53963 : n36798;
  assign n53965 = pi18 ? n53964 : n53466;
  assign n53966 = pi17 ? n53965 : n53475;
  assign n53967 = pi16 ? n32 : n53966;
  assign n53968 = pi20 ? n32 : n49845;
  assign n53969 = pi19 ? n53968 : n53482;
  assign n53970 = pi18 ? n53969 : n53487;
  assign n53971 = pi17 ? n53970 : n53492;
  assign n53972 = pi16 ? n32 : n53971;
  assign n53973 = pi15 ? n53967 : n53972;
  assign n53974 = pi14 ? n53962 : n53973;
  assign n53975 = pi22 ? n36659 : n50792;
  assign n53976 = pi21 ? n53975 : n36659;
  assign n53977 = pi22 ? n43198 : n50339;
  assign n53978 = pi21 ? n53977 : n50796;
  assign n53979 = pi20 ? n53976 : n53978;
  assign n53980 = pi19 ? n53968 : n53979;
  assign n53981 = pi18 ? n53980 : n36659;
  assign n53982 = pi23 ? n51565 : n32;
  assign n53983 = pi22 ? n53982 : n32;
  assign n53984 = pi21 ? n53983 : n32;
  assign n53985 = pi20 ? n53984 : n32;
  assign n53986 = pi19 ? n53502 : n53985;
  assign n53987 = pi18 ? n36659 : n53986;
  assign n53988 = pi17 ? n53981 : n53987;
  assign n53989 = pi16 ? n32 : n53988;
  assign n53990 = pi22 ? n46789 : n36659;
  assign n53991 = pi21 ? n32 : n53990;
  assign n53992 = pi20 ? n32 : n53991;
  assign n53993 = pi21 ? n37878 : n36659;
  assign n53994 = pi20 ? n37878 : n53993;
  assign n53995 = pi19 ? n53992 : n53994;
  assign n53996 = pi18 ? n53995 : n53518;
  assign n53997 = pi17 ? n53996 : n53531;
  assign n53998 = pi16 ? n32 : n53997;
  assign n53999 = pi15 ? n53989 : n53998;
  assign n54000 = pi22 ? n46275 : n36781;
  assign n54001 = pi21 ? n32 : n54000;
  assign n54002 = pi20 ? n32 : n54001;
  assign n54003 = pi19 ? n54002 : n36781;
  assign n54004 = pi18 ? n54003 : n36781;
  assign n54005 = pi17 ? n54004 : n53546;
  assign n54006 = pi16 ? n32 : n54005;
  assign n54007 = pi21 ? n32 : n47902;
  assign n54008 = pi20 ? n32 : n54007;
  assign n54009 = pi21 ? n47397 : n43198;
  assign n54010 = pi20 ? n54009 : n47396;
  assign n54011 = pi19 ? n54008 : n54010;
  assign n54012 = pi18 ? n54011 : n53557;
  assign n54013 = pi17 ? n54012 : n53563;
  assign n54014 = pi16 ? n32 : n54013;
  assign n54015 = pi15 ? n54006 : n54014;
  assign n54016 = pi14 ? n53999 : n54015;
  assign n54017 = pi13 ? n53974 : n54016;
  assign n54018 = pi12 ? n53951 : n54017;
  assign n54019 = pi11 ? n53905 : n54018;
  assign n54020 = pi10 ? n53784 : n54019;
  assign n54021 = pi09 ? n53588 : n54020;
  assign n54022 = pi08 ? n53572 : n54021;
  assign n54023 = pi20 ? n46815 : n30096;
  assign n54024 = pi21 ? n297 : n8015;
  assign n54025 = pi20 ? n37 : n54024;
  assign n54026 = pi19 ? n54023 : n54025;
  assign n54027 = pi18 ? n20563 : n54026;
  assign n54028 = pi17 ? n46447 : n54027;
  assign n54029 = pi16 ? n32 : n54028;
  assign n54030 = pi15 ? n32 : n54029;
  assign n54031 = pi21 ? n297 : n8557;
  assign n54032 = pi20 ? n37 : n54031;
  assign n54033 = pi19 ? n32898 : n54032;
  assign n54034 = pi18 ? n20563 : n54033;
  assign n54035 = pi17 ? n39374 : n54034;
  assign n54036 = pi16 ? n32 : n54035;
  assign n54037 = pi21 ? n30867 : n31889;
  assign n54038 = pi20 ? n54037 : n20563;
  assign n54039 = pi19 ? n20563 : n54038;
  assign n54040 = pi21 ? n35230 : n20563;
  assign n54041 = pi20 ? n54040 : n30096;
  assign n54042 = pi21 ? n569 : n8557;
  assign n54043 = pi20 ? n37 : n54042;
  assign n54044 = pi19 ? n54041 : n54043;
  assign n54045 = pi18 ? n54039 : n54044;
  assign n54046 = pi17 ? n39374 : n54045;
  assign n54047 = pi16 ? n32 : n54046;
  assign n54048 = pi15 ? n54036 : n54047;
  assign n54049 = pi14 ? n54030 : n54048;
  assign n54050 = pi13 ? n32 : n54049;
  assign n54051 = pi12 ? n32 : n54050;
  assign n54052 = pi11 ? n32 : n54051;
  assign n54053 = pi10 ? n32 : n54052;
  assign n54054 = pi19 ? n40531 : n38962;
  assign n54055 = pi18 ? n32 : n54054;
  assign n54056 = pi21 ? n37 : n31294;
  assign n54057 = pi20 ? n54056 : n20563;
  assign n54058 = pi19 ? n32294 : n54057;
  assign n54059 = pi21 ? n20228 : n8044;
  assign n54060 = pi20 ? n3086 : n54059;
  assign n54061 = pi19 ? n37 : n54060;
  assign n54062 = pi18 ? n54058 : n54061;
  assign n54063 = pi17 ? n54055 : n54062;
  assign n54064 = pi16 ? n32 : n54063;
  assign n54065 = pi20 ? n20563 : n47432;
  assign n54066 = pi19 ? n41707 : n54065;
  assign n54067 = pi18 ? n32 : n54066;
  assign n54068 = pi21 ? n31885 : n20563;
  assign n54069 = pi20 ? n54068 : n31266;
  assign n54070 = pi21 ? n36249 : n31294;
  assign n54071 = pi20 ? n54070 : n31266;
  assign n54072 = pi19 ? n54069 : n54071;
  assign n54073 = pi21 ? n29838 : n2469;
  assign n54074 = pi20 ? n37 : n54073;
  assign n54075 = pi19 ? n37 : n54074;
  assign n54076 = pi18 ? n54072 : n54075;
  assign n54077 = pi17 ? n54067 : n54076;
  assign n54078 = pi16 ? n32 : n54077;
  assign n54079 = pi15 ? n54064 : n54078;
  assign n54080 = pi20 ? n20563 : n38966;
  assign n54081 = pi19 ? n54080 : n35854;
  assign n54082 = pi20 ? n36250 : n37;
  assign n54083 = pi19 ? n54082 : n26630;
  assign n54084 = pi18 ? n54081 : n54083;
  assign n54085 = pi17 ? n38949 : n54084;
  assign n54086 = pi16 ? n32 : n54085;
  assign n54087 = pi22 ? n37 : n3935;
  assign n54088 = pi21 ? n54087 : n32;
  assign n54089 = pi20 ? n37 : n54088;
  assign n54090 = pi19 ? n38522 : n54089;
  assign n54091 = pi18 ? n48972 : n54090;
  assign n54092 = pi17 ? n40046 : n54091;
  assign n54093 = pi16 ? n32 : n54092;
  assign n54094 = pi15 ? n54086 : n54093;
  assign n54095 = pi14 ? n54079 : n54094;
  assign n54096 = pi20 ? n37 : n22814;
  assign n54097 = pi19 ? n31267 : n54096;
  assign n54098 = pi18 ? n20563 : n54097;
  assign n54099 = pi17 ? n40046 : n54098;
  assign n54100 = pi16 ? n32 : n54099;
  assign n54101 = pi19 ? n20563 : n51932;
  assign n54102 = pi18 ? n37928 : n54101;
  assign n54103 = pi20 ? n20563 : n47433;
  assign n54104 = pi20 ? n54068 : n36929;
  assign n54105 = pi19 ? n54103 : n54104;
  assign n54106 = pi20 ? n37 : n11200;
  assign n54107 = pi19 ? n31280 : n54106;
  assign n54108 = pi18 ? n54105 : n54107;
  assign n54109 = pi17 ? n54102 : n54108;
  assign n54110 = pi16 ? n32 : n54109;
  assign n54111 = pi15 ? n54100 : n54110;
  assign n54112 = pi19 ? n37 : n54106;
  assign n54113 = pi18 ? n53013 : n54112;
  assign n54114 = pi17 ? n38984 : n54113;
  assign n54115 = pi16 ? n32 : n54114;
  assign n54116 = pi21 ? n30843 : n31877;
  assign n54117 = pi20 ? n54116 : n38966;
  assign n54118 = pi19 ? n20563 : n54117;
  assign n54119 = pi18 ? n40056 : n54118;
  assign n54120 = pi21 ? n31885 : n31294;
  assign n54121 = pi20 ? n54120 : n37;
  assign n54122 = pi19 ? n50854 : n54121;
  assign n54123 = pi20 ? n37 : n22836;
  assign n54124 = pi19 ? n37 : n54123;
  assign n54125 = pi18 ? n54122 : n54124;
  assign n54126 = pi17 ? n54119 : n54125;
  assign n54127 = pi16 ? n32 : n54126;
  assign n54128 = pi15 ? n54115 : n54127;
  assign n54129 = pi14 ? n54111 : n54128;
  assign n54130 = pi13 ? n54095 : n54129;
  assign n54131 = pi19 ? n50906 : n31267;
  assign n54132 = pi22 ? n37 : n6365;
  assign n54133 = pi21 ? n54132 : n32;
  assign n54134 = pi20 ? n37 : n54133;
  assign n54135 = pi19 ? n37 : n54134;
  assign n54136 = pi18 ? n54131 : n54135;
  assign n54137 = pi17 ? n37936 : n54136;
  assign n54138 = pi16 ? n32 : n54137;
  assign n54139 = pi20 ? n37 : n49916;
  assign n54140 = pi22 ? n99 : n1475;
  assign n54141 = pi21 ? n54140 : n32;
  assign n54142 = pi20 ? n30096 : n54141;
  assign n54143 = pi19 ? n54139 : n54142;
  assign n54144 = pi18 ? n37441 : n54143;
  assign n54145 = pi17 ? n37958 : n54144;
  assign n54146 = pi16 ? n32 : n54145;
  assign n54147 = pi15 ? n54138 : n54146;
  assign n54148 = pi20 ? n30096 : n24850;
  assign n54149 = pi19 ? n51953 : n54148;
  assign n54150 = pi18 ? n20563 : n54149;
  assign n54151 = pi17 ? n36162 : n54150;
  assign n54152 = pi16 ? n32 : n54151;
  assign n54153 = pi21 ? n30195 : n20563;
  assign n54154 = pi20 ? n31925 : n54153;
  assign n54155 = pi21 ? n31877 : n20563;
  assign n54156 = pi20 ? n31913 : n54155;
  assign n54157 = pi19 ? n54154 : n54156;
  assign n54158 = pi21 ? n37 : n31877;
  assign n54159 = pi20 ? n37 : n54158;
  assign n54160 = pi23 ? n685 : n1149;
  assign n54161 = pi22 ? n37 : n54160;
  assign n54162 = pi21 ? n54161 : n32;
  assign n54163 = pi20 ? n30096 : n54162;
  assign n54164 = pi19 ? n54159 : n54163;
  assign n54165 = pi18 ? n54157 : n54164;
  assign n54166 = pi17 ? n36162 : n54165;
  assign n54167 = pi16 ? n32 : n54166;
  assign n54168 = pi15 ? n54152 : n54167;
  assign n54169 = pi14 ? n54147 : n54168;
  assign n54170 = pi20 ? n54068 : n20563;
  assign n54171 = pi19 ? n20563 : n54170;
  assign n54172 = pi18 ? n28159 : n54171;
  assign n54173 = pi22 ? n37 : n730;
  assign n54174 = pi21 ? n54173 : n32;
  assign n54175 = pi20 ? n37 : n54174;
  assign n54176 = pi19 ? n37 : n54175;
  assign n54177 = pi18 ? n54131 : n54176;
  assign n54178 = pi17 ? n54172 : n54177;
  assign n54179 = pi16 ? n32 : n54178;
  assign n54180 = pi19 ? n32876 : n20563;
  assign n54181 = pi18 ? n31265 : n54180;
  assign n54182 = pi20 ? n31903 : n52962;
  assign n54183 = pi19 ? n54182 : n32287;
  assign n54184 = pi21 ? n17806 : n32;
  assign n54185 = pi20 ? n37 : n54184;
  assign n54186 = pi19 ? n37 : n54185;
  assign n54187 = pi18 ? n54183 : n54186;
  assign n54188 = pi17 ? n54181 : n54187;
  assign n54189 = pi16 ? n32 : n54188;
  assign n54190 = pi15 ? n54179 : n54189;
  assign n54191 = pi18 ? n34295 : n54186;
  assign n54192 = pi17 ? n36215 : n54191;
  assign n54193 = pi16 ? n32 : n54192;
  assign n54194 = pi20 ? n37 : n11215;
  assign n54195 = pi19 ? n51953 : n54194;
  assign n54196 = pi18 ? n34258 : n54195;
  assign n54197 = pi17 ? n36215 : n54196;
  assign n54198 = pi16 ? n32 : n54197;
  assign n54199 = pi15 ? n54193 : n54198;
  assign n54200 = pi14 ? n54190 : n54199;
  assign n54201 = pi13 ? n54169 : n54200;
  assign n54202 = pi12 ? n54130 : n54201;
  assign n54203 = pi22 ? n5011 : n316;
  assign n54204 = pi21 ? n54203 : n32;
  assign n54205 = pi20 ? n30096 : n54204;
  assign n54206 = pi19 ? n53104 : n54205;
  assign n54207 = pi18 ? n20563 : n54206;
  assign n54208 = pi17 ? n36215 : n54207;
  assign n54209 = pi16 ? n32 : n54208;
  assign n54210 = pi20 ? n33845 : n20563;
  assign n54211 = pi20 ? n36929 : n31220;
  assign n54212 = pi19 ? n54210 : n54211;
  assign n54213 = pi20 ? n37 : n53577;
  assign n54214 = pi22 ? n112 : n1511;
  assign n54215 = pi21 ? n54214 : n32;
  assign n54216 = pi20 ? n37 : n54215;
  assign n54217 = pi19 ? n54213 : n54216;
  assign n54218 = pi18 ? n54212 : n54217;
  assign n54219 = pi17 ? n50390 : n54218;
  assign n54220 = pi16 ? n32 : n54219;
  assign n54221 = pi15 ? n54209 : n54220;
  assign n54222 = pi19 ? n32294 : n20563;
  assign n54223 = pi18 ? n44686 : n54222;
  assign n54224 = pi19 ? n53051 : n32933;
  assign n54225 = pi22 ? n893 : n430;
  assign n54226 = pi21 ? n54225 : n32;
  assign n54227 = pi20 ? n37 : n54226;
  assign n54228 = pi19 ? n37 : n54227;
  assign n54229 = pi18 ? n54224 : n54228;
  assign n54230 = pi17 ? n54223 : n54229;
  assign n54231 = pi16 ? n32 : n54230;
  assign n54232 = pi18 ? n43217 : n34865;
  assign n54233 = pi21 ? n30843 : n20563;
  assign n54234 = pi20 ? n54233 : n20563;
  assign n54235 = pi19 ? n54234 : n31280;
  assign n54236 = pi20 ? n6434 : n25822;
  assign n54237 = pi19 ? n37 : n54236;
  assign n54238 = pi18 ? n54235 : n54237;
  assign n54239 = pi17 ? n54232 : n54238;
  assign n54240 = pi16 ? n32 : n54239;
  assign n54241 = pi15 ? n54231 : n54240;
  assign n54242 = pi14 ? n54221 : n54241;
  assign n54243 = pi20 ? n48905 : n31925;
  assign n54244 = pi22 ? n157 : n664;
  assign n54245 = pi21 ? n54244 : n32;
  assign n54246 = pi20 ? n24493 : n54245;
  assign n54247 = pi19 ? n54243 : n54246;
  assign n54248 = pi18 ? n34869 : n54247;
  assign n54249 = pi17 ? n49888 : n54248;
  assign n54250 = pi16 ? n32 : n54249;
  assign n54251 = pi20 ? n5077 : n5667;
  assign n54252 = pi19 ? n53104 : n54251;
  assign n54253 = pi18 ? n34869 : n54252;
  assign n54254 = pi17 ? n49888 : n54253;
  assign n54255 = pi16 ? n32 : n54254;
  assign n54256 = pi15 ? n54250 : n54255;
  assign n54257 = pi20 ? n24493 : n5667;
  assign n54258 = pi19 ? n53104 : n54257;
  assign n54259 = pi18 ? n20563 : n54258;
  assign n54260 = pi17 ? n49888 : n54259;
  assign n54261 = pi16 ? n32 : n54260;
  assign n54262 = pi20 ? n36872 : n20563;
  assign n54263 = pi20 ? n54040 : n20563;
  assign n54264 = pi19 ? n54262 : n54263;
  assign n54265 = pi20 ? n48905 : n37439;
  assign n54266 = pi19 ? n54265 : n53722;
  assign n54267 = pi18 ? n54264 : n54266;
  assign n54268 = pi17 ? n49888 : n54267;
  assign n54269 = pi16 ? n32 : n54268;
  assign n54270 = pi15 ? n54261 : n54269;
  assign n54271 = pi14 ? n54256 : n54270;
  assign n54272 = pi13 ? n54242 : n54271;
  assign n54273 = pi18 ? n44273 : n20563;
  assign n54274 = pi19 ? n53104 : n32348;
  assign n54275 = pi21 ? n37 : n15305;
  assign n54276 = pi20 ? n54275 : n5667;
  assign n54277 = pi19 ? n37 : n54276;
  assign n54278 = pi18 ? n54274 : n54277;
  assign n54279 = pi17 ? n54273 : n54278;
  assign n54280 = pi16 ? n32 : n54279;
  assign n54281 = pi21 ? n181 : n22940;
  assign n54282 = pi20 ? n54281 : n24937;
  assign n54283 = pi19 ? n51996 : n54282;
  assign n54284 = pi18 ? n34869 : n54283;
  assign n54285 = pi17 ? n49900 : n54284;
  assign n54286 = pi16 ? n32 : n54285;
  assign n54287 = pi15 ? n54280 : n54286;
  assign n54288 = pi19 ? n53344 : n53159;
  assign n54289 = pi18 ? n20563 : n54288;
  assign n54290 = pi17 ? n49900 : n54289;
  assign n54291 = pi16 ? n32 : n54290;
  assign n54292 = pi20 ? n22941 : n3210;
  assign n54293 = pi19 ? n32294 : n54292;
  assign n54294 = pi18 ? n20563 : n54293;
  assign n54295 = pi17 ? n49900 : n54294;
  assign n54296 = pi16 ? n32 : n54295;
  assign n54297 = pi15 ? n54291 : n54296;
  assign n54298 = pi14 ? n54287 : n54297;
  assign n54299 = pi20 ? n14927 : n6417;
  assign n54300 = pi19 ? n32294 : n54299;
  assign n54301 = pi18 ? n20563 : n54300;
  assign n54302 = pi17 ? n49900 : n54301;
  assign n54303 = pi16 ? n32 : n54302;
  assign n54304 = pi20 ? n14927 : n4116;
  assign n54305 = pi19 ? n51069 : n54304;
  assign n54306 = pi18 ? n20563 : n54305;
  assign n54307 = pi17 ? n49900 : n54306;
  assign n54308 = pi16 ? n32 : n54307;
  assign n54309 = pi15 ? n54303 : n54308;
  assign n54310 = pi20 ? n21732 : n5830;
  assign n54311 = pi19 ? n32294 : n54310;
  assign n54312 = pi18 ? n20563 : n54311;
  assign n54313 = pi17 ? n50426 : n54312;
  assign n54314 = pi16 ? n32 : n54313;
  assign n54315 = pi21 ? n37 : n11808;
  assign n54316 = pi20 ? n54315 : n10011;
  assign n54317 = pi19 ? n32294 : n54316;
  assign n54318 = pi18 ? n20563 : n54317;
  assign n54319 = pi17 ? n50426 : n54318;
  assign n54320 = pi16 ? n32 : n54319;
  assign n54321 = pi15 ? n54314 : n54320;
  assign n54322 = pi14 ? n54309 : n54321;
  assign n54323 = pi13 ? n54298 : n54322;
  assign n54324 = pi12 ? n54272 : n54323;
  assign n54325 = pi11 ? n54202 : n54324;
  assign n54326 = pi21 ? n37 : n29992;
  assign n54327 = pi20 ? n54326 : n2653;
  assign n54328 = pi19 ? n32294 : n54327;
  assign n54329 = pi18 ? n20563 : n54328;
  assign n54330 = pi17 ? n50426 : n54329;
  assign n54331 = pi16 ? n32 : n54330;
  assign n54332 = pi20 ? n51634 : n2701;
  assign n54333 = pi19 ? n32294 : n54332;
  assign n54334 = pi18 ? n20563 : n54333;
  assign n54335 = pi17 ? n50426 : n54334;
  assign n54336 = pi16 ? n32 : n54335;
  assign n54337 = pi15 ? n54331 : n54336;
  assign n54338 = pi22 ? n4537 : n2299;
  assign n54339 = pi21 ? n139 : n54338;
  assign n54340 = pi20 ? n54339 : n1822;
  assign n54341 = pi19 ? n32294 : n54340;
  assign n54342 = pi18 ? n20563 : n54341;
  assign n54343 = pi17 ? n50426 : n54342;
  assign n54344 = pi16 ? n32 : n54343;
  assign n54345 = pi22 ? n51509 : n316;
  assign n54346 = pi21 ? n37 : n54345;
  assign n54347 = pi20 ? n54346 : n1822;
  assign n54348 = pi19 ? n31221 : n54347;
  assign n54349 = pi18 ? n20563 : n54348;
  assign n54350 = pi17 ? n48904 : n54349;
  assign n54351 = pi16 ? n32 : n54350;
  assign n54352 = pi15 ? n54344 : n54351;
  assign n54353 = pi14 ? n54337 : n54352;
  assign n54354 = pi21 ? n20563 : n99;
  assign n54355 = pi20 ? n20563 : n54354;
  assign n54356 = pi23 ? n3491 : n157;
  assign n54357 = pi22 ? n54356 : n233;
  assign n54358 = pi21 ? n37 : n54357;
  assign n54359 = pi20 ? n54358 : n32;
  assign n54360 = pi19 ? n54355 : n54359;
  assign n54361 = pi18 ? n20563 : n54360;
  assign n54362 = pi17 ? n48904 : n54361;
  assign n54363 = pi16 ? n32 : n54362;
  assign n54364 = pi23 ? n11962 : n233;
  assign n54365 = pi22 ? n54364 : n6365;
  assign n54366 = pi21 ? n139 : n54365;
  assign n54367 = pi20 ? n54366 : n32;
  assign n54368 = pi19 ? n32294 : n54367;
  assign n54369 = pi18 ? n20563 : n54368;
  assign n54370 = pi17 ? n48904 : n54369;
  assign n54371 = pi16 ? n32 : n54370;
  assign n54372 = pi15 ? n54363 : n54371;
  assign n54373 = pi23 ? n3134 : n233;
  assign n54374 = pi22 ? n54373 : n1070;
  assign n54375 = pi21 ? n4247 : n54374;
  assign n54376 = pi20 ? n54375 : n32;
  assign n54377 = pi19 ? n32294 : n54376;
  assign n54378 = pi18 ? n20563 : n54377;
  assign n54379 = pi17 ? n48904 : n54378;
  assign n54380 = pi16 ? n32 : n54379;
  assign n54381 = pi22 ? n673 : n3338;
  assign n54382 = pi21 ? n335 : n54381;
  assign n54383 = pi20 ? n54382 : n32;
  assign n54384 = pi19 ? n32294 : n54383;
  assign n54385 = pi18 ? n20563 : n54384;
  assign n54386 = pi17 ? n48904 : n54385;
  assign n54387 = pi16 ? n32 : n54386;
  assign n54388 = pi15 ? n54380 : n54387;
  assign n54389 = pi14 ? n54372 : n54388;
  assign n54390 = pi13 ? n54353 : n54389;
  assign n54391 = pi18 ? n41630 : n20563;
  assign n54392 = pi21 ? n45016 : n29133;
  assign n54393 = pi20 ? n20563 : n54392;
  assign n54394 = pi21 ? n335 : n53398;
  assign n54395 = pi20 ? n54394 : n32;
  assign n54396 = pi19 ? n54393 : n54395;
  assign n54397 = pi18 ? n20563 : n54396;
  assign n54398 = pi17 ? n54391 : n54397;
  assign n54399 = pi16 ? n32 : n54398;
  assign n54400 = pi22 ? n46165 : n20563;
  assign n54401 = pi21 ? n32 : n54400;
  assign n54402 = pi20 ? n32 : n54401;
  assign n54403 = pi19 ? n54402 : n20563;
  assign n54404 = pi18 ? n54403 : n20563;
  assign n54405 = pi22 ? n1457 : n1407;
  assign n54406 = pi21 ? n363 : n54405;
  assign n54407 = pi20 ? n54406 : n32;
  assign n54408 = pi19 ? n32294 : n54407;
  assign n54409 = pi18 ? n20563 : n54408;
  assign n54410 = pi17 ? n54404 : n54409;
  assign n54411 = pi16 ? n32 : n54410;
  assign n54412 = pi15 ? n54399 : n54411;
  assign n54413 = pi21 ? n48173 : n39801;
  assign n54414 = pi21 ? n20563 : n40913;
  assign n54415 = pi20 ? n54413 : n54414;
  assign n54416 = pi19 ? n46062 : n54415;
  assign n54417 = pi21 ? n45049 : n20563;
  assign n54418 = pi20 ? n54417 : n20563;
  assign n54419 = pi19 ? n54418 : n20563;
  assign n54420 = pi18 ? n54416 : n54419;
  assign n54421 = pi21 ? n14865 : n8916;
  assign n54422 = pi20 ? n54421 : n32;
  assign n54423 = pi19 ? n20563 : n54422;
  assign n54424 = pi18 ? n20563 : n54423;
  assign n54425 = pi17 ? n54420 : n54424;
  assign n54426 = pi16 ? n32 : n54425;
  assign n54427 = pi22 ? n45516 : n30868;
  assign n54428 = pi21 ? n32 : n54427;
  assign n54429 = pi20 ? n32 : n54428;
  assign n54430 = pi19 ? n54429 : n30868;
  assign n54431 = pi20 ? n40915 : n30868;
  assign n54432 = pi19 ? n30868 : n54431;
  assign n54433 = pi18 ? n54430 : n54432;
  assign n54434 = pi19 ? n54431 : n20563;
  assign n54435 = pi20 ? n38754 : n31220;
  assign n54436 = pi21 ? n157 : n2230;
  assign n54437 = pi20 ? n54436 : n32;
  assign n54438 = pi19 ? n54435 : n54437;
  assign n54439 = pi18 ? n54434 : n54438;
  assign n54440 = pi17 ? n54433 : n54439;
  assign n54441 = pi16 ? n32 : n54440;
  assign n54442 = pi15 ? n54426 : n54441;
  assign n54443 = pi14 ? n54412 : n54442;
  assign n54444 = pi21 ? n32 : n52259;
  assign n54445 = pi20 ? n32 : n54444;
  assign n54446 = pi22 ? n37173 : n33792;
  assign n54447 = pi21 ? n54446 : n40957;
  assign n54448 = pi20 ? n54447 : n41486;
  assign n54449 = pi19 ? n54445 : n54448;
  assign n54450 = pi21 ? n40954 : n20563;
  assign n54451 = pi20 ? n54450 : n20563;
  assign n54452 = pi19 ? n54451 : n20563;
  assign n54453 = pi18 ? n54449 : n54452;
  assign n54454 = pi21 ? n7986 : n8486;
  assign n54455 = pi20 ? n54454 : n32;
  assign n54456 = pi19 ? n53312 : n54455;
  assign n54457 = pi18 ? n20563 : n54456;
  assign n54458 = pi17 ? n54453 : n54457;
  assign n54459 = pi16 ? n32 : n54458;
  assign n54460 = pi22 ? n36615 : n37173;
  assign n54461 = pi21 ? n45008 : n54460;
  assign n54462 = pi21 ? n51744 : n40957;
  assign n54463 = pi20 ? n54461 : n54462;
  assign n54464 = pi19 ? n54445 : n54463;
  assign n54465 = pi21 ? n40955 : n37173;
  assign n54466 = pi21 ? n40954 : n45526;
  assign n54467 = pi20 ? n54465 : n54466;
  assign n54468 = pi21 ? n20563 : n40957;
  assign n54469 = pi21 ? n33792 : n37173;
  assign n54470 = pi20 ? n54468 : n54469;
  assign n54471 = pi19 ? n54467 : n54470;
  assign n54472 = pi18 ? n54464 : n54471;
  assign n54473 = pi21 ? n36615 : n37768;
  assign n54474 = pi21 ? n37768 : n33792;
  assign n54475 = pi20 ? n54473 : n54474;
  assign n54476 = pi19 ? n54475 : n20563;
  assign n54477 = pi21 ? n36837 : n3523;
  assign n54478 = pi20 ? n54477 : n32;
  assign n54479 = pi19 ? n53327 : n54478;
  assign n54480 = pi18 ? n54476 : n54479;
  assign n54481 = pi17 ? n54472 : n54480;
  assign n54482 = pi16 ? n32 : n54481;
  assign n54483 = pi15 ? n54459 : n54482;
  assign n54484 = pi21 ? n5054 : n2320;
  assign n54485 = pi20 ? n54484 : n32;
  assign n54486 = pi19 ? n31221 : n54485;
  assign n54487 = pi18 ? n20563 : n54486;
  assign n54488 = pi17 ? n48469 : n54487;
  assign n54489 = pi16 ? n32 : n54488;
  assign n54490 = pi22 ? n52307 : n204;
  assign n54491 = pi21 ? n54490 : n882;
  assign n54492 = pi20 ? n54491 : n32;
  assign n54493 = pi19 ? n53344 : n54492;
  assign n54494 = pi18 ? n20563 : n54493;
  assign n54495 = pi17 ? n48466 : n54494;
  assign n54496 = pi16 ? n32 : n54495;
  assign n54497 = pi15 ? n54489 : n54496;
  assign n54498 = pi14 ? n54483 : n54497;
  assign n54499 = pi13 ? n54443 : n54498;
  assign n54500 = pi12 ? n54390 : n54499;
  assign n54501 = pi21 ? n53359 : n882;
  assign n54502 = pi20 ? n54501 : n32;
  assign n54503 = pi19 ? n53357 : n54502;
  assign n54504 = pi18 ? n20563 : n54503;
  assign n54505 = pi17 ? n48466 : n54504;
  assign n54506 = pi16 ? n32 : n54505;
  assign n54507 = pi21 ? n53370 : n53983;
  assign n54508 = pi20 ? n54507 : n32;
  assign n54509 = pi19 ? n53368 : n54508;
  assign n54510 = pi18 ? n20563 : n54509;
  assign n54511 = pi17 ? n48466 : n54510;
  assign n54512 = pi16 ? n32 : n54511;
  assign n54513 = pi15 ? n54506 : n54512;
  assign n54514 = pi17 ? n48460 : n53382;
  assign n54515 = pi16 ? n32 : n54514;
  assign n54516 = pi17 ? n53151 : n53390;
  assign n54517 = pi16 ? n32 : n54516;
  assign n54518 = pi15 ? n54515 : n54517;
  assign n54519 = pi14 ? n54513 : n54518;
  assign n54520 = pi23 ? n685 : n51565;
  assign n54521 = pi22 ? n1457 : n54520;
  assign n54522 = pi21 ? n54521 : n32;
  assign n54523 = pi20 ? n54522 : n32;
  assign n54524 = pi19 ? n53397 : n54523;
  assign n54525 = pi18 ? n20563 : n54524;
  assign n54526 = pi17 ? n53151 : n54525;
  assign n54527 = pi16 ? n32 : n54526;
  assign n54528 = pi18 ? n48805 : n43012;
  assign n54529 = pi22 ? n14626 : n396;
  assign n54530 = pi21 ? n54529 : n32;
  assign n54531 = pi20 ? n54530 : n32;
  assign n54532 = pi19 ? n53410 : n54531;
  assign n54533 = pi18 ? n20563 : n54532;
  assign n54534 = pi17 ? n54528 : n54533;
  assign n54535 = pi16 ? n32 : n54534;
  assign n54536 = pi15 ? n54527 : n54535;
  assign n54537 = pi20 ? n30868 : n42005;
  assign n54538 = pi19 ? n46168 : n54537;
  assign n54539 = pi19 ? n51203 : n20563;
  assign n54540 = pi18 ? n54538 : n54539;
  assign n54541 = pi17 ? n54540 : n53425;
  assign n54542 = pi16 ? n32 : n54541;
  assign n54543 = pi20 ? n50735 : n20563;
  assign n54544 = pi19 ? n40055 : n54543;
  assign n54545 = pi18 ? n54544 : n20563;
  assign n54546 = pi22 ? n316 : n53982;
  assign n54547 = pi21 ? n54546 : n32;
  assign n54548 = pi20 ? n54547 : n32;
  assign n54549 = pi19 ? n53434 : n54548;
  assign n54550 = pi18 ? n20563 : n54549;
  assign n54551 = pi17 ? n54545 : n54550;
  assign n54552 = pi16 ? n32 : n54551;
  assign n54553 = pi15 ? n54542 : n54552;
  assign n54554 = pi14 ? n54536 : n54553;
  assign n54555 = pi13 ? n54519 : n54554;
  assign n54556 = pi19 ? n51815 : n30868;
  assign n54557 = pi18 ? n54556 : n30868;
  assign n54558 = pi17 ? n54557 : n53447;
  assign n54559 = pi16 ? n32 : n54558;
  assign n54560 = pi22 ? n30868 : n49800;
  assign n54561 = pi21 ? n54560 : n51564;
  assign n54562 = pi20 ? n30868 : n54561;
  assign n54563 = pi23 ? n51564 : n395;
  assign n54564 = pi22 ? n54563 : n32;
  assign n54565 = pi21 ? n54564 : n32;
  assign n54566 = pi20 ? n54565 : n32;
  assign n54567 = pi19 ? n54562 : n54566;
  assign n54568 = pi18 ? n30868 : n54567;
  assign n54569 = pi17 ? n54557 : n54568;
  assign n54570 = pi16 ? n32 : n54569;
  assign n54571 = pi15 ? n54559 : n54570;
  assign n54572 = pi20 ? n32 : n52918;
  assign n54573 = pi19 ? n54572 : n36798;
  assign n54574 = pi23 ? n33792 : n36798;
  assign n54575 = pi22 ? n36798 : n54574;
  assign n54576 = pi21 ? n53463 : n54575;
  assign n54577 = pi20 ? n50300 : n54576;
  assign n54578 = pi19 ? n36798 : n54577;
  assign n54579 = pi18 ? n54573 : n54578;
  assign n54580 = pi23 ? n36798 : n33792;
  assign n54581 = pi22 ? n33792 : n54580;
  assign n54582 = pi21 ? n54581 : n33792;
  assign n54583 = pi20 ? n36798 : n54582;
  assign n54584 = pi19 ? n54583 : n33792;
  assign n54585 = pi18 ? n54584 : n53474;
  assign n54586 = pi17 ? n54579 : n54585;
  assign n54587 = pi16 ? n32 : n54586;
  assign n54588 = pi19 ? n46278 : n43198;
  assign n54589 = pi21 ? n43198 : n53471;
  assign n54590 = pi20 ? n54589 : n43198;
  assign n54591 = pi21 ? n43198 : n33792;
  assign n54592 = pi22 ? n33792 : n52875;
  assign n54593 = pi21 ? n33792 : n54592;
  assign n54594 = pi20 ? n54591 : n54593;
  assign n54595 = pi19 ? n54590 : n54594;
  assign n54596 = pi18 ? n54588 : n54595;
  assign n54597 = pi22 ? n33792 : n52873;
  assign n54598 = pi21 ? n54597 : n33792;
  assign n54599 = pi20 ? n43198 : n54598;
  assign n54600 = pi19 ? n54599 : n33792;
  assign n54601 = pi19 ? n53490 : n37641;
  assign n54602 = pi18 ? n54600 : n54601;
  assign n54603 = pi17 ? n54596 : n54602;
  assign n54604 = pi16 ? n32 : n54603;
  assign n54605 = pi15 ? n54587 : n54604;
  assign n54606 = pi14 ? n54571 : n54605;
  assign n54607 = pi21 ? n36659 : n50795;
  assign n54608 = pi20 ? n51354 : n54607;
  assign n54609 = pi19 ? n46278 : n54608;
  assign n54610 = pi21 ? n50795 : n36659;
  assign n54611 = pi20 ? n54610 : n36659;
  assign n54612 = pi19 ? n54611 : n36659;
  assign n54613 = pi18 ? n54609 : n54612;
  assign n54614 = pi17 ? n54613 : n53987;
  assign n54615 = pi16 ? n32 : n54614;
  assign n54616 = pi21 ? n52416 : n36781;
  assign n54617 = pi22 ? n36781 : n49412;
  assign n54618 = pi21 ? n38285 : n54617;
  assign n54619 = pi20 ? n54616 : n54618;
  assign n54620 = pi19 ? n32 : n54619;
  assign n54621 = pi22 ? n37288 : n36781;
  assign n54622 = pi21 ? n54621 : n40002;
  assign n54623 = pi21 ? n36781 : n54621;
  assign n54624 = pi20 ? n54622 : n54623;
  assign n54625 = pi21 ? n53520 : n54621;
  assign n54626 = pi21 ? n37288 : n36781;
  assign n54627 = pi20 ? n54625 : n54626;
  assign n54628 = pi19 ? n54624 : n54627;
  assign n54629 = pi18 ? n54620 : n54628;
  assign n54630 = pi21 ? n36781 : n40002;
  assign n54631 = pi21 ? n36781 : n37288;
  assign n54632 = pi20 ? n54630 : n54631;
  assign n54633 = pi19 ? n54632 : n36781;
  assign n54634 = pi21 ? n53520 : n37288;
  assign n54635 = pi21 ? n36781 : n13481;
  assign n54636 = pi20 ? n54634 : n54635;
  assign n54637 = pi19 ? n54636 : n35482;
  assign n54638 = pi18 ? n54633 : n54637;
  assign n54639 = pi17 ? n54629 : n54638;
  assign n54640 = pi16 ? n32 : n54639;
  assign n54641 = pi15 ? n54615 : n54640;
  assign n54642 = pi22 ? n51366 : n36781;
  assign n54643 = pi21 ? n54642 : n36781;
  assign n54644 = pi21 ? n36781 : n43200;
  assign n54645 = pi20 ? n54643 : n54644;
  assign n54646 = pi19 ? n32 : n54645;
  assign n54647 = pi18 ? n54646 : n36781;
  assign n54648 = pi22 ? n13481 : n54563;
  assign n54649 = pi21 ? n39972 : n54648;
  assign n54650 = pi20 ? n36781 : n54649;
  assign n54651 = pi19 ? n54650 : n32;
  assign n54652 = pi18 ? n36781 : n54651;
  assign n54653 = pi17 ? n54647 : n54652;
  assign n54654 = pi16 ? n32 : n54653;
  assign n54655 = pi21 ? n47396 : n43198;
  assign n54656 = pi20 ? n43198 : n54655;
  assign n54657 = pi19 ? n32 : n54656;
  assign n54658 = pi20 ? n49401 : n36798;
  assign n54659 = pi19 ? n54658 : n36798;
  assign n54660 = pi18 ? n54657 : n54659;
  assign n54661 = pi21 ? n36798 : n47397;
  assign n54662 = pi20 ? n54661 : n36798;
  assign n54663 = pi19 ? n54662 : n36798;
  assign n54664 = pi23 ? n43198 : n685;
  assign n54665 = pi22 ? n54664 : n21502;
  assign n54666 = pi21 ? n43198 : n54665;
  assign n54667 = pi20 ? n36798 : n54666;
  assign n54668 = pi19 ? n54667 : n32;
  assign n54669 = pi18 ? n54663 : n54668;
  assign n54670 = pi17 ? n54660 : n54669;
  assign n54671 = pi16 ? n32 : n54670;
  assign n54672 = pi15 ? n54654 : n54671;
  assign n54673 = pi14 ? n54641 : n54672;
  assign n54674 = pi13 ? n54606 : n54673;
  assign n54675 = pi12 ? n54555 : n54674;
  assign n54676 = pi11 ? n54500 : n54675;
  assign n54677 = pi10 ? n54325 : n54676;
  assign n54678 = pi09 ? n54053 : n54677;
  assign n54679 = pi17 ? n41158 : n54027;
  assign n54680 = pi16 ? n32 : n54679;
  assign n54681 = pi15 ? n32 : n54680;
  assign n54682 = pi17 ? n46447 : n54034;
  assign n54683 = pi16 ? n32 : n54682;
  assign n54684 = pi20 ? n37308 : n38961;
  assign n54685 = pi19 ? n43672 : n54684;
  assign n54686 = pi18 ? n32 : n54685;
  assign n54687 = pi21 ? n31890 : n31200;
  assign n54688 = pi21 ? n30867 : n20563;
  assign n54689 = pi20 ? n54687 : n54688;
  assign n54690 = pi19 ? n54065 : n54689;
  assign n54691 = pi19 ? n53106 : n54043;
  assign n54692 = pi18 ? n54690 : n54691;
  assign n54693 = pi17 ? n54686 : n54692;
  assign n54694 = pi16 ? n32 : n54693;
  assign n54695 = pi15 ? n54683 : n54694;
  assign n54696 = pi14 ? n54681 : n54695;
  assign n54697 = pi13 ? n32 : n54696;
  assign n54698 = pi12 ? n32 : n54697;
  assign n54699 = pi11 ? n32 : n54698;
  assign n54700 = pi10 ? n32 : n54699;
  assign n54701 = pi21 ? n20563 : n31885;
  assign n54702 = pi20 ? n54701 : n38961;
  assign n54703 = pi19 ? n40496 : n54702;
  assign n54704 = pi18 ? n32 : n54703;
  assign n54705 = pi20 ? n30120 : n20563;
  assign n54706 = pi19 ? n32294 : n54705;
  assign n54707 = pi18 ? n54706 : n54061;
  assign n54708 = pi17 ? n54704 : n54707;
  assign n54709 = pi16 ? n32 : n54708;
  assign n54710 = pi21 ? n31294 : n31877;
  assign n54711 = pi20 ? n54710 : n38477;
  assign n54712 = pi19 ? n41681 : n54711;
  assign n54713 = pi18 ? n32 : n54712;
  assign n54714 = pi20 ? n52962 : n31266;
  assign n54715 = pi20 ? n37439 : n31266;
  assign n54716 = pi19 ? n54714 : n54715;
  assign n54717 = pi18 ? n54716 : n54075;
  assign n54718 = pi17 ? n54713 : n54717;
  assign n54719 = pi16 ? n32 : n54718;
  assign n54720 = pi15 ? n54709 : n54719;
  assign n54721 = pi21 ? n36249 : n31200;
  assign n54722 = pi20 ? n54721 : n37;
  assign n54723 = pi19 ? n54722 : n26630;
  assign n54724 = pi18 ? n34258 : n54723;
  assign n54725 = pi17 ? n39374 : n54724;
  assign n54726 = pi16 ? n32 : n54725;
  assign n54727 = pi17 ? n40533 : n54091;
  assign n54728 = pi16 ? n32 : n54727;
  assign n54729 = pi15 ? n54726 : n54728;
  assign n54730 = pi14 ? n54720 : n54729;
  assign n54731 = pi20 ? n37 : n23828;
  assign n54732 = pi19 ? n31267 : n54731;
  assign n54733 = pi18 ? n20563 : n54732;
  assign n54734 = pi17 ? n40046 : n54733;
  assign n54735 = pi16 ? n32 : n54734;
  assign n54736 = pi20 ? n38376 : n31925;
  assign n54737 = pi24 ? n20563 : n37;
  assign n54738 = pi23 ? n54737 : n37;
  assign n54739 = pi22 ? n20563 : n54738;
  assign n54740 = pi21 ? n20563 : n54739;
  assign n54741 = pi20 ? n54740 : n20563;
  assign n54742 = pi19 ? n54736 : n54741;
  assign n54743 = pi18 ? n32 : n54742;
  assign n54744 = pi20 ? n47432 : n30096;
  assign n54745 = pi19 ? n54744 : n51465;
  assign n54746 = pi21 ? n11199 : n2678;
  assign n54747 = pi20 ? n37 : n54746;
  assign n54748 = pi19 ? n31280 : n54747;
  assign n54749 = pi18 ? n54745 : n54748;
  assign n54750 = pi17 ? n54743 : n54749;
  assign n54751 = pi16 ? n32 : n54750;
  assign n54752 = pi15 ? n54735 : n54751;
  assign n54753 = pi20 ? n39395 : n31913;
  assign n54754 = pi19 ? n54753 : n20563;
  assign n54755 = pi18 ? n32 : n54754;
  assign n54756 = pi19 ? n37 : n54747;
  assign n54757 = pi18 ? n53013 : n54756;
  assign n54758 = pi17 ? n54755 : n54757;
  assign n54759 = pi16 ? n32 : n54758;
  assign n54760 = pi20 ? n28157 : n36929;
  assign n54761 = pi20 ? n46815 : n38477;
  assign n54762 = pi19 ? n54760 : n54761;
  assign n54763 = pi18 ? n32 : n54762;
  assign n54764 = pi20 ? n54070 : n37;
  assign n54765 = pi19 ? n50854 : n54764;
  assign n54766 = pi20 ? n37 : n23859;
  assign n54767 = pi19 ? n37 : n54766;
  assign n54768 = pi18 ? n54765 : n54767;
  assign n54769 = pi17 ? n54763 : n54768;
  assign n54770 = pi16 ? n32 : n54769;
  assign n54771 = pi15 ? n54759 : n54770;
  assign n54772 = pi14 ? n54752 : n54771;
  assign n54773 = pi13 ? n54730 : n54772;
  assign n54774 = pi20 ? n35316 : n20563;
  assign n54775 = pi19 ? n54774 : n31926;
  assign n54776 = pi21 ? n54132 : n2700;
  assign n54777 = pi20 ? n37 : n54776;
  assign n54778 = pi19 ? n37 : n54777;
  assign n54779 = pi18 ? n54775 : n54778;
  assign n54780 = pi17 ? n45393 : n54779;
  assign n54781 = pi16 ? n32 : n54780;
  assign n54782 = pi20 ? n20563 : n54070;
  assign n54783 = pi19 ? n20563 : n54782;
  assign n54784 = pi21 ? n54140 : n1009;
  assign n54785 = pi20 ? n30096 : n54784;
  assign n54786 = pi19 ? n54139 : n54785;
  assign n54787 = pi18 ? n54783 : n54786;
  assign n54788 = pi17 ? n37929 : n54787;
  assign n54789 = pi16 ? n32 : n54788;
  assign n54790 = pi15 ? n54781 : n54789;
  assign n54791 = pi20 ? n30096 : n24844;
  assign n54792 = pi19 ? n51953 : n54791;
  assign n54793 = pi18 ? n20563 : n54792;
  assign n54794 = pi17 ? n37958 : n54793;
  assign n54795 = pi16 ? n32 : n54794;
  assign n54796 = pi20 ? n31266 : n49916;
  assign n54797 = pi20 ? n31266 : n52962;
  assign n54798 = pi19 ? n54796 : n54797;
  assign n54799 = pi22 ? n37 : n7780;
  assign n54800 = pi21 ? n54799 : n32;
  assign n54801 = pi20 ? n30096 : n54800;
  assign n54802 = pi19 ? n54139 : n54801;
  assign n54803 = pi18 ? n54798 : n54802;
  assign n54804 = pi17 ? n37958 : n54803;
  assign n54805 = pi16 ? n32 : n54804;
  assign n54806 = pi15 ? n54795 : n54805;
  assign n54807 = pi14 ? n54790 : n54806;
  assign n54808 = pi18 ? n38999 : n54171;
  assign n54809 = pi20 ? n37 : n54800;
  assign n54810 = pi19 ? n37 : n54809;
  assign n54811 = pi18 ? n54131 : n54810;
  assign n54812 = pi17 ? n54808 : n54811;
  assign n54813 = pi16 ? n32 : n54812;
  assign n54814 = pi20 ? n31205 : n52962;
  assign n54815 = pi19 ? n54814 : n32871;
  assign n54816 = pi18 ? n54815 : n54186;
  assign n54817 = pi17 ? n37336 : n54816;
  assign n54818 = pi16 ? n32 : n54817;
  assign n54819 = pi15 ? n54813 : n54818;
  assign n54820 = pi21 ? n37 : n31200;
  assign n54821 = pi20 ? n20563 : n54820;
  assign n54822 = pi19 ? n20563 : n54821;
  assign n54823 = pi20 ? n37 : n49441;
  assign n54824 = pi20 ? n31903 : n54184;
  assign n54825 = pi19 ? n54823 : n54824;
  assign n54826 = pi18 ? n54822 : n54825;
  assign n54827 = pi17 ? n37336 : n54826;
  assign n54828 = pi16 ? n32 : n54827;
  assign n54829 = pi20 ? n31903 : n11215;
  assign n54830 = pi19 ? n51953 : n54829;
  assign n54831 = pi18 ? n34258 : n54830;
  assign n54832 = pi17 ? n36162 : n54831;
  assign n54833 = pi16 ? n32 : n54832;
  assign n54834 = pi15 ? n54828 : n54833;
  assign n54835 = pi14 ? n54819 : n54834;
  assign n54836 = pi13 ? n54807 : n54835;
  assign n54837 = pi12 ? n54773 : n54836;
  assign n54838 = pi17 ? n36162 : n54207;
  assign n54839 = pi16 ? n32 : n54838;
  assign n54840 = pi19 ? n51932 : n20563;
  assign n54841 = pi18 ? n28159 : n54840;
  assign n54842 = pi20 ? n30096 : n54040;
  assign n54843 = pi20 ? n33821 : n31220;
  assign n54844 = pi19 ? n54842 : n54843;
  assign n54845 = pi20 ? n37 : n54820;
  assign n54846 = pi19 ? n54845 : n54216;
  assign n54847 = pi18 ? n54844 : n54846;
  assign n54848 = pi17 ? n54841 : n54847;
  assign n54849 = pi16 ? n32 : n54848;
  assign n54850 = pi15 ? n54839 : n54849;
  assign n54851 = pi18 ? n30119 : n54222;
  assign n54852 = pi19 ? n53051 : n30097;
  assign n54853 = pi18 ? n54852 : n54228;
  assign n54854 = pi17 ? n54851 : n54853;
  assign n54855 = pi16 ? n32 : n54854;
  assign n54856 = pi17 ? n35194 : n54238;
  assign n54857 = pi16 ? n32 : n54856;
  assign n54858 = pi15 ? n54855 : n54857;
  assign n54859 = pi14 ? n54850 : n54858;
  assign n54860 = pi20 ? n24493 : n40749;
  assign n54861 = pi19 ? n54243 : n54860;
  assign n54862 = pi18 ? n34869 : n54861;
  assign n54863 = pi17 ? n35764 : n54862;
  assign n54864 = pi16 ? n32 : n54863;
  assign n54865 = pi20 ? n5077 : n6935;
  assign n54866 = pi19 ? n53104 : n54865;
  assign n54867 = pi18 ? n34869 : n54866;
  assign n54868 = pi17 ? n35764 : n54867;
  assign n54869 = pi16 ? n32 : n54868;
  assign n54870 = pi15 ? n54864 : n54869;
  assign n54871 = pi20 ? n24493 : n6935;
  assign n54872 = pi19 ? n53104 : n54871;
  assign n54873 = pi18 ? n20563 : n54872;
  assign n54874 = pi17 ? n50386 : n54873;
  assign n54875 = pi16 ? n32 : n54874;
  assign n54876 = pi20 ? n31220 : n54155;
  assign n54877 = pi19 ? n54876 : n53104;
  assign n54878 = pi20 ? n53138 : n6935;
  assign n54879 = pi19 ? n54265 : n54878;
  assign n54880 = pi18 ? n54877 : n54879;
  assign n54881 = pi17 ? n50386 : n54880;
  assign n54882 = pi16 ? n32 : n54881;
  assign n54883 = pi15 ? n54875 : n54882;
  assign n54884 = pi14 ? n54870 : n54883;
  assign n54885 = pi13 ? n54859 : n54884;
  assign n54886 = pi17 ? n50390 : n54278;
  assign n54887 = pi16 ? n32 : n54886;
  assign n54888 = pi17 ? n50393 : n54284;
  assign n54889 = pi16 ? n32 : n54888;
  assign n54890 = pi15 ? n54887 : n54889;
  assign n54891 = pi20 ? n1665 : n24937;
  assign n54892 = pi19 ? n53344 : n54891;
  assign n54893 = pi18 ? n20563 : n54892;
  assign n54894 = pi17 ? n50393 : n54893;
  assign n54895 = pi16 ? n32 : n54894;
  assign n54896 = pi19 ? n32294 : n22942;
  assign n54897 = pi18 ? n20563 : n54896;
  assign n54898 = pi17 ? n50393 : n54897;
  assign n54899 = pi16 ? n32 : n54898;
  assign n54900 = pi15 ? n54895 : n54899;
  assign n54901 = pi14 ? n54890 : n54900;
  assign n54902 = pi20 ? n14927 : n3176;
  assign n54903 = pi19 ? n32294 : n54902;
  assign n54904 = pi18 ? n20563 : n54903;
  assign n54905 = pi17 ? n50393 : n54904;
  assign n54906 = pi16 ? n32 : n54905;
  assign n54907 = pi19 ? n51069 : n54902;
  assign n54908 = pi18 ? n20563 : n54907;
  assign n54909 = pi17 ? n50905 : n54908;
  assign n54910 = pi16 ? n32 : n54909;
  assign n54911 = pi15 ? n54906 : n54910;
  assign n54912 = pi18 ? n43247 : n20563;
  assign n54913 = pi20 ? n21732 : n3176;
  assign n54914 = pi19 ? n32294 : n54913;
  assign n54915 = pi18 ? n20563 : n54914;
  assign n54916 = pi17 ? n54912 : n54915;
  assign n54917 = pi16 ? n32 : n54916;
  assign n54918 = pi20 ? n54315 : n4110;
  assign n54919 = pi19 ? n32294 : n54918;
  assign n54920 = pi18 ? n20563 : n54919;
  assign n54921 = pi17 ? n54912 : n54920;
  assign n54922 = pi16 ? n32 : n54921;
  assign n54923 = pi15 ? n54917 : n54922;
  assign n54924 = pi14 ? n54911 : n54923;
  assign n54925 = pi13 ? n54901 : n54924;
  assign n54926 = pi12 ? n54885 : n54925;
  assign n54927 = pi11 ? n54837 : n54926;
  assign n54928 = pi20 ? n54326 : n3210;
  assign n54929 = pi19 ? n32294 : n54928;
  assign n54930 = pi18 ? n20563 : n54929;
  assign n54931 = pi17 ? n54912 : n54930;
  assign n54932 = pi16 ? n32 : n54931;
  assign n54933 = pi20 ? n51634 : n4116;
  assign n54934 = pi19 ? n32294 : n54933;
  assign n54935 = pi18 ? n20563 : n54934;
  assign n54936 = pi17 ? n54912 : n54935;
  assign n54937 = pi16 ? n32 : n54936;
  assign n54938 = pi15 ? n54932 : n54937;
  assign n54939 = pi23 ? n20627 : n363;
  assign n54940 = pi22 ? n54939 : n2299;
  assign n54941 = pi21 ? n139 : n54940;
  assign n54942 = pi20 ? n54941 : n10011;
  assign n54943 = pi19 ? n32294 : n54942;
  assign n54944 = pi18 ? n20563 : n54943;
  assign n54945 = pi17 ? n54912 : n54944;
  assign n54946 = pi16 ? n32 : n54945;
  assign n54947 = pi20 ? n54346 : n10011;
  assign n54948 = pi19 ? n31221 : n54947;
  assign n54949 = pi18 ? n20563 : n54948;
  assign n54950 = pi17 ? n49448 : n54949;
  assign n54951 = pi16 ? n32 : n54950;
  assign n54952 = pi15 ? n54946 : n54951;
  assign n54953 = pi14 ? n54938 : n54952;
  assign n54954 = pi24 ? n99 : n33792;
  assign n54955 = pi23 ? n54954 : n157;
  assign n54956 = pi22 ? n54955 : n233;
  assign n54957 = pi21 ? n37 : n54956;
  assign n54958 = pi20 ? n54957 : n32;
  assign n54959 = pi19 ? n54355 : n54958;
  assign n54960 = pi18 ? n20563 : n54959;
  assign n54961 = pi17 ? n49448 : n54960;
  assign n54962 = pi16 ? n32 : n54961;
  assign n54963 = pi17 ? n49448 : n54369;
  assign n54964 = pi16 ? n32 : n54963;
  assign n54965 = pi15 ? n54962 : n54964;
  assign n54966 = pi17 ? n49448 : n54378;
  assign n54967 = pi16 ? n32 : n54966;
  assign n54968 = pi22 ? n35902 : n3338;
  assign n54969 = pi21 ? n335 : n54968;
  assign n54970 = pi20 ? n54969 : n32;
  assign n54971 = pi19 ? n32294 : n54970;
  assign n54972 = pi18 ? n20563 : n54971;
  assign n54973 = pi17 ? n49448 : n54972;
  assign n54974 = pi16 ? n32 : n54973;
  assign n54975 = pi15 ? n54967 : n54974;
  assign n54976 = pi14 ? n54965 : n54975;
  assign n54977 = pi13 ? n54953 : n54976;
  assign n54978 = pi18 ? n43254 : n20563;
  assign n54979 = pi22 ? n15294 : n2192;
  assign n54980 = pi21 ? n335 : n54979;
  assign n54981 = pi20 ? n54980 : n32;
  assign n54982 = pi19 ? n54393 : n54981;
  assign n54983 = pi18 ? n20563 : n54982;
  assign n54984 = pi17 ? n54978 : n54983;
  assign n54985 = pi16 ? n32 : n54984;
  assign n54986 = pi22 ? n18448 : n1407;
  assign n54987 = pi21 ? n363 : n54986;
  assign n54988 = pi20 ? n54987 : n32;
  assign n54989 = pi19 ? n32294 : n54988;
  assign n54990 = pi18 ? n20563 : n54989;
  assign n54991 = pi17 ? n54978 : n54990;
  assign n54992 = pi16 ? n32 : n54991;
  assign n54993 = pi15 ? n54985 : n54992;
  assign n54994 = pi21 ? n46187 : n40913;
  assign n54995 = pi20 ? n54994 : n40791;
  assign n54996 = pi19 ? n32 : n54995;
  assign n54997 = pi18 ? n54996 : n54419;
  assign n54998 = pi21 ? n20563 : n45049;
  assign n54999 = pi20 ? n54998 : n20563;
  assign n55000 = pi19 ? n54999 : n20563;
  assign n55001 = pi18 ? n55000 : n54423;
  assign n55002 = pi17 ? n54997 : n55001;
  assign n55003 = pi16 ? n32 : n55002;
  assign n55004 = pi19 ? n32 : n46715;
  assign n55005 = pi18 ? n55004 : n54432;
  assign n55006 = pi17 ? n55005 : n54439;
  assign n55007 = pi16 ? n32 : n55006;
  assign n55008 = pi15 ? n55003 : n55007;
  assign n55009 = pi14 ? n54993 : n55008;
  assign n55010 = pi21 ? n52742 : n40955;
  assign n55011 = pi20 ? n55010 : n53307;
  assign n55012 = pi19 ? n32 : n55011;
  assign n55013 = pi18 ? n55012 : n54452;
  assign n55014 = pi21 ? n20563 : n40954;
  assign n55015 = pi20 ? n55014 : n20563;
  assign n55016 = pi19 ? n55015 : n20563;
  assign n55017 = pi18 ? n55016 : n54456;
  assign n55018 = pi17 ? n55013 : n55017;
  assign n55019 = pi16 ? n32 : n55018;
  assign n55020 = pi21 ? n20563 : n41489;
  assign n55021 = pi20 ? n55020 : n40961;
  assign n55022 = pi19 ? n38982 : n55021;
  assign n55023 = pi21 ? n40957 : n37768;
  assign n55024 = pi21 ? n40954 : n40957;
  assign n55025 = pi20 ? n55023 : n55024;
  assign n55026 = pi21 ? n33792 : n37768;
  assign n55027 = pi20 ? n54468 : n55026;
  assign n55028 = pi19 ? n55025 : n55027;
  assign n55029 = pi18 ? n55022 : n55028;
  assign n55030 = pi21 ? n40954 : n37768;
  assign n55031 = pi20 ? n55030 : n53326;
  assign n55032 = pi19 ? n55031 : n20563;
  assign n55033 = pi18 ? n55032 : n54479;
  assign n55034 = pi17 ? n55029 : n55033;
  assign n55035 = pi16 ? n32 : n55034;
  assign n55036 = pi15 ? n55019 : n55035;
  assign n55037 = pi17 ? n48912 : n54487;
  assign n55038 = pi16 ? n32 : n55037;
  assign n55039 = pi23 ? n54954 : n363;
  assign n55040 = pi22 ? n55039 : n204;
  assign n55041 = pi21 ? n55040 : n882;
  assign n55042 = pi20 ? n55041 : n32;
  assign n55043 = pi19 ? n53344 : n55042;
  assign n55044 = pi18 ? n20563 : n55043;
  assign n55045 = pi17 ? n48912 : n55044;
  assign n55046 = pi16 ? n32 : n55045;
  assign n55047 = pi15 ? n55038 : n55046;
  assign n55048 = pi14 ? n55036 : n55047;
  assign n55049 = pi13 ? n55009 : n55048;
  assign n55050 = pi12 ? n54977 : n55049;
  assign n55051 = pi17 ? n48904 : n54504;
  assign n55052 = pi16 ? n32 : n55051;
  assign n55053 = pi24 ? n33792 : n363;
  assign n55054 = pi23 ? n55053 : n157;
  assign n55055 = pi22 ? n55054 : n685;
  assign n55056 = pi21 ? n55055 : n53983;
  assign n55057 = pi20 ? n55056 : n32;
  assign n55058 = pi19 ? n53368 : n55057;
  assign n55059 = pi18 ? n20563 : n55058;
  assign n55060 = pi17 ? n48904 : n55059;
  assign n55061 = pi16 ? n32 : n55060;
  assign n55062 = pi15 ? n55052 : n55061;
  assign n55063 = pi17 ? n53727 : n53382;
  assign n55064 = pi16 ? n32 : n55063;
  assign n55065 = pi17 ? n53727 : n53390;
  assign n55066 = pi16 ? n32 : n55065;
  assign n55067 = pi15 ? n55064 : n55066;
  assign n55068 = pi14 ? n55062 : n55067;
  assign n55069 = pi17 ? n53727 : n53402;
  assign n55070 = pi16 ? n32 : n55069;
  assign n55071 = pi18 ? n49219 : n43012;
  assign n55072 = pi17 ? n55071 : n54533;
  assign n55073 = pi16 ? n32 : n55072;
  assign n55074 = pi15 ? n55070 : n55073;
  assign n55075 = pi20 ? n37806 : n42005;
  assign n55076 = pi19 ? n32 : n55075;
  assign n55077 = pi18 ? n55076 : n54539;
  assign n55078 = pi17 ? n55077 : n53425;
  assign n55079 = pi16 ? n32 : n55078;
  assign n55080 = pi21 ? n51232 : n20563;
  assign n55081 = pi20 ? n55080 : n20563;
  assign n55082 = pi19 ? n32 : n55081;
  assign n55083 = pi18 ? n55082 : n20563;
  assign n55084 = pi17 ? n55083 : n53436;
  assign n55085 = pi16 ? n32 : n55084;
  assign n55086 = pi15 ? n55079 : n55085;
  assign n55087 = pi14 ? n55074 : n55086;
  assign n55088 = pi13 ? n55068 : n55087;
  assign n55089 = pi19 ? n32 : n46700;
  assign n55090 = pi18 ? n55089 : n30868;
  assign n55091 = pi17 ? n55090 : n53447;
  assign n55092 = pi16 ? n32 : n55091;
  assign n55093 = pi17 ? n55090 : n54568;
  assign n55094 = pi16 ? n32 : n55093;
  assign n55095 = pi15 ? n55092 : n55094;
  assign n55096 = pi20 ? n50768 : n36798;
  assign n55097 = pi19 ? n32 : n55096;
  assign n55098 = pi22 ? n54580 : n33792;
  assign n55099 = pi21 ? n36798 : n55098;
  assign n55100 = pi21 ? n53463 : n45142;
  assign n55101 = pi20 ? n55099 : n55100;
  assign n55102 = pi19 ? n36798 : n55101;
  assign n55103 = pi18 ? n55097 : n55102;
  assign n55104 = pi20 ? n36798 : n54581;
  assign n55105 = pi19 ? n55104 : n33792;
  assign n55106 = pi18 ? n55105 : n53474;
  assign n55107 = pi17 ? n55103 : n55106;
  assign n55108 = pi16 ? n32 : n55107;
  assign n55109 = pi20 ? n50787 : n43198;
  assign n55110 = pi19 ? n32 : n55109;
  assign n55111 = pi20 ? n53481 : n33792;
  assign n55112 = pi19 ? n54590 : n55111;
  assign n55113 = pi18 ? n55110 : n55112;
  assign n55114 = pi20 ? n43198 : n54597;
  assign n55115 = pi19 ? n55114 : n33792;
  assign n55116 = pi18 ? n55115 : n54601;
  assign n55117 = pi17 ? n55113 : n55116;
  assign n55118 = pi16 ? n32 : n55117;
  assign n55119 = pi15 ? n55108 : n55118;
  assign n55120 = pi14 ? n55095 : n55119;
  assign n55121 = pi21 ? n50786 : n53977;
  assign n55122 = pi21 ? n50796 : n50795;
  assign n55123 = pi20 ? n55121 : n55122;
  assign n55124 = pi19 ? n32 : n55123;
  assign n55125 = pi22 ? n50339 : n43198;
  assign n55126 = pi21 ? n55125 : n36659;
  assign n55127 = pi20 ? n55126 : n36659;
  assign n55128 = pi19 ? n55127 : n36659;
  assign n55129 = pi18 ? n55124 : n55128;
  assign n55130 = pi23 ? n36659 : n363;
  assign n55131 = pi22 ? n36659 : n55130;
  assign n55132 = pi21 ? n55131 : n13481;
  assign n55133 = pi20 ? n36659 : n55132;
  assign n55134 = pi19 ? n55133 : n1823;
  assign n55135 = pi18 ? n36659 : n55134;
  assign n55136 = pi17 ? n55129 : n55135;
  assign n55137 = pi16 ? n32 : n55136;
  assign n55138 = pi21 ? n46790 : n36781;
  assign n55139 = pi21 ? n36781 : n54617;
  assign n55140 = pi20 ? n55138 : n55139;
  assign n55141 = pi19 ? n32 : n55140;
  assign n55142 = pi18 ? n55141 : n36781;
  assign n55143 = pi22 ? n36781 : n51895;
  assign n55144 = pi21 ? n55143 : n51895;
  assign n55145 = pi20 ? n55144 : n54635;
  assign n55146 = pi19 ? n55145 : n35482;
  assign n55147 = pi18 ? n36781 : n55146;
  assign n55148 = pi17 ? n55142 : n55147;
  assign n55149 = pi16 ? n32 : n55148;
  assign n55150 = pi15 ? n55137 : n55149;
  assign n55151 = pi21 ? n46276 : n36781;
  assign n55152 = pi20 ? n55151 : n54644;
  assign n55153 = pi19 ? n32 : n55152;
  assign n55154 = pi18 ? n55153 : n36781;
  assign n55155 = pi17 ? n55154 : n54652;
  assign n55156 = pi16 ? n32 : n55155;
  assign n55157 = pi20 ? n46791 : n54655;
  assign n55158 = pi19 ? n32 : n55157;
  assign n55159 = pi18 ? n55158 : n54659;
  assign n55160 = pi17 ? n55159 : n54669;
  assign n55161 = pi16 ? n32 : n55160;
  assign n55162 = pi15 ? n55156 : n55161;
  assign n55163 = pi14 ? n55150 : n55162;
  assign n55164 = pi13 ? n55120 : n55163;
  assign n55165 = pi12 ? n55088 : n55164;
  assign n55166 = pi11 ? n55050 : n55165;
  assign n55167 = pi10 ? n54927 : n55166;
  assign n55168 = pi09 ? n54700 : n55167;
  assign n55169 = pi08 ? n54678 : n55168;
  assign n55170 = pi07 ? n54022 : n55169;
  assign n55171 = pi06 ? n52935 : n55170;
  assign n55172 = pi05 ? n50853 : n55171;
  assign n55173 = pi04 ? n46814 : n55172;
  assign n55174 = pi03 ? n38314 : n55173;
  assign n55175 = pi02 ? n22600 : n55174;
  assign n55176 = pi01 ? n32 : n55175;
  assign n55177 = pi21 ? n297 : n3022;
  assign n55178 = pi20 ? n37 : n55177;
  assign n55179 = pi19 ? n20563 : n55178;
  assign n55180 = pi18 ? n20563 : n55179;
  assign n55181 = pi17 ? n41169 : n55180;
  assign n55182 = pi16 ? n32 : n55181;
  assign n55183 = pi15 ? n32 : n55182;
  assign n55184 = pi20 ? n31220 : n10158;
  assign n55185 = pi19 ? n20563 : n55184;
  assign n55186 = pi18 ? n20563 : n55185;
  assign n55187 = pi17 ? n41169 : n55186;
  assign n55188 = pi16 ? n32 : n55187;
  assign n55189 = pi17 ? n40024 : n55186;
  assign n55190 = pi16 ? n32 : n55189;
  assign n55191 = pi15 ? n55188 : n55190;
  assign n55192 = pi14 ? n55183 : n55191;
  assign n55193 = pi13 ? n32 : n55192;
  assign n55194 = pi12 ? n32 : n55193;
  assign n55195 = pi11 ? n32 : n55194;
  assign n55196 = pi10 ? n32 : n55195;
  assign n55197 = pi21 ? n297 : n9238;
  assign n55198 = pi20 ? n20563 : n55197;
  assign n55199 = pi19 ? n20563 : n55198;
  assign n55200 = pi18 ? n20563 : n55199;
  assign n55201 = pi17 ? n41182 : n55200;
  assign n55202 = pi16 ? n32 : n55201;
  assign n55203 = pi21 ? n297 : n9246;
  assign n55204 = pi20 ? n31220 : n55203;
  assign n55205 = pi19 ? n20563 : n55204;
  assign n55206 = pi18 ? n20563 : n55205;
  assign n55207 = pi17 ? n46447 : n55206;
  assign n55208 = pi16 ? n32 : n55207;
  assign n55209 = pi15 ? n55202 : n55208;
  assign n55210 = pi21 ? n569 : n2565;
  assign n55211 = pi20 ? n31220 : n55210;
  assign n55212 = pi19 ? n20563 : n55211;
  assign n55213 = pi18 ? n20563 : n55212;
  assign n55214 = pi17 ? n40498 : n55213;
  assign n55215 = pi16 ? n32 : n55214;
  assign n55216 = pi21 ? n569 : n2469;
  assign n55217 = pi20 ? n31220 : n55216;
  assign n55218 = pi19 ? n20563 : n55217;
  assign n55219 = pi18 ? n20563 : n55218;
  assign n55220 = pi17 ? n40533 : n55219;
  assign n55221 = pi16 ? n32 : n55220;
  assign n55222 = pi15 ? n55215 : n55221;
  assign n55223 = pi14 ? n55209 : n55222;
  assign n55224 = pi21 ? n335 : n2553;
  assign n55225 = pi20 ? n31220 : n55224;
  assign n55226 = pi19 ? n20563 : n55225;
  assign n55227 = pi18 ? n20563 : n55226;
  assign n55228 = pi17 ? n40533 : n55227;
  assign n55229 = pi16 ? n32 : n55228;
  assign n55230 = pi20 ? n31220 : n38437;
  assign n55231 = pi19 ? n20563 : n55230;
  assign n55232 = pi18 ? n20563 : n55231;
  assign n55233 = pi17 ? n41709 : n55232;
  assign n55234 = pi16 ? n32 : n55233;
  assign n55235 = pi15 ? n55229 : n55234;
  assign n55236 = pi21 ? n569 : n2678;
  assign n55237 = pi20 ? n31220 : n55236;
  assign n55238 = pi19 ? n20563 : n55237;
  assign n55239 = pi18 ? n20563 : n55238;
  assign n55240 = pi17 ? n45367 : n55239;
  assign n55241 = pi16 ? n32 : n55240;
  assign n55242 = pi21 ? n569 : n2700;
  assign n55243 = pi20 ? n31220 : n55242;
  assign n55244 = pi19 ? n20563 : n55243;
  assign n55245 = pi18 ? n20563 : n55244;
  assign n55246 = pi17 ? n38949 : n55245;
  assign n55247 = pi16 ? n32 : n55246;
  assign n55248 = pi15 ? n55241 : n55247;
  assign n55249 = pi14 ? n55235 : n55248;
  assign n55250 = pi13 ? n55223 : n55249;
  assign n55251 = pi17 ? n40046 : n55245;
  assign n55252 = pi16 ? n32 : n55251;
  assign n55253 = pi20 ? n31220 : n25766;
  assign n55254 = pi19 ? n20563 : n55253;
  assign n55255 = pi18 ? n20563 : n55254;
  assign n55256 = pi17 ? n40046 : n55255;
  assign n55257 = pi16 ? n32 : n55256;
  assign n55258 = pi15 ? n55252 : n55257;
  assign n55259 = pi17 ? n37929 : n55255;
  assign n55260 = pi16 ? n32 : n55259;
  assign n55261 = pi20 ? n31220 : n11665;
  assign n55262 = pi19 ? n20563 : n55261;
  assign n55263 = pi18 ? n20563 : n55262;
  assign n55264 = pi17 ? n38984 : n55263;
  assign n55265 = pi16 ? n32 : n55264;
  assign n55266 = pi15 ? n55260 : n55265;
  assign n55267 = pi14 ? n55258 : n55266;
  assign n55268 = pi20 ? n31220 : n11215;
  assign n55269 = pi19 ? n20563 : n55268;
  assign n55270 = pi18 ? n20563 : n55269;
  assign n55271 = pi17 ? n40057 : n55270;
  assign n55272 = pi16 ? n32 : n55271;
  assign n55273 = pi20 ? n31220 : n12486;
  assign n55274 = pi19 ? n20563 : n55273;
  assign n55275 = pi18 ? n20563 : n55274;
  assign n55276 = pi17 ? n37936 : n55275;
  assign n55277 = pi16 ? n32 : n55276;
  assign n55278 = pi15 ? n55272 : n55277;
  assign n55279 = pi20 ? n31220 : n12101;
  assign n55280 = pi19 ? n20563 : n55279;
  assign n55281 = pi18 ? n20563 : n55280;
  assign n55282 = pi17 ? n37958 : n55281;
  assign n55283 = pi16 ? n32 : n55282;
  assign n55284 = pi14 ? n55278 : n55283;
  assign n55285 = pi13 ? n55267 : n55284;
  assign n55286 = pi12 ? n55250 : n55285;
  assign n55287 = pi20 ? n31220 : n24844;
  assign n55288 = pi19 ? n20563 : n55287;
  assign n55289 = pi18 ? n20563 : n55288;
  assign n55290 = pi17 ? n37958 : n55289;
  assign n55291 = pi16 ? n32 : n55290;
  assign n55292 = pi20 ? n37 : n48905;
  assign n55293 = pi21 ? n20563 : n3392;
  assign n55294 = pi20 ? n55293 : n24850;
  assign n55295 = pi19 ? n55292 : n55294;
  assign n55296 = pi18 ? n20563 : n55295;
  assign n55297 = pi17 ? n39000 : n55296;
  assign n55298 = pi16 ? n32 : n55297;
  assign n55299 = pi15 ? n55291 : n55298;
  assign n55300 = pi21 ? n29319 : n32;
  assign n55301 = pi20 ? n31220 : n55300;
  assign n55302 = pi19 ? n54170 : n55301;
  assign n55303 = pi18 ? n20563 : n55302;
  assign n55304 = pi17 ? n37323 : n55303;
  assign n55305 = pi16 ? n32 : n55304;
  assign n55306 = pi22 ? n37 : n1388;
  assign n55307 = pi21 ? n55306 : n32;
  assign n55308 = pi20 ? n31220 : n55307;
  assign n55309 = pi19 ? n20563 : n55308;
  assign n55310 = pi18 ? n20563 : n55309;
  assign n55311 = pi17 ? n37323 : n55310;
  assign n55312 = pi16 ? n32 : n55311;
  assign n55313 = pi15 ? n55305 : n55312;
  assign n55314 = pi14 ? n55299 : n55313;
  assign n55315 = pi22 ? n157 : n6415;
  assign n55316 = pi21 ? n55315 : n32;
  assign n55317 = pi20 ? n31220 : n55316;
  assign n55318 = pi19 ? n20563 : n55317;
  assign n55319 = pi18 ? n20563 : n55318;
  assign n55320 = pi17 ? n39456 : n55319;
  assign n55321 = pi16 ? n32 : n55320;
  assign n55322 = pi20 ? n31220 : n39589;
  assign n55323 = pi19 ? n20563 : n55322;
  assign n55324 = pi18 ? n20563 : n55323;
  assign n55325 = pi17 ? n39456 : n55324;
  assign n55326 = pi16 ? n32 : n55325;
  assign n55327 = pi15 ? n55321 : n55326;
  assign n55328 = pi20 ? n31220 : n6935;
  assign n55329 = pi19 ? n53012 : n55328;
  assign n55330 = pi18 ? n20563 : n55329;
  assign n55331 = pi17 ? n39456 : n55330;
  assign n55332 = pi16 ? n32 : n55331;
  assign n55333 = pi22 ? n37 : n19177;
  assign n55334 = pi21 ? n36249 : n55333;
  assign n55335 = pi20 ? n55334 : n6935;
  assign n55336 = pi19 ? n55292 : n55335;
  assign n55337 = pi18 ? n38951 : n55336;
  assign n55338 = pi17 ? n36162 : n55337;
  assign n55339 = pi16 ? n32 : n55338;
  assign n55340 = pi15 ? n55332 : n55339;
  assign n55341 = pi14 ? n55327 : n55340;
  assign n55342 = pi13 ? n55314 : n55341;
  assign n55343 = pi21 ? n20563 : n6433;
  assign n55344 = pi20 ? n55343 : n5667;
  assign n55345 = pi19 ? n53104 : n55344;
  assign n55346 = pi18 ? n20563 : n55345;
  assign n55347 = pi17 ? n34859 : n55346;
  assign n55348 = pi16 ? n32 : n55347;
  assign n55349 = pi21 ? n20563 : n55333;
  assign n55350 = pi20 ? n55349 : n26293;
  assign n55351 = pi19 ? n20563 : n55350;
  assign n55352 = pi18 ? n20563 : n55351;
  assign n55353 = pi17 ? n34859 : n55352;
  assign n55354 = pi16 ? n32 : n55353;
  assign n55355 = pi15 ? n55348 : n55354;
  assign n55356 = pi20 ? n55349 : n12149;
  assign n55357 = pi19 ? n20563 : n55356;
  assign n55358 = pi18 ? n20563 : n55357;
  assign n55359 = pi17 ? n34859 : n55358;
  assign n55360 = pi16 ? n32 : n55359;
  assign n55361 = pi18 ? n43673 : n20563;
  assign n55362 = pi21 ? n29133 : n4451;
  assign n55363 = pi20 ? n55362 : n4008;
  assign n55364 = pi19 ? n20563 : n55363;
  assign n55365 = pi18 ? n20563 : n55364;
  assign n55366 = pi17 ? n55361 : n55365;
  assign n55367 = pi16 ? n32 : n55366;
  assign n55368 = pi15 ? n55360 : n55367;
  assign n55369 = pi14 ? n55355 : n55368;
  assign n55370 = pi21 ? n29133 : n6706;
  assign n55371 = pi20 ? n55370 : n7035;
  assign n55372 = pi19 ? n20563 : n55371;
  assign n55373 = pi18 ? n20563 : n55372;
  assign n55374 = pi17 ? n55361 : n55373;
  assign n55375 = pi16 ? n32 : n55374;
  assign n55376 = pi21 ? n30843 : n30195;
  assign n55377 = pi20 ? n55376 : n52962;
  assign n55378 = pi21 ? n31294 : n36249;
  assign n55379 = pi20 ? n55378 : n37;
  assign n55380 = pi19 ? n55377 : n55379;
  assign n55381 = pi21 ? n36249 : n35230;
  assign n55382 = pi20 ? n37 : n55381;
  assign n55383 = pi21 ? n2957 : n6706;
  assign n55384 = pi20 ? n55383 : n7724;
  assign n55385 = pi19 ? n55382 : n55384;
  assign n55386 = pi18 ? n55380 : n55385;
  assign n55387 = pi17 ? n55361 : n55386;
  assign n55388 = pi16 ? n32 : n55387;
  assign n55389 = pi15 ? n55375 : n55388;
  assign n55390 = pi21 ? n31294 : n1056;
  assign n55391 = pi20 ? n55390 : n7724;
  assign n55392 = pi19 ? n53104 : n55391;
  assign n55393 = pi18 ? n20563 : n55392;
  assign n55394 = pi17 ? n50386 : n55393;
  assign n55395 = pi16 ? n32 : n55394;
  assign n55396 = pi21 ? n29133 : n3759;
  assign n55397 = pi20 ? n55396 : n3210;
  assign n55398 = pi19 ? n20563 : n55397;
  assign n55399 = pi18 ? n20563 : n55398;
  assign n55400 = pi17 ? n50386 : n55399;
  assign n55401 = pi16 ? n32 : n55400;
  assign n55402 = pi15 ? n55395 : n55401;
  assign n55403 = pi14 ? n55389 : n55402;
  assign n55404 = pi13 ? n55369 : n55403;
  assign n55405 = pi12 ? n55342 : n55404;
  assign n55406 = pi11 ? n55286 : n55405;
  assign n55407 = pi21 ? n20563 : n916;
  assign n55408 = pi20 ? n55407 : n3210;
  assign n55409 = pi19 ? n20563 : n55408;
  assign n55410 = pi18 ? n20563 : n55409;
  assign n55411 = pi17 ? n50386 : n55410;
  assign n55412 = pi16 ? n32 : n55411;
  assign n55413 = pi23 ? n20627 : n139;
  assign n55414 = pi22 ? n55413 : n204;
  assign n55415 = pi21 ? n20563 : n55414;
  assign n55416 = pi20 ? n55415 : n6417;
  assign n55417 = pi19 ? n20563 : n55416;
  assign n55418 = pi18 ? n20563 : n55417;
  assign n55419 = pi17 ? n50386 : n55418;
  assign n55420 = pi16 ? n32 : n55419;
  assign n55421 = pi15 ? n55412 : n55420;
  assign n55422 = pi22 ? n52290 : n204;
  assign n55423 = pi21 ? n20563 : n55422;
  assign n55424 = pi20 ? n55423 : n5830;
  assign n55425 = pi19 ? n50906 : n55424;
  assign n55426 = pi18 ? n20563 : n55425;
  assign n55427 = pi17 ? n49888 : n55426;
  assign n55428 = pi16 ? n32 : n55427;
  assign n55429 = pi23 ? n5612 : n335;
  assign n55430 = pi22 ? n55429 : n233;
  assign n55431 = pi21 ? n29133 : n55430;
  assign n55432 = pi20 ? n55431 : n5830;
  assign n55433 = pi19 ? n55292 : n55432;
  assign n55434 = pi18 ? n33245 : n55433;
  assign n55435 = pi17 ? n49894 : n55434;
  assign n55436 = pi16 ? n32 : n55435;
  assign n55437 = pi15 ? n55428 : n55436;
  assign n55438 = pi14 ? n55421 : n55437;
  assign n55439 = pi20 ? n20563 : n43935;
  assign n55440 = pi22 ? n55039 : n233;
  assign n55441 = pi21 ? n29133 : n55440;
  assign n55442 = pi20 ? n55441 : n2653;
  assign n55443 = pi19 ? n55439 : n55442;
  assign n55444 = pi18 ? n20563 : n55443;
  assign n55445 = pi17 ? n49894 : n55444;
  assign n55446 = pi16 ? n32 : n55445;
  assign n55447 = pi23 ? n11962 : n363;
  assign n55448 = pi22 ? n55447 : n685;
  assign n55449 = pi21 ? n20563 : n55448;
  assign n55450 = pi20 ? n55449 : n2653;
  assign n55451 = pi19 ? n40792 : n55450;
  assign n55452 = pi18 ? n20563 : n55451;
  assign n55453 = pi17 ? n49894 : n55452;
  assign n55454 = pi16 ? n32 : n55453;
  assign n55455 = pi15 ? n55446 : n55454;
  assign n55456 = pi22 ? n30867 : n30868;
  assign n55457 = pi21 ? n20563 : n55456;
  assign n55458 = pi20 ? n20563 : n55457;
  assign n55459 = pi21 ? n30868 : n53370;
  assign n55460 = pi20 ? n55459 : n1822;
  assign n55461 = pi19 ? n55458 : n55460;
  assign n55462 = pi18 ? n20563 : n55461;
  assign n55463 = pi17 ? n49894 : n55462;
  assign n55464 = pi16 ? n32 : n55463;
  assign n55465 = pi22 ? n35902 : n316;
  assign n55466 = pi21 ? n30868 : n55465;
  assign n55467 = pi20 ? n55466 : n32;
  assign n55468 = pi19 ? n47159 : n55467;
  assign n55469 = pi18 ? n20563 : n55468;
  assign n55470 = pi17 ? n49894 : n55469;
  assign n55471 = pi16 ? n32 : n55470;
  assign n55472 = pi15 ? n55464 : n55471;
  assign n55473 = pi14 ? n55455 : n55472;
  assign n55474 = pi13 ? n55438 : n55473;
  assign n55475 = pi21 ? n20563 : n40986;
  assign n55476 = pi20 ? n20563 : n55475;
  assign n55477 = pi21 ? n36659 : n42178;
  assign n55478 = pi20 ? n55477 : n32;
  assign n55479 = pi19 ? n55476 : n55478;
  assign n55480 = pi18 ? n20563 : n55479;
  assign n55481 = pi17 ? n54273 : n55480;
  assign n55482 = pi16 ? n32 : n55481;
  assign n55483 = pi21 ? n47321 : n20563;
  assign n55484 = pi20 ? n55483 : n20563;
  assign n55485 = pi19 ? n32 : n55484;
  assign n55486 = pi18 ? n55485 : n20563;
  assign n55487 = pi20 ? n37 : n55475;
  assign n55488 = pi23 ? n157 : n35938;
  assign n55489 = pi22 ? n55488 : n1407;
  assign n55490 = pi21 ? n36659 : n55489;
  assign n55491 = pi20 ? n55490 : n32;
  assign n55492 = pi19 ? n55487 : n55491;
  assign n55493 = pi18 ? n20563 : n55492;
  assign n55494 = pi17 ? n55486 : n55493;
  assign n55495 = pi16 ? n32 : n55494;
  assign n55496 = pi15 ? n55482 : n55495;
  assign n55497 = pi21 ? n32 : n52822;
  assign n55498 = pi21 ? n30868 : n46116;
  assign n55499 = pi20 ? n55497 : n55498;
  assign n55500 = pi19 ? n32 : n55499;
  assign n55501 = pi24 ? n30868 : n20563;
  assign n55502 = pi23 ? n30868 : n55501;
  assign n55503 = pi22 ? n39190 : n55502;
  assign n55504 = pi21 ? n55503 : n40386;
  assign n55505 = pi20 ? n55504 : n51187;
  assign n55506 = pi19 ? n55505 : n54418;
  assign n55507 = pi18 ? n55500 : n55506;
  assign n55508 = pi20 ? n38754 : n50735;
  assign n55509 = pi19 ? n55508 : n20563;
  assign n55510 = pi21 ? n36781 : n8916;
  assign n55511 = pi20 ? n55510 : n32;
  assign n55512 = pi19 ? n20563 : n55511;
  assign n55513 = pi18 ? n55509 : n55512;
  assign n55514 = pi17 ? n55507 : n55513;
  assign n55515 = pi16 ? n32 : n55514;
  assign n55516 = pi22 ? n32 : n45516;
  assign n55517 = pi21 ? n55516 : n40249;
  assign n55518 = pi20 ? n55517 : n30868;
  assign n55519 = pi19 ? n32 : n55518;
  assign n55520 = pi18 ? n55519 : n30868;
  assign n55521 = pi20 ? n30868 : n43010;
  assign n55522 = pi19 ? n30868 : n55521;
  assign n55523 = pi21 ? n36781 : n2230;
  assign n55524 = pi20 ? n55523 : n32;
  assign n55525 = pi19 ? n50101 : n55524;
  assign n55526 = pi18 ? n55522 : n55525;
  assign n55527 = pi17 ? n55520 : n55526;
  assign n55528 = pi16 ? n32 : n55527;
  assign n55529 = pi15 ? n55515 : n55528;
  assign n55530 = pi14 ? n55496 : n55529;
  assign n55531 = pi21 ? n32 : n54460;
  assign n55532 = pi20 ? n55531 : n55026;
  assign n55533 = pi19 ? n32 : n55532;
  assign n55534 = pi24 ? n33792 : n20563;
  assign n55535 = pi23 ? n33792 : n55534;
  assign n55536 = pi22 ? n37173 : n55535;
  assign n55537 = pi21 ? n55536 : n36615;
  assign n55538 = pi20 ? n55537 : n51220;
  assign n55539 = pi22 ? n36615 : n30868;
  assign n55540 = pi21 ? n55539 : n30868;
  assign n55541 = pi20 ? n55540 : n20563;
  assign n55542 = pi19 ? n55538 : n55541;
  assign n55543 = pi18 ? n55533 : n55542;
  assign n55544 = pi21 ? n30868 : n45016;
  assign n55545 = pi20 ? n55544 : n47280;
  assign n55546 = pi19 ? n55545 : n43010;
  assign n55547 = pi21 ? n36781 : n8486;
  assign n55548 = pi20 ? n55547 : n32;
  assign n55549 = pi19 ? n50101 : n55548;
  assign n55550 = pi18 ? n55546 : n55549;
  assign n55551 = pi17 ? n55543 : n55550;
  assign n55552 = pi16 ? n32 : n55551;
  assign n55553 = pi21 ? n36798 : n3523;
  assign n55554 = pi20 ? n55553 : n32;
  assign n55555 = pi19 ? n20563 : n55554;
  assign n55556 = pi18 ? n20563 : n55555;
  assign n55557 = pi17 ? n49451 : n55556;
  assign n55558 = pi16 ? n32 : n55557;
  assign n55559 = pi15 ? n55552 : n55558;
  assign n55560 = pi22 ? n13481 : n32;
  assign n55561 = pi21 ? n43198 : n55560;
  assign n55562 = pi20 ? n55561 : n32;
  assign n55563 = pi19 ? n20563 : n55562;
  assign n55564 = pi18 ? n20563 : n55563;
  assign n55565 = pi17 ? n49451 : n55564;
  assign n55566 = pi16 ? n32 : n55565;
  assign n55567 = pi24 ? n30868 : n33792;
  assign n55568 = pi23 ? n55567 : n363;
  assign n55569 = pi22 ? n55568 : n43198;
  assign n55570 = pi21 ? n55569 : n882;
  assign n55571 = pi20 ? n55570 : n32;
  assign n55572 = pi19 ? n42915 : n55571;
  assign n55573 = pi18 ? n20563 : n55572;
  assign n55574 = pi17 ? n49448 : n55573;
  assign n55575 = pi16 ? n32 : n55574;
  assign n55576 = pi15 ? n55566 : n55575;
  assign n55577 = pi14 ? n55559 : n55576;
  assign n55578 = pi13 ? n55530 : n55577;
  assign n55579 = pi12 ? n55474 : n55578;
  assign n55580 = pi24 ? n33792 : n36659;
  assign n55581 = pi23 ? n55580 : n157;
  assign n55582 = pi22 ? n55581 : n14626;
  assign n55583 = pi21 ? n55582 : n882;
  assign n55584 = pi20 ? n55583 : n32;
  assign n55585 = pi19 ? n47159 : n55584;
  assign n55586 = pi18 ? n20563 : n55585;
  assign n55587 = pi17 ? n49448 : n55586;
  assign n55588 = pi16 ? n32 : n55587;
  assign n55589 = pi22 ? n55054 : n51564;
  assign n55590 = pi21 ? n55589 : n53983;
  assign n55591 = pi20 ? n55590 : n32;
  assign n55592 = pi19 ? n55476 : n55591;
  assign n55593 = pi18 ? n20563 : n55592;
  assign n55594 = pi17 ? n49448 : n55593;
  assign n55595 = pi16 ? n32 : n55594;
  assign n55596 = pi15 ? n55588 : n55595;
  assign n55597 = pi22 ? n43199 : n13481;
  assign n55598 = pi21 ? n55597 : n32;
  assign n55599 = pi20 ? n55598 : n32;
  assign n55600 = pi19 ? n55476 : n55599;
  assign n55601 = pi18 ? n20563 : n55600;
  assign n55602 = pi17 ? n49440 : n55601;
  assign n55603 = pi16 ? n32 : n55602;
  assign n55604 = pi21 ? n20563 : n37878;
  assign n55605 = pi20 ? n20563 : n55604;
  assign n55606 = pi22 ? n53550 : n13481;
  assign n55607 = pi21 ? n55606 : n32;
  assign n55608 = pi20 ? n55607 : n32;
  assign n55609 = pi19 ? n55605 : n55608;
  assign n55610 = pi18 ? n20563 : n55609;
  assign n55611 = pi17 ? n49900 : n55610;
  assign n55612 = pi16 ? n32 : n55611;
  assign n55613 = pi15 ? n55603 : n55612;
  assign n55614 = pi14 ? n55596 : n55613;
  assign n55615 = pi20 ? n53943 : n38754;
  assign n55616 = pi19 ? n32 : n55615;
  assign n55617 = pi19 ? n55521 : n30868;
  assign n55618 = pi18 ? n55616 : n55617;
  assign n55619 = pi19 ? n51301 : n42014;
  assign n55620 = pi21 ? n30868 : n51313;
  assign n55621 = pi20 ? n20563 : n55620;
  assign n55622 = pi23 ? n36798 : n14626;
  assign n55623 = pi22 ? n55622 : n2192;
  assign n55624 = pi21 ? n55623 : n32;
  assign n55625 = pi20 ? n55624 : n32;
  assign n55626 = pi19 ? n55621 : n55625;
  assign n55627 = pi18 ? n55619 : n55626;
  assign n55628 = pi17 ? n55618 : n55627;
  assign n55629 = pi16 ? n32 : n55628;
  assign n55630 = pi21 ? n47321 : n40249;
  assign n55631 = pi20 ? n55630 : n43010;
  assign n55632 = pi19 ? n32 : n55631;
  assign n55633 = pi20 ? n30868 : n36489;
  assign n55634 = pi20 ? n30868 : n39805;
  assign n55635 = pi19 ? n55633 : n55634;
  assign n55636 = pi18 ? n55632 : n55635;
  assign n55637 = pi20 ? n38754 : n43010;
  assign n55638 = pi19 ? n55637 : n43011;
  assign n55639 = pi21 ? n30868 : n39972;
  assign n55640 = pi20 ? n20563 : n55639;
  assign n55641 = pi23 ? n43198 : n14626;
  assign n55642 = pi22 ? n55641 : n396;
  assign n55643 = pi21 ? n55642 : n32;
  assign n55644 = pi20 ? n55643 : n32;
  assign n55645 = pi19 ? n55640 : n55644;
  assign n55646 = pi18 ? n55638 : n55645;
  assign n55647 = pi17 ? n55636 : n55646;
  assign n55648 = pi16 ? n32 : n55647;
  assign n55649 = pi15 ? n55629 : n55648;
  assign n55650 = pi20 ? n40915 : n36489;
  assign n55651 = pi19 ? n55650 : n43011;
  assign n55652 = pi18 ? n55632 : n55651;
  assign n55653 = pi20 ? n38754 : n49241;
  assign n55654 = pi19 ? n55653 : n20563;
  assign n55655 = pi21 ? n36489 : n36798;
  assign n55656 = pi20 ? n20563 : n55655;
  assign n55657 = pi21 ? n53559 : n32;
  assign n55658 = pi20 ? n55657 : n32;
  assign n55659 = pi19 ? n55656 : n55658;
  assign n55660 = pi18 ? n55654 : n55659;
  assign n55661 = pi17 ? n55652 : n55660;
  assign n55662 = pi16 ? n32 : n55661;
  assign n55663 = pi21 ? n32 : n49206;
  assign n55664 = pi20 ? n55663 : n20563;
  assign n55665 = pi19 ? n32 : n55664;
  assign n55666 = pi18 ? n55665 : n20563;
  assign n55667 = pi22 ? n13481 : n706;
  assign n55668 = pi21 ? n55667 : n32;
  assign n55669 = pi20 ? n55668 : n32;
  assign n55670 = pi19 ? n55656 : n55669;
  assign n55671 = pi18 ? n20563 : n55670;
  assign n55672 = pi17 ? n55666 : n55671;
  assign n55673 = pi16 ? n32 : n55672;
  assign n55674 = pi15 ? n55662 : n55673;
  assign n55675 = pi14 ? n55649 : n55674;
  assign n55676 = pi13 ? n55614 : n55675;
  assign n55677 = pi19 ? n32 : n52835;
  assign n55678 = pi18 ? n55677 : n30868;
  assign n55679 = pi21 ? n30868 : n46283;
  assign n55680 = pi20 ? n30868 : n55679;
  assign n55681 = pi19 ? n55680 : n55669;
  assign n55682 = pi18 ? n30868 : n55681;
  assign n55683 = pi17 ? n55678 : n55682;
  assign n55684 = pi16 ? n32 : n55683;
  assign n55685 = pi22 ? n30868 : n36659;
  assign n55686 = pi21 ? n55685 : n53551;
  assign n55687 = pi20 ? n30868 : n55686;
  assign n55688 = pi23 ? n13481 : n395;
  assign n55689 = pi22 ? n55688 : n32;
  assign n55690 = pi21 ? n55689 : n32;
  assign n55691 = pi20 ? n55690 : n32;
  assign n55692 = pi19 ? n55687 : n55691;
  assign n55693 = pi18 ? n30868 : n55692;
  assign n55694 = pi17 ? n55678 : n55693;
  assign n55695 = pi16 ? n32 : n55694;
  assign n55696 = pi15 ? n55684 : n55695;
  assign n55697 = pi22 ? n46789 : n36798;
  assign n55698 = pi21 ? n32 : n55697;
  assign n55699 = pi20 ? n55698 : n36798;
  assign n55700 = pi19 ? n32 : n55699;
  assign n55701 = pi21 ? n36798 : n43198;
  assign n55702 = pi20 ? n49401 : n55701;
  assign n55703 = pi20 ? n55701 : n53555;
  assign n55704 = pi19 ? n55702 : n55703;
  assign n55705 = pi18 ? n55700 : n55704;
  assign n55706 = pi20 ? n54655 : n49401;
  assign n55707 = pi19 ? n55702 : n55706;
  assign n55708 = pi22 ? n36798 : n14626;
  assign n55709 = pi21 ? n43198 : n55708;
  assign n55710 = pi20 ? n33792 : n55709;
  assign n55711 = pi19 ? n55710 : n37641;
  assign n55712 = pi18 ? n55707 : n55711;
  assign n55713 = pi17 ? n55705 : n55712;
  assign n55714 = pi16 ? n32 : n55713;
  assign n55715 = pi22 ? n43199 : n43198;
  assign n55716 = pi21 ? n55715 : n43198;
  assign n55717 = pi22 ? n43198 : n43199;
  assign n55718 = pi21 ? n43198 : n55717;
  assign n55719 = pi20 ? n55716 : n55718;
  assign n55720 = pi21 ? n43198 : n52874;
  assign n55721 = pi20 ? n43198 : n55720;
  assign n55722 = pi19 ? n55719 : n55721;
  assign n55723 = pi18 ? n49868 : n55722;
  assign n55724 = pi21 ? n43198 : n52875;
  assign n55725 = pi21 ? n43198 : n53484;
  assign n55726 = pi20 ? n55724 : n55725;
  assign n55727 = pi22 ? n52875 : n43198;
  assign n55728 = pi21 ? n55727 : n43198;
  assign n55729 = pi21 ? n33792 : n43198;
  assign n55730 = pi20 ? n55728 : n55729;
  assign n55731 = pi19 ? n55726 : n55730;
  assign n55732 = pi22 ? n43198 : n54664;
  assign n55733 = pi21 ? n39952 : n55732;
  assign n55734 = pi20 ? n55725 : n55733;
  assign n55735 = pi19 ? n55734 : n37641;
  assign n55736 = pi18 ? n55731 : n55735;
  assign n55737 = pi17 ? n55723 : n55736;
  assign n55738 = pi16 ? n32 : n55737;
  assign n55739 = pi15 ? n55714 : n55738;
  assign n55740 = pi14 ? n55696 : n55739;
  assign n55741 = pi21 ? n55125 : n50338;
  assign n55742 = pi20 ? n47411 : n55741;
  assign n55743 = pi19 ? n32 : n55742;
  assign n55744 = pi21 ? n50795 : n53977;
  assign n55745 = pi20 ? n55744 : n36659;
  assign n55746 = pi20 ? n50338 : n50342;
  assign n55747 = pi19 ? n55745 : n55746;
  assign n55748 = pi18 ? n55743 : n55747;
  assign n55749 = pi19 ? n53498 : n54611;
  assign n55750 = pi23 ? n13481 : n685;
  assign n55751 = pi22 ? n43198 : n55750;
  assign n55752 = pi21 ? n55131 : n55751;
  assign n55753 = pi20 ? n36659 : n55752;
  assign n55754 = pi19 ? n55753 : n35482;
  assign n55755 = pi18 ? n55749 : n55754;
  assign n55756 = pi17 ? n55748 : n55755;
  assign n55757 = pi16 ? n32 : n55756;
  assign n55758 = pi22 ? n43199 : n49412;
  assign n55759 = pi21 ? n55758 : n36781;
  assign n55760 = pi20 ? n51368 : n55759;
  assign n55761 = pi19 ? n32 : n55760;
  assign n55762 = pi20 ? n49414 : n36781;
  assign n55763 = pi19 ? n55762 : n36781;
  assign n55764 = pi18 ? n55761 : n55763;
  assign n55765 = pi22 ? n363 : n36781;
  assign n55766 = pi23 ? n43198 : n233;
  assign n55767 = pi22 ? n55766 : n13481;
  assign n55768 = pi21 ? n55765 : n55767;
  assign n55769 = pi20 ? n36781 : n55768;
  assign n55770 = pi19 ? n55769 : n35482;
  assign n55771 = pi18 ? n36781 : n55770;
  assign n55772 = pi17 ? n55764 : n55771;
  assign n55773 = pi16 ? n32 : n55772;
  assign n55774 = pi15 ? n55757 : n55773;
  assign n55775 = pi20 ? n51368 : n52435;
  assign n55776 = pi19 ? n32 : n55775;
  assign n55777 = pi21 ? n36781 : n53537;
  assign n55778 = pi20 ? n55777 : n36781;
  assign n55779 = pi20 ? n42170 : n36781;
  assign n55780 = pi19 ? n55778 : n55779;
  assign n55781 = pi18 ? n55776 : n55780;
  assign n55782 = pi19 ? n55779 : n40001;
  assign n55783 = pi24 ? n36798 : n43198;
  assign n55784 = pi23 ? n55783 : n685;
  assign n55785 = pi22 ? n55784 : n55688;
  assign n55786 = pi21 ? n39972 : n55785;
  assign n55787 = pi20 ? n36781 : n55786;
  assign n55788 = pi19 ? n55787 : n32;
  assign n55789 = pi18 ? n55782 : n55788;
  assign n55790 = pi17 ? n55781 : n55789;
  assign n55791 = pi16 ? n32 : n55790;
  assign n55792 = pi22 ? n53550 : n43198;
  assign n55793 = pi21 ? n55792 : n47396;
  assign n55794 = pi20 ? n48857 : n55793;
  assign n55795 = pi19 ? n32 : n55794;
  assign n55796 = pi20 ? n43198 : n53555;
  assign n55797 = pi19 ? n55796 : n54658;
  assign n55798 = pi18 ? n55795 : n55797;
  assign n55799 = pi23 ? n43198 : n36798;
  assign n55800 = pi22 ? n55799 : n36798;
  assign n55801 = pi21 ? n43198 : n55800;
  assign n55802 = pi20 ? n36798 : n55801;
  assign n55803 = pi19 ? n55802 : n36798;
  assign n55804 = pi18 ? n55803 : n54668;
  assign n55805 = pi17 ? n55798 : n55804;
  assign n55806 = pi16 ? n32 : n55805;
  assign n55807 = pi15 ? n55791 : n55806;
  assign n55808 = pi14 ? n55774 : n55807;
  assign n55809 = pi13 ? n55740 : n55808;
  assign n55810 = pi12 ? n55676 : n55809;
  assign n55811 = pi11 ? n55579 : n55810;
  assign n55812 = pi10 ? n55406 : n55811;
  assign n55813 = pi09 ? n55196 : n55812;
  assign n55814 = pi17 ? n41631 : n55180;
  assign n55815 = pi16 ? n32 : n55814;
  assign n55816 = pi15 ? n32 : n55815;
  assign n55817 = pi17 ? n41631 : n55186;
  assign n55818 = pi16 ? n32 : n55817;
  assign n55819 = pi17 ? n41642 : n55186;
  assign n55820 = pi16 ? n32 : n55819;
  assign n55821 = pi15 ? n55818 : n55820;
  assign n55822 = pi14 ? n55816 : n55821;
  assign n55823 = pi13 ? n32 : n55822;
  assign n55824 = pi12 ? n32 : n55823;
  assign n55825 = pi11 ? n32 : n55824;
  assign n55826 = pi10 ? n32 : n55825;
  assign n55827 = pi17 ? n42700 : n55200;
  assign n55828 = pi16 ? n32 : n55827;
  assign n55829 = pi17 ? n41158 : n55206;
  assign n55830 = pi16 ? n32 : n55829;
  assign n55831 = pi15 ? n55828 : n55830;
  assign n55832 = pi17 ? n41169 : n55213;
  assign n55833 = pi16 ? n32 : n55832;
  assign n55834 = pi17 ? n40498 : n55219;
  assign n55835 = pi16 ? n32 : n55834;
  assign n55836 = pi15 ? n55833 : n55835;
  assign n55837 = pi14 ? n55831 : n55836;
  assign n55838 = pi20 ? n31220 : n24781;
  assign n55839 = pi19 ? n20563 : n55838;
  assign n55840 = pi18 ? n20563 : n55839;
  assign n55841 = pi17 ? n40498 : n55840;
  assign n55842 = pi16 ? n32 : n55841;
  assign n55843 = pi17 ? n41683 : n55840;
  assign n55844 = pi16 ? n32 : n55843;
  assign n55845 = pi15 ? n55842 : n55844;
  assign n55846 = pi21 ? n569 : n2578;
  assign n55847 = pi20 ? n36872 : n55846;
  assign n55848 = pi19 ? n20563 : n55847;
  assign n55849 = pi18 ? n20563 : n55848;
  assign n55850 = pi17 ? n40511 : n55849;
  assign n55851 = pi16 ? n32 : n55850;
  assign n55852 = pi20 ? n31220 : n55846;
  assign n55853 = pi19 ? n20563 : n55852;
  assign n55854 = pi18 ? n20563 : n55853;
  assign n55855 = pi17 ? n39374 : n55854;
  assign n55856 = pi16 ? n32 : n55855;
  assign n55857 = pi15 ? n55851 : n55856;
  assign n55858 = pi14 ? n55845 : n55857;
  assign n55859 = pi13 ? n55837 : n55858;
  assign n55860 = pi21 ? n569 : n2637;
  assign n55861 = pi20 ? n31220 : n55860;
  assign n55862 = pi19 ? n20563 : n55861;
  assign n55863 = pi18 ? n20563 : n55862;
  assign n55864 = pi17 ? n40533 : n55863;
  assign n55865 = pi16 ? n32 : n55864;
  assign n55866 = pi20 ? n31220 : n40649;
  assign n55867 = pi19 ? n20563 : n55866;
  assign n55868 = pi18 ? n20563 : n55867;
  assign n55869 = pi17 ? n40046 : n55868;
  assign n55870 = pi16 ? n32 : n55869;
  assign n55871 = pi15 ? n55865 : n55870;
  assign n55872 = pi20 ? n31220 : n25760;
  assign n55873 = pi19 ? n20563 : n55872;
  assign n55874 = pi18 ? n20563 : n55873;
  assign n55875 = pi17 ? n40046 : n55874;
  assign n55876 = pi16 ? n32 : n55875;
  assign n55877 = pi21 ? n2106 : n928;
  assign n55878 = pi20 ? n31220 : n55877;
  assign n55879 = pi19 ? n20563 : n55878;
  assign n55880 = pi18 ? n20563 : n55879;
  assign n55881 = pi17 ? n39398 : n55880;
  assign n55882 = pi16 ? n32 : n55881;
  assign n55883 = pi15 ? n55876 : n55882;
  assign n55884 = pi14 ? n55871 : n55883;
  assign n55885 = pi20 ? n31220 : n40142;
  assign n55886 = pi19 ? n20563 : n55885;
  assign n55887 = pi18 ? n20563 : n55886;
  assign n55888 = pi17 ? n40551 : n55887;
  assign n55889 = pi16 ? n32 : n55888;
  assign n55890 = pi21 ? n11208 : n2678;
  assign n55891 = pi20 ? n31220 : n55890;
  assign n55892 = pi19 ? n20563 : n55891;
  assign n55893 = pi18 ? n20563 : n55892;
  assign n55894 = pi17 ? n45393 : n55893;
  assign n55895 = pi16 ? n32 : n55894;
  assign n55896 = pi15 ? n55889 : n55895;
  assign n55897 = pi17 ? n37929 : n55281;
  assign n55898 = pi16 ? n32 : n55897;
  assign n55899 = pi14 ? n55896 : n55898;
  assign n55900 = pi13 ? n55884 : n55899;
  assign n55901 = pi12 ? n55859 : n55900;
  assign n55902 = pi17 ? n37929 : n55289;
  assign n55903 = pi16 ? n32 : n55902;
  assign n55904 = pi20 ? n33964 : n48905;
  assign n55905 = pi19 ? n55904 : n55294;
  assign n55906 = pi18 ? n20563 : n55905;
  assign n55907 = pi17 ? n38984 : n55906;
  assign n55908 = pi16 ? n32 : n55907;
  assign n55909 = pi15 ? n55903 : n55908;
  assign n55910 = pi19 ? n20563 : n55301;
  assign n55911 = pi18 ? n20563 : n55910;
  assign n55912 = pi17 ? n40057 : n55911;
  assign n55913 = pi16 ? n32 : n55912;
  assign n55914 = pi17 ? n40057 : n55310;
  assign n55915 = pi16 ? n32 : n55914;
  assign n55916 = pi15 ? n55913 : n55915;
  assign n55917 = pi14 ? n55909 : n55916;
  assign n55918 = pi17 ? n36870 : n55319;
  assign n55919 = pi16 ? n32 : n55918;
  assign n55920 = pi17 ? n36870 : n55324;
  assign n55921 = pi16 ? n32 : n55920;
  assign n55922 = pi15 ? n55919 : n55921;
  assign n55923 = pi20 ? n31220 : n13398;
  assign n55924 = pi19 ? n53012 : n55923;
  assign n55925 = pi18 ? n20563 : n55924;
  assign n55926 = pi17 ? n36870 : n55925;
  assign n55927 = pi16 ? n32 : n55926;
  assign n55928 = pi20 ? n31903 : n48905;
  assign n55929 = pi21 ? n31885 : n55333;
  assign n55930 = pi20 ? n55929 : n13398;
  assign n55931 = pi19 ? n55928 : n55930;
  assign n55932 = pi18 ? n20563 : n55931;
  assign n55933 = pi17 ? n37958 : n55932;
  assign n55934 = pi16 ? n32 : n55933;
  assign n55935 = pi15 ? n55927 : n55934;
  assign n55936 = pi14 ? n55922 : n55935;
  assign n55937 = pi13 ? n55917 : n55936;
  assign n55938 = pi20 ? n55343 : n13398;
  assign n55939 = pi19 ? n54234 : n55938;
  assign n55940 = pi18 ? n20563 : n55939;
  assign n55941 = pi17 ? n39000 : n55940;
  assign n55942 = pi16 ? n32 : n55941;
  assign n55943 = pi20 ? n55349 : n6935;
  assign n55944 = pi19 ? n20563 : n55943;
  assign n55945 = pi18 ? n20563 : n55944;
  assign n55946 = pi17 ? n39000 : n55945;
  assign n55947 = pi16 ? n32 : n55946;
  assign n55948 = pi15 ? n55942 : n55947;
  assign n55949 = pi17 ? n38379 : n55945;
  assign n55950 = pi16 ? n32 : n55949;
  assign n55951 = pi20 ? n55362 : n6935;
  assign n55952 = pi19 ? n20563 : n55951;
  assign n55953 = pi18 ? n20563 : n55952;
  assign n55954 = pi17 ? n38379 : n55953;
  assign n55955 = pi16 ? n32 : n55954;
  assign n55956 = pi15 ? n55950 : n55955;
  assign n55957 = pi14 ? n55948 : n55956;
  assign n55958 = pi21 ? n31294 : n6706;
  assign n55959 = pi20 ? n55958 : n7035;
  assign n55960 = pi19 ? n20563 : n55959;
  assign n55961 = pi18 ? n20563 : n55960;
  assign n55962 = pi17 ? n38379 : n55961;
  assign n55963 = pi16 ? n32 : n55962;
  assign n55964 = pi21 ? n31294 : n30195;
  assign n55965 = pi20 ? n55964 : n54068;
  assign n55966 = pi20 ? n54701 : n40358;
  assign n55967 = pi19 ? n55965 : n55966;
  assign n55968 = pi20 ? n37 : n36249;
  assign n55969 = pi22 ? n37 : n43579;
  assign n55970 = pi21 ? n55969 : n6706;
  assign n55971 = pi20 ? n55970 : n7724;
  assign n55972 = pi19 ? n55968 : n55971;
  assign n55973 = pi18 ? n55967 : n55972;
  assign n55974 = pi17 ? n39456 : n55973;
  assign n55975 = pi16 ? n32 : n55974;
  assign n55976 = pi15 ? n55963 : n55975;
  assign n55977 = pi21 ? n20563 : n1056;
  assign n55978 = pi20 ? n55977 : n7724;
  assign n55979 = pi19 ? n53104 : n55978;
  assign n55980 = pi18 ? n20563 : n55979;
  assign n55981 = pi17 ? n39456 : n55980;
  assign n55982 = pi16 ? n32 : n55981;
  assign n55983 = pi17 ? n39456 : n55399;
  assign n55984 = pi16 ? n32 : n55983;
  assign n55985 = pi15 ? n55982 : n55984;
  assign n55986 = pi14 ? n55976 : n55985;
  assign n55987 = pi13 ? n55957 : n55986;
  assign n55988 = pi12 ? n55937 : n55987;
  assign n55989 = pi11 ? n55901 : n55988;
  assign n55990 = pi17 ? n39456 : n55410;
  assign n55991 = pi16 ? n32 : n55990;
  assign n55992 = pi17 ? n35764 : n55418;
  assign n55993 = pi16 ? n32 : n55992;
  assign n55994 = pi15 ? n55991 : n55993;
  assign n55995 = pi17 ? n35764 : n55426;
  assign n55996 = pi16 ? n32 : n55995;
  assign n55997 = pi18 ? n39432 : n55433;
  assign n55998 = pi17 ? n36215 : n55997;
  assign n55999 = pi16 ? n32 : n55998;
  assign n56000 = pi15 ? n55996 : n55999;
  assign n56001 = pi14 ? n55994 : n56000;
  assign n56002 = pi22 ? n55447 : n233;
  assign n56003 = pi21 ? n29133 : n56002;
  assign n56004 = pi20 ? n56003 : n2653;
  assign n56005 = pi19 ? n55439 : n56004;
  assign n56006 = pi18 ? n20563 : n56005;
  assign n56007 = pi17 ? n36215 : n56006;
  assign n56008 = pi16 ? n32 : n56007;
  assign n56009 = pi17 ? n36215 : n55452;
  assign n56010 = pi16 ? n32 : n56009;
  assign n56011 = pi15 ? n56008 : n56010;
  assign n56012 = pi22 ? n36617 : n30868;
  assign n56013 = pi21 ? n20563 : n56012;
  assign n56014 = pi20 ? n20563 : n56013;
  assign n56015 = pi19 ? n56014 : n55460;
  assign n56016 = pi18 ? n20563 : n56015;
  assign n56017 = pi17 ? n36215 : n56016;
  assign n56018 = pi16 ? n32 : n56017;
  assign n56019 = pi17 ? n50390 : n55469;
  assign n56020 = pi16 ? n32 : n56019;
  assign n56021 = pi15 ? n56018 : n56020;
  assign n56022 = pi14 ? n56011 : n56021;
  assign n56023 = pi13 ? n56001 : n56022;
  assign n56024 = pi17 ? n50390 : n55480;
  assign n56025 = pi16 ? n32 : n56024;
  assign n56026 = pi23 ? n157 : n43198;
  assign n56027 = pi22 ? n56026 : n1407;
  assign n56028 = pi21 ? n36659 : n56027;
  assign n56029 = pi20 ? n56028 : n32;
  assign n56030 = pi19 ? n55487 : n56029;
  assign n56031 = pi18 ? n20563 : n56030;
  assign n56032 = pi17 ? n50390 : n56031;
  assign n56033 = pi16 ? n32 : n56032;
  assign n56034 = pi15 ? n56025 : n56033;
  assign n56035 = pi20 ? n47848 : n40915;
  assign n56036 = pi19 ? n32 : n56035;
  assign n56037 = pi22 ? n39190 : n39174;
  assign n56038 = pi21 ? n56037 : n40913;
  assign n56039 = pi20 ? n56038 : n51187;
  assign n56040 = pi19 ? n56039 : n54418;
  assign n56041 = pi18 ? n56036 : n56040;
  assign n56042 = pi17 ? n56041 : n55513;
  assign n56043 = pi16 ? n32 : n56042;
  assign n56044 = pi19 ? n32 : n47849;
  assign n56045 = pi18 ? n56044 : n30868;
  assign n56046 = pi17 ? n56045 : n55526;
  assign n56047 = pi16 ? n32 : n56046;
  assign n56048 = pi15 ? n56043 : n56047;
  assign n56049 = pi14 ? n56034 : n56048;
  assign n56050 = pi20 ? n51731 : n40958;
  assign n56051 = pi19 ? n32 : n56050;
  assign n56052 = pi22 ? n37173 : n39291;
  assign n56053 = pi21 ? n56052 : n40955;
  assign n56054 = pi20 ? n56053 : n51220;
  assign n56055 = pi19 ? n56054 : n55541;
  assign n56056 = pi18 ? n56051 : n56055;
  assign n56057 = pi17 ? n56056 : n55550;
  assign n56058 = pi16 ? n32 : n56057;
  assign n56059 = pi17 ? n50905 : n55556;
  assign n56060 = pi16 ? n32 : n56059;
  assign n56061 = pi15 ? n56058 : n56060;
  assign n56062 = pi17 ? n50905 : n55564;
  assign n56063 = pi16 ? n32 : n56062;
  assign n56064 = pi24 ? n30868 : n36659;
  assign n56065 = pi23 ? n56064 : n363;
  assign n56066 = pi22 ? n56065 : n43198;
  assign n56067 = pi21 ? n56066 : n882;
  assign n56068 = pi20 ? n56067 : n32;
  assign n56069 = pi19 ? n42915 : n56068;
  assign n56070 = pi18 ? n20563 : n56069;
  assign n56071 = pi17 ? n50905 : n56070;
  assign n56072 = pi16 ? n32 : n56071;
  assign n56073 = pi15 ? n56063 : n56072;
  assign n56074 = pi14 ? n56061 : n56073;
  assign n56075 = pi13 ? n56049 : n56074;
  assign n56076 = pi12 ? n56023 : n56075;
  assign n56077 = pi17 ? n49894 : n55586;
  assign n56078 = pi16 ? n32 : n56077;
  assign n56079 = pi24 ? n36659 : n36781;
  assign n56080 = pi23 ? n56079 : n157;
  assign n56081 = pi22 ? n56080 : n51564;
  assign n56082 = pi21 ? n56081 : n53983;
  assign n56083 = pi20 ? n56082 : n32;
  assign n56084 = pi19 ? n55476 : n56083;
  assign n56085 = pi18 ? n20563 : n56084;
  assign n56086 = pi17 ? n49894 : n56085;
  assign n56087 = pi16 ? n32 : n56086;
  assign n56088 = pi15 ? n56078 : n56087;
  assign n56089 = pi17 ? n50393 : n55601;
  assign n56090 = pi16 ? n32 : n56089;
  assign n56091 = pi17 ? n50393 : n55610;
  assign n56092 = pi16 ? n32 : n56091;
  assign n56093 = pi15 ? n56090 : n56092;
  assign n56094 = pi14 ? n56088 : n56093;
  assign n56095 = pi20 ? n40054 : n38754;
  assign n56096 = pi19 ? n32 : n56095;
  assign n56097 = pi18 ? n56096 : n55617;
  assign n56098 = pi17 ? n56097 : n55627;
  assign n56099 = pi16 ? n32 : n56098;
  assign n56100 = pi20 ? n47746 : n43010;
  assign n56101 = pi19 ? n32 : n56100;
  assign n56102 = pi18 ? n56101 : n55635;
  assign n56103 = pi22 ? n54664 : n19696;
  assign n56104 = pi21 ? n56103 : n32;
  assign n56105 = pi20 ? n56104 : n32;
  assign n56106 = pi19 ? n55640 : n56105;
  assign n56107 = pi18 ? n55638 : n56106;
  assign n56108 = pi17 ? n56102 : n56107;
  assign n56109 = pi16 ? n32 : n56108;
  assign n56110 = pi15 ? n56099 : n56109;
  assign n56111 = pi23 ? n55501 : n20563;
  assign n56112 = pi22 ? n30868 : n56111;
  assign n56113 = pi21 ? n30868 : n56112;
  assign n56114 = pi20 ? n56113 : n36489;
  assign n56115 = pi19 ? n56114 : n43011;
  assign n56116 = pi18 ? n56101 : n56115;
  assign n56117 = pi17 ? n56116 : n55660;
  assign n56118 = pi16 ? n32 : n56117;
  assign n56119 = pi20 ? n47848 : n20563;
  assign n56120 = pi19 ? n32 : n56119;
  assign n56121 = pi18 ? n56120 : n20563;
  assign n56122 = pi17 ? n56121 : n55671;
  assign n56123 = pi16 ? n32 : n56122;
  assign n56124 = pi15 ? n56118 : n56123;
  assign n56125 = pi14 ? n56110 : n56124;
  assign n56126 = pi13 ? n56094 : n56125;
  assign n56127 = pi19 ? n32 : n47836;
  assign n56128 = pi18 ? n56127 : n30868;
  assign n56129 = pi22 ? n13481 : n14363;
  assign n56130 = pi21 ? n56129 : n32;
  assign n56131 = pi20 ? n56130 : n32;
  assign n56132 = pi19 ? n55680 : n56131;
  assign n56133 = pi18 ? n30868 : n56132;
  assign n56134 = pi17 ? n56128 : n56133;
  assign n56135 = pi16 ? n32 : n56134;
  assign n56136 = pi17 ? n56128 : n55693;
  assign n56137 = pi16 ? n32 : n56136;
  assign n56138 = pi15 ? n56135 : n56137;
  assign n56139 = pi18 ? n41603 : n55704;
  assign n56140 = pi17 ? n56139 : n55712;
  assign n56141 = pi16 ? n32 : n56140;
  assign n56142 = pi21 ? n49844 : n43198;
  assign n56143 = pi20 ? n32 : n56142;
  assign n56144 = pi19 ? n32 : n56143;
  assign n56145 = pi22 ? n38271 : n43198;
  assign n56146 = pi21 ? n56145 : n43198;
  assign n56147 = pi22 ? n43198 : n52875;
  assign n56148 = pi22 ? n43198 : n38271;
  assign n56149 = pi21 ? n56147 : n56148;
  assign n56150 = pi20 ? n56146 : n56149;
  assign n56151 = pi20 ? n43198 : n55725;
  assign n56152 = pi19 ? n56150 : n56151;
  assign n56153 = pi18 ? n56144 : n56152;
  assign n56154 = pi21 ? n53471 : n43198;
  assign n56155 = pi20 ? n56154 : n55729;
  assign n56156 = pi19 ? n55726 : n56155;
  assign n56157 = pi19 ? n55734 : n35482;
  assign n56158 = pi18 ? n56156 : n56157;
  assign n56159 = pi17 ? n56153 : n56158;
  assign n56160 = pi16 ? n32 : n56159;
  assign n56161 = pi15 ? n56141 : n56160;
  assign n56162 = pi14 ? n56138 : n56161;
  assign n56163 = pi20 ? n32 : n51870;
  assign n56164 = pi19 ? n32 : n56163;
  assign n56165 = pi21 ? n50795 : n43198;
  assign n56166 = pi24 ? n43198 : n36659;
  assign n56167 = pi23 ? n56166 : n36659;
  assign n56168 = pi22 ? n56167 : n36659;
  assign n56169 = pi21 ? n56168 : n36659;
  assign n56170 = pi20 ? n56165 : n56169;
  assign n56171 = pi19 ? n56170 : n55746;
  assign n56172 = pi18 ? n56164 : n56171;
  assign n56173 = pi23 ? n51564 : n685;
  assign n56174 = pi22 ? n43198 : n56173;
  assign n56175 = pi21 ? n55131 : n56174;
  assign n56176 = pi20 ? n36659 : n56175;
  assign n56177 = pi19 ? n56176 : n35482;
  assign n56178 = pi18 ? n55749 : n56177;
  assign n56179 = pi17 ? n56172 : n56178;
  assign n56180 = pi16 ? n32 : n56179;
  assign n56181 = pi22 ? n46789 : n36781;
  assign n56182 = pi21 ? n56181 : n36781;
  assign n56183 = pi20 ? n32 : n56182;
  assign n56184 = pi19 ? n32 : n56183;
  assign n56185 = pi18 ? n56184 : n36781;
  assign n56186 = pi23 ? n51564 : n13481;
  assign n56187 = pi22 ? n55766 : n56186;
  assign n56188 = pi21 ? n55765 : n56187;
  assign n56189 = pi20 ? n36781 : n56188;
  assign n56190 = pi19 ? n56189 : n32;
  assign n56191 = pi18 ? n36781 : n56190;
  assign n56192 = pi17 ? n56185 : n56191;
  assign n56193 = pi16 ? n32 : n56192;
  assign n56194 = pi15 ? n56180 : n56193;
  assign n56195 = pi21 ? n54000 : n36781;
  assign n56196 = pi20 ? n32 : n56195;
  assign n56197 = pi19 ? n32 : n56196;
  assign n56198 = pi19 ? n36781 : n55779;
  assign n56199 = pi18 ? n56197 : n56198;
  assign n56200 = pi22 ? n54664 : n55688;
  assign n56201 = pi21 ? n39972 : n56200;
  assign n56202 = pi20 ? n36781 : n56201;
  assign n56203 = pi19 ? n56202 : n32;
  assign n56204 = pi18 ? n55782 : n56203;
  assign n56205 = pi17 ? n56199 : n56204;
  assign n56206 = pi16 ? n32 : n56205;
  assign n56207 = pi22 ? n43198 : n53550;
  assign n56208 = pi21 ? n47902 : n56207;
  assign n56209 = pi20 ? n32 : n56208;
  assign n56210 = pi19 ? n32 : n56209;
  assign n56211 = pi22 ? n55799 : n43198;
  assign n56212 = pi22 ? n53550 : n36798;
  assign n56213 = pi21 ? n56211 : n56212;
  assign n56214 = pi20 ? n43198 : n56213;
  assign n56215 = pi19 ? n56214 : n54658;
  assign n56216 = pi18 ? n56210 : n56215;
  assign n56217 = pi17 ? n56216 : n55804;
  assign n56218 = pi16 ? n32 : n56217;
  assign n56219 = pi15 ? n56206 : n56218;
  assign n56220 = pi14 ? n56194 : n56219;
  assign n56221 = pi13 ? n56162 : n56220;
  assign n56222 = pi12 ? n56126 : n56221;
  assign n56223 = pi11 ? n56076 : n56222;
  assign n56224 = pi10 ? n55989 : n56223;
  assign n56225 = pi09 ? n55826 : n56224;
  assign n56226 = pi08 ? n55813 : n56225;
  assign n56227 = pi21 ? n297 : n18039;
  assign n56228 = pi20 ? n37 : n56227;
  assign n56229 = pi19 ? n20563 : n56228;
  assign n56230 = pi18 ? n20563 : n56229;
  assign n56231 = pi17 ? n42201 : n56230;
  assign n56232 = pi16 ? n32 : n56231;
  assign n56233 = pi15 ? n32 : n56232;
  assign n56234 = pi21 ? n37 : n18039;
  assign n56235 = pi20 ? n31220 : n56234;
  assign n56236 = pi19 ? n20563 : n56235;
  assign n56237 = pi18 ? n20563 : n56236;
  assign n56238 = pi17 ? n42201 : n56237;
  assign n56239 = pi16 ? n32 : n56238;
  assign n56240 = pi20 ? n31220 : n39419;
  assign n56241 = pi19 ? n20563 : n56240;
  assign n56242 = pi18 ? n20563 : n56241;
  assign n56243 = pi17 ? n48121 : n56242;
  assign n56244 = pi16 ? n32 : n56243;
  assign n56245 = pi15 ? n56239 : n56244;
  assign n56246 = pi14 ? n56233 : n56245;
  assign n56247 = pi13 ? n32 : n56246;
  assign n56248 = pi12 ? n32 : n56247;
  assign n56249 = pi11 ? n32 : n56248;
  assign n56250 = pi10 ? n32 : n56249;
  assign n56251 = pi21 ? n297 : n12003;
  assign n56252 = pi20 ? n20563 : n56251;
  assign n56253 = pi19 ? n20563 : n56252;
  assign n56254 = pi18 ? n20563 : n56253;
  assign n56255 = pi17 ? n47593 : n56254;
  assign n56256 = pi16 ? n32 : n56255;
  assign n56257 = pi21 ? n297 : n33397;
  assign n56258 = pi20 ? n31220 : n56257;
  assign n56259 = pi19 ? n20563 : n56258;
  assign n56260 = pi18 ? n20563 : n56259;
  assign n56261 = pi17 ? n41631 : n56260;
  assign n56262 = pi16 ? n32 : n56261;
  assign n56263 = pi15 ? n56256 : n56262;
  assign n56264 = pi21 ? n569 : n28467;
  assign n56265 = pi20 ? n31220 : n56264;
  assign n56266 = pi19 ? n20563 : n56265;
  assign n56267 = pi18 ? n20563 : n56266;
  assign n56268 = pi17 ? n42688 : n56267;
  assign n56269 = pi16 ? n32 : n56268;
  assign n56270 = pi21 ? n569 : n9246;
  assign n56271 = pi20 ? n31220 : n56270;
  assign n56272 = pi19 ? n20563 : n56271;
  assign n56273 = pi18 ? n20563 : n56272;
  assign n56274 = pi17 ? n40024 : n56273;
  assign n56275 = pi16 ? n32 : n56274;
  assign n56276 = pi15 ? n56269 : n56275;
  assign n56277 = pi14 ? n56263 : n56276;
  assign n56278 = pi17 ? n40024 : n55840;
  assign n56279 = pi16 ? n32 : n56278;
  assign n56280 = pi21 ? n4938 : n2578;
  assign n56281 = pi20 ? n31220 : n56280;
  assign n56282 = pi19 ? n20563 : n56281;
  assign n56283 = pi18 ? n20563 : n56282;
  assign n56284 = pi17 ? n41182 : n56283;
  assign n56285 = pi16 ? n32 : n56284;
  assign n56286 = pi15 ? n56279 : n56285;
  assign n56287 = pi17 ? n42240 : n55849;
  assign n56288 = pi16 ? n32 : n56287;
  assign n56289 = pi17 ? n40498 : n55854;
  assign n56290 = pi16 ? n32 : n56289;
  assign n56291 = pi15 ? n56288 : n56290;
  assign n56292 = pi14 ? n56286 : n56291;
  assign n56293 = pi13 ? n56277 : n56292;
  assign n56294 = pi17 ? n40498 : n55863;
  assign n56295 = pi16 ? n32 : n56294;
  assign n56296 = pi17 ? n40533 : n55868;
  assign n56297 = pi16 ? n32 : n56296;
  assign n56298 = pi15 ? n56295 : n56297;
  assign n56299 = pi22 ? n686 : n685;
  assign n56300 = pi21 ? n56299 : n2637;
  assign n56301 = pi20 ? n31220 : n56300;
  assign n56302 = pi19 ? n20563 : n56301;
  assign n56303 = pi18 ? n20563 : n56302;
  assign n56304 = pi17 ? n41709 : n56303;
  assign n56305 = pi16 ? n32 : n56304;
  assign n56306 = pi15 ? n56297 : n56305;
  assign n56307 = pi14 ? n56298 : n56306;
  assign n56308 = pi20 ? n36872 : n56300;
  assign n56309 = pi19 ? n20563 : n56308;
  assign n56310 = pi18 ? n20563 : n56309;
  assign n56311 = pi17 ? n45367 : n56310;
  assign n56312 = pi16 ? n32 : n56311;
  assign n56313 = pi20 ? n31220 : n12894;
  assign n56314 = pi19 ? n20563 : n56313;
  assign n56315 = pi18 ? n20563 : n56314;
  assign n56316 = pi17 ? n38949 : n56315;
  assign n56317 = pi16 ? n32 : n56316;
  assign n56318 = pi15 ? n56312 : n56317;
  assign n56319 = pi17 ? n40046 : n56315;
  assign n56320 = pi16 ? n32 : n56319;
  assign n56321 = pi21 ? n11208 : n928;
  assign n56322 = pi20 ? n31220 : n56321;
  assign n56323 = pi19 ? n20563 : n56322;
  assign n56324 = pi18 ? n20563 : n56323;
  assign n56325 = pi17 ? n40046 : n56324;
  assign n56326 = pi16 ? n32 : n56325;
  assign n56327 = pi15 ? n56320 : n56326;
  assign n56328 = pi14 ? n56318 : n56327;
  assign n56329 = pi13 ? n56307 : n56328;
  assign n56330 = pi12 ? n56293 : n56329;
  assign n56331 = pi21 ? n3436 : n928;
  assign n56332 = pi20 ? n31220 : n56331;
  assign n56333 = pi19 ? n20563 : n56332;
  assign n56334 = pi18 ? n20563 : n56333;
  assign n56335 = pi17 ? n40046 : n56334;
  assign n56336 = pi16 ? n32 : n56335;
  assign n56337 = pi20 ? n31220 : n12508;
  assign n56338 = pi19 ? n38478 : n56337;
  assign n56339 = pi18 ? n20563 : n56338;
  assign n56340 = pi17 ? n39398 : n56339;
  assign n56341 = pi16 ? n32 : n56340;
  assign n56342 = pi15 ? n56336 : n56341;
  assign n56343 = pi21 ? n20563 : n2957;
  assign n56344 = pi21 ? n10021 : n32;
  assign n56345 = pi20 ? n56343 : n56344;
  assign n56346 = pi19 ? n20563 : n56345;
  assign n56347 = pi18 ? n20563 : n56346;
  assign n56348 = pi17 ? n40551 : n56347;
  assign n56349 = pi16 ? n32 : n56348;
  assign n56350 = pi21 ? n20563 : n3073;
  assign n56351 = pi21 ? n52373 : n32;
  assign n56352 = pi20 ? n56350 : n56351;
  assign n56353 = pi19 ? n20563 : n56352;
  assign n56354 = pi18 ? n20563 : n56353;
  assign n56355 = pi17 ? n40551 : n56354;
  assign n56356 = pi16 ? n32 : n56355;
  assign n56357 = pi15 ? n56349 : n56356;
  assign n56358 = pi14 ? n56342 : n56357;
  assign n56359 = pi17 ? n38330 : n56354;
  assign n56360 = pi16 ? n32 : n56359;
  assign n56361 = pi21 ? n20563 : n584;
  assign n56362 = pi21 ? n41982 : n32;
  assign n56363 = pi20 ? n56361 : n56362;
  assign n56364 = pi19 ? n20563 : n56363;
  assign n56365 = pi18 ? n20563 : n56364;
  assign n56366 = pi17 ? n38330 : n56365;
  assign n56367 = pi16 ? n32 : n56366;
  assign n56368 = pi15 ? n56360 : n56367;
  assign n56369 = pi19 ? n53012 : n56363;
  assign n56370 = pi18 ? n20563 : n56369;
  assign n56371 = pi17 ? n38330 : n56370;
  assign n56372 = pi16 ? n32 : n56371;
  assign n56373 = pi20 ? n31266 : n48905;
  assign n56374 = pi21 ? n20563 : n6401;
  assign n56375 = pi20 ? n56374 : n13398;
  assign n56376 = pi19 ? n56373 : n56375;
  assign n56377 = pi18 ? n20563 : n56376;
  assign n56378 = pi17 ? n37929 : n56377;
  assign n56379 = pi16 ? n32 : n56378;
  assign n56380 = pi15 ? n56372 : n56379;
  assign n56381 = pi14 ? n56368 : n56380;
  assign n56382 = pi13 ? n56358 : n56381;
  assign n56383 = pi21 ? n3990 : n32;
  assign n56384 = pi20 ? n55343 : n56383;
  assign n56385 = pi19 ? n20563 : n56384;
  assign n56386 = pi18 ? n20563 : n56385;
  assign n56387 = pi17 ? n38984 : n56386;
  assign n56388 = pi16 ? n32 : n56387;
  assign n56389 = pi21 ? n20563 : n214;
  assign n56390 = pi21 ? n8454 : n32;
  assign n56391 = pi20 ? n56389 : n56390;
  assign n56392 = pi19 ? n20563 : n56391;
  assign n56393 = pi18 ? n20563 : n56392;
  assign n56394 = pi17 ? n38984 : n56393;
  assign n56395 = pi16 ? n32 : n56394;
  assign n56396 = pi15 ? n56388 : n56395;
  assign n56397 = pi21 ? n20563 : n7195;
  assign n56398 = pi21 ? n8464 : n32;
  assign n56399 = pi20 ? n56397 : n56398;
  assign n56400 = pi19 ? n20563 : n56399;
  assign n56401 = pi18 ? n20563 : n56400;
  assign n56402 = pi17 ? n37936 : n56401;
  assign n56403 = pi16 ? n32 : n56402;
  assign n56404 = pi20 ? n56397 : n15407;
  assign n56405 = pi19 ? n20563 : n56404;
  assign n56406 = pi18 ? n20563 : n56405;
  assign n56407 = pi17 ? n37936 : n56406;
  assign n56408 = pi16 ? n32 : n56407;
  assign n56409 = pi15 ? n56403 : n56408;
  assign n56410 = pi14 ? n56396 : n56409;
  assign n56411 = pi21 ? n20563 : n2074;
  assign n56412 = pi20 ? n56411 : n16519;
  assign n56413 = pi19 ? n20563 : n56412;
  assign n56414 = pi18 ? n20563 : n56413;
  assign n56415 = pi17 ? n37936 : n56414;
  assign n56416 = pi16 ? n32 : n56415;
  assign n56417 = pi20 ? n31220 : n36249;
  assign n56418 = pi20 ? n56411 : n9963;
  assign n56419 = pi19 ? n56417 : n56418;
  assign n56420 = pi18 ? n20563 : n56419;
  assign n56421 = pi17 ? n36870 : n56420;
  assign n56422 = pi16 ? n32 : n56421;
  assign n56423 = pi15 ? n56416 : n56422;
  assign n56424 = pi21 ? n20563 : n17764;
  assign n56425 = pi20 ? n56424 : n9963;
  assign n56426 = pi19 ? n20563 : n56425;
  assign n56427 = pi18 ? n20563 : n56426;
  assign n56428 = pi17 ? n36870 : n56427;
  assign n56429 = pi16 ? n32 : n56428;
  assign n56430 = pi21 ? n20563 : n767;
  assign n56431 = pi20 ? n56430 : n12149;
  assign n56432 = pi19 ? n20563 : n56431;
  assign n56433 = pi18 ? n20563 : n56432;
  assign n56434 = pi17 ? n36870 : n56433;
  assign n56435 = pi16 ? n32 : n56434;
  assign n56436 = pi15 ? n56429 : n56435;
  assign n56437 = pi14 ? n56423 : n56436;
  assign n56438 = pi13 ? n56410 : n56437;
  assign n56439 = pi12 ? n56382 : n56438;
  assign n56440 = pi11 ? n56330 : n56439;
  assign n56441 = pi21 ? n20563 : n7468;
  assign n56442 = pi20 ? n56441 : n4008;
  assign n56443 = pi19 ? n20563 : n56442;
  assign n56444 = pi18 ? n20563 : n56443;
  assign n56445 = pi17 ? n37323 : n56444;
  assign n56446 = pi16 ? n32 : n56445;
  assign n56447 = pi22 ? n55413 : n316;
  assign n56448 = pi21 ? n20563 : n56447;
  assign n56449 = pi20 ? n56448 : n4008;
  assign n56450 = pi19 ? n20563 : n56449;
  assign n56451 = pi18 ? n20563 : n56450;
  assign n56452 = pi17 ? n37323 : n56451;
  assign n56453 = pi16 ? n32 : n56452;
  assign n56454 = pi15 ? n56446 : n56453;
  assign n56455 = pi20 ? n42006 : n43935;
  assign n56456 = pi19 ? n56455 : n20563;
  assign n56457 = pi18 ? n37322 : n56456;
  assign n56458 = pi24 ? n37 : n30868;
  assign n56459 = pi23 ? n56458 : n335;
  assign n56460 = pi22 ? n56459 : n204;
  assign n56461 = pi21 ? n20563 : n56460;
  assign n56462 = pi20 ? n56461 : n3340;
  assign n56463 = pi19 ? n50906 : n56462;
  assign n56464 = pi18 ? n20563 : n56463;
  assign n56465 = pi17 ? n56457 : n56464;
  assign n56466 = pi16 ? n32 : n56465;
  assign n56467 = pi24 ? n20563 : n139;
  assign n56468 = pi23 ? n56467 : n335;
  assign n56469 = pi22 ? n56468 : n233;
  assign n56470 = pi21 ? n29133 : n56469;
  assign n56471 = pi20 ? n56470 : n5830;
  assign n56472 = pi19 ? n50854 : n56471;
  assign n56473 = pi18 ? n20563 : n56472;
  assign n56474 = pi17 ? n37336 : n56473;
  assign n56475 = pi16 ? n32 : n56474;
  assign n56476 = pi15 ? n56466 : n56475;
  assign n56477 = pi14 ? n56454 : n56476;
  assign n56478 = pi24 ? n30868 : n335;
  assign n56479 = pi23 ? n56478 : n363;
  assign n56480 = pi22 ? n56479 : n233;
  assign n56481 = pi21 ? n20563 : n56480;
  assign n56482 = pi20 ? n56481 : n2653;
  assign n56483 = pi19 ? n20563 : n56482;
  assign n56484 = pi18 ? n20563 : n56483;
  assign n56485 = pi17 ? n37336 : n56484;
  assign n56486 = pi16 ? n32 : n56485;
  assign n56487 = pi22 ? n37 : n30868;
  assign n56488 = pi21 ? n20563 : n56487;
  assign n56489 = pi20 ? n20563 : n56488;
  assign n56490 = pi22 ? n56479 : n685;
  assign n56491 = pi21 ? n20563 : n56490;
  assign n56492 = pi20 ? n56491 : n37640;
  assign n56493 = pi19 ? n56489 : n56492;
  assign n56494 = pi18 ? n20563 : n56493;
  assign n56495 = pi17 ? n37336 : n56494;
  assign n56496 = pi16 ? n32 : n56495;
  assign n56497 = pi15 ? n56486 : n56496;
  assign n56498 = pi21 ? n30868 : n55055;
  assign n56499 = pi20 ? n56498 : n2653;
  assign n56500 = pi19 ? n56489 : n56499;
  assign n56501 = pi18 ? n20563 : n56500;
  assign n56502 = pi17 ? n37336 : n56501;
  assign n56503 = pi16 ? n32 : n56502;
  assign n56504 = pi22 ? n35902 : n685;
  assign n56505 = pi21 ? n30868 : n56504;
  assign n56506 = pi20 ? n56505 : n32;
  assign n56507 = pi19 ? n47159 : n56506;
  assign n56508 = pi18 ? n20563 : n56507;
  assign n56509 = pi17 ? n36162 : n56508;
  assign n56510 = pi16 ? n32 : n56509;
  assign n56511 = pi15 ? n56503 : n56510;
  assign n56512 = pi14 ? n56497 : n56511;
  assign n56513 = pi13 ? n56477 : n56512;
  assign n56514 = pi22 ? n15294 : n13481;
  assign n56515 = pi21 ? n36659 : n56514;
  assign n56516 = pi20 ? n56515 : n32;
  assign n56517 = pi19 ? n55476 : n56516;
  assign n56518 = pi18 ? n20563 : n56517;
  assign n56519 = pi17 ? n36162 : n56518;
  assign n56520 = pi16 ? n32 : n56519;
  assign n56521 = pi22 ? n53550 : n316;
  assign n56522 = pi21 ? n36659 : n56521;
  assign n56523 = pi20 ? n56522 : n32;
  assign n56524 = pi19 ? n55487 : n56523;
  assign n56525 = pi18 ? n20563 : n56524;
  assign n56526 = pi17 ? n36162 : n56525;
  assign n56527 = pi16 ? n32 : n56526;
  assign n56528 = pi15 ? n56520 : n56527;
  assign n56529 = pi22 ? n32 : n40386;
  assign n56530 = pi21 ? n56529 : n40917;
  assign n56531 = pi20 ? n32 : n56530;
  assign n56532 = pi19 ? n32 : n56531;
  assign n56533 = pi23 ? n20563 : n55501;
  assign n56534 = pi22 ? n56533 : n20563;
  assign n56535 = pi21 ? n56534 : n45049;
  assign n56536 = pi20 ? n39192 : n56535;
  assign n56537 = pi19 ? n56536 : n20563;
  assign n56538 = pi18 ? n56532 : n56537;
  assign n56539 = pi21 ? n20563 : n51270;
  assign n56540 = pi20 ? n20563 : n56539;
  assign n56541 = pi22 ? n233 : n21502;
  assign n56542 = pi21 ? n36781 : n56541;
  assign n56543 = pi20 ? n56542 : n32;
  assign n56544 = pi19 ? n56540 : n56543;
  assign n56545 = pi18 ? n20563 : n56544;
  assign n56546 = pi17 ? n56538 : n56545;
  assign n56547 = pi16 ? n32 : n56546;
  assign n56548 = pi21 ? n56529 : n36489;
  assign n56549 = pi20 ? n32 : n56548;
  assign n56550 = pi19 ? n32 : n56549;
  assign n56551 = pi18 ? n56550 : n30868;
  assign n56552 = pi21 ? n30868 : n51270;
  assign n56553 = pi20 ? n20563 : n56552;
  assign n56554 = pi22 ? n685 : n21502;
  assign n56555 = pi21 ? n36781 : n56554;
  assign n56556 = pi20 ? n56555 : n32;
  assign n56557 = pi19 ? n56553 : n56556;
  assign n56558 = pi18 ? n55522 : n56557;
  assign n56559 = pi17 ? n56551 : n56558;
  assign n56560 = pi16 ? n32 : n56559;
  assign n56561 = pi15 ? n56547 : n56560;
  assign n56562 = pi14 ? n56528 : n56561;
  assign n56563 = pi22 ? n32 : n36615;
  assign n56564 = pi21 ? n56563 : n40960;
  assign n56565 = pi20 ? n32 : n56564;
  assign n56566 = pi19 ? n32 : n56565;
  assign n56567 = pi21 ? n20563 : n52246;
  assign n56568 = pi23 ? n20563 : n55534;
  assign n56569 = pi22 ? n56568 : n40386;
  assign n56570 = pi22 ? n42106 : n20563;
  assign n56571 = pi21 ? n56569 : n56570;
  assign n56572 = pi20 ? n56567 : n56571;
  assign n56573 = pi20 ? n48184 : n20563;
  assign n56574 = pi19 ? n56572 : n56573;
  assign n56575 = pi18 ? n56566 : n56574;
  assign n56576 = pi20 ? n39805 : n20563;
  assign n56577 = pi19 ? n56576 : n43010;
  assign n56578 = pi18 ? n56577 : n55549;
  assign n56579 = pi17 ? n56575 : n56578;
  assign n56580 = pi16 ? n32 : n56579;
  assign n56581 = pi17 ? n55361 : n55556;
  assign n56582 = pi16 ? n32 : n56581;
  assign n56583 = pi15 ? n56580 : n56582;
  assign n56584 = pi17 ? n55361 : n55564;
  assign n56585 = pi16 ? n32 : n56584;
  assign n56586 = pi20 ? n20563 : n46587;
  assign n56587 = pi21 ? n46283 : n882;
  assign n56588 = pi20 ? n56587 : n32;
  assign n56589 = pi19 ? n56586 : n56588;
  assign n56590 = pi18 ? n20563 : n56589;
  assign n56591 = pi17 ? n36215 : n56590;
  assign n56592 = pi16 ? n32 : n56591;
  assign n56593 = pi15 ? n56585 : n56592;
  assign n56594 = pi14 ? n56583 : n56593;
  assign n56595 = pi13 ? n56562 : n56594;
  assign n56596 = pi12 ? n56513 : n56595;
  assign n56597 = pi21 ? n55708 : n55689;
  assign n56598 = pi20 ? n56597 : n32;
  assign n56599 = pi19 ? n42915 : n56598;
  assign n56600 = pi18 ? n20563 : n56599;
  assign n56601 = pi17 ? n36215 : n56600;
  assign n56602 = pi16 ? n32 : n56601;
  assign n56603 = pi22 ? n20563 : n42109;
  assign n56604 = pi21 ? n20563 : n56603;
  assign n56605 = pi20 ? n20563 : n56604;
  assign n56606 = pi23 ? n56079 : n36798;
  assign n56607 = pi23 ? n43198 : n51564;
  assign n56608 = pi22 ? n56606 : n56607;
  assign n56609 = pi21 ? n56608 : n53983;
  assign n56610 = pi20 ? n56609 : n32;
  assign n56611 = pi19 ? n56605 : n56610;
  assign n56612 = pi18 ? n20563 : n56611;
  assign n56613 = pi17 ? n36215 : n56612;
  assign n56614 = pi16 ? n32 : n56613;
  assign n56615 = pi15 ? n56602 : n56614;
  assign n56616 = pi23 ? n33792 : n335;
  assign n56617 = pi22 ? n20563 : n56616;
  assign n56618 = pi21 ? n20563 : n56617;
  assign n56619 = pi20 ? n20563 : n56618;
  assign n56620 = pi24 ? n36781 : n36798;
  assign n56621 = pi23 ? n56620 : n43198;
  assign n56622 = pi23 ? n14626 : n13481;
  assign n56623 = pi22 ? n56621 : n56622;
  assign n56624 = pi21 ? n56623 : n32;
  assign n56625 = pi20 ? n56624 : n32;
  assign n56626 = pi19 ? n56619 : n56625;
  assign n56627 = pi18 ? n20563 : n56626;
  assign n56628 = pi17 ? n35764 : n56627;
  assign n56629 = pi16 ? n32 : n56628;
  assign n56630 = pi21 ? n20563 : n36659;
  assign n56631 = pi20 ? n20563 : n56630;
  assign n56632 = pi22 ? n55622 : n56186;
  assign n56633 = pi21 ? n56632 : n32;
  assign n56634 = pi20 ? n56633 : n32;
  assign n56635 = pi19 ? n56631 : n56634;
  assign n56636 = pi18 ? n20563 : n56635;
  assign n56637 = pi17 ? n34859 : n56636;
  assign n56638 = pi16 ? n32 : n56637;
  assign n56639 = pi15 ? n56629 : n56638;
  assign n56640 = pi14 ? n56615 : n56639;
  assign n56641 = pi21 ? n51232 : n48173;
  assign n56642 = pi20 ? n32 : n56641;
  assign n56643 = pi19 ? n32 : n56642;
  assign n56644 = pi18 ? n56643 : n55617;
  assign n56645 = pi22 ? n30868 : n55130;
  assign n56646 = pi21 ? n30868 : n56645;
  assign n56647 = pi20 ? n20563 : n56646;
  assign n56648 = pi22 ? n55784 : n54563;
  assign n56649 = pi21 ? n56648 : n32;
  assign n56650 = pi20 ? n56649 : n32;
  assign n56651 = pi19 ? n56647 : n56650;
  assign n56652 = pi18 ? n55619 : n56651;
  assign n56653 = pi17 ? n56644 : n56652;
  assign n56654 = pi16 ? n32 : n56653;
  assign n56655 = pi22 ? n46165 : n40386;
  assign n56656 = pi21 ? n56655 : n48173;
  assign n56657 = pi20 ? n32 : n56656;
  assign n56658 = pi19 ? n32 : n56657;
  assign n56659 = pi18 ? n56658 : n30868;
  assign n56660 = pi20 ? n38754 : n30868;
  assign n56661 = pi19 ? n56660 : n56576;
  assign n56662 = pi21 ? n30868 : n36781;
  assign n56663 = pi20 ? n20563 : n56662;
  assign n56664 = pi23 ? n55783 : n51564;
  assign n56665 = pi23 ? n13481 : n14362;
  assign n56666 = pi22 ? n56664 : n56665;
  assign n56667 = pi21 ? n56666 : n32;
  assign n56668 = pi20 ? n56667 : n32;
  assign n56669 = pi19 ? n56663 : n56668;
  assign n56670 = pi18 ? n56661 : n56669;
  assign n56671 = pi17 ? n56659 : n56670;
  assign n56672 = pi16 ? n32 : n56671;
  assign n56673 = pi15 ? n56654 : n56672;
  assign n56674 = pi19 ? n30868 : n43011;
  assign n56675 = pi18 ? n56658 : n56674;
  assign n56676 = pi20 ? n38754 : n43935;
  assign n56677 = pi19 ? n56676 : n20563;
  assign n56678 = pi23 ? n14626 : n316;
  assign n56679 = pi22 ? n56678 : n21502;
  assign n56680 = pi21 ? n56679 : n32;
  assign n56681 = pi20 ? n56680 : n32;
  assign n56682 = pi19 ? n55656 : n56681;
  assign n56683 = pi18 ? n56677 : n56682;
  assign n56684 = pi17 ? n56675 : n56683;
  assign n56685 = pi16 ? n32 : n56684;
  assign n56686 = pi21 ? n39394 : n46116;
  assign n56687 = pi20 ? n32 : n56686;
  assign n56688 = pi19 ? n32 : n56687;
  assign n56689 = pi18 ? n56688 : n20563;
  assign n56690 = pi17 ? n56689 : n55671;
  assign n56691 = pi16 ? n32 : n56690;
  assign n56692 = pi15 ? n56685 : n56691;
  assign n56693 = pi14 ? n56673 : n56692;
  assign n56694 = pi13 ? n56640 : n56693;
  assign n56695 = pi22 ? n36781 : n53550;
  assign n56696 = pi21 ? n30868 : n56695;
  assign n56697 = pi20 ? n30868 : n56696;
  assign n56698 = pi22 ? n56186 : n14363;
  assign n56699 = pi21 ? n56698 : n32;
  assign n56700 = pi20 ? n56699 : n32;
  assign n56701 = pi19 ? n56697 : n56700;
  assign n56702 = pi18 ? n30868 : n56701;
  assign n56703 = pi17 ? n45624 : n56702;
  assign n56704 = pi16 ? n32 : n56703;
  assign n56705 = pi21 ? n55685 : n47397;
  assign n56706 = pi20 ? n30868 : n56705;
  assign n56707 = pi19 ? n56706 : n10012;
  assign n56708 = pi18 ? n30868 : n56707;
  assign n56709 = pi17 ? n45624 : n56708;
  assign n56710 = pi16 ? n32 : n56709;
  assign n56711 = pi15 ? n56704 : n56710;
  assign n56712 = pi23 ? n36798 : n36781;
  assign n56713 = pi22 ? n56712 : n52875;
  assign n56714 = pi21 ? n46790 : n56713;
  assign n56715 = pi20 ? n32 : n56714;
  assign n56716 = pi19 ? n32 : n56715;
  assign n56717 = pi21 ? n43198 : n47396;
  assign n56718 = pi20 ? n56717 : n55701;
  assign n56719 = pi20 ? n54009 : n47397;
  assign n56720 = pi19 ? n56718 : n56719;
  assign n56721 = pi18 ? n56716 : n56720;
  assign n56722 = pi20 ? n43198 : n49401;
  assign n56723 = pi19 ? n55702 : n56722;
  assign n56724 = pi22 ? n36798 : n55641;
  assign n56725 = pi21 ? n43198 : n56724;
  assign n56726 = pi20 ? n33792 : n56725;
  assign n56727 = pi19 ? n56726 : n37641;
  assign n56728 = pi18 ? n56723 : n56727;
  assign n56729 = pi17 ? n56721 : n56728;
  assign n56730 = pi16 ? n32 : n56729;
  assign n56731 = pi22 ? n55799 : n50339;
  assign n56732 = pi21 ? n46276 : n56731;
  assign n56733 = pi20 ? n32 : n56732;
  assign n56734 = pi19 ? n32 : n56733;
  assign n56735 = pi18 ? n56734 : n43198;
  assign n56736 = pi21 ? n50338 : n43198;
  assign n56737 = pi20 ? n43198 : n56736;
  assign n56738 = pi19 ? n51355 : n56737;
  assign n56739 = pi22 ? n43198 : n335;
  assign n56740 = pi21 ? n43198 : n56739;
  assign n56741 = pi22 ? n335 : n36781;
  assign n56742 = pi22 ? n43198 : n685;
  assign n56743 = pi21 ? n56741 : n56742;
  assign n56744 = pi20 ? n56740 : n56743;
  assign n56745 = pi19 ? n56744 : n1823;
  assign n56746 = pi18 ? n56738 : n56745;
  assign n56747 = pi17 ? n56735 : n56746;
  assign n56748 = pi16 ? n32 : n56747;
  assign n56749 = pi15 ? n56730 : n56748;
  assign n56750 = pi14 ? n56711 : n56749;
  assign n56751 = pi21 ? n50338 : n47396;
  assign n56752 = pi20 ? n50338 : n56751;
  assign n56753 = pi19 ? n43198 : n56752;
  assign n56754 = pi18 ? n56734 : n56753;
  assign n56755 = pi20 ? n50338 : n56736;
  assign n56756 = pi21 ? n43198 : n46260;
  assign n56757 = pi20 ? n56756 : n50338;
  assign n56758 = pi19 ? n56755 : n56757;
  assign n56759 = pi21 ? n38926 : n335;
  assign n56760 = pi22 ? n43198 : n51564;
  assign n56761 = pi21 ? n56741 : n56760;
  assign n56762 = pi20 ? n56759 : n56761;
  assign n56763 = pi19 ? n56762 : n35482;
  assign n56764 = pi18 ? n56758 : n56763;
  assign n56765 = pi17 ? n56754 : n56764;
  assign n56766 = pi16 ? n32 : n56765;
  assign n56767 = pi22 ? n52431 : n43199;
  assign n56768 = pi21 ? n32 : n56767;
  assign n56769 = pi20 ? n32 : n56768;
  assign n56770 = pi19 ? n32 : n56769;
  assign n56771 = pi21 ? n49413 : n36781;
  assign n56772 = pi21 ? n46283 : n36781;
  assign n56773 = pi20 ? n56771 : n56772;
  assign n56774 = pi19 ? n56773 : n36781;
  assign n56775 = pi18 ? n56770 : n56774;
  assign n56776 = pi23 ? n36781 : n157;
  assign n56777 = pi22 ? n363 : n56776;
  assign n56778 = pi22 ? n14626 : n316;
  assign n56779 = pi21 ? n56777 : n56778;
  assign n56780 = pi20 ? n36781 : n56779;
  assign n56781 = pi19 ? n56780 : n32;
  assign n56782 = pi18 ? n36781 : n56781;
  assign n56783 = pi17 ? n56775 : n56782;
  assign n56784 = pi16 ? n32 : n56783;
  assign n56785 = pi15 ? n56766 : n56784;
  assign n56786 = pi21 ? n32 : n54642;
  assign n56787 = pi20 ? n32 : n56786;
  assign n56788 = pi19 ? n32 : n56787;
  assign n56789 = pi20 ? n53538 : n56772;
  assign n56790 = pi19 ? n56789 : n55779;
  assign n56791 = pi18 ? n56788 : n56790;
  assign n56792 = pi21 ? n36798 : n55143;
  assign n56793 = pi20 ? n56792 : n36781;
  assign n56794 = pi19 ? n55779 : n56793;
  assign n56795 = pi22 ? n685 : n56665;
  assign n56796 = pi21 ? n39972 : n56795;
  assign n56797 = pi20 ? n40442 : n56796;
  assign n56798 = pi19 ? n56797 : n32;
  assign n56799 = pi18 ? n56794 : n56798;
  assign n56800 = pi17 ? n56791 : n56799;
  assign n56801 = pi16 ? n32 : n56800;
  assign n56802 = pi23 ? n46274 : n36798;
  assign n56803 = pi22 ? n56802 : n53550;
  assign n56804 = pi21 ? n32 : n56803;
  assign n56805 = pi20 ? n32 : n56804;
  assign n56806 = pi19 ? n32 : n56805;
  assign n56807 = pi18 ? n56806 : n55797;
  assign n56808 = pi20 ? n36798 : n49401;
  assign n56809 = pi19 ? n56808 : n36798;
  assign n56810 = pi22 ? n56607 : n21502;
  assign n56811 = pi21 ? n43198 : n56810;
  assign n56812 = pi20 ? n36798 : n56811;
  assign n56813 = pi19 ? n56812 : n32;
  assign n56814 = pi18 ? n56809 : n56813;
  assign n56815 = pi17 ? n56807 : n56814;
  assign n56816 = pi16 ? n32 : n56815;
  assign n56817 = pi15 ? n56801 : n56816;
  assign n56818 = pi14 ? n56785 : n56817;
  assign n56819 = pi13 ? n56750 : n56818;
  assign n56820 = pi12 ? n56694 : n56819;
  assign n56821 = pi11 ? n56596 : n56820;
  assign n56822 = pi10 ? n56440 : n56821;
  assign n56823 = pi09 ? n56250 : n56822;
  assign n56824 = pi17 ? n44274 : n56230;
  assign n56825 = pi16 ? n32 : n56824;
  assign n56826 = pi15 ? n32 : n56825;
  assign n56827 = pi17 ? n48624 : n56237;
  assign n56828 = pi16 ? n32 : n56827;
  assign n56829 = pi17 ? n42645 : n56242;
  assign n56830 = pi16 ? n32 : n56829;
  assign n56831 = pi15 ? n56828 : n56830;
  assign n56832 = pi14 ? n56826 : n56831;
  assign n56833 = pi13 ? n32 : n56832;
  assign n56834 = pi12 ? n32 : n56833;
  assign n56835 = pi11 ? n32 : n56834;
  assign n56836 = pi10 ? n32 : n56835;
  assign n56837 = pi17 ? n42655 : n56254;
  assign n56838 = pi16 ? n32 : n56837;
  assign n56839 = pi17 ? n42201 : n56260;
  assign n56840 = pi16 ? n32 : n56839;
  assign n56841 = pi15 ? n56838 : n56840;
  assign n56842 = pi21 ? n569 : n11569;
  assign n56843 = pi20 ? n31220 : n56842;
  assign n56844 = pi19 ? n20563 : n56843;
  assign n56845 = pi18 ? n20563 : n56844;
  assign n56846 = pi17 ? n43262 : n56845;
  assign n56847 = pi16 ? n32 : n56846;
  assign n56848 = pi21 ? n4938 : n3066;
  assign n56849 = pi20 ? n31220 : n56848;
  assign n56850 = pi19 ? n20563 : n56849;
  assign n56851 = pi18 ? n20563 : n56850;
  assign n56852 = pi17 ? n42688 : n56851;
  assign n56853 = pi16 ? n32 : n56852;
  assign n56854 = pi15 ? n56847 : n56853;
  assign n56855 = pi14 ? n56841 : n56854;
  assign n56856 = pi21 ? n4938 : n4109;
  assign n56857 = pi20 ? n31220 : n56856;
  assign n56858 = pi19 ? n20563 : n56857;
  assign n56859 = pi18 ? n20563 : n56858;
  assign n56860 = pi17 ? n42688 : n56859;
  assign n56861 = pi16 ? n32 : n56860;
  assign n56862 = pi17 ? n42700 : n56859;
  assign n56863 = pi16 ? n32 : n56862;
  assign n56864 = pi15 ? n56861 : n56863;
  assign n56865 = pi20 ? n36872 : n11602;
  assign n56866 = pi19 ? n20563 : n56865;
  assign n56867 = pi18 ? n20563 : n56866;
  assign n56868 = pi17 ? n46998 : n56867;
  assign n56869 = pi16 ? n32 : n56868;
  assign n56870 = pi20 ? n31220 : n12448;
  assign n56871 = pi19 ? n20563 : n56870;
  assign n56872 = pi18 ? n20563 : n56871;
  assign n56873 = pi17 ? n41169 : n56872;
  assign n56874 = pi16 ? n32 : n56873;
  assign n56875 = pi15 ? n56869 : n56874;
  assign n56876 = pi14 ? n56864 : n56875;
  assign n56877 = pi13 ? n56855 : n56876;
  assign n56878 = pi20 ? n31220 : n11610;
  assign n56879 = pi19 ? n20563 : n56878;
  assign n56880 = pi18 ? n20563 : n56879;
  assign n56881 = pi17 ? n41169 : n56880;
  assign n56882 = pi16 ? n32 : n56881;
  assign n56883 = pi21 ? n3392 : n5829;
  assign n56884 = pi20 ? n31220 : n56883;
  assign n56885 = pi19 ? n20563 : n56884;
  assign n56886 = pi18 ? n20563 : n56885;
  assign n56887 = pi17 ? n40498 : n56886;
  assign n56888 = pi16 ? n32 : n56887;
  assign n56889 = pi15 ? n56882 : n56888;
  assign n56890 = pi17 ? n40498 : n55868;
  assign n56891 = pi16 ? n32 : n56890;
  assign n56892 = pi17 ? n41683 : n56303;
  assign n56893 = pi16 ? n32 : n56892;
  assign n56894 = pi15 ? n56891 : n56893;
  assign n56895 = pi14 ? n56889 : n56894;
  assign n56896 = pi17 ? n40511 : n56310;
  assign n56897 = pi16 ? n32 : n56896;
  assign n56898 = pi17 ? n39374 : n56315;
  assign n56899 = pi16 ? n32 : n56898;
  assign n56900 = pi15 ? n56897 : n56899;
  assign n56901 = pi17 ? n40533 : n56315;
  assign n56902 = pi16 ? n32 : n56901;
  assign n56903 = pi17 ? n40533 : n56324;
  assign n56904 = pi16 ? n32 : n56903;
  assign n56905 = pi15 ? n56902 : n56904;
  assign n56906 = pi14 ? n56900 : n56905;
  assign n56907 = pi13 ? n56895 : n56906;
  assign n56908 = pi12 ? n56877 : n56907;
  assign n56909 = pi21 ? n3436 : n1009;
  assign n56910 = pi20 ? n31220 : n56909;
  assign n56911 = pi19 ? n20563 : n56910;
  assign n56912 = pi18 ? n20563 : n56911;
  assign n56913 = pi17 ? n40533 : n56912;
  assign n56914 = pi16 ? n32 : n56913;
  assign n56915 = pi17 ? n41709 : n56339;
  assign n56916 = pi16 ? n32 : n56915;
  assign n56917 = pi15 ? n56914 : n56916;
  assign n56918 = pi17 ? n45367 : n56347;
  assign n56919 = pi16 ? n32 : n56918;
  assign n56920 = pi17 ? n45367 : n56354;
  assign n56921 = pi16 ? n32 : n56920;
  assign n56922 = pi15 ? n56919 : n56921;
  assign n56923 = pi14 ? n56917 : n56922;
  assign n56924 = pi17 ? n38958 : n56354;
  assign n56925 = pi16 ? n32 : n56924;
  assign n56926 = pi17 ? n38958 : n56365;
  assign n56927 = pi16 ? n32 : n56926;
  assign n56928 = pi15 ? n56925 : n56927;
  assign n56929 = pi17 ? n38958 : n56370;
  assign n56930 = pi16 ? n32 : n56929;
  assign n56931 = pi17 ? n40046 : n56377;
  assign n56932 = pi16 ? n32 : n56931;
  assign n56933 = pi15 ? n56930 : n56932;
  assign n56934 = pi14 ? n56928 : n56933;
  assign n56935 = pi13 ? n56923 : n56934;
  assign n56936 = pi23 ? n204 : n13481;
  assign n56937 = pi22 ? n316 : n56936;
  assign n56938 = pi21 ? n56937 : n32;
  assign n56939 = pi20 ? n55343 : n56938;
  assign n56940 = pi19 ? n20563 : n56939;
  assign n56941 = pi18 ? n20563 : n56940;
  assign n56942 = pi17 ? n39398 : n56941;
  assign n56943 = pi16 ? n32 : n56942;
  assign n56944 = pi17 ? n39398 : n56393;
  assign n56945 = pi16 ? n32 : n56944;
  assign n56946 = pi15 ? n56943 : n56945;
  assign n56947 = pi17 ? n38317 : n56401;
  assign n56948 = pi16 ? n32 : n56947;
  assign n56949 = pi17 ? n38317 : n56406;
  assign n56950 = pi16 ? n32 : n56949;
  assign n56951 = pi15 ? n56948 : n56950;
  assign n56952 = pi14 ? n56946 : n56951;
  assign n56953 = pi17 ? n38317 : n56414;
  assign n56954 = pi16 ? n32 : n56953;
  assign n56955 = pi17 ? n38330 : n56420;
  assign n56956 = pi16 ? n32 : n56955;
  assign n56957 = pi15 ? n56954 : n56956;
  assign n56958 = pi20 ? n56424 : n8295;
  assign n56959 = pi19 ? n20563 : n56958;
  assign n56960 = pi18 ? n20563 : n56959;
  assign n56961 = pi17 ? n38330 : n56960;
  assign n56962 = pi16 ? n32 : n56961;
  assign n56963 = pi17 ? n38330 : n56433;
  assign n56964 = pi16 ? n32 : n56963;
  assign n56965 = pi15 ? n56962 : n56964;
  assign n56966 = pi14 ? n56957 : n56965;
  assign n56967 = pi13 ? n56952 : n56966;
  assign n56968 = pi12 ? n56935 : n56967;
  assign n56969 = pi11 ? n56908 : n56968;
  assign n56970 = pi21 ? n20563 : n15007;
  assign n56971 = pi20 ? n56970 : n4008;
  assign n56972 = pi19 ? n20563 : n56971;
  assign n56973 = pi18 ? n20563 : n56972;
  assign n56974 = pi17 ? n38984 : n56973;
  assign n56975 = pi16 ? n32 : n56974;
  assign n56976 = pi24 ? n20563 : n99;
  assign n56977 = pi23 ? n56976 : n139;
  assign n56978 = pi22 ? n56977 : n316;
  assign n56979 = pi21 ? n20563 : n56978;
  assign n56980 = pi20 ? n56979 : n12192;
  assign n56981 = pi19 ? n20563 : n56980;
  assign n56982 = pi18 ? n20563 : n56981;
  assign n56983 = pi17 ? n38984 : n56982;
  assign n56984 = pi16 ? n32 : n56983;
  assign n56985 = pi15 ? n56975 : n56984;
  assign n56986 = pi18 ? n38983 : n56456;
  assign n56987 = pi24 ? n20563 : n30868;
  assign n56988 = pi23 ? n56987 : n335;
  assign n56989 = pi22 ? n56988 : n204;
  assign n56990 = pi21 ? n20563 : n56989;
  assign n56991 = pi20 ? n56990 : n3340;
  assign n56992 = pi19 ? n50906 : n56991;
  assign n56993 = pi18 ? n20563 : n56992;
  assign n56994 = pi17 ? n56986 : n56993;
  assign n56995 = pi16 ? n32 : n56994;
  assign n56996 = pi21 ? n52252 : n32;
  assign n56997 = pi20 ? n56470 : n56996;
  assign n56998 = pi19 ? n50854 : n56997;
  assign n56999 = pi18 ? n20563 : n56998;
  assign n57000 = pi17 ? n40057 : n56999;
  assign n57001 = pi16 ? n32 : n57000;
  assign n57002 = pi15 ? n56995 : n57001;
  assign n57003 = pi14 ? n56985 : n57002;
  assign n57004 = pi17 ? n40057 : n56484;
  assign n57005 = pi16 ? n32 : n57004;
  assign n57006 = pi17 ? n40057 : n56494;
  assign n57007 = pi16 ? n32 : n57006;
  assign n57008 = pi15 ? n57005 : n57007;
  assign n57009 = pi20 ? n56498 : n1822;
  assign n57010 = pi19 ? n56489 : n57009;
  assign n57011 = pi18 ? n20563 : n57010;
  assign n57012 = pi17 ? n37958 : n57011;
  assign n57013 = pi16 ? n32 : n57012;
  assign n57014 = pi24 ? n363 : n36798;
  assign n57015 = pi23 ? n363 : n57014;
  assign n57016 = pi22 ? n57015 : n685;
  assign n57017 = pi21 ? n30868 : n57016;
  assign n57018 = pi20 ? n57017 : n32;
  assign n57019 = pi19 ? n47159 : n57018;
  assign n57020 = pi18 ? n20563 : n57019;
  assign n57021 = pi17 ? n37958 : n57020;
  assign n57022 = pi16 ? n32 : n57021;
  assign n57023 = pi15 ? n57013 : n57022;
  assign n57024 = pi14 ? n57008 : n57023;
  assign n57025 = pi13 ? n57003 : n57024;
  assign n57026 = pi17 ? n37958 : n56518;
  assign n57027 = pi16 ? n32 : n57026;
  assign n57028 = pi18 ? n51235 : n20563;
  assign n57029 = pi24 ? n36798 : n233;
  assign n57030 = pi23 ? n36798 : n57029;
  assign n57031 = pi22 ? n57030 : n317;
  assign n57032 = pi21 ? n36659 : n57031;
  assign n57033 = pi20 ? n57032 : n32;
  assign n57034 = pi19 ? n55487 : n57033;
  assign n57035 = pi18 ? n20563 : n57034;
  assign n57036 = pi17 ? n57028 : n57035;
  assign n57037 = pi16 ? n32 : n57036;
  assign n57038 = pi15 ? n57027 : n57037;
  assign n57039 = pi22 ? n45597 : n40386;
  assign n57040 = pi21 ? n32 : n57039;
  assign n57041 = pi20 ? n32 : n57040;
  assign n57042 = pi19 ? n32 : n57041;
  assign n57043 = pi21 ? n40917 : n39191;
  assign n57044 = pi22 ? n30195 : n39190;
  assign n57045 = pi21 ? n57044 : n45049;
  assign n57046 = pi20 ? n57043 : n57045;
  assign n57047 = pi19 ? n57046 : n20563;
  assign n57048 = pi18 ? n57042 : n57047;
  assign n57049 = pi17 ? n57048 : n56545;
  assign n57050 = pi16 ? n32 : n57049;
  assign n57051 = pi22 ? n49720 : n30868;
  assign n57052 = pi21 ? n32 : n57051;
  assign n57053 = pi20 ? n32 : n57052;
  assign n57054 = pi19 ? n32 : n57053;
  assign n57055 = pi18 ? n57054 : n30868;
  assign n57056 = pi17 ? n57055 : n56558;
  assign n57057 = pi16 ? n32 : n57056;
  assign n57058 = pi15 ? n57050 : n57057;
  assign n57059 = pi14 ? n57038 : n57058;
  assign n57060 = pi22 ? n51754 : n36615;
  assign n57061 = pi21 ? n32 : n57060;
  assign n57062 = pi20 ? n32 : n57061;
  assign n57063 = pi19 ? n32 : n57062;
  assign n57064 = pi21 ? n40960 : n52246;
  assign n57065 = pi22 ? n30195 : n42109;
  assign n57066 = pi21 ? n57065 : n56570;
  assign n57067 = pi20 ? n57064 : n57066;
  assign n57068 = pi19 ? n57067 : n56573;
  assign n57069 = pi18 ? n57063 : n57068;
  assign n57070 = pi21 ? n36781 : n37547;
  assign n57071 = pi20 ? n57070 : n32;
  assign n57072 = pi19 ? n50101 : n57071;
  assign n57073 = pi18 ? n56577 : n57072;
  assign n57074 = pi17 ? n57069 : n57073;
  assign n57075 = pi16 ? n32 : n57074;
  assign n57076 = pi21 ? n36798 : n33095;
  assign n57077 = pi20 ? n57076 : n32;
  assign n57078 = pi19 ? n20563 : n57077;
  assign n57079 = pi18 ? n20563 : n57078;
  assign n57080 = pi17 ? n38379 : n57079;
  assign n57081 = pi16 ? n32 : n57080;
  assign n57082 = pi15 ? n57075 : n57081;
  assign n57083 = pi17 ? n37336 : n55564;
  assign n57084 = pi16 ? n32 : n57083;
  assign n57085 = pi23 ? n20563 : n56987;
  assign n57086 = pi22 ? n20563 : n57085;
  assign n57087 = pi21 ? n20563 : n57086;
  assign n57088 = pi20 ? n20563 : n57087;
  assign n57089 = pi19 ? n57088 : n56588;
  assign n57090 = pi18 ? n20563 : n57089;
  assign n57091 = pi17 ? n38379 : n57090;
  assign n57092 = pi16 ? n32 : n57091;
  assign n57093 = pi15 ? n57084 : n57092;
  assign n57094 = pi14 ? n57082 : n57093;
  assign n57095 = pi13 ? n57059 : n57094;
  assign n57096 = pi12 ? n57025 : n57095;
  assign n57097 = pi22 ? n56665 : n32;
  assign n57098 = pi21 ? n55708 : n57097;
  assign n57099 = pi20 ? n57098 : n32;
  assign n57100 = pi19 ? n42915 : n57099;
  assign n57101 = pi18 ? n20563 : n57100;
  assign n57102 = pi17 ? n37336 : n57101;
  assign n57103 = pi16 ? n32 : n57102;
  assign n57104 = pi22 ? n49412 : n56607;
  assign n57105 = pi21 ? n57104 : n1009;
  assign n57106 = pi20 ? n57105 : n32;
  assign n57107 = pi19 ? n56605 : n57106;
  assign n57108 = pi18 ? n20563 : n57107;
  assign n57109 = pi17 ? n37336 : n57108;
  assign n57110 = pi16 ? n32 : n57109;
  assign n57111 = pi15 ? n57103 : n57110;
  assign n57112 = pi22 ? n53550 : n56622;
  assign n57113 = pi21 ? n57112 : n32;
  assign n57114 = pi20 ? n57113 : n32;
  assign n57115 = pi19 ? n56619 : n57114;
  assign n57116 = pi18 ? n20563 : n57115;
  assign n57117 = pi17 ? n39000 : n57116;
  assign n57118 = pi16 ? n32 : n57117;
  assign n57119 = pi22 ? n55622 : n54563;
  assign n57120 = pi21 ? n57119 : n32;
  assign n57121 = pi20 ? n57120 : n32;
  assign n57122 = pi19 ? n56631 : n57121;
  assign n57123 = pi18 ? n20563 : n57122;
  assign n57124 = pi17 ? n39000 : n57123;
  assign n57125 = pi16 ? n32 : n57124;
  assign n57126 = pi15 ? n57118 : n57125;
  assign n57127 = pi14 ? n57111 : n57126;
  assign n57128 = pi18 ? n51323 : n55617;
  assign n57129 = pi22 ? n54664 : n54563;
  assign n57130 = pi21 ? n57129 : n32;
  assign n57131 = pi20 ? n57130 : n32;
  assign n57132 = pi19 ? n56647 : n57131;
  assign n57133 = pi18 ? n55619 : n57132;
  assign n57134 = pi17 ? n57128 : n57133;
  assign n57135 = pi16 ? n32 : n57134;
  assign n57136 = pi18 ? n51323 : n30868;
  assign n57137 = pi21 ? n56810 : n32;
  assign n57138 = pi20 ? n57137 : n32;
  assign n57139 = pi19 ? n56663 : n57138;
  assign n57140 = pi18 ? n56661 : n57139;
  assign n57141 = pi17 ? n57136 : n57140;
  assign n57142 = pi16 ? n32 : n57141;
  assign n57143 = pi15 ? n57135 : n57142;
  assign n57144 = pi18 ? n46190 : n56674;
  assign n57145 = pi17 ? n57144 : n56683;
  assign n57146 = pi16 ? n32 : n57145;
  assign n57147 = pi19 ? n55656 : n56131;
  assign n57148 = pi18 ? n20563 : n57147;
  assign n57149 = pi17 ? n57028 : n57148;
  assign n57150 = pi16 ? n32 : n57149;
  assign n57151 = pi15 ? n57146 : n57150;
  assign n57152 = pi14 ? n57143 : n57151;
  assign n57153 = pi13 ? n57127 : n57152;
  assign n57154 = pi19 ? n56697 : n54566;
  assign n57155 = pi18 ? n30868 : n57154;
  assign n57156 = pi17 ? n46170 : n57155;
  assign n57157 = pi16 ? n32 : n57156;
  assign n57158 = pi17 ? n46170 : n56708;
  assign n57159 = pi16 ? n32 : n57158;
  assign n57160 = pi15 ? n57157 : n57159;
  assign n57161 = pi20 ? n32 : n52872;
  assign n57162 = pi19 ? n32 : n57161;
  assign n57163 = pi18 ? n57162 : n56720;
  assign n57164 = pi17 ? n57163 : n56728;
  assign n57165 = pi16 ? n32 : n57164;
  assign n57166 = pi18 ? n57162 : n43198;
  assign n57167 = pi17 ? n57166 : n56746;
  assign n57168 = pi16 ? n32 : n57167;
  assign n57169 = pi15 ? n57165 : n57168;
  assign n57170 = pi14 ? n57160 : n57169;
  assign n57171 = pi19 ? n32 : n54572;
  assign n57172 = pi18 ? n57171 : n56753;
  assign n57173 = pi17 ? n57172 : n56764;
  assign n57174 = pi16 ? n32 : n57173;
  assign n57175 = pi20 ? n36781 : n56772;
  assign n57176 = pi19 ? n57175 : n36781;
  assign n57177 = pi18 ? n57171 : n57176;
  assign n57178 = pi21 ? n5054 : n56778;
  assign n57179 = pi20 ? n36781 : n57178;
  assign n57180 = pi19 ? n57179 : n32;
  assign n57181 = pi18 ? n36781 : n57180;
  assign n57182 = pi17 ? n57177 : n57181;
  assign n57183 = pi16 ? n32 : n57182;
  assign n57184 = pi15 ? n57174 : n57183;
  assign n57185 = pi22 ? n36781 : n49406;
  assign n57186 = pi21 ? n57185 : n36781;
  assign n57187 = pi20 ? n36781 : n57186;
  assign n57188 = pi19 ? n57187 : n55779;
  assign n57189 = pi18 ? n46227 : n57188;
  assign n57190 = pi21 ? n55143 : n363;
  assign n57191 = pi20 ? n57190 : n56796;
  assign n57192 = pi19 ? n57191 : n32;
  assign n57193 = pi18 ? n55782 : n57192;
  assign n57194 = pi17 ? n57189 : n57193;
  assign n57195 = pi16 ? n32 : n57194;
  assign n57196 = pi18 ? n57171 : n55797;
  assign n57197 = pi23 ? n14626 : n51564;
  assign n57198 = pi22 ? n57197 : n32;
  assign n57199 = pi21 ? n43198 : n57198;
  assign n57200 = pi20 ? n36798 : n57199;
  assign n57201 = pi19 ? n57200 : n32;
  assign n57202 = pi18 ? n56809 : n57201;
  assign n57203 = pi17 ? n57196 : n57202;
  assign n57204 = pi16 ? n32 : n57203;
  assign n57205 = pi15 ? n57195 : n57204;
  assign n57206 = pi14 ? n57184 : n57205;
  assign n57207 = pi13 ? n57170 : n57206;
  assign n57208 = pi12 ? n57153 : n57207;
  assign n57209 = pi11 ? n57096 : n57208;
  assign n57210 = pi10 ? n56969 : n57209;
  assign n57211 = pi09 ? n56836 : n57210;
  assign n57212 = pi08 ? n56823 : n57211;
  assign n57213 = pi07 ? n56226 : n57212;
  assign n57214 = pi21 ? n297 : n10453;
  assign n57215 = pi20 ? n31220 : n57214;
  assign n57216 = pi19 ? n20563 : n57215;
  assign n57217 = pi18 ? n20563 : n57216;
  assign n57218 = pi17 ? n44247 : n57217;
  assign n57219 = pi16 ? n32 : n57218;
  assign n57220 = pi15 ? n32 : n57219;
  assign n57221 = pi20 ? n31220 : n11394;
  assign n57222 = pi19 ? n20563 : n57221;
  assign n57223 = pi18 ? n20563 : n57222;
  assign n57224 = pi17 ? n44247 : n57223;
  assign n57225 = pi16 ? n32 : n57224;
  assign n57226 = pi17 ? n43223 : n57223;
  assign n57227 = pi16 ? n32 : n57226;
  assign n57228 = pi15 ? n57225 : n57227;
  assign n57229 = pi14 ? n57220 : n57228;
  assign n57230 = pi13 ? n32 : n57229;
  assign n57231 = pi12 ? n32 : n57230;
  assign n57232 = pi11 ? n32 : n57231;
  assign n57233 = pi10 ? n32 : n57232;
  assign n57234 = pi21 ? n37 : n11015;
  assign n57235 = pi20 ? n20563 : n57234;
  assign n57236 = pi19 ? n20563 : n57235;
  assign n57237 = pi18 ? n20563 : n57236;
  assign n57238 = pi17 ? n43227 : n57237;
  assign n57239 = pi16 ? n32 : n57238;
  assign n57240 = pi21 ? n37 : n11026;
  assign n57241 = pi20 ? n20563 : n57240;
  assign n57242 = pi19 ? n20563 : n57241;
  assign n57243 = pi18 ? n20563 : n57242;
  assign n57244 = pi17 ? n44274 : n57243;
  assign n57245 = pi16 ? n32 : n57244;
  assign n57246 = pi15 ? n57239 : n57245;
  assign n57247 = pi21 ? n37 : n12404;
  assign n57248 = pi20 ? n20563 : n57247;
  assign n57249 = pi19 ? n20563 : n57248;
  assign n57250 = pi18 ? n20563 : n57249;
  assign n57251 = pi17 ? n43262 : n57250;
  assign n57252 = pi16 ? n32 : n57251;
  assign n57253 = pi21 ? n4938 : n7034;
  assign n57254 = pi20 ? n20563 : n57253;
  assign n57255 = pi19 ? n20563 : n57254;
  assign n57256 = pi18 ? n20563 : n57255;
  assign n57257 = pi17 ? n43262 : n57256;
  assign n57258 = pi16 ? n32 : n57257;
  assign n57259 = pi15 ? n57252 : n57258;
  assign n57260 = pi14 ? n57246 : n57259;
  assign n57261 = pi21 ? n11199 : n11569;
  assign n57262 = pi20 ? n31220 : n57261;
  assign n57263 = pi19 ? n20563 : n57262;
  assign n57264 = pi18 ? n20563 : n57263;
  assign n57265 = pi17 ? n43262 : n57264;
  assign n57266 = pi16 ? n32 : n57265;
  assign n57267 = pi21 ? n11199 : n17630;
  assign n57268 = pi20 ? n31220 : n57267;
  assign n57269 = pi19 ? n20563 : n57268;
  assign n57270 = pi18 ? n20563 : n57269;
  assign n57271 = pi17 ? n47593 : n57270;
  assign n57272 = pi16 ? n32 : n57271;
  assign n57273 = pi15 ? n57266 : n57272;
  assign n57274 = pi21 ? n11199 : n6406;
  assign n57275 = pi20 ? n31220 : n57274;
  assign n57276 = pi19 ? n20563 : n57275;
  assign n57277 = pi18 ? n20563 : n57276;
  assign n57278 = pi17 ? n42207 : n57277;
  assign n57279 = pi16 ? n32 : n57278;
  assign n57280 = pi21 ? n22842 : n20889;
  assign n57281 = pi20 ? n31266 : n57280;
  assign n57282 = pi19 ? n20563 : n57281;
  assign n57283 = pi18 ? n20563 : n57282;
  assign n57284 = pi17 ? n42688 : n57283;
  assign n57285 = pi16 ? n32 : n57284;
  assign n57286 = pi15 ? n57279 : n57285;
  assign n57287 = pi14 ? n57273 : n57286;
  assign n57288 = pi13 ? n57260 : n57287;
  assign n57289 = pi21 ? n22842 : n1512;
  assign n57290 = pi20 ? n31220 : n57289;
  assign n57291 = pi19 ? n20563 : n57290;
  assign n57292 = pi18 ? n20563 : n57291;
  assign n57293 = pi17 ? n42688 : n57292;
  assign n57294 = pi16 ? n32 : n57293;
  assign n57295 = pi21 ? n11208 : n16358;
  assign n57296 = pi20 ? n31220 : n57295;
  assign n57297 = pi19 ? n20563 : n57296;
  assign n57298 = pi18 ? n20563 : n57297;
  assign n57299 = pi17 ? n40024 : n57298;
  assign n57300 = pi16 ? n32 : n57299;
  assign n57301 = pi15 ? n57294 : n57300;
  assign n57302 = pi21 ? n11208 : n2565;
  assign n57303 = pi20 ? n31220 : n57302;
  assign n57304 = pi19 ? n20563 : n57303;
  assign n57305 = pi18 ? n20563 : n57304;
  assign n57306 = pi17 ? n40024 : n57305;
  assign n57307 = pi16 ? n32 : n57306;
  assign n57308 = pi21 ? n11208 : n2578;
  assign n57309 = pi20 ? n31220 : n57308;
  assign n57310 = pi19 ? n20563 : n57309;
  assign n57311 = pi18 ? n20563 : n57310;
  assign n57312 = pi17 ? n41182 : n57311;
  assign n57313 = pi16 ? n32 : n57312;
  assign n57314 = pi15 ? n57307 : n57313;
  assign n57315 = pi14 ? n57301 : n57314;
  assign n57316 = pi21 ? n17806 : n760;
  assign n57317 = pi20 ? n20563 : n57316;
  assign n57318 = pi19 ? n20563 : n57317;
  assign n57319 = pi18 ? n20563 : n57318;
  assign n57320 = pi17 ? n42240 : n57319;
  assign n57321 = pi16 ? n32 : n57320;
  assign n57322 = pi20 ? n31220 : n57316;
  assign n57323 = pi19 ? n20563 : n57322;
  assign n57324 = pi18 ? n20563 : n57323;
  assign n57325 = pi17 ? n40498 : n57324;
  assign n57326 = pi16 ? n32 : n57325;
  assign n57327 = pi15 ? n57321 : n57326;
  assign n57328 = pi14 ? n57327 : n57326;
  assign n57329 = pi13 ? n57315 : n57328;
  assign n57330 = pi12 ? n57288 : n57329;
  assign n57331 = pi21 ? n52795 : n5829;
  assign n57332 = pi20 ? n54354 : n57331;
  assign n57333 = pi19 ? n20563 : n57332;
  assign n57334 = pi18 ? n20563 : n57333;
  assign n57335 = pi17 ? n40498 : n57334;
  assign n57336 = pi16 ? n32 : n57335;
  assign n57337 = pi20 ? n54354 : n8644;
  assign n57338 = pi19 ? n20563 : n57337;
  assign n57339 = pi18 ? n20563 : n57338;
  assign n57340 = pi17 ? n41683 : n57339;
  assign n57341 = pi16 ? n32 : n57340;
  assign n57342 = pi15 ? n57336 : n57341;
  assign n57343 = pi21 ? n20563 : n55969;
  assign n57344 = pi20 ? n57343 : n8644;
  assign n57345 = pi19 ? n20563 : n57344;
  assign n57346 = pi18 ? n20563 : n57345;
  assign n57347 = pi17 ? n40511 : n57346;
  assign n57348 = pi16 ? n32 : n57347;
  assign n57349 = pi23 ? n8160 : n316;
  assign n57350 = pi22 ? n57349 : n316;
  assign n57351 = pi21 ? n57350 : n928;
  assign n57352 = pi20 ? n56350 : n57351;
  assign n57353 = pi19 ? n20563 : n57352;
  assign n57354 = pi18 ? n20563 : n57353;
  assign n57355 = pi17 ? n40511 : n57354;
  assign n57356 = pi16 ? n32 : n57355;
  assign n57357 = pi15 ? n57348 : n57356;
  assign n57358 = pi14 ? n57342 : n57357;
  assign n57359 = pi17 ? n39374 : n57354;
  assign n57360 = pi16 ? n32 : n57359;
  assign n57361 = pi20 ? n56361 : n980;
  assign n57362 = pi19 ? n20563 : n57361;
  assign n57363 = pi18 ? n20563 : n57362;
  assign n57364 = pi17 ? n39374 : n57363;
  assign n57365 = pi16 ? n32 : n57364;
  assign n57366 = pi15 ? n57360 : n57365;
  assign n57367 = pi20 ? n3299 : n980;
  assign n57368 = pi19 ? n20563 : n57367;
  assign n57369 = pi18 ? n20563 : n57368;
  assign n57370 = pi17 ? n39374 : n57369;
  assign n57371 = pi16 ? n32 : n57370;
  assign n57372 = pi20 ? n6402 : n1010;
  assign n57373 = pi19 ? n20563 : n57372;
  assign n57374 = pi18 ? n20563 : n57373;
  assign n57375 = pi17 ? n40533 : n57374;
  assign n57376 = pi16 ? n32 : n57375;
  assign n57377 = pi15 ? n57371 : n57376;
  assign n57378 = pi14 ? n57366 : n57377;
  assign n57379 = pi13 ? n57358 : n57378;
  assign n57380 = pi23 ? n20563 : n363;
  assign n57381 = pi22 ? n37 : n57380;
  assign n57382 = pi21 ? n20563 : n57381;
  assign n57383 = pi20 ? n57382 : n1010;
  assign n57384 = pi19 ? n20563 : n57383;
  assign n57385 = pi18 ? n20563 : n57384;
  assign n57386 = pi17 ? n41709 : n57385;
  assign n57387 = pi16 ? n32 : n57386;
  assign n57388 = pi20 ? n55343 : n1010;
  assign n57389 = pi19 ? n20563 : n57388;
  assign n57390 = pi18 ? n20563 : n57389;
  assign n57391 = pi17 ? n41709 : n57390;
  assign n57392 = pi16 ? n32 : n57391;
  assign n57393 = pi15 ? n57387 : n57392;
  assign n57394 = pi23 ? n139 : n36798;
  assign n57395 = pi22 ? n37 : n57394;
  assign n57396 = pi21 ? n37 : n57395;
  assign n57397 = pi22 ? n13481 : n6415;
  assign n57398 = pi21 ? n57397 : n32;
  assign n57399 = pi20 ? n57396 : n57398;
  assign n57400 = pi19 ? n20563 : n57399;
  assign n57401 = pi18 ? n20563 : n57400;
  assign n57402 = pi17 ? n38949 : n57401;
  assign n57403 = pi16 ? n32 : n57402;
  assign n57404 = pi21 ? n37 : n7195;
  assign n57405 = pi20 ? n57404 : n44443;
  assign n57406 = pi19 ? n20563 : n57405;
  assign n57407 = pi18 ? n20563 : n57406;
  assign n57408 = pi17 ? n38949 : n57407;
  assign n57409 = pi16 ? n32 : n57408;
  assign n57410 = pi15 ? n57403 : n57409;
  assign n57411 = pi14 ? n57393 : n57410;
  assign n57412 = pi20 ? n31410 : n16519;
  assign n57413 = pi19 ? n31221 : n57412;
  assign n57414 = pi18 ? n20563 : n57413;
  assign n57415 = pi17 ? n38949 : n57414;
  assign n57416 = pi16 ? n32 : n57415;
  assign n57417 = pi20 ? n31410 : n8917;
  assign n57418 = pi19 ? n31221 : n57417;
  assign n57419 = pi18 ? n20563 : n57418;
  assign n57420 = pi17 ? n38958 : n57419;
  assign n57421 = pi16 ? n32 : n57420;
  assign n57422 = pi15 ? n57416 : n57421;
  assign n57423 = pi22 ? n20563 : n5782;
  assign n57424 = pi21 ? n20563 : n57423;
  assign n57425 = pi21 ? n56554 : n32;
  assign n57426 = pi20 ? n57424 : n57425;
  assign n57427 = pi19 ? n20563 : n57426;
  assign n57428 = pi18 ? n20563 : n57427;
  assign n57429 = pi17 ? n38958 : n57428;
  assign n57430 = pi16 ? n32 : n57429;
  assign n57431 = pi22 ? n99 : n51564;
  assign n57432 = pi21 ? n20563 : n57431;
  assign n57433 = pi22 ? n51564 : n688;
  assign n57434 = pi21 ? n57433 : n32;
  assign n57435 = pi20 ? n57432 : n57434;
  assign n57436 = pi19 ? n20563 : n57435;
  assign n57437 = pi18 ? n20563 : n57436;
  assign n57438 = pi17 ? n38958 : n57437;
  assign n57439 = pi16 ? n32 : n57438;
  assign n57440 = pi15 ? n57430 : n57439;
  assign n57441 = pi14 ? n57422 : n57440;
  assign n57442 = pi13 ? n57411 : n57441;
  assign n57443 = pi12 ? n57379 : n57442;
  assign n57444 = pi11 ? n57330 : n57443;
  assign n57445 = pi17 ? n45393 : n56444;
  assign n57446 = pi16 ? n32 : n57445;
  assign n57447 = pi22 ? n56977 : n13481;
  assign n57448 = pi21 ? n20563 : n57447;
  assign n57449 = pi20 ? n57448 : n56130;
  assign n57450 = pi19 ? n20563 : n57449;
  assign n57451 = pi18 ? n20563 : n57450;
  assign n57452 = pi17 ? n45393 : n57451;
  assign n57453 = pi16 ? n32 : n57452;
  assign n57454 = pi15 ? n57446 : n57453;
  assign n57455 = pi22 ? n56468 : n204;
  assign n57456 = pi21 ? n20563 : n57455;
  assign n57457 = pi23 ? n14626 : n395;
  assign n57458 = pi22 ? n57457 : n32;
  assign n57459 = pi21 ? n57458 : n32;
  assign n57460 = pi20 ? n57456 : n57459;
  assign n57461 = pi19 ? n20563 : n57460;
  assign n57462 = pi18 ? n20563 : n57461;
  assign n57463 = pi17 ? n45393 : n57462;
  assign n57464 = pi16 ? n32 : n57463;
  assign n57465 = pi24 ? n30868 : n139;
  assign n57466 = pi23 ? n57465 : n335;
  assign n57467 = pi22 ? n57466 : n233;
  assign n57468 = pi21 ? n36249 : n57467;
  assign n57469 = pi20 ? n57468 : n56996;
  assign n57470 = pi19 ? n20563 : n57469;
  assign n57471 = pi18 ? n20563 : n57470;
  assign n57472 = pi17 ? n45414 : n57471;
  assign n57473 = pi16 ? n32 : n57472;
  assign n57474 = pi15 ? n57464 : n57473;
  assign n57475 = pi14 ? n57454 : n57474;
  assign n57476 = pi21 ? n36249 : n233;
  assign n57477 = pi20 ? n57476 : n2653;
  assign n57478 = pi19 ? n20563 : n57477;
  assign n57479 = pi18 ? n20563 : n57478;
  assign n57480 = pi17 ? n45414 : n57479;
  assign n57481 = pi16 ? n32 : n57480;
  assign n57482 = pi23 ? n8184 : n363;
  assign n57483 = pi22 ? n57482 : n685;
  assign n57484 = pi21 ? n56487 : n57483;
  assign n57485 = pi20 ? n57484 : n37640;
  assign n57486 = pi19 ? n20563 : n57485;
  assign n57487 = pi18 ? n20563 : n57486;
  assign n57488 = pi17 ? n45414 : n57487;
  assign n57489 = pi16 ? n32 : n57488;
  assign n57490 = pi15 ? n57481 : n57489;
  assign n57491 = pi22 ? n37 : n37173;
  assign n57492 = pi23 ? n19714 : n157;
  assign n57493 = pi22 ? n57492 : n51564;
  assign n57494 = pi21 ? n57491 : n57493;
  assign n57495 = pi20 ? n57494 : n37640;
  assign n57496 = pi19 ? n20563 : n57495;
  assign n57497 = pi18 ? n20563 : n57496;
  assign n57498 = pi17 ? n38330 : n57497;
  assign n57499 = pi16 ? n32 : n57498;
  assign n57500 = pi22 ? n37 : n33792;
  assign n57501 = pi23 ? n36781 : n57014;
  assign n57502 = pi22 ? n57501 : n316;
  assign n57503 = pi21 ? n57500 : n57502;
  assign n57504 = pi20 ? n57503 : n32;
  assign n57505 = pi19 ? n20563 : n57504;
  assign n57506 = pi18 ? n20563 : n57505;
  assign n57507 = pi17 ? n38330 : n57506;
  assign n57508 = pi16 ? n32 : n57507;
  assign n57509 = pi15 ? n57499 : n57508;
  assign n57510 = pi14 ? n57490 : n57509;
  assign n57511 = pi13 ? n57475 : n57510;
  assign n57512 = pi20 ? n43935 : n40791;
  assign n57513 = pi20 ? n40791 : n20563;
  assign n57514 = pi19 ? n57512 : n57513;
  assign n57515 = pi18 ? n32 : n57514;
  assign n57516 = pi22 ? n99 : n56616;
  assign n57517 = pi24 ? n36798 : n204;
  assign n57518 = pi23 ? n36798 : n57517;
  assign n57519 = pi22 ? n57518 : n13481;
  assign n57520 = pi21 ? n57516 : n57519;
  assign n57521 = pi20 ? n57520 : n32;
  assign n57522 = pi19 ? n20563 : n57521;
  assign n57523 = pi18 ? n52168 : n57522;
  assign n57524 = pi17 ? n57515 : n57523;
  assign n57525 = pi16 ? n32 : n57524;
  assign n57526 = pi22 ? n39190 : n56533;
  assign n57527 = pi21 ? n20563 : n57526;
  assign n57528 = pi20 ? n54998 : n57527;
  assign n57529 = pi19 ? n57528 : n20563;
  assign n57530 = pi18 ? n32 : n57529;
  assign n57531 = pi22 ? n99 : n36659;
  assign n57532 = pi22 ? n57030 : n13481;
  assign n57533 = pi21 ? n57531 : n57532;
  assign n57534 = pi20 ? n57533 : n32;
  assign n57535 = pi19 ? n20563 : n57534;
  assign n57536 = pi18 ? n20563 : n57535;
  assign n57537 = pi17 ? n57530 : n57536;
  assign n57538 = pi16 ? n32 : n57537;
  assign n57539 = pi15 ? n57525 : n57538;
  assign n57540 = pi21 ? n20563 : n55536;
  assign n57541 = pi20 ? n55014 : n57540;
  assign n57542 = pi19 ? n57541 : n20563;
  assign n57543 = pi18 ? n32 : n57542;
  assign n57544 = pi19 ? n20563 : n56543;
  assign n57545 = pi18 ? n20563 : n57544;
  assign n57546 = pi17 ? n57543 : n57545;
  assign n57547 = pi16 ? n32 : n57546;
  assign n57548 = pi22 ? n37173 : n56568;
  assign n57549 = pi21 ? n20563 : n57548;
  assign n57550 = pi20 ? n55014 : n57549;
  assign n57551 = pi19 ? n57550 : n20563;
  assign n57552 = pi18 ? n32 : n57551;
  assign n57553 = pi22 ? n139 : n36781;
  assign n57554 = pi21 ? n57553 : n56554;
  assign n57555 = pi20 ? n57554 : n32;
  assign n57556 = pi19 ? n20563 : n57555;
  assign n57557 = pi18 ? n20563 : n57556;
  assign n57558 = pi17 ? n57552 : n57557;
  assign n57559 = pi16 ? n32 : n57558;
  assign n57560 = pi15 ? n57547 : n57559;
  assign n57561 = pi14 ? n57539 : n57560;
  assign n57562 = pi22 ? n335 : n36798;
  assign n57563 = pi22 ? n51564 : n14363;
  assign n57564 = pi21 ? n57562 : n57563;
  assign n57565 = pi20 ? n57564 : n32;
  assign n57566 = pi19 ? n20563 : n57565;
  assign n57567 = pi18 ? n20563 : n57566;
  assign n57568 = pi17 ? n37936 : n57567;
  assign n57569 = pi16 ? n32 : n57568;
  assign n57570 = pi22 ? n363 : n49412;
  assign n57571 = pi21 ? n57570 : n33095;
  assign n57572 = pi20 ? n57571 : n32;
  assign n57573 = pi19 ? n56489 : n57572;
  assign n57574 = pi18 ? n20563 : n57573;
  assign n57575 = pi17 ? n37936 : n57574;
  assign n57576 = pi16 ? n32 : n57575;
  assign n57577 = pi15 ? n57569 : n57576;
  assign n57578 = pi21 ? n20563 : n297;
  assign n57579 = pi20 ? n20563 : n57578;
  assign n57580 = pi22 ? n157 : n43198;
  assign n57581 = pi21 ? n57580 : n55560;
  assign n57582 = pi20 ? n57581 : n32;
  assign n57583 = pi19 ? n57579 : n57582;
  assign n57584 = pi18 ? n20563 : n57583;
  assign n57585 = pi17 ? n40057 : n57584;
  assign n57586 = pi16 ? n32 : n57585;
  assign n57587 = pi22 ? n37 : n57085;
  assign n57588 = pi21 ? n20563 : n57587;
  assign n57589 = pi20 ? n20563 : n57588;
  assign n57590 = pi21 ? n14626 : n57097;
  assign n57591 = pi20 ? n57590 : n32;
  assign n57592 = pi19 ? n57589 : n57591;
  assign n57593 = pi18 ? n20563 : n57592;
  assign n57594 = pi17 ? n40057 : n57593;
  assign n57595 = pi16 ? n32 : n57594;
  assign n57596 = pi15 ? n57586 : n57595;
  assign n57597 = pi14 ? n57577 : n57596;
  assign n57598 = pi13 ? n57561 : n57597;
  assign n57599 = pi12 ? n57511 : n57598;
  assign n57600 = pi22 ? n233 : n14626;
  assign n57601 = pi21 ? n57600 : n57097;
  assign n57602 = pi20 ? n57601 : n32;
  assign n57603 = pi19 ? n47159 : n57602;
  assign n57604 = pi18 ? n20563 : n57603;
  assign n57605 = pi17 ? n40057 : n57604;
  assign n57606 = pi16 ? n32 : n57605;
  assign n57607 = pi21 ? n51564 : n20952;
  assign n57608 = pi20 ? n57607 : n32;
  assign n57609 = pi19 ? n56631 : n57608;
  assign n57610 = pi18 ? n20563 : n57609;
  assign n57611 = pi17 ? n38984 : n57610;
  assign n57612 = pi16 ? n32 : n57611;
  assign n57613 = pi15 ? n57606 : n57612;
  assign n57614 = pi21 ? n20563 : n57553;
  assign n57615 = pi20 ? n20563 : n57614;
  assign n57616 = pi22 ? n685 : n13481;
  assign n57617 = pi21 ? n57616 : n32;
  assign n57618 = pi20 ? n57617 : n32;
  assign n57619 = pi19 ? n57615 : n57618;
  assign n57620 = pi18 ? n20563 : n57619;
  assign n57621 = pi17 ? n38984 : n57620;
  assign n57622 = pi16 ? n32 : n57621;
  assign n57623 = pi20 ? n47801 : n38754;
  assign n57624 = pi19 ? n50091 : n57623;
  assign n57625 = pi18 ? n37928 : n57624;
  assign n57626 = pi20 ? n40918 : n40791;
  assign n57627 = pi21 ? n40917 : n48173;
  assign n57628 = pi20 ? n57627 : n39801;
  assign n57629 = pi19 ? n57626 : n57628;
  assign n57630 = pi21 ? n20563 : n36781;
  assign n57631 = pi20 ? n43010 : n57630;
  assign n57632 = pi23 ? n36798 : n685;
  assign n57633 = pi22 ? n57632 : n56665;
  assign n57634 = pi21 ? n57633 : n32;
  assign n57635 = pi20 ? n57634 : n32;
  assign n57636 = pi19 ? n57631 : n57635;
  assign n57637 = pi18 ? n57629 : n57636;
  assign n57638 = pi17 ? n57625 : n57637;
  assign n57639 = pi16 ? n32 : n57638;
  assign n57640 = pi15 ? n57622 : n57639;
  assign n57641 = pi14 ? n57613 : n57640;
  assign n57642 = pi20 ? n42006 : n30868;
  assign n57643 = pi19 ? n57642 : n30868;
  assign n57644 = pi18 ? n37928 : n57643;
  assign n57645 = pi21 ? n30868 : n57562;
  assign n57646 = pi20 ? n20563 : n57645;
  assign n57647 = pi23 ? n51564 : n14362;
  assign n57648 = pi22 ? n316 : n57647;
  assign n57649 = pi21 ? n57648 : n32;
  assign n57650 = pi20 ? n57649 : n32;
  assign n57651 = pi19 ? n57646 : n57650;
  assign n57652 = pi18 ? n55521 : n57651;
  assign n57653 = pi17 ? n57644 : n57652;
  assign n57654 = pi16 ? n32 : n57653;
  assign n57655 = pi19 ? n51301 : n30868;
  assign n57656 = pi18 ? n51823 : n57655;
  assign n57657 = pi21 ? n30868 : n53432;
  assign n57658 = pi20 ? n20563 : n57657;
  assign n57659 = pi23 ? n233 : n13481;
  assign n57660 = pi22 ? n57659 : n21502;
  assign n57661 = pi21 ? n57660 : n32;
  assign n57662 = pi20 ? n57661 : n32;
  assign n57663 = pi19 ? n57658 : n57662;
  assign n57664 = pi18 ? n55521 : n57663;
  assign n57665 = pi17 ? n57656 : n57664;
  assign n57666 = pi16 ? n32 : n57665;
  assign n57667 = pi15 ? n57654 : n57666;
  assign n57668 = pi20 ? n54417 : n43010;
  assign n57669 = pi19 ? n57668 : n20563;
  assign n57670 = pi18 ? n32 : n57669;
  assign n57671 = pi22 ? n36781 : n233;
  assign n57672 = pi21 ? n36659 : n57671;
  assign n57673 = pi20 ? n20563 : n57672;
  assign n57674 = pi23 ? n685 : n13481;
  assign n57675 = pi22 ? n57674 : n21502;
  assign n57676 = pi21 ? n57675 : n32;
  assign n57677 = pi20 ? n57676 : n32;
  assign n57678 = pi19 ? n57673 : n57677;
  assign n57679 = pi18 ? n40793 : n57678;
  assign n57680 = pi17 ? n57670 : n57679;
  assign n57681 = pi16 ? n32 : n57680;
  assign n57682 = pi20 ? n31313 : n38754;
  assign n57683 = pi20 ? n50735 : n43935;
  assign n57684 = pi19 ? n57682 : n57683;
  assign n57685 = pi18 ? n32 : n57684;
  assign n57686 = pi22 ? n57674 : n14363;
  assign n57687 = pi21 ? n57686 : n32;
  assign n57688 = pi20 ? n57687 : n32;
  assign n57689 = pi19 ? n57673 : n57688;
  assign n57690 = pi18 ? n20563 : n57689;
  assign n57691 = pi17 ? n57685 : n57690;
  assign n57692 = pi16 ? n32 : n57691;
  assign n57693 = pi15 ? n57681 : n57692;
  assign n57694 = pi14 ? n57667 : n57693;
  assign n57695 = pi13 ? n57641 : n57694;
  assign n57696 = pi19 ? n49218 : n30868;
  assign n57697 = pi18 ? n32 : n57696;
  assign n57698 = pi22 ? n36798 : n685;
  assign n57699 = pi21 ? n36781 : n57698;
  assign n57700 = pi20 ? n30868 : n57699;
  assign n57701 = pi19 ? n57700 : n52867;
  assign n57702 = pi18 ? n30868 : n57701;
  assign n57703 = pi17 ? n57697 : n57702;
  assign n57704 = pi16 ? n32 : n57703;
  assign n57705 = pi22 ? n45160 : n36781;
  assign n57706 = pi21 ? n57705 : n47396;
  assign n57707 = pi20 ? n57706 : n55701;
  assign n57708 = pi19 ? n57707 : n56722;
  assign n57709 = pi18 ? n32 : n57708;
  assign n57710 = pi20 ? n36798 : n38923;
  assign n57711 = pi19 ? n57710 : n56808;
  assign n57712 = pi21 ? n36781 : n43198;
  assign n57713 = pi22 ? n204 : n51564;
  assign n57714 = pi21 ? n36781 : n57713;
  assign n57715 = pi20 ? n57712 : n57714;
  assign n57716 = pi21 ? n57097 : n32;
  assign n57717 = pi20 ? n57716 : n32;
  assign n57718 = pi19 ? n57715 : n57717;
  assign n57719 = pi18 ? n57711 : n57718;
  assign n57720 = pi17 ? n57709 : n57719;
  assign n57721 = pi16 ? n32 : n57720;
  assign n57722 = pi15 ? n57704 : n57721;
  assign n57723 = pi22 ? n46789 : n49412;
  assign n57724 = pi21 ? n57723 : n43198;
  assign n57725 = pi20 ? n57724 : n43198;
  assign n57726 = pi20 ? n52447 : n56717;
  assign n57727 = pi19 ? n57725 : n57726;
  assign n57728 = pi18 ? n32 : n57727;
  assign n57729 = pi21 ? n53484 : n47397;
  assign n57730 = pi20 ? n43198 : n57729;
  assign n57731 = pi19 ? n43198 : n57730;
  assign n57732 = pi21 ? n36798 : n53484;
  assign n57733 = pi22 ? n43198 : n316;
  assign n57734 = pi21 ? n43198 : n57733;
  assign n57735 = pi20 ? n57732 : n57734;
  assign n57736 = pi19 ? n57735 : n35482;
  assign n57737 = pi18 ? n57731 : n57736;
  assign n57738 = pi17 ? n57728 : n57737;
  assign n57739 = pi16 ? n32 : n57738;
  assign n57740 = pi21 ? n47341 : n47396;
  assign n57741 = pi20 ? n57740 : n54009;
  assign n57742 = pi19 ? n57741 : n43198;
  assign n57743 = pi18 ? n32 : n57742;
  assign n57744 = pi20 ? n55701 : n43198;
  assign n57745 = pi19 ? n43198 : n57744;
  assign n57746 = pi22 ? n14626 : n13481;
  assign n57747 = pi21 ? n43198 : n57746;
  assign n57748 = pi20 ? n49369 : n57747;
  assign n57749 = pi19 ? n57748 : n35482;
  assign n57750 = pi18 ? n57745 : n57749;
  assign n57751 = pi17 ? n57743 : n57750;
  assign n57752 = pi16 ? n32 : n57751;
  assign n57753 = pi15 ? n57739 : n57752;
  assign n57754 = pi14 ? n57722 : n57753;
  assign n57755 = pi22 ? n46275 : n53550;
  assign n57756 = pi21 ? n57755 : n55125;
  assign n57757 = pi20 ? n57756 : n43198;
  assign n57758 = pi19 ? n57757 : n43198;
  assign n57759 = pi18 ? n32 : n57758;
  assign n57760 = pi22 ? n51564 : n13481;
  assign n57761 = pi21 ? n43198 : n57760;
  assign n57762 = pi20 ? n51356 : n57761;
  assign n57763 = pi19 ? n57762 : n32;
  assign n57764 = pi18 ? n43198 : n57763;
  assign n57765 = pi17 ? n57759 : n57764;
  assign n57766 = pi16 ? n32 : n57765;
  assign n57767 = pi22 ? n32 : n49406;
  assign n57768 = pi21 ? n57767 : n36781;
  assign n57769 = pi20 ? n57768 : n36781;
  assign n57770 = pi21 ? n54617 : n36781;
  assign n57771 = pi20 ? n57770 : n36781;
  assign n57772 = pi19 ? n57769 : n57771;
  assign n57773 = pi18 ? n32 : n57772;
  assign n57774 = pi22 ? n36781 : n14626;
  assign n57775 = pi21 ? n57774 : n57760;
  assign n57776 = pi20 ? n36781 : n57775;
  assign n57777 = pi19 ? n57776 : n32;
  assign n57778 = pi18 ? n36781 : n57777;
  assign n57779 = pi17 ? n57773 : n57778;
  assign n57780 = pi16 ? n32 : n57779;
  assign n57781 = pi15 ? n57766 : n57780;
  assign n57782 = pi23 ? n56620 : n36798;
  assign n57783 = pi22 ? n36781 : n57782;
  assign n57784 = pi21 ? n45211 : n57783;
  assign n57785 = pi21 ? n36781 : n39972;
  assign n57786 = pi20 ? n57784 : n57785;
  assign n57787 = pi21 ? n49858 : n36781;
  assign n57788 = pi20 ? n57787 : n36781;
  assign n57789 = pi19 ? n57786 : n57788;
  assign n57790 = pi18 ? n32 : n57789;
  assign n57791 = pi21 ? n56695 : n55560;
  assign n57792 = pi20 ? n36781 : n57791;
  assign n57793 = pi19 ? n57792 : n32;
  assign n57794 = pi18 ? n36781 : n57793;
  assign n57795 = pi17 ? n57790 : n57794;
  assign n57796 = pi16 ? n32 : n57795;
  assign n57797 = pi20 ? n50768 : n55701;
  assign n57798 = pi19 ? n57797 : n56808;
  assign n57799 = pi18 ? n32 : n57798;
  assign n57800 = pi22 ? n36798 : n53930;
  assign n57801 = pi21 ? n57800 : n55560;
  assign n57802 = pi20 ? n36798 : n57801;
  assign n57803 = pi19 ? n57802 : n32;
  assign n57804 = pi18 ? n36798 : n57803;
  assign n57805 = pi17 ? n57799 : n57804;
  assign n57806 = pi16 ? n32 : n57805;
  assign n57807 = pi15 ? n57796 : n57806;
  assign n57808 = pi14 ? n57781 : n57807;
  assign n57809 = pi13 ? n57754 : n57808;
  assign n57810 = pi12 ? n57695 : n57809;
  assign n57811 = pi11 ? n57599 : n57810;
  assign n57812 = pi10 ? n57444 : n57811;
  assign n57813 = pi09 ? n57233 : n57812;
  assign n57814 = pi17 ? n44670 : n57217;
  assign n57815 = pi16 ? n32 : n57814;
  assign n57816 = pi15 ? n32 : n57815;
  assign n57817 = pi17 ? n44670 : n57223;
  assign n57818 = pi16 ? n32 : n57817;
  assign n57819 = pi17 ? n43684 : n57223;
  assign n57820 = pi16 ? n32 : n57819;
  assign n57821 = pi15 ? n57818 : n57820;
  assign n57822 = pi14 ? n57816 : n57821;
  assign n57823 = pi13 ? n32 : n57822;
  assign n57824 = pi12 ? n32 : n57823;
  assign n57825 = pi11 ? n32 : n57824;
  assign n57826 = pi10 ? n32 : n57825;
  assign n57827 = pi17 ? n43218 : n57237;
  assign n57828 = pi16 ? n32 : n57827;
  assign n57829 = pi17 ? n44247 : n57243;
  assign n57830 = pi16 ? n32 : n57829;
  assign n57831 = pi15 ? n57828 : n57830;
  assign n57832 = pi17 ? n48624 : n57250;
  assign n57833 = pi16 ? n32 : n57832;
  assign n57834 = pi21 ? n4938 : n650;
  assign n57835 = pi20 ? n20563 : n57834;
  assign n57836 = pi19 ? n20563 : n57835;
  assign n57837 = pi18 ? n20563 : n57836;
  assign n57838 = pi17 ? n48624 : n57837;
  assign n57839 = pi16 ? n32 : n57838;
  assign n57840 = pi15 ? n57833 : n57839;
  assign n57841 = pi14 ? n57831 : n57840;
  assign n57842 = pi21 ? n11199 : n5771;
  assign n57843 = pi20 ? n31220 : n57842;
  assign n57844 = pi19 ? n20563 : n57843;
  assign n57845 = pi18 ? n20563 : n57844;
  assign n57846 = pi17 ? n42645 : n57845;
  assign n57847 = pi16 ? n32 : n57846;
  assign n57848 = pi17 ? n42655 : n57845;
  assign n57849 = pi16 ? n32 : n57848;
  assign n57850 = pi15 ? n57847 : n57849;
  assign n57851 = pi21 ? n11199 : n21387;
  assign n57852 = pi20 ? n31220 : n57851;
  assign n57853 = pi19 ? n20563 : n57852;
  assign n57854 = pi18 ? n20563 : n57853;
  assign n57855 = pi17 ? n42681 : n57854;
  assign n57856 = pi16 ? n32 : n57855;
  assign n57857 = pi21 ? n22842 : n21387;
  assign n57858 = pi20 ? n31266 : n57857;
  assign n57859 = pi19 ? n20563 : n57858;
  assign n57860 = pi18 ? n20563 : n57859;
  assign n57861 = pi17 ? n43262 : n57860;
  assign n57862 = pi16 ? n32 : n57861;
  assign n57863 = pi15 ? n57856 : n57862;
  assign n57864 = pi14 ? n57850 : n57863;
  assign n57865 = pi13 ? n57841 : n57864;
  assign n57866 = pi22 ? n13278 : n685;
  assign n57867 = pi21 ? n57866 : n1485;
  assign n57868 = pi20 ? n31220 : n57867;
  assign n57869 = pi19 ? n20563 : n57868;
  assign n57870 = pi18 ? n20563 : n57869;
  assign n57871 = pi17 ? n43262 : n57870;
  assign n57872 = pi16 ? n32 : n57871;
  assign n57873 = pi23 ? n204 : n5630;
  assign n57874 = pi22 ? n57873 : n32;
  assign n57875 = pi21 ? n11208 : n57874;
  assign n57876 = pi20 ? n31220 : n57875;
  assign n57877 = pi19 ? n20563 : n57876;
  assign n57878 = pi18 ? n20563 : n57877;
  assign n57879 = pi17 ? n42688 : n57878;
  assign n57880 = pi16 ? n32 : n57879;
  assign n57881 = pi15 ? n57872 : n57880;
  assign n57882 = pi23 ? n1432 : n363;
  assign n57883 = pi22 ? n57882 : n685;
  assign n57884 = pi21 ? n57883 : n57874;
  assign n57885 = pi20 ? n31220 : n57884;
  assign n57886 = pi19 ? n20563 : n57885;
  assign n57887 = pi18 ? n20563 : n57886;
  assign n57888 = pi17 ? n42688 : n57887;
  assign n57889 = pi16 ? n32 : n57888;
  assign n57890 = pi23 ? n233 : n5630;
  assign n57891 = pi22 ? n57890 : n32;
  assign n57892 = pi21 ? n57883 : n57891;
  assign n57893 = pi20 ? n31220 : n57892;
  assign n57894 = pi19 ? n20563 : n57893;
  assign n57895 = pi18 ? n20563 : n57894;
  assign n57896 = pi17 ? n42700 : n57895;
  assign n57897 = pi16 ? n32 : n57896;
  assign n57898 = pi15 ? n57889 : n57897;
  assign n57899 = pi14 ? n57881 : n57898;
  assign n57900 = pi22 ? n48052 : n685;
  assign n57901 = pi22 ? n54160 : n32;
  assign n57902 = pi21 ? n57900 : n57901;
  assign n57903 = pi20 ? n20563 : n57902;
  assign n57904 = pi19 ? n20563 : n57903;
  assign n57905 = pi18 ? n20563 : n57904;
  assign n57906 = pi17 ? n46998 : n57905;
  assign n57907 = pi16 ? n32 : n57906;
  assign n57908 = pi21 ? n57900 : n731;
  assign n57909 = pi20 ? n31220 : n57908;
  assign n57910 = pi19 ? n20563 : n57909;
  assign n57911 = pi18 ? n20563 : n57910;
  assign n57912 = pi17 ? n41169 : n57911;
  assign n57913 = pi16 ? n32 : n57912;
  assign n57914 = pi15 ? n57907 : n57913;
  assign n57915 = pi21 ? n57900 : n33622;
  assign n57916 = pi20 ? n31220 : n57915;
  assign n57917 = pi19 ? n20563 : n57916;
  assign n57918 = pi18 ? n20563 : n57917;
  assign n57919 = pi17 ? n41169 : n57918;
  assign n57920 = pi16 ? n32 : n57919;
  assign n57921 = pi21 ? n57900 : n760;
  assign n57922 = pi20 ? n31220 : n57921;
  assign n57923 = pi19 ? n20563 : n57922;
  assign n57924 = pi18 ? n20563 : n57923;
  assign n57925 = pi17 ? n40024 : n57924;
  assign n57926 = pi16 ? n32 : n57925;
  assign n57927 = pi15 ? n57920 : n57926;
  assign n57928 = pi14 ? n57914 : n57927;
  assign n57929 = pi13 ? n57899 : n57928;
  assign n57930 = pi12 ? n57865 : n57929;
  assign n57931 = pi17 ? n40024 : n57334;
  assign n57932 = pi16 ? n32 : n57931;
  assign n57933 = pi17 ? n41182 : n57339;
  assign n57934 = pi16 ? n32 : n57933;
  assign n57935 = pi15 ? n57932 : n57934;
  assign n57936 = pi17 ? n42240 : n57346;
  assign n57937 = pi16 ? n32 : n57936;
  assign n57938 = pi21 ? n2412 : n928;
  assign n57939 = pi20 ? n56350 : n57938;
  assign n57940 = pi19 ? n20563 : n57939;
  assign n57941 = pi18 ? n20563 : n57940;
  assign n57942 = pi17 ? n46447 : n57941;
  assign n57943 = pi16 ? n32 : n57942;
  assign n57944 = pi15 ? n57937 : n57943;
  assign n57945 = pi14 ? n57935 : n57944;
  assign n57946 = pi17 ? n46447 : n57363;
  assign n57947 = pi16 ? n32 : n57946;
  assign n57948 = pi15 ? n57943 : n57947;
  assign n57949 = pi17 ? n46447 : n57369;
  assign n57950 = pi16 ? n32 : n57949;
  assign n57951 = pi20 ? n6402 : n43905;
  assign n57952 = pi19 ? n20563 : n57951;
  assign n57953 = pi18 ? n20563 : n57952;
  assign n57954 = pi17 ? n40498 : n57953;
  assign n57955 = pi16 ? n32 : n57954;
  assign n57956 = pi15 ? n57950 : n57955;
  assign n57957 = pi14 ? n57948 : n57956;
  assign n57958 = pi13 ? n57945 : n57957;
  assign n57959 = pi20 ? n57382 : n43905;
  assign n57960 = pi19 ? n20563 : n57959;
  assign n57961 = pi18 ? n20563 : n57960;
  assign n57962 = pi17 ? n41683 : n57961;
  assign n57963 = pi16 ? n32 : n57962;
  assign n57964 = pi20 ? n56389 : n1010;
  assign n57965 = pi19 ? n20563 : n57964;
  assign n57966 = pi18 ? n20563 : n57965;
  assign n57967 = pi17 ? n41683 : n57966;
  assign n57968 = pi16 ? n32 : n57967;
  assign n57969 = pi15 ? n57963 : n57968;
  assign n57970 = pi17 ? n40511 : n57401;
  assign n57971 = pi16 ? n32 : n57970;
  assign n57972 = pi17 ? n40511 : n57407;
  assign n57973 = pi16 ? n32 : n57972;
  assign n57974 = pi15 ? n57971 : n57973;
  assign n57975 = pi14 ? n57969 : n57974;
  assign n57976 = pi17 ? n40511 : n57414;
  assign n57977 = pi16 ? n32 : n57976;
  assign n57978 = pi17 ? n39374 : n57419;
  assign n57979 = pi16 ? n32 : n57978;
  assign n57980 = pi15 ? n57977 : n57979;
  assign n57981 = pi23 ? n36659 : n685;
  assign n57982 = pi22 ? n20563 : n57981;
  assign n57983 = pi21 ? n20563 : n57982;
  assign n57984 = pi20 ? n57983 : n57425;
  assign n57985 = pi19 ? n20563 : n57984;
  assign n57986 = pi18 ? n20563 : n57985;
  assign n57987 = pi17 ? n39374 : n57986;
  assign n57988 = pi16 ? n32 : n57987;
  assign n57989 = pi17 ? n39374 : n57437;
  assign n57990 = pi16 ? n32 : n57989;
  assign n57991 = pi15 ? n57988 : n57990;
  assign n57992 = pi14 ? n57980 : n57991;
  assign n57993 = pi13 ? n57975 : n57992;
  assign n57994 = pi12 ? n57958 : n57993;
  assign n57995 = pi11 ? n57930 : n57994;
  assign n57996 = pi23 ? n36781 : n316;
  assign n57997 = pi22 ? n139 : n57996;
  assign n57998 = pi21 ? n20563 : n57997;
  assign n57999 = pi20 ? n57998 : n4008;
  assign n58000 = pi19 ? n20563 : n57999;
  assign n58001 = pi18 ? n20563 : n58000;
  assign n58002 = pi17 ? n45367 : n58001;
  assign n58003 = pi16 ? n32 : n58002;
  assign n58004 = pi22 ? n49800 : n13481;
  assign n58005 = pi21 ? n20563 : n58004;
  assign n58006 = pi20 ? n58005 : n56130;
  assign n58007 = pi19 ? n20563 : n58006;
  assign n58008 = pi18 ? n20563 : n58007;
  assign n58009 = pi17 ? n41709 : n58008;
  assign n58010 = pi16 ? n32 : n58009;
  assign n58011 = pi15 ? n58003 : n58010;
  assign n58012 = pi22 ? n9827 : n42172;
  assign n58013 = pi21 ? n20563 : n58012;
  assign n58014 = pi20 ? n58013 : n57459;
  assign n58015 = pi19 ? n20563 : n58014;
  assign n58016 = pi18 ? n20563 : n58015;
  assign n58017 = pi17 ? n41709 : n58016;
  assign n58018 = pi16 ? n32 : n58017;
  assign n58019 = pi22 ? n56616 : n233;
  assign n58020 = pi21 ? n36249 : n58019;
  assign n58021 = pi20 ? n58020 : n56996;
  assign n58022 = pi19 ? n20563 : n58021;
  assign n58023 = pi18 ? n20563 : n58022;
  assign n58024 = pi17 ? n45367 : n58023;
  assign n58025 = pi16 ? n32 : n58024;
  assign n58026 = pi15 ? n58018 : n58025;
  assign n58027 = pi14 ? n58011 : n58026;
  assign n58028 = pi17 ? n45367 : n57479;
  assign n58029 = pi16 ? n32 : n58028;
  assign n58030 = pi23 ? n55580 : n363;
  assign n58031 = pi22 ? n58030 : n685;
  assign n58032 = pi21 ? n56487 : n58031;
  assign n58033 = pi20 ? n58032 : n37640;
  assign n58034 = pi19 ? n20563 : n58033;
  assign n58035 = pi18 ? n20563 : n58034;
  assign n58036 = pi17 ? n45367 : n58035;
  assign n58037 = pi16 ? n32 : n58036;
  assign n58038 = pi15 ? n58029 : n58037;
  assign n58039 = pi20 ? n57494 : n1822;
  assign n58040 = pi19 ? n20563 : n58039;
  assign n58041 = pi18 ? n20563 : n58040;
  assign n58042 = pi17 ? n39398 : n58041;
  assign n58043 = pi16 ? n32 : n58042;
  assign n58044 = pi23 ? n36781 : n56620;
  assign n58045 = pi22 ? n58044 : n316;
  assign n58046 = pi21 ? n57500 : n58045;
  assign n58047 = pi20 ? n58046 : n32;
  assign n58048 = pi19 ? n20563 : n58047;
  assign n58049 = pi18 ? n20563 : n58048;
  assign n58050 = pi17 ? n39398 : n58049;
  assign n58051 = pi16 ? n32 : n58050;
  assign n58052 = pi15 ? n58043 : n58051;
  assign n58053 = pi14 ? n58038 : n58052;
  assign n58054 = pi13 ? n58027 : n58053;
  assign n58055 = pi21 ? n39394 : n39801;
  assign n58056 = pi20 ? n58055 : n40791;
  assign n58057 = pi19 ? n58056 : n57513;
  assign n58058 = pi18 ? n32 : n58057;
  assign n58059 = pi17 ? n58058 : n57523;
  assign n58060 = pi16 ? n32 : n58059;
  assign n58061 = pi21 ? n39394 : n45049;
  assign n58062 = pi20 ? n58061 : n43946;
  assign n58063 = pi19 ? n58062 : n20563;
  assign n58064 = pi18 ? n32 : n58063;
  assign n58065 = pi22 ? n57030 : n21502;
  assign n58066 = pi21 ? n57531 : n58065;
  assign n58067 = pi20 ? n58066 : n32;
  assign n58068 = pi19 ? n20563 : n58067;
  assign n58069 = pi18 ? n20563 : n58068;
  assign n58070 = pi17 ? n58064 : n58069;
  assign n58071 = pi16 ? n32 : n58070;
  assign n58072 = pi15 ? n58060 : n58071;
  assign n58073 = pi21 ? n45620 : n40954;
  assign n58074 = pi21 ? n20563 : n37174;
  assign n58075 = pi20 ? n58073 : n58074;
  assign n58076 = pi19 ? n58075 : n20563;
  assign n58077 = pi18 ? n32 : n58076;
  assign n58078 = pi17 ? n58077 : n57545;
  assign n58079 = pi16 ? n32 : n58078;
  assign n58080 = pi21 ? n47768 : n40954;
  assign n58081 = pi22 ? n37173 : n30195;
  assign n58082 = pi21 ? n20563 : n58081;
  assign n58083 = pi20 ? n58080 : n58082;
  assign n58084 = pi19 ? n58083 : n20563;
  assign n58085 = pi18 ? n32 : n58084;
  assign n58086 = pi22 ? n685 : n53982;
  assign n58087 = pi21 ? n57553 : n58086;
  assign n58088 = pi20 ? n58087 : n32;
  assign n58089 = pi19 ? n20563 : n58088;
  assign n58090 = pi18 ? n20563 : n58089;
  assign n58091 = pi17 ? n58085 : n58090;
  assign n58092 = pi16 ? n32 : n58091;
  assign n58093 = pi15 ? n58079 : n58092;
  assign n58094 = pi14 ? n58072 : n58093;
  assign n58095 = pi17 ? n38317 : n57567;
  assign n58096 = pi16 ? n32 : n58095;
  assign n58097 = pi21 ? n57570 : n2320;
  assign n58098 = pi20 ? n58097 : n32;
  assign n58099 = pi19 ? n56489 : n58098;
  assign n58100 = pi18 ? n20563 : n58099;
  assign n58101 = pi17 ? n45393 : n58100;
  assign n58102 = pi16 ? n32 : n58101;
  assign n58103 = pi15 ? n58096 : n58102;
  assign n58104 = pi17 ? n45393 : n57584;
  assign n58105 = pi16 ? n32 : n58104;
  assign n58106 = pi19 ? n57579 : n57591;
  assign n58107 = pi18 ? n20563 : n58106;
  assign n58108 = pi17 ? n45414 : n58107;
  assign n58109 = pi16 ? n32 : n58108;
  assign n58110 = pi15 ? n58105 : n58109;
  assign n58111 = pi14 ? n58103 : n58110;
  assign n58112 = pi13 ? n58094 : n58111;
  assign n58113 = pi12 ? n58054 : n58112;
  assign n58114 = pi21 ? n57600 : n53983;
  assign n58115 = pi20 ? n58114 : n32;
  assign n58116 = pi19 ? n47159 : n58115;
  assign n58117 = pi18 ? n20563 : n58116;
  assign n58118 = pi17 ? n45414 : n58117;
  assign n58119 = pi16 ? n32 : n58118;
  assign n58120 = pi17 ? n45393 : n57610;
  assign n58121 = pi16 ? n32 : n58120;
  assign n58122 = pi15 ? n58119 : n58121;
  assign n58123 = pi17 ? n45393 : n57620;
  assign n58124 = pi16 ? n32 : n58123;
  assign n58125 = pi22 ? n46165 : n39190;
  assign n58126 = pi21 ? n58125 : n51714;
  assign n58127 = pi21 ? n40912 : n20563;
  assign n58128 = pi20 ? n58126 : n58127;
  assign n58129 = pi22 ? n20563 : n39174;
  assign n58130 = pi21 ? n39801 : n58129;
  assign n58131 = pi21 ? n39191 : n36489;
  assign n58132 = pi20 ? n58130 : n58131;
  assign n58133 = pi19 ? n58128 : n58132;
  assign n58134 = pi18 ? n32 : n58133;
  assign n58135 = pi22 ? n3762 : n56665;
  assign n58136 = pi21 ? n58135 : n32;
  assign n58137 = pi20 ? n58136 : n32;
  assign n58138 = pi19 ? n57631 : n58137;
  assign n58139 = pi18 ? n57629 : n58138;
  assign n58140 = pi17 ? n58134 : n58139;
  assign n58141 = pi16 ? n32 : n58140;
  assign n58142 = pi15 ? n58124 : n58141;
  assign n58143 = pi14 ? n58122 : n58142;
  assign n58144 = pi21 ? n46060 : n20563;
  assign n58145 = pi20 ? n58144 : n30868;
  assign n58146 = pi19 ? n58145 : n30868;
  assign n58147 = pi18 ? n32 : n58146;
  assign n58148 = pi17 ? n58147 : n57652;
  assign n58149 = pi16 ? n32 : n58148;
  assign n58150 = pi20 ? n38376 : n30868;
  assign n58151 = pi19 ? n58150 : n30868;
  assign n58152 = pi18 ? n32 : n58151;
  assign n58153 = pi17 ? n58152 : n57664;
  assign n58154 = pi16 ? n32 : n58153;
  assign n58155 = pi15 ? n58149 : n58154;
  assign n58156 = pi20 ? n38376 : n43010;
  assign n58157 = pi19 ? n58156 : n20563;
  assign n58158 = pi18 ? n32 : n58157;
  assign n58159 = pi17 ? n58158 : n57679;
  assign n58160 = pi16 ? n32 : n58159;
  assign n58161 = pi21 ? n38375 : n39191;
  assign n58162 = pi20 ? n58161 : n38754;
  assign n58163 = pi21 ? n56112 : n20563;
  assign n58164 = pi20 ? n58163 : n43935;
  assign n58165 = pi19 ? n58162 : n58164;
  assign n58166 = pi18 ? n32 : n58165;
  assign n58167 = pi22 ? n54520 : n32;
  assign n58168 = pi21 ? n58167 : n32;
  assign n58169 = pi20 ? n58168 : n32;
  assign n58170 = pi19 ? n57673 : n58169;
  assign n58171 = pi18 ? n20563 : n58170;
  assign n58172 = pi17 ? n58166 : n58171;
  assign n58173 = pi16 ? n32 : n58172;
  assign n58174 = pi15 ? n58160 : n58173;
  assign n58175 = pi14 ? n58155 : n58174;
  assign n58176 = pi13 ? n58143 : n58175;
  assign n58177 = pi19 ? n49709 : n30868;
  assign n58178 = pi18 ? n32 : n58177;
  assign n58179 = pi17 ? n58178 : n57702;
  assign n58180 = pi16 ? n32 : n58179;
  assign n58181 = pi21 ? n45653 : n47396;
  assign n58182 = pi20 ? n58181 : n55701;
  assign n58183 = pi19 ? n58182 : n56722;
  assign n58184 = pi18 ? n32 : n58183;
  assign n58185 = pi17 ? n58184 : n57719;
  assign n58186 = pi16 ? n32 : n58185;
  assign n58187 = pi15 ? n58180 : n58186;
  assign n58188 = pi19 ? n52406 : n57726;
  assign n58189 = pi18 ? n32 : n58188;
  assign n58190 = pi17 ? n58189 : n57737;
  assign n58191 = pi16 ? n32 : n58190;
  assign n58192 = pi21 ? n32 : n47396;
  assign n58193 = pi20 ? n58192 : n54009;
  assign n58194 = pi19 ? n58193 : n43198;
  assign n58195 = pi18 ? n32 : n58194;
  assign n58196 = pi17 ? n58195 : n57750;
  assign n58197 = pi16 ? n32 : n58196;
  assign n58198 = pi15 ? n58191 : n58197;
  assign n58199 = pi14 ? n58187 : n58198;
  assign n58200 = pi20 ? n54007 : n43198;
  assign n58201 = pi19 ? n58200 : n43198;
  assign n58202 = pi18 ? n32 : n58201;
  assign n58203 = pi17 ? n58202 : n57764;
  assign n58204 = pi16 ? n32 : n58203;
  assign n58205 = pi20 ? n45663 : n56771;
  assign n58206 = pi24 ? n36798 : n36781;
  assign n58207 = pi23 ? n58206 : n36781;
  assign n58208 = pi22 ? n58207 : n36781;
  assign n58209 = pi21 ? n39972 : n58208;
  assign n58210 = pi20 ? n58209 : n36781;
  assign n58211 = pi19 ? n58205 : n58210;
  assign n58212 = pi18 ? n32 : n58211;
  assign n58213 = pi17 ? n58212 : n57778;
  assign n58214 = pi16 ? n32 : n58213;
  assign n58215 = pi15 ? n58204 : n58214;
  assign n58216 = pi22 ? n45135 : n49412;
  assign n58217 = pi21 ? n32 : n58216;
  assign n58218 = pi21 ? n53537 : n39972;
  assign n58219 = pi20 ? n58217 : n58218;
  assign n58220 = pi24 ? n43198 : n36781;
  assign n58221 = pi23 ? n58220 : n36781;
  assign n58222 = pi22 ? n58221 : n36781;
  assign n58223 = pi21 ? n47397 : n58222;
  assign n58224 = pi20 ? n58223 : n36781;
  assign n58225 = pi19 ? n58219 : n58224;
  assign n58226 = pi18 ? n32 : n58225;
  assign n58227 = pi17 ? n58226 : n57794;
  assign n58228 = pi16 ? n32 : n58227;
  assign n58229 = pi20 ? n45670 : n55701;
  assign n58230 = pi19 ? n58229 : n56808;
  assign n58231 = pi18 ? n32 : n58230;
  assign n58232 = pi17 ? n58231 : n57804;
  assign n58233 = pi16 ? n32 : n58232;
  assign n58234 = pi15 ? n58228 : n58233;
  assign n58235 = pi14 ? n58215 : n58234;
  assign n58236 = pi13 ? n58199 : n58235;
  assign n58237 = pi12 ? n58176 : n58236;
  assign n58238 = pi11 ? n58113 : n58237;
  assign n58239 = pi10 ? n57995 : n58238;
  assign n58240 = pi09 ? n57826 : n58239;
  assign n58241 = pi08 ? n57813 : n58240;
  assign n58242 = pi22 ? n13624 : n139;
  assign n58243 = pi21 ? n58242 : n5623;
  assign n58244 = pi20 ? n31220 : n58243;
  assign n58245 = pi19 ? n20563 : n58244;
  assign n58246 = pi18 ? n20563 : n58245;
  assign n58247 = pi17 ? n44652 : n58246;
  assign n58248 = pi16 ? n32 : n58247;
  assign n58249 = pi15 ? n32 : n58248;
  assign n58250 = pi20 ? n31220 : n12252;
  assign n58251 = pi19 ? n20563 : n58250;
  assign n58252 = pi18 ? n20563 : n58251;
  assign n58253 = pi17 ? n44222 : n58252;
  assign n58254 = pi16 ? n32 : n58253;
  assign n58255 = pi21 ? n37 : n5640;
  assign n58256 = pi20 ? n31220 : n58255;
  assign n58257 = pi19 ? n20563 : n58256;
  assign n58258 = pi18 ? n20563 : n58257;
  assign n58259 = pi17 ? n45242 : n58258;
  assign n58260 = pi16 ? n32 : n58259;
  assign n58261 = pi15 ? n58254 : n58260;
  assign n58262 = pi14 ? n58249 : n58261;
  assign n58263 = pi13 ? n32 : n58262;
  assign n58264 = pi12 ? n32 : n58263;
  assign n58265 = pi11 ? n32 : n58264;
  assign n58266 = pi10 ? n32 : n58265;
  assign n58267 = pi21 ? n37 : n22885;
  assign n58268 = pi20 ? n20563 : n58267;
  assign n58269 = pi19 ? n20563 : n58268;
  assign n58270 = pi18 ? n20563 : n58269;
  assign n58271 = pi17 ? n43663 : n58270;
  assign n58272 = pi16 ? n32 : n58271;
  assign n58273 = pi21 ? n37 : n11928;
  assign n58274 = pi20 ? n20563 : n58273;
  assign n58275 = pi19 ? n20563 : n58274;
  assign n58276 = pi18 ? n20563 : n58275;
  assign n58277 = pi17 ? n44670 : n58276;
  assign n58278 = pi16 ? n32 : n58277;
  assign n58279 = pi15 ? n58272 : n58278;
  assign n58280 = pi21 ? n37 : n4748;
  assign n58281 = pi20 ? n20563 : n58280;
  assign n58282 = pi19 ? n20563 : n58281;
  assign n58283 = pi18 ? n20563 : n58282;
  assign n58284 = pi17 ? n43223 : n58283;
  assign n58285 = pi16 ? n32 : n58284;
  assign n58286 = pi20 ? n20563 : n12042;
  assign n58287 = pi19 ? n20563 : n58286;
  assign n58288 = pi18 ? n20563 : n58287;
  assign n58289 = pi17 ? n43223 : n58288;
  assign n58290 = pi16 ? n32 : n58289;
  assign n58291 = pi15 ? n58285 : n58290;
  assign n58292 = pi14 ? n58279 : n58291;
  assign n58293 = pi21 ? n2091 : n7034;
  assign n58294 = pi20 ? n31220 : n58293;
  assign n58295 = pi19 ? n20563 : n58294;
  assign n58296 = pi18 ? n20563 : n58295;
  assign n58297 = pi17 ? n43223 : n58296;
  assign n58298 = pi16 ? n32 : n58297;
  assign n58299 = pi17 ? n43227 : n58296;
  assign n58300 = pi16 ? n32 : n58299;
  assign n58301 = pi15 ? n58298 : n58300;
  assign n58302 = pi21 ? n2091 : n7723;
  assign n58303 = pi20 ? n31220 : n58302;
  assign n58304 = pi19 ? n20563 : n58303;
  assign n58305 = pi18 ? n20563 : n58304;
  assign n58306 = pi17 ? n43248 : n58305;
  assign n58307 = pi16 ? n32 : n58306;
  assign n58308 = pi21 ? n2106 : n7048;
  assign n58309 = pi20 ? n31266 : n58308;
  assign n58310 = pi19 ? n20563 : n58309;
  assign n58311 = pi18 ? n20563 : n58310;
  assign n58312 = pi17 ? n48624 : n58311;
  assign n58313 = pi16 ? n32 : n58312;
  assign n58314 = pi15 ? n58307 : n58313;
  assign n58315 = pi14 ? n58301 : n58314;
  assign n58316 = pi13 ? n58292 : n58315;
  assign n58317 = pi21 ? n2106 : n2320;
  assign n58318 = pi20 ? n31220 : n58317;
  assign n58319 = pi19 ? n20563 : n58318;
  assign n58320 = pi18 ? n20563 : n58319;
  assign n58321 = pi17 ? n43262 : n58320;
  assign n58322 = pi16 ? n32 : n58321;
  assign n58323 = pi23 ? n685 : n260;
  assign n58324 = pi22 ? n58323 : n32;
  assign n58325 = pi21 ? n17806 : n58324;
  assign n58326 = pi20 ? n31220 : n58325;
  assign n58327 = pi19 ? n20563 : n58326;
  assign n58328 = pi18 ? n20563 : n58327;
  assign n58329 = pi17 ? n43262 : n58328;
  assign n58330 = pi16 ? n32 : n58329;
  assign n58331 = pi15 ? n58322 : n58330;
  assign n58332 = pi23 ? n20627 : n685;
  assign n58333 = pi22 ? n58332 : n685;
  assign n58334 = pi23 ? n685 : n586;
  assign n58335 = pi22 ? n58334 : n32;
  assign n58336 = pi21 ? n58333 : n58335;
  assign n58337 = pi20 ? n31220 : n58336;
  assign n58338 = pi19 ? n20563 : n58337;
  assign n58339 = pi18 ? n20563 : n58338;
  assign n58340 = pi17 ? n43262 : n58339;
  assign n58341 = pi16 ? n32 : n58340;
  assign n58342 = pi23 ? n685 : n5630;
  assign n58343 = pi22 ? n58342 : n32;
  assign n58344 = pi21 ? n58333 : n58343;
  assign n58345 = pi20 ? n31220 : n58344;
  assign n58346 = pi19 ? n20563 : n58345;
  assign n58347 = pi18 ? n20563 : n58346;
  assign n58348 = pi17 ? n47593 : n58347;
  assign n58349 = pi16 ? n32 : n58348;
  assign n58350 = pi15 ? n58341 : n58349;
  assign n58351 = pi14 ? n58331 : n58350;
  assign n58352 = pi23 ? n5612 : n685;
  assign n58353 = pi22 ? n58352 : n685;
  assign n58354 = pi21 ? n58353 : n57901;
  assign n58355 = pi20 ? n20563 : n58354;
  assign n58356 = pi19 ? n20563 : n58355;
  assign n58357 = pi18 ? n20563 : n58356;
  assign n58358 = pi17 ? n42207 : n58357;
  assign n58359 = pi16 ? n32 : n58358;
  assign n58360 = pi21 ? n58353 : n731;
  assign n58361 = pi20 ? n31220 : n58360;
  assign n58362 = pi19 ? n20563 : n58361;
  assign n58363 = pi18 ? n20563 : n58362;
  assign n58364 = pi17 ? n42688 : n58363;
  assign n58365 = pi16 ? n32 : n58364;
  assign n58366 = pi15 ? n58359 : n58365;
  assign n58367 = pi22 ? n48040 : n685;
  assign n58368 = pi21 ? n58367 : n33622;
  assign n58369 = pi20 ? n31220 : n58368;
  assign n58370 = pi19 ? n20563 : n58369;
  assign n58371 = pi18 ? n20563 : n58370;
  assign n58372 = pi17 ? n42688 : n58371;
  assign n58373 = pi16 ? n32 : n58372;
  assign n58374 = pi22 ? n5782 : n685;
  assign n58375 = pi21 ? n58374 : n760;
  assign n58376 = pi20 ? n31220 : n58375;
  assign n58377 = pi19 ? n20563 : n58376;
  assign n58378 = pi18 ? n20563 : n58377;
  assign n58379 = pi17 ? n42688 : n58378;
  assign n58380 = pi16 ? n32 : n58379;
  assign n58381 = pi15 ? n58373 : n58380;
  assign n58382 = pi14 ? n58366 : n58381;
  assign n58383 = pi13 ? n58351 : n58382;
  assign n58384 = pi12 ? n58316 : n58383;
  assign n58385 = pi22 ? n705 : n316;
  assign n58386 = pi21 ? n58385 : n882;
  assign n58387 = pi20 ? n54354 : n58386;
  assign n58388 = pi19 ? n20563 : n58387;
  assign n58389 = pi18 ? n20563 : n58388;
  assign n58390 = pi17 ? n42688 : n58389;
  assign n58391 = pi16 ? n32 : n58390;
  assign n58392 = pi17 ? n42700 : n57339;
  assign n58393 = pi16 ? n32 : n58392;
  assign n58394 = pi15 ? n58391 : n58393;
  assign n58395 = pi21 ? n20563 : n181;
  assign n58396 = pi20 ? n58395 : n8644;
  assign n58397 = pi19 ? n20563 : n58396;
  assign n58398 = pi18 ? n20563 : n58397;
  assign n58399 = pi17 ? n46998 : n58398;
  assign n58400 = pi16 ? n32 : n58399;
  assign n58401 = pi21 ? n1027 : n2578;
  assign n58402 = pi20 ? n56350 : n58401;
  assign n58403 = pi19 ? n20563 : n58402;
  assign n58404 = pi18 ? n20563 : n58403;
  assign n58405 = pi17 ? n41158 : n58404;
  assign n58406 = pi16 ? n32 : n58405;
  assign n58407 = pi15 ? n58400 : n58406;
  assign n58408 = pi14 ? n58394 : n58407;
  assign n58409 = pi21 ? n1027 : n2637;
  assign n58410 = pi20 ? n56350 : n58409;
  assign n58411 = pi19 ? n20563 : n58410;
  assign n58412 = pi18 ? n20563 : n58411;
  assign n58413 = pi17 ? n41158 : n58412;
  assign n58414 = pi16 ? n32 : n58413;
  assign n58415 = pi17 ? n41169 : n57363;
  assign n58416 = pi16 ? n32 : n58415;
  assign n58417 = pi15 ? n58414 : n58416;
  assign n58418 = pi17 ? n41169 : n57369;
  assign n58419 = pi16 ? n32 : n58418;
  assign n58420 = pi20 ? n6402 : n980;
  assign n58421 = pi19 ? n20563 : n58420;
  assign n58422 = pi18 ? n20563 : n58421;
  assign n58423 = pi17 ? n40024 : n58422;
  assign n58424 = pi16 ? n32 : n58423;
  assign n58425 = pi15 ? n58419 : n58424;
  assign n58426 = pi14 ? n58417 : n58425;
  assign n58427 = pi13 ? n58408 : n58426;
  assign n58428 = pi23 ? n20563 : n36781;
  assign n58429 = pi22 ? n37 : n58428;
  assign n58430 = pi21 ? n20563 : n58429;
  assign n58431 = pi20 ? n58430 : n1010;
  assign n58432 = pi19 ? n20563 : n58431;
  assign n58433 = pi18 ? n20563 : n58432;
  assign n58434 = pi17 ? n41182 : n58433;
  assign n58435 = pi16 ? n32 : n58434;
  assign n58436 = pi17 ? n47057 : n57966;
  assign n58437 = pi16 ? n32 : n58436;
  assign n58438 = pi15 ? n58435 : n58437;
  assign n58439 = pi21 ? n13481 : n20952;
  assign n58440 = pi20 ? n57404 : n58439;
  assign n58441 = pi19 ? n20563 : n58440;
  assign n58442 = pi18 ? n20563 : n58441;
  assign n58443 = pi17 ? n47057 : n58442;
  assign n58444 = pi16 ? n32 : n58443;
  assign n58445 = pi20 ? n57404 : n15407;
  assign n58446 = pi19 ? n20563 : n58445;
  assign n58447 = pi18 ? n20563 : n58446;
  assign n58448 = pi17 ? n47057 : n58447;
  assign n58449 = pi16 ? n32 : n58448;
  assign n58450 = pi15 ? n58444 : n58449;
  assign n58451 = pi14 ? n58438 : n58450;
  assign n58452 = pi23 ? n51564 : n32;
  assign n58453 = pi22 ? n233 : n58452;
  assign n58454 = pi21 ? n58453 : n32;
  assign n58455 = pi20 ? n31410 : n58454;
  assign n58456 = pi19 ? n31221 : n58455;
  assign n58457 = pi18 ? n20563 : n58456;
  assign n58458 = pi17 ? n47057 : n58457;
  assign n58459 = pi16 ? n32 : n58458;
  assign n58460 = pi17 ? n46447 : n57419;
  assign n58461 = pi16 ? n32 : n58460;
  assign n58462 = pi15 ? n58459 : n58461;
  assign n58463 = pi22 ? n20563 : n686;
  assign n58464 = pi21 ? n20563 : n58463;
  assign n58465 = pi20 ? n58464 : n57425;
  assign n58466 = pi19 ? n20563 : n58465;
  assign n58467 = pi18 ? n20563 : n58466;
  assign n58468 = pi17 ? n46447 : n58467;
  assign n58469 = pi16 ? n32 : n58468;
  assign n58470 = pi22 ? n51564 : n21502;
  assign n58471 = pi21 ? n58470 : n32;
  assign n58472 = pi20 ? n57432 : n58471;
  assign n58473 = pi19 ? n20563 : n58472;
  assign n58474 = pi18 ? n20563 : n58473;
  assign n58475 = pi17 ? n46447 : n58474;
  assign n58476 = pi16 ? n32 : n58475;
  assign n58477 = pi15 ? n58469 : n58476;
  assign n58478 = pi14 ? n58462 : n58477;
  assign n58479 = pi13 ? n58451 : n58478;
  assign n58480 = pi12 ? n58427 : n58479;
  assign n58481 = pi11 ? n58384 : n58480;
  assign n58482 = pi21 ? n20563 : n346;
  assign n58483 = pi20 ? n58482 : n4008;
  assign n58484 = pi19 ? n20563 : n58483;
  assign n58485 = pi18 ? n20563 : n58484;
  assign n58486 = pi17 ? n40498 : n58485;
  assign n58487 = pi16 ? n32 : n58486;
  assign n58488 = pi22 ? n139 : n13481;
  assign n58489 = pi21 ? n20563 : n58488;
  assign n58490 = pi20 ? n58489 : n56130;
  assign n58491 = pi19 ? n20563 : n58490;
  assign n58492 = pi18 ? n20563 : n58491;
  assign n58493 = pi17 ? n40498 : n58492;
  assign n58494 = pi16 ? n32 : n58493;
  assign n58495 = pi15 ? n58487 : n58494;
  assign n58496 = pi21 ? n20563 : n1079;
  assign n58497 = pi20 ? n58496 : n5830;
  assign n58498 = pi19 ? n20563 : n58497;
  assign n58499 = pi18 ? n20563 : n58498;
  assign n58500 = pi17 ? n40498 : n58499;
  assign n58501 = pi16 ? n32 : n58500;
  assign n58502 = pi21 ? n31890 : n6376;
  assign n58503 = pi22 ? n57647 : n32;
  assign n58504 = pi21 ? n58503 : n32;
  assign n58505 = pi20 ? n58502 : n58504;
  assign n58506 = pi19 ? n20563 : n58505;
  assign n58507 = pi18 ? n20563 : n58506;
  assign n58508 = pi17 ? n41683 : n58507;
  assign n58509 = pi16 ? n32 : n58508;
  assign n58510 = pi15 ? n58501 : n58509;
  assign n58511 = pi14 ? n58495 : n58510;
  assign n58512 = pi21 ? n31890 : n233;
  assign n58513 = pi20 ? n58512 : n2653;
  assign n58514 = pi19 ? n20563 : n58513;
  assign n58515 = pi18 ? n20563 : n58514;
  assign n58516 = pi17 ? n41683 : n58515;
  assign n58517 = pi16 ? n32 : n58516;
  assign n58518 = pi22 ? n37 : n37240;
  assign n58519 = pi23 ? n55580 : n36781;
  assign n58520 = pi22 ? n58519 : n685;
  assign n58521 = pi21 ? n58518 : n58520;
  assign n58522 = pi20 ? n58521 : n37640;
  assign n58523 = pi19 ? n20563 : n58522;
  assign n58524 = pi18 ? n20563 : n58523;
  assign n58525 = pi17 ? n41683 : n58524;
  assign n58526 = pi16 ? n32 : n58525;
  assign n58527 = pi15 ? n58517 : n58526;
  assign n58528 = pi24 ? n335 : n36781;
  assign n58529 = pi23 ? n58528 : n157;
  assign n58530 = pi22 ? n58529 : n51564;
  assign n58531 = pi21 ? n57500 : n58530;
  assign n58532 = pi20 ? n58531 : n1822;
  assign n58533 = pi19 ? n20563 : n58532;
  assign n58534 = pi18 ? n20563 : n58533;
  assign n58535 = pi17 ? n41709 : n58534;
  assign n58536 = pi16 ? n32 : n58535;
  assign n58537 = pi22 ? n37 : n40428;
  assign n58538 = pi24 ? n36781 : n204;
  assign n58539 = pi23 ? n36781 : n58538;
  assign n58540 = pi22 ? n58539 : n316;
  assign n58541 = pi21 ? n58537 : n58540;
  assign n58542 = pi20 ? n58541 : n32;
  assign n58543 = pi19 ? n20563 : n58542;
  assign n58544 = pi18 ? n20563 : n58543;
  assign n58545 = pi17 ? n40533 : n58544;
  assign n58546 = pi16 ? n32 : n58545;
  assign n58547 = pi15 ? n58536 : n58546;
  assign n58548 = pi14 ? n58527 : n58547;
  assign n58549 = pi13 ? n58511 : n58548;
  assign n58550 = pi20 ? n54401 : n40791;
  assign n58551 = pi19 ? n58550 : n57513;
  assign n58552 = pi18 ? n32 : n58551;
  assign n58553 = pi23 ? n58538 : n204;
  assign n58554 = pi22 ? n58553 : n13481;
  assign n58555 = pi21 ? n57531 : n58554;
  assign n58556 = pi20 ? n58555 : n32;
  assign n58557 = pi19 ? n20563 : n58556;
  assign n58558 = pi18 ? n52168 : n58557;
  assign n58559 = pi17 ? n58552 : n58558;
  assign n58560 = pi16 ? n32 : n58559;
  assign n58561 = pi20 ? n37933 : n39192;
  assign n58562 = pi20 ? n51188 : n20563;
  assign n58563 = pi19 ? n58561 : n58562;
  assign n58564 = pi18 ? n32 : n58563;
  assign n58565 = pi22 ? n99 : n38926;
  assign n58566 = pi24 ? n43198 : n233;
  assign n58567 = pi23 ? n43198 : n58566;
  assign n58568 = pi22 ? n58567 : n317;
  assign n58569 = pi21 ? n58565 : n58568;
  assign n58570 = pi20 ? n58569 : n32;
  assign n58571 = pi19 ? n20563 : n58570;
  assign n58572 = pi18 ? n20563 : n58571;
  assign n58573 = pi17 ? n58564 : n58572;
  assign n58574 = pi16 ? n32 : n58573;
  assign n58575 = pi15 ? n58560 : n58574;
  assign n58576 = pi22 ? n45516 : n20563;
  assign n58577 = pi21 ? n32 : n58576;
  assign n58578 = pi21 ? n40917 : n51214;
  assign n58579 = pi20 ? n58577 : n58578;
  assign n58580 = pi22 ? n55502 : n40386;
  assign n58581 = pi21 ? n52632 : n58580;
  assign n58582 = pi20 ? n58581 : n20563;
  assign n58583 = pi19 ? n58579 : n58582;
  assign n58584 = pi18 ? n32 : n58583;
  assign n58585 = pi21 ? n40957 : n20563;
  assign n58586 = pi20 ? n20563 : n58585;
  assign n58587 = pi19 ? n20563 : n58586;
  assign n58588 = pi18 ? n58587 : n57544;
  assign n58589 = pi17 ? n58584 : n58588;
  assign n58590 = pi16 ? n32 : n58589;
  assign n58591 = pi22 ? n43571 : n37173;
  assign n58592 = pi21 ? n40960 : n58591;
  assign n58593 = pi20 ? n37933 : n58592;
  assign n58594 = pi22 ? n55535 : n20563;
  assign n58595 = pi21 ? n52758 : n58594;
  assign n58596 = pi20 ? n58595 : n20563;
  assign n58597 = pi19 ? n58593 : n58596;
  assign n58598 = pi18 ? n32 : n58597;
  assign n58599 = pi22 ? n139 : n40004;
  assign n58600 = pi21 ? n58599 : n8486;
  assign n58601 = pi20 ? n58600 : n32;
  assign n58602 = pi19 ? n20563 : n58601;
  assign n58603 = pi18 ? n20563 : n58602;
  assign n58604 = pi17 ? n58598 : n58603;
  assign n58605 = pi16 ? n32 : n58604;
  assign n58606 = pi15 ? n58590 : n58605;
  assign n58607 = pi14 ? n58575 : n58606;
  assign n58608 = pi21 ? n1079 : n57563;
  assign n58609 = pi20 ? n58608 : n32;
  assign n58610 = pi19 ? n20563 : n58609;
  assign n58611 = pi18 ? n20563 : n58610;
  assign n58612 = pi17 ? n38949 : n58611;
  assign n58613 = pi16 ? n32 : n58612;
  assign n58614 = pi22 ? n363 : n43198;
  assign n58615 = pi21 ? n58614 : n2320;
  assign n58616 = pi20 ? n58615 : n32;
  assign n58617 = pi19 ? n56489 : n58616;
  assign n58618 = pi18 ? n20563 : n58617;
  assign n58619 = pi17 ? n38949 : n58618;
  assign n58620 = pi16 ? n32 : n58619;
  assign n58621 = pi15 ? n58613 : n58620;
  assign n58622 = pi21 ? n52373 : n55560;
  assign n58623 = pi20 ? n58622 : n32;
  assign n58624 = pi19 ? n57579 : n58623;
  assign n58625 = pi18 ? n20563 : n58624;
  assign n58626 = pi17 ? n38949 : n58625;
  assign n58627 = pi16 ? n32 : n58626;
  assign n58628 = pi21 ? n20563 : n57500;
  assign n58629 = pi20 ? n20563 : n58628;
  assign n58630 = pi19 ? n58629 : n57591;
  assign n58631 = pi18 ? n20563 : n58630;
  assign n58632 = pi17 ? n38958 : n58631;
  assign n58633 = pi16 ? n32 : n58632;
  assign n58634 = pi15 ? n58627 : n58633;
  assign n58635 = pi14 ? n58621 : n58634;
  assign n58636 = pi13 ? n58607 : n58635;
  assign n58637 = pi12 ? n58549 : n58636;
  assign n58638 = pi23 ? n335 : n33792;
  assign n58639 = pi22 ? n20563 : n58638;
  assign n58640 = pi21 ? n20563 : n58639;
  assign n58641 = pi20 ? n20563 : n58640;
  assign n58642 = pi22 ? n233 : n51564;
  assign n58643 = pi21 ? n58642 : n1009;
  assign n58644 = pi20 ? n58643 : n32;
  assign n58645 = pi19 ? n58641 : n58644;
  assign n58646 = pi18 ? n20563 : n58645;
  assign n58647 = pi17 ? n38958 : n58646;
  assign n58648 = pi16 ? n32 : n58647;
  assign n58649 = pi17 ? n38949 : n57610;
  assign n58650 = pi16 ? n32 : n58649;
  assign n58651 = pi15 ? n58648 : n58650;
  assign n58652 = pi22 ? n685 : n57647;
  assign n58653 = pi21 ? n58652 : n32;
  assign n58654 = pi20 ? n58653 : n32;
  assign n58655 = pi19 ? n57615 : n58654;
  assign n58656 = pi18 ? n20563 : n58655;
  assign n58657 = pi17 ? n41709 : n58656;
  assign n58658 = pi16 ? n32 : n58657;
  assign n58659 = pi20 ? n51233 : n48184;
  assign n58660 = pi20 ? n42005 : n36489;
  assign n58661 = pi19 ? n58659 : n58660;
  assign n58662 = pi18 ? n32 : n58661;
  assign n58663 = pi20 ? n38754 : n39801;
  assign n58664 = pi19 ? n40791 : n58663;
  assign n58665 = pi22 ? n51564 : n57647;
  assign n58666 = pi21 ? n58665 : n32;
  assign n58667 = pi20 ? n58666 : n32;
  assign n58668 = pi19 ? n57631 : n58667;
  assign n58669 = pi18 ? n58664 : n58668;
  assign n58670 = pi17 ? n58662 : n58669;
  assign n58671 = pi16 ? n32 : n58670;
  assign n58672 = pi15 ? n58658 : n58671;
  assign n58673 = pi14 ? n58651 : n58672;
  assign n58674 = pi19 ? n52840 : n30868;
  assign n58675 = pi18 ? n32 : n58674;
  assign n58676 = pi22 ? n316 : n21502;
  assign n58677 = pi21 ? n58676 : n32;
  assign n58678 = pi20 ? n58677 : n32;
  assign n58679 = pi19 ? n57646 : n58678;
  assign n58680 = pi18 ? n55521 : n58679;
  assign n58681 = pi17 ? n58675 : n58680;
  assign n58682 = pi16 ? n32 : n58681;
  assign n58683 = pi17 ? n58675 : n57664;
  assign n58684 = pi16 ? n32 : n58683;
  assign n58685 = pi15 ? n58682 : n58684;
  assign n58686 = pi20 ? n36867 : n43010;
  assign n58687 = pi19 ? n58686 : n20563;
  assign n58688 = pi18 ? n32 : n58687;
  assign n58689 = pi19 ? n57673 : n4117;
  assign n58690 = pi18 ? n40793 : n58689;
  assign n58691 = pi17 ? n58688 : n58690;
  assign n58692 = pi16 ? n32 : n58691;
  assign n58693 = pi21 ? n30868 : n40249;
  assign n58694 = pi20 ? n30868 : n58693;
  assign n58695 = pi20 ? n30868 : n41463;
  assign n58696 = pi19 ? n58694 : n58695;
  assign n58697 = pi20 ? n30868 : n57672;
  assign n58698 = pi19 ? n58697 : n54566;
  assign n58699 = pi18 ? n58696 : n58698;
  assign n58700 = pi17 ? n58675 : n58699;
  assign n58701 = pi16 ? n32 : n58700;
  assign n58702 = pi15 ? n58692 : n58701;
  assign n58703 = pi14 ? n58685 : n58702;
  assign n58704 = pi13 ? n58673 : n58703;
  assign n58705 = pi18 ? n32 : n52852;
  assign n58706 = pi17 ? n58705 : n57702;
  assign n58707 = pi16 ? n32 : n58706;
  assign n58708 = pi22 ? n32 : n55799;
  assign n58709 = pi21 ? n32 : n58708;
  assign n58710 = pi23 ? n33792 : n36659;
  assign n58711 = pi22 ? n58710 : n36798;
  assign n58712 = pi21 ? n58711 : n43198;
  assign n58713 = pi20 ? n58709 : n58712;
  assign n58714 = pi19 ? n58713 : n56722;
  assign n58715 = pi18 ? n32 : n58714;
  assign n58716 = pi19 ? n57715 : n37641;
  assign n58717 = pi18 ? n57711 : n58716;
  assign n58718 = pi17 ? n58715 : n58717;
  assign n58719 = pi16 ? n32 : n58718;
  assign n58720 = pi15 ? n58707 : n58719;
  assign n58721 = pi22 ? n38284 : n43198;
  assign n58722 = pi22 ? n54580 : n43198;
  assign n58723 = pi21 ? n58721 : n58722;
  assign n58724 = pi20 ? n52918 : n58723;
  assign n58725 = pi22 ? n36798 : n56712;
  assign n58726 = pi21 ? n43198 : n58725;
  assign n58727 = pi21 ? n53471 : n53484;
  assign n58728 = pi20 ? n58726 : n58727;
  assign n58729 = pi19 ? n58724 : n58728;
  assign n58730 = pi18 ? n32 : n58729;
  assign n58731 = pi21 ? n53484 : n43198;
  assign n58732 = pi22 ? n43198 : n52395;
  assign n58733 = pi21 ? n58732 : n43198;
  assign n58734 = pi20 ? n58731 : n58733;
  assign n58735 = pi22 ? n43198 : n49406;
  assign n58736 = pi23 ? n36659 : n33792;
  assign n58737 = pi22 ? n58736 : n43198;
  assign n58738 = pi21 ? n58735 : n58737;
  assign n58739 = pi20 ? n58731 : n58738;
  assign n58740 = pi19 ? n58734 : n58739;
  assign n58741 = pi19 ? n57735 : n32;
  assign n58742 = pi18 ? n58740 : n58741;
  assign n58743 = pi17 ? n58730 : n58742;
  assign n58744 = pi16 ? n32 : n58743;
  assign n58745 = pi21 ? n58721 : n43198;
  assign n58746 = pi20 ? n46201 : n58745;
  assign n58747 = pi19 ? n58746 : n43198;
  assign n58748 = pi18 ? n32 : n58747;
  assign n58749 = pi19 ? n57748 : n32;
  assign n58750 = pi18 ? n57745 : n58749;
  assign n58751 = pi17 ? n58748 : n58750;
  assign n58752 = pi16 ? n32 : n58751;
  assign n58753 = pi15 ? n58744 : n58752;
  assign n58754 = pi14 ? n58720 : n58753;
  assign n58755 = pi22 ? n49412 : n43198;
  assign n58756 = pi21 ? n58755 : n43198;
  assign n58757 = pi20 ? n46225 : n58756;
  assign n58758 = pi19 ? n58757 : n43198;
  assign n58759 = pi18 ? n32 : n58758;
  assign n58760 = pi17 ? n58759 : n57764;
  assign n58761 = pi16 ? n32 : n58760;
  assign n58762 = pi21 ? n58755 : n36798;
  assign n58763 = pi20 ? n46225 : n58762;
  assign n58764 = pi21 ? n36781 : n38901;
  assign n58765 = pi20 ? n57785 : n58764;
  assign n58766 = pi19 ? n58763 : n58765;
  assign n58767 = pi18 ? n32 : n58766;
  assign n58768 = pi21 ? n36798 : n46280;
  assign n58769 = pi20 ? n46280 : n58768;
  assign n58770 = pi22 ? n40004 : n36781;
  assign n58771 = pi21 ? n58770 : n55765;
  assign n58772 = pi22 ? n363 : n36798;
  assign n58773 = pi21 ? n58772 : n43198;
  assign n58774 = pi20 ? n58771 : n58773;
  assign n58775 = pi19 ? n58769 : n58774;
  assign n58776 = pi21 ? n51895 : n55765;
  assign n58777 = pi22 ? n43198 : n14626;
  assign n58778 = pi22 ? n51564 : n706;
  assign n58779 = pi21 ? n58777 : n58778;
  assign n58780 = pi20 ? n58776 : n58779;
  assign n58781 = pi19 ? n58780 : n32;
  assign n58782 = pi18 ? n58775 : n58781;
  assign n58783 = pi17 ? n58767 : n58782;
  assign n58784 = pi16 ? n32 : n58783;
  assign n58785 = pi15 ? n58761 : n58784;
  assign n58786 = pi22 ? n56712 : n49406;
  assign n58787 = pi21 ? n58786 : n39972;
  assign n58788 = pi20 ? n46225 : n58787;
  assign n58789 = pi19 ? n58788 : n38902;
  assign n58790 = pi18 ? n32 : n58789;
  assign n58791 = pi21 ? n39972 : n57185;
  assign n58792 = pi20 ? n36781 : n58791;
  assign n58793 = pi19 ? n36781 : n58792;
  assign n58794 = pi22 ? n36781 : n55622;
  assign n58795 = pi21 ? n58794 : n55560;
  assign n58796 = pi20 ? n36781 : n58795;
  assign n58797 = pi19 ? n58796 : n32;
  assign n58798 = pi18 ? n58793 : n58797;
  assign n58799 = pi17 ? n58790 : n58798;
  assign n58800 = pi16 ? n32 : n58799;
  assign n58801 = pi20 ? n46225 : n55701;
  assign n58802 = pi19 ? n58801 : n56808;
  assign n58803 = pi18 ? n32 : n58802;
  assign n58804 = pi22 ? n36798 : n56607;
  assign n58805 = pi21 ? n58804 : n55560;
  assign n58806 = pi20 ? n36798 : n58805;
  assign n58807 = pi19 ? n58806 : n32;
  assign n58808 = pi18 ? n36798 : n58807;
  assign n58809 = pi17 ? n58803 : n58808;
  assign n58810 = pi16 ? n32 : n58809;
  assign n58811 = pi15 ? n58800 : n58810;
  assign n58812 = pi14 ? n58785 : n58811;
  assign n58813 = pi13 ? n58754 : n58812;
  assign n58814 = pi12 ? n58704 : n58813;
  assign n58815 = pi11 ? n58637 : n58814;
  assign n58816 = pi10 ? n58481 : n58815;
  assign n58817 = pi09 ? n58266 : n58816;
  assign n58818 = pi21 ? n297 : n5623;
  assign n58819 = pi20 ? n31220 : n58818;
  assign n58820 = pi19 ? n20563 : n58819;
  assign n58821 = pi18 ? n20563 : n58820;
  assign n58822 = pi17 ? n45739 : n58821;
  assign n58823 = pi16 ? n32 : n58822;
  assign n58824 = pi15 ? n32 : n58823;
  assign n58825 = pi17 ? n45739 : n58252;
  assign n58826 = pi16 ? n32 : n58825;
  assign n58827 = pi17 ? n50066 : n58258;
  assign n58828 = pi16 ? n32 : n58827;
  assign n58829 = pi15 ? n58826 : n58828;
  assign n58830 = pi14 ? n58824 : n58829;
  assign n58831 = pi13 ? n32 : n58830;
  assign n58832 = pi12 ? n32 : n58831;
  assign n58833 = pi11 ? n32 : n58832;
  assign n58834 = pi10 ? n32 : n58833;
  assign n58835 = pi17 ? n44643 : n58270;
  assign n58836 = pi16 ? n32 : n58835;
  assign n58837 = pi17 ? n44652 : n58276;
  assign n58838 = pi16 ? n32 : n58837;
  assign n58839 = pi15 ? n58836 : n58838;
  assign n58840 = pi17 ? n43674 : n58283;
  assign n58841 = pi16 ? n32 : n58840;
  assign n58842 = pi17 ? n43674 : n58288;
  assign n58843 = pi16 ? n32 : n58842;
  assign n58844 = pi15 ? n58841 : n58843;
  assign n58845 = pi14 ? n58839 : n58844;
  assign n58846 = pi21 ? n4920 : n650;
  assign n58847 = pi20 ? n31220 : n58846;
  assign n58848 = pi19 ? n20563 : n58847;
  assign n58849 = pi18 ? n20563 : n58848;
  assign n58850 = pi17 ? n43674 : n58849;
  assign n58851 = pi16 ? n32 : n58850;
  assign n58852 = pi17 ? n44687 : n58849;
  assign n58853 = pi16 ? n32 : n58852;
  assign n58854 = pi15 ? n58851 : n58853;
  assign n58855 = pi21 ? n4920 : n22919;
  assign n58856 = pi20 ? n31220 : n58855;
  assign n58857 = pi19 ? n20563 : n58856;
  assign n58858 = pi18 ? n20563 : n58857;
  assign n58859 = pi17 ? n44247 : n58858;
  assign n58860 = pi16 ? n32 : n58859;
  assign n58861 = pi21 ? n17806 : n696;
  assign n58862 = pi20 ? n31266 : n58861;
  assign n58863 = pi19 ? n20563 : n58862;
  assign n58864 = pi18 ? n20563 : n58863;
  assign n58865 = pi17 ? n43223 : n58864;
  assign n58866 = pi16 ? n32 : n58865;
  assign n58867 = pi15 ? n58860 : n58866;
  assign n58868 = pi14 ? n58854 : n58867;
  assign n58869 = pi13 ? n58845 : n58868;
  assign n58870 = pi21 ? n17806 : n3494;
  assign n58871 = pi20 ? n31220 : n58870;
  assign n58872 = pi19 ? n20563 : n58871;
  assign n58873 = pi18 ? n20563 : n58872;
  assign n58874 = pi17 ? n48624 : n58873;
  assign n58875 = pi16 ? n32 : n58874;
  assign n58876 = pi24 ? n37 : n685;
  assign n58877 = pi23 ? n58876 : n685;
  assign n58878 = pi22 ? n58877 : n685;
  assign n58879 = pi21 ? n58878 : n696;
  assign n58880 = pi20 ? n31220 : n58879;
  assign n58881 = pi19 ? n20563 : n58880;
  assign n58882 = pi18 ? n20563 : n58881;
  assign n58883 = pi17 ? n48624 : n58882;
  assign n58884 = pi16 ? n32 : n58883;
  assign n58885 = pi15 ? n58875 : n58884;
  assign n58886 = pi17 ? n42645 : n58882;
  assign n58887 = pi16 ? n32 : n58886;
  assign n58888 = pi17 ? n42655 : n58882;
  assign n58889 = pi16 ? n32 : n58888;
  assign n58890 = pi15 ? n58887 : n58889;
  assign n58891 = pi14 ? n58885 : n58890;
  assign n58892 = pi20 ? n20563 : n58879;
  assign n58893 = pi19 ? n20563 : n58892;
  assign n58894 = pi18 ? n20563 : n58893;
  assign n58895 = pi17 ? n42681 : n58894;
  assign n58896 = pi16 ? n32 : n58895;
  assign n58897 = pi17 ? n43262 : n58882;
  assign n58898 = pi16 ? n32 : n58897;
  assign n58899 = pi15 ? n58896 : n58898;
  assign n58900 = pi14 ? n58899 : n58898;
  assign n58901 = pi13 ? n58891 : n58900;
  assign n58902 = pi12 ? n58869 : n58901;
  assign n58903 = pi23 ? n10750 : n316;
  assign n58904 = pi22 ? n58903 : n316;
  assign n58905 = pi21 ? n58904 : n2320;
  assign n58906 = pi20 ? n54354 : n58905;
  assign n58907 = pi19 ? n20563 : n58906;
  assign n58908 = pi18 ? n20563 : n58907;
  assign n58909 = pi17 ? n43262 : n58908;
  assign n58910 = pi16 ? n32 : n58909;
  assign n58911 = pi24 ? n36781 : n316;
  assign n58912 = pi23 ? n58911 : n316;
  assign n58913 = pi22 ? n58912 : n316;
  assign n58914 = pi21 ? n58913 : n2320;
  assign n58915 = pi20 ? n54354 : n58914;
  assign n58916 = pi19 ? n20563 : n58915;
  assign n58917 = pi18 ? n20563 : n58916;
  assign n58918 = pi17 ? n47593 : n58917;
  assign n58919 = pi16 ? n32 : n58918;
  assign n58920 = pi15 ? n58910 : n58919;
  assign n58921 = pi22 ? n22383 : n316;
  assign n58922 = pi21 ? n58921 : n2320;
  assign n58923 = pi20 ? n58395 : n58922;
  assign n58924 = pi19 ? n20563 : n58923;
  assign n58925 = pi18 ? n20563 : n58924;
  assign n58926 = pi17 ? n42207 : n58925;
  assign n58927 = pi16 ? n32 : n58926;
  assign n58928 = pi17 ? n41631 : n58404;
  assign n58929 = pi16 ? n32 : n58928;
  assign n58930 = pi15 ? n58927 : n58929;
  assign n58931 = pi14 ? n58920 : n58930;
  assign n58932 = pi17 ? n41631 : n58412;
  assign n58933 = pi16 ? n32 : n58932;
  assign n58934 = pi17 ? n41631 : n57363;
  assign n58935 = pi16 ? n32 : n58934;
  assign n58936 = pi15 ? n58933 : n58935;
  assign n58937 = pi17 ? n41631 : n57369;
  assign n58938 = pi16 ? n32 : n58937;
  assign n58939 = pi17 ? n41642 : n58422;
  assign n58940 = pi16 ? n32 : n58939;
  assign n58941 = pi15 ? n58938 : n58940;
  assign n58942 = pi14 ? n58936 : n58941;
  assign n58943 = pi13 ? n58931 : n58942;
  assign n58944 = pi21 ? n316 : n53983;
  assign n58945 = pi20 ? n58430 : n58944;
  assign n58946 = pi19 ? n20563 : n58945;
  assign n58947 = pi18 ? n20563 : n58946;
  assign n58948 = pi17 ? n42700 : n58947;
  assign n58949 = pi16 ? n32 : n58948;
  assign n58950 = pi17 ? n40486 : n57966;
  assign n58951 = pi16 ? n32 : n58950;
  assign n58952 = pi15 ? n58949 : n58951;
  assign n58953 = pi17 ? n40486 : n58442;
  assign n58954 = pi16 ? n32 : n58953;
  assign n58955 = pi17 ? n41158 : n58447;
  assign n58956 = pi16 ? n32 : n58955;
  assign n58957 = pi15 ? n58954 : n58956;
  assign n58958 = pi14 ? n58952 : n58957;
  assign n58959 = pi17 ? n41158 : n58457;
  assign n58960 = pi16 ? n32 : n58959;
  assign n58961 = pi17 ? n41169 : n57419;
  assign n58962 = pi16 ? n32 : n58961;
  assign n58963 = pi15 ? n58960 : n58962;
  assign n58964 = pi17 ? n41169 : n58467;
  assign n58965 = pi16 ? n32 : n58964;
  assign n58966 = pi22 ? n51564 : n53982;
  assign n58967 = pi21 ? n58966 : n32;
  assign n58968 = pi20 ? n57432 : n58967;
  assign n58969 = pi19 ? n20563 : n58968;
  assign n58970 = pi18 ? n20563 : n58969;
  assign n58971 = pi17 ? n41182 : n58970;
  assign n58972 = pi16 ? n32 : n58971;
  assign n58973 = pi15 ? n58965 : n58972;
  assign n58974 = pi14 ? n58963 : n58973;
  assign n58975 = pi13 ? n58958 : n58974;
  assign n58976 = pi12 ? n58943 : n58975;
  assign n58977 = pi11 ? n58902 : n58976;
  assign n58978 = pi17 ? n41182 : n58485;
  assign n58979 = pi16 ? n32 : n58978;
  assign n58980 = pi17 ? n41182 : n58492;
  assign n58981 = pi16 ? n32 : n58980;
  assign n58982 = pi15 ? n58979 : n58981;
  assign n58983 = pi17 ? n41182 : n58499;
  assign n58984 = pi16 ? n32 : n58983;
  assign n58985 = pi21 ? n2957 : n6376;
  assign n58986 = pi20 ? n58985 : n58504;
  assign n58987 = pi19 ? n20563 : n58986;
  assign n58988 = pi18 ? n20563 : n58987;
  assign n58989 = pi17 ? n42240 : n58988;
  assign n58990 = pi16 ? n32 : n58989;
  assign n58991 = pi15 ? n58984 : n58990;
  assign n58992 = pi14 ? n58982 : n58991;
  assign n58993 = pi21 ? n50596 : n233;
  assign n58994 = pi20 ? n58993 : n2653;
  assign n58995 = pi19 ? n20563 : n58994;
  assign n58996 = pi18 ? n20563 : n58995;
  assign n58997 = pi17 ? n42240 : n58996;
  assign n58998 = pi16 ? n32 : n58997;
  assign n58999 = pi22 ? n36781 : n685;
  assign n59000 = pi21 ? n47664 : n58999;
  assign n59001 = pi20 ? n59000 : n37640;
  assign n59002 = pi19 ? n20563 : n59001;
  assign n59003 = pi18 ? n20563 : n59002;
  assign n59004 = pi17 ? n42240 : n59003;
  assign n59005 = pi16 ? n32 : n59004;
  assign n59006 = pi15 ? n58998 : n59005;
  assign n59007 = pi17 ? n47057 : n58534;
  assign n59008 = pi16 ? n32 : n59007;
  assign n59009 = pi23 ? n57014 : n204;
  assign n59010 = pi22 ? n59009 : n316;
  assign n59011 = pi21 ? n15050 : n59010;
  assign n59012 = pi20 ? n59011 : n32;
  assign n59013 = pi19 ? n20563 : n59012;
  assign n59014 = pi18 ? n20563 : n59013;
  assign n59015 = pi17 ? n47057 : n59014;
  assign n59016 = pi16 ? n32 : n59015;
  assign n59017 = pi15 ? n59008 : n59016;
  assign n59018 = pi14 ? n59006 : n59017;
  assign n59019 = pi13 ? n58992 : n59018;
  assign n59020 = pi21 ? n30866 : n30868;
  assign n59021 = pi20 ? n32 : n59020;
  assign n59022 = pi19 ? n59021 : n57513;
  assign n59023 = pi18 ? n32 : n59022;
  assign n59024 = pi17 ? n59023 : n58558;
  assign n59025 = pi16 ? n32 : n59024;
  assign n59026 = pi22 ? n56533 : n39190;
  assign n59027 = pi21 ? n30866 : n59026;
  assign n59028 = pi20 ? n32 : n59027;
  assign n59029 = pi20 ? n38754 : n20563;
  assign n59030 = pi19 ? n59028 : n59029;
  assign n59031 = pi18 ? n32 : n59030;
  assign n59032 = pi22 ? n99 : n39976;
  assign n59033 = pi21 ? n59032 : n58568;
  assign n59034 = pi20 ? n59033 : n32;
  assign n59035 = pi19 ? n20563 : n59034;
  assign n59036 = pi18 ? n20563 : n59035;
  assign n59037 = pi17 ? n59031 : n59036;
  assign n59038 = pi16 ? n32 : n59037;
  assign n59039 = pi15 ? n59025 : n59038;
  assign n59040 = pi22 ? n30865 : n40386;
  assign n59041 = pi23 ? n33792 : n55501;
  assign n59042 = pi22 ? n59041 : n39190;
  assign n59043 = pi21 ? n59040 : n59042;
  assign n59044 = pi20 ? n32 : n59043;
  assign n59045 = pi22 ? n36617 : n42109;
  assign n59046 = pi21 ? n52632 : n59045;
  assign n59047 = pi20 ? n59046 : n20563;
  assign n59048 = pi19 ? n59044 : n59047;
  assign n59049 = pi18 ? n32 : n59048;
  assign n59050 = pi17 ? n59049 : n58588;
  assign n59051 = pi16 ? n32 : n59050;
  assign n59052 = pi23 ? n36659 : n55534;
  assign n59053 = pi22 ? n59052 : n37173;
  assign n59054 = pi21 ? n36616 : n59053;
  assign n59055 = pi20 ? n32 : n59054;
  assign n59056 = pi23 ? n37 : n36659;
  assign n59057 = pi22 ? n59056 : n36659;
  assign n59058 = pi21 ? n52758 : n59057;
  assign n59059 = pi20 ? n59058 : n20563;
  assign n59060 = pi19 ? n59055 : n59059;
  assign n59061 = pi18 ? n32 : n59060;
  assign n59062 = pi22 ? n139 : n46796;
  assign n59063 = pi21 ? n59062 : n8486;
  assign n59064 = pi20 ? n59063 : n32;
  assign n59065 = pi19 ? n20563 : n59064;
  assign n59066 = pi18 ? n20563 : n59065;
  assign n59067 = pi17 ? n59061 : n59066;
  assign n59068 = pi16 ? n32 : n59067;
  assign n59069 = pi15 ? n59051 : n59068;
  assign n59070 = pi14 ? n59039 : n59069;
  assign n59071 = pi17 ? n39374 : n58611;
  assign n59072 = pi16 ? n32 : n59071;
  assign n59073 = pi17 ? n40511 : n58618;
  assign n59074 = pi16 ? n32 : n59073;
  assign n59075 = pi15 ? n59072 : n59074;
  assign n59076 = pi17 ? n40511 : n58625;
  assign n59077 = pi16 ? n32 : n59076;
  assign n59078 = pi21 ? n14626 : n53983;
  assign n59079 = pi20 ? n59078 : n32;
  assign n59080 = pi19 ? n58629 : n59079;
  assign n59081 = pi18 ? n20563 : n59080;
  assign n59082 = pi17 ? n41683 : n59081;
  assign n59083 = pi16 ? n32 : n59082;
  assign n59084 = pi15 ? n59077 : n59083;
  assign n59085 = pi14 ? n59075 : n59084;
  assign n59086 = pi13 ? n59070 : n59085;
  assign n59087 = pi12 ? n59019 : n59086;
  assign n59088 = pi19 ? n53368 : n58644;
  assign n59089 = pi18 ? n20563 : n59088;
  assign n59090 = pi17 ? n40498 : n59089;
  assign n59091 = pi16 ? n32 : n59090;
  assign n59092 = pi17 ? n40498 : n57610;
  assign n59093 = pi16 ? n32 : n59092;
  assign n59094 = pi15 ? n59091 : n59093;
  assign n59095 = pi17 ? n40498 : n58656;
  assign n59096 = pi16 ? n32 : n59095;
  assign n59097 = pi20 ? n37926 : n48184;
  assign n59098 = pi19 ? n59097 : n58660;
  assign n59099 = pi18 ? n32 : n59098;
  assign n59100 = pi17 ? n59099 : n58669;
  assign n59101 = pi16 ? n32 : n59100;
  assign n59102 = pi15 ? n59096 : n59101;
  assign n59103 = pi14 ? n59094 : n59102;
  assign n59104 = pi17 ? n47838 : n58680;
  assign n59105 = pi16 ? n32 : n59104;
  assign n59106 = pi17 ? n47838 : n57664;
  assign n59107 = pi16 ? n32 : n59106;
  assign n59108 = pi15 ? n59105 : n59107;
  assign n59109 = pi20 ? n32 : n43010;
  assign n59110 = pi19 ? n59109 : n20563;
  assign n59111 = pi18 ? n32 : n59110;
  assign n59112 = pi18 ? n40793 : n58170;
  assign n59113 = pi17 ? n59111 : n59112;
  assign n59114 = pi16 ? n32 : n59113;
  assign n59115 = pi19 ? n53290 : n30868;
  assign n59116 = pi18 ? n32 : n59115;
  assign n59117 = pi19 ? n41566 : n30868;
  assign n59118 = pi18 ? n59117 : n58698;
  assign n59119 = pi17 ? n59116 : n59118;
  assign n59120 = pi16 ? n32 : n59119;
  assign n59121 = pi15 ? n59114 : n59120;
  assign n59122 = pi14 ? n59108 : n59121;
  assign n59123 = pi13 ? n59103 : n59122;
  assign n59124 = pi20 ? n32 : n46714;
  assign n59125 = pi19 ? n59124 : n30868;
  assign n59126 = pi18 ? n32 : n59125;
  assign n59127 = pi17 ? n59126 : n57702;
  assign n59128 = pi16 ? n32 : n59127;
  assign n59129 = pi22 ? n45634 : n36798;
  assign n59130 = pi21 ? n59129 : n43198;
  assign n59131 = pi20 ? n32 : n59130;
  assign n59132 = pi19 ? n59131 : n56722;
  assign n59133 = pi18 ? n32 : n59132;
  assign n59134 = pi17 ? n59133 : n58717;
  assign n59135 = pi16 ? n32 : n59134;
  assign n59136 = pi15 ? n59128 : n59135;
  assign n59137 = pi22 ? n49720 : n43198;
  assign n59138 = pi21 ? n59137 : n58722;
  assign n59139 = pi20 ? n32 : n59138;
  assign n59140 = pi21 ? n43198 : n55098;
  assign n59141 = pi20 ? n59140 : n58727;
  assign n59142 = pi19 ? n59139 : n59141;
  assign n59143 = pi18 ? n32 : n59142;
  assign n59144 = pi21 ? n52874 : n53471;
  assign n59145 = pi20 ? n58731 : n59144;
  assign n59146 = pi19 ? n58731 : n59145;
  assign n59147 = pi18 ? n59146 : n58741;
  assign n59148 = pi17 ? n59143 : n59147;
  assign n59149 = pi16 ? n32 : n59148;
  assign n59150 = pi19 ? n53479 : n43198;
  assign n59151 = pi18 ? n32 : n59150;
  assign n59152 = pi17 ? n59151 : n58750;
  assign n59153 = pi16 ? n32 : n59152;
  assign n59154 = pi15 ? n59149 : n59153;
  assign n59155 = pi14 ? n59136 : n59154;
  assign n59156 = pi21 ? n43198 : n58470;
  assign n59157 = pi20 ? n51356 : n59156;
  assign n59158 = pi19 ? n59157 : n32;
  assign n59159 = pi18 ? n43198 : n59158;
  assign n59160 = pi17 ? n59151 : n59159;
  assign n59161 = pi16 ? n32 : n59160;
  assign n59162 = pi21 ? n48856 : n36798;
  assign n59163 = pi20 ? n32 : n59162;
  assign n59164 = pi22 ? n36781 : n42171;
  assign n59165 = pi21 ? n36781 : n59164;
  assign n59166 = pi20 ? n59165 : n58764;
  assign n59167 = pi19 ? n59163 : n59166;
  assign n59168 = pi18 ? n32 : n59167;
  assign n59169 = pi21 ? n55143 : n55765;
  assign n59170 = pi20 ? n59169 : n58779;
  assign n59171 = pi19 ? n59170 : n32;
  assign n59172 = pi18 ? n58775 : n59171;
  assign n59173 = pi17 ? n59168 : n59172;
  assign n59174 = pi16 ? n32 : n59173;
  assign n59175 = pi15 ? n59161 : n59174;
  assign n59176 = pi21 ? n57767 : n39972;
  assign n59177 = pi20 ? n32 : n59176;
  assign n59178 = pi19 ? n59177 : n38902;
  assign n59179 = pi18 ? n32 : n59178;
  assign n59180 = pi22 ? n36781 : n53930;
  assign n59181 = pi21 ? n59180 : n55560;
  assign n59182 = pi20 ? n36781 : n59181;
  assign n59183 = pi19 ? n59182 : n32;
  assign n59184 = pi18 ? n58793 : n59183;
  assign n59185 = pi17 ? n59179 : n59184;
  assign n59186 = pi16 ? n32 : n59185;
  assign n59187 = pi21 ? n46772 : n43198;
  assign n59188 = pi20 ? n32 : n59187;
  assign n59189 = pi19 ? n59188 : n56808;
  assign n59190 = pi18 ? n32 : n59189;
  assign n59191 = pi17 ? n59190 : n58808;
  assign n59192 = pi16 ? n32 : n59191;
  assign n59193 = pi15 ? n59186 : n59192;
  assign n59194 = pi14 ? n59175 : n59193;
  assign n59195 = pi13 ? n59155 : n59194;
  assign n59196 = pi12 ? n59123 : n59195;
  assign n59197 = pi11 ? n59087 : n59196;
  assign n59198 = pi10 ? n58977 : n59197;
  assign n59199 = pi09 ? n58834 : n59198;
  assign n59200 = pi08 ? n58817 : n59199;
  assign n59201 = pi07 ? n58241 : n59200;
  assign n59202 = pi06 ? n57213 : n59201;
  assign n59203 = pi21 ? n1721 : n12243;
  assign n59204 = pi20 ? n31220 : n59203;
  assign n59205 = pi19 ? n38478 : n59204;
  assign n59206 = pi18 ? n38316 : n59205;
  assign n59207 = pi17 ? n32 : n59206;
  assign n59208 = pi16 ? n32 : n59207;
  assign n59209 = pi15 ? n32 : n59208;
  assign n59210 = pi19 ? n20563 : n59204;
  assign n59211 = pi18 ? n20563 : n59210;
  assign n59212 = pi17 ? n46325 : n59211;
  assign n59213 = pi16 ? n32 : n59212;
  assign n59214 = pi21 ? n1721 : n19777;
  assign n59215 = pi20 ? n30096 : n59214;
  assign n59216 = pi19 ? n38478 : n59215;
  assign n59217 = pi18 ? n20563 : n59216;
  assign n59218 = pi17 ? n46325 : n59217;
  assign n59219 = pi16 ? n32 : n59218;
  assign n59220 = pi15 ? n59213 : n59219;
  assign n59221 = pi14 ? n59209 : n59220;
  assign n59222 = pi13 ? n32 : n59221;
  assign n59223 = pi12 ? n32 : n59222;
  assign n59224 = pi11 ? n32 : n59223;
  assign n59225 = pi10 ? n32 : n59224;
  assign n59226 = pi22 ? n335 : n1370;
  assign n59227 = pi21 ? n4938 : n59226;
  assign n59228 = pi20 ? n31220 : n59227;
  assign n59229 = pi19 ? n20563 : n59228;
  assign n59230 = pi18 ? n20563 : n59229;
  assign n59231 = pi17 ? n45232 : n59230;
  assign n59232 = pi16 ? n32 : n59231;
  assign n59233 = pi22 ? n335 : n1378;
  assign n59234 = pi21 ? n4938 : n59233;
  assign n59235 = pi20 ? n31220 : n59234;
  assign n59236 = pi19 ? n20563 : n59235;
  assign n59237 = pi18 ? n20563 : n59236;
  assign n59238 = pi17 ? n44634 : n59237;
  assign n59239 = pi16 ? n32 : n59238;
  assign n59240 = pi15 ? n59232 : n59239;
  assign n59241 = pi21 ? n4938 : n20793;
  assign n59242 = pi20 ? n20563 : n59241;
  assign n59243 = pi19 ? n20563 : n59242;
  assign n59244 = pi18 ? n20563 : n59243;
  assign n59245 = pi17 ? n44222 : n59244;
  assign n59246 = pi16 ? n32 : n59245;
  assign n59247 = pi22 ? n1656 : n335;
  assign n59248 = pi21 ? n59247 : n588;
  assign n59249 = pi20 ? n20563 : n59248;
  assign n59250 = pi19 ? n20563 : n59249;
  assign n59251 = pi18 ? n20563 : n59250;
  assign n59252 = pi17 ? n44222 : n59251;
  assign n59253 = pi16 ? n32 : n59252;
  assign n59254 = pi15 ? n59246 : n59253;
  assign n59255 = pi14 ? n59240 : n59254;
  assign n59256 = pi22 ? n13278 : n335;
  assign n59257 = pi21 ? n59256 : n588;
  assign n59258 = pi20 ? n31220 : n59257;
  assign n59259 = pi19 ? n20563 : n59258;
  assign n59260 = pi18 ? n20563 : n59259;
  assign n59261 = pi17 ? n45242 : n59260;
  assign n59262 = pi16 ? n32 : n59261;
  assign n59263 = pi17 ? n46348 : n59260;
  assign n59264 = pi16 ? n32 : n59263;
  assign n59265 = pi15 ? n59262 : n59264;
  assign n59266 = pi17 ? n44670 : n59260;
  assign n59267 = pi16 ? n32 : n59266;
  assign n59268 = pi17 ? n43674 : n59260;
  assign n59269 = pi16 ? n32 : n59268;
  assign n59270 = pi15 ? n59267 : n59269;
  assign n59271 = pi14 ? n59265 : n59270;
  assign n59272 = pi13 ? n59255 : n59271;
  assign n59273 = pi22 ? n57882 : n363;
  assign n59274 = pi22 ? n363 : n5631;
  assign n59275 = pi21 ? n59273 : n59274;
  assign n59276 = pi20 ? n20563 : n59275;
  assign n59277 = pi19 ? n20563 : n59276;
  assign n59278 = pi18 ? n20563 : n59277;
  assign n59279 = pi17 ? n43223 : n59278;
  assign n59280 = pi16 ? n32 : n59279;
  assign n59281 = pi23 ? n31328 : n157;
  assign n59282 = pi22 ? n59281 : n157;
  assign n59283 = pi21 ? n59282 : n11928;
  assign n59284 = pi20 ? n31220 : n59283;
  assign n59285 = pi19 ? n20563 : n59284;
  assign n59286 = pi18 ? n20563 : n59285;
  assign n59287 = pi17 ? n43223 : n59286;
  assign n59288 = pi16 ? n32 : n59287;
  assign n59289 = pi17 ? n43227 : n59286;
  assign n59290 = pi16 ? n32 : n59289;
  assign n59291 = pi15 ? n59288 : n59290;
  assign n59292 = pi14 ? n59280 : n59291;
  assign n59293 = pi22 ? n32905 : n204;
  assign n59294 = pi21 ? n59293 : n4748;
  assign n59295 = pi20 ? n20563 : n59294;
  assign n59296 = pi19 ? n20563 : n59295;
  assign n59297 = pi18 ? n20563 : n59296;
  assign n59298 = pi17 ? n43248 : n59297;
  assign n59299 = pi16 ? n32 : n59298;
  assign n59300 = pi17 ? n48624 : n59297;
  assign n59301 = pi16 ? n32 : n59300;
  assign n59302 = pi15 ? n59299 : n59301;
  assign n59303 = pi23 ? n11127 : n233;
  assign n59304 = pi22 ? n59303 : n233;
  assign n59305 = pi21 ? n59304 : n650;
  assign n59306 = pi20 ? n20563 : n59305;
  assign n59307 = pi19 ? n20563 : n59306;
  assign n59308 = pi18 ? n20563 : n59307;
  assign n59309 = pi17 ? n48624 : n59308;
  assign n59310 = pi16 ? n32 : n59309;
  assign n59311 = pi23 ? n11127 : n685;
  assign n59312 = pi22 ? n59311 : n685;
  assign n59313 = pi21 ? n59312 : n696;
  assign n59314 = pi20 ? n20563 : n59313;
  assign n59315 = pi19 ? n20563 : n59314;
  assign n59316 = pi18 ? n20563 : n59315;
  assign n59317 = pi17 ? n48624 : n59316;
  assign n59318 = pi16 ? n32 : n59317;
  assign n59319 = pi15 ? n59310 : n59318;
  assign n59320 = pi14 ? n59302 : n59319;
  assign n59321 = pi13 ? n59292 : n59320;
  assign n59322 = pi12 ? n59272 : n59321;
  assign n59323 = pi23 ? n7420 : n685;
  assign n59324 = pi22 ? n59323 : n685;
  assign n59325 = pi21 ? n59324 : n7723;
  assign n59326 = pi20 ? n54354 : n59325;
  assign n59327 = pi19 ? n20563 : n59326;
  assign n59328 = pi18 ? n20563 : n59327;
  assign n59329 = pi17 ? n42645 : n59328;
  assign n59330 = pi16 ? n32 : n59329;
  assign n59331 = pi20 ? n54354 : n58922;
  assign n59332 = pi19 ? n20563 : n59331;
  assign n59333 = pi18 ? n20563 : n59332;
  assign n59334 = pi17 ? n42655 : n59333;
  assign n59335 = pi16 ? n32 : n59334;
  assign n59336 = pi15 ? n59330 : n59335;
  assign n59337 = pi17 ? n42681 : n58925;
  assign n59338 = pi16 ? n32 : n59337;
  assign n59339 = pi22 ? n37 : n37218;
  assign n59340 = pi21 ? n20563 : n59339;
  assign n59341 = pi23 ? n14626 : n32;
  assign n59342 = pi22 ? n59341 : n32;
  assign n59343 = pi21 ? n204 : n59342;
  assign n59344 = pi20 ? n59340 : n59343;
  assign n59345 = pi19 ? n20563 : n59344;
  assign n59346 = pi18 ? n20563 : n59345;
  assign n59347 = pi17 ? n42201 : n59346;
  assign n59348 = pi16 ? n32 : n59347;
  assign n59349 = pi15 ? n59338 : n59348;
  assign n59350 = pi14 ? n59336 : n59349;
  assign n59351 = pi21 ? n14626 : n2637;
  assign n59352 = pi20 ? n56350 : n59351;
  assign n59353 = pi19 ? n20563 : n59352;
  assign n59354 = pi18 ? n20563 : n59353;
  assign n59355 = pi17 ? n42201 : n59354;
  assign n59356 = pi16 ? n32 : n59355;
  assign n59357 = pi22 ? n58452 : n32;
  assign n59358 = pi21 ? n14626 : n59357;
  assign n59359 = pi20 ? n56361 : n59358;
  assign n59360 = pi19 ? n20563 : n59359;
  assign n59361 = pi18 ? n20563 : n59360;
  assign n59362 = pi17 ? n42201 : n59361;
  assign n59363 = pi16 ? n32 : n59362;
  assign n59364 = pi15 ? n59356 : n59363;
  assign n59365 = pi22 ? n37 : n59056;
  assign n59366 = pi21 ? n20563 : n59365;
  assign n59367 = pi21 ? n51564 : n928;
  assign n59368 = pi20 ? n59366 : n59367;
  assign n59369 = pi19 ? n20563 : n59368;
  assign n59370 = pi18 ? n20563 : n59369;
  assign n59371 = pi17 ? n42201 : n59370;
  assign n59372 = pi16 ? n32 : n59371;
  assign n59373 = pi21 ? n51564 : n37639;
  assign n59374 = pi20 ? n56374 : n59373;
  assign n59375 = pi19 ? n20563 : n59374;
  assign n59376 = pi18 ? n20563 : n59375;
  assign n59377 = pi17 ? n48121 : n59376;
  assign n59378 = pi16 ? n32 : n59377;
  assign n59379 = pi15 ? n59372 : n59378;
  assign n59380 = pi14 ? n59364 : n59379;
  assign n59381 = pi13 ? n59350 : n59380;
  assign n59382 = pi21 ? n13481 : n53983;
  assign n59383 = pi20 ? n55343 : n59382;
  assign n59384 = pi19 ? n20563 : n59383;
  assign n59385 = pi18 ? n20563 : n59384;
  assign n59386 = pi17 ? n47593 : n59385;
  assign n59387 = pi16 ? n32 : n59386;
  assign n59388 = pi21 ? n13481 : n1009;
  assign n59389 = pi20 ? n56389 : n59388;
  assign n59390 = pi19 ? n20563 : n59389;
  assign n59391 = pi18 ? n20563 : n59390;
  assign n59392 = pi17 ? n42207 : n59391;
  assign n59393 = pi16 ? n32 : n59392;
  assign n59394 = pi15 ? n59387 : n59393;
  assign n59395 = pi23 ? n14626 : n687;
  assign n59396 = pi22 ? n204 : n59395;
  assign n59397 = pi21 ? n59396 : n32;
  assign n59398 = pi20 ? n56397 : n59397;
  assign n59399 = pi19 ? n20563 : n59398;
  assign n59400 = pi18 ? n20563 : n59399;
  assign n59401 = pi17 ? n42207 : n59400;
  assign n59402 = pi16 ? n32 : n59401;
  assign n59403 = pi17 ? n42207 : n56406;
  assign n59404 = pi16 ? n32 : n59403;
  assign n59405 = pi15 ? n59402 : n59404;
  assign n59406 = pi14 ? n59394 : n59405;
  assign n59407 = pi20 ? n56411 : n58454;
  assign n59408 = pi19 ? n20563 : n59407;
  assign n59409 = pi18 ? n20563 : n59408;
  assign n59410 = pi17 ? n42207 : n59409;
  assign n59411 = pi16 ? n32 : n59410;
  assign n59412 = pi23 ? n36659 : n14626;
  assign n59413 = pi22 ? n20563 : n59412;
  assign n59414 = pi21 ? n20563 : n59413;
  assign n59415 = pi22 ? n14626 : n317;
  assign n59416 = pi21 ? n59415 : n32;
  assign n59417 = pi20 ? n59414 : n59416;
  assign n59418 = pi19 ? n20563 : n59417;
  assign n59419 = pi18 ? n20563 : n59418;
  assign n59420 = pi17 ? n42688 : n59419;
  assign n59421 = pi16 ? n32 : n59420;
  assign n59422 = pi15 ? n59411 : n59421;
  assign n59423 = pi23 ? n36781 : n685;
  assign n59424 = pi22 ? n99 : n59423;
  assign n59425 = pi21 ? n20563 : n59424;
  assign n59426 = pi20 ? n59425 : n57434;
  assign n59427 = pi19 ? n20563 : n59426;
  assign n59428 = pi18 ? n20563 : n59427;
  assign n59429 = pi17 ? n42688 : n59428;
  assign n59430 = pi16 ? n32 : n59429;
  assign n59431 = pi22 ? n30868 : n51564;
  assign n59432 = pi21 ? n20563 : n59431;
  assign n59433 = pi20 ? n59432 : n54547;
  assign n59434 = pi19 ? n20563 : n59433;
  assign n59435 = pi18 ? n20563 : n59434;
  assign n59436 = pi17 ? n42700 : n59435;
  assign n59437 = pi16 ? n32 : n59436;
  assign n59438 = pi15 ? n59430 : n59437;
  assign n59439 = pi14 ? n59422 : n59438;
  assign n59440 = pi13 ? n59406 : n59439;
  assign n59441 = pi12 ? n59381 : n59440;
  assign n59442 = pi11 ? n59322 : n59441;
  assign n59443 = pi20 ? n58489 : n55668;
  assign n59444 = pi19 ? n40792 : n59443;
  assign n59445 = pi18 ? n20563 : n59444;
  assign n59446 = pi17 ? n42700 : n59445;
  assign n59447 = pi16 ? n32 : n59446;
  assign n59448 = pi21 ? n20563 : n204;
  assign n59449 = pi23 ? n14626 : n51565;
  assign n59450 = pi22 ? n59449 : n32;
  assign n59451 = pi21 ? n59450 : n32;
  assign n59452 = pi20 ? n59448 : n59451;
  assign n59453 = pi19 ? n40792 : n59452;
  assign n59454 = pi18 ? n20563 : n59453;
  assign n59455 = pi17 ? n46998 : n59454;
  assign n59456 = pi16 ? n32 : n59455;
  assign n59457 = pi15 ? n59447 : n59456;
  assign n59458 = pi20 ? n20563 : n53326;
  assign n59459 = pi21 ? n36489 : n14626;
  assign n59460 = pi20 ? n59459 : n5830;
  assign n59461 = pi19 ? n59458 : n59460;
  assign n59462 = pi18 ? n20563 : n59461;
  assign n59463 = pi17 ? n46998 : n59462;
  assign n59464 = pi16 ? n32 : n59463;
  assign n59465 = pi21 ? n2957 : n14626;
  assign n59466 = pi21 ? n59357 : n32;
  assign n59467 = pi20 ? n59465 : n59466;
  assign n59468 = pi19 ? n20563 : n59467;
  assign n59469 = pi18 ? n20563 : n59468;
  assign n59470 = pi17 ? n40486 : n59469;
  assign n59471 = pi16 ? n32 : n59470;
  assign n59472 = pi15 ? n59464 : n59471;
  assign n59473 = pi14 ? n59457 : n59472;
  assign n59474 = pi21 ? n59339 : n685;
  assign n59475 = pi20 ? n59474 : n2653;
  assign n59476 = pi19 ? n20563 : n59475;
  assign n59477 = pi18 ? n20563 : n59476;
  assign n59478 = pi17 ? n40486 : n59477;
  assign n59479 = pi16 ? n32 : n59478;
  assign n59480 = pi21 ? n33792 : n13481;
  assign n59481 = pi20 ? n59480 : n2701;
  assign n59482 = pi19 ? n47159 : n59481;
  assign n59483 = pi18 ? n20563 : n59482;
  assign n59484 = pi17 ? n41169 : n59483;
  assign n59485 = pi16 ? n32 : n59484;
  assign n59486 = pi15 ? n59479 : n59485;
  assign n59487 = pi22 ? n58529 : n316;
  assign n59488 = pi21 ? n36659 : n59487;
  assign n59489 = pi20 ? n59488 : n1822;
  assign n59490 = pi19 ? n56631 : n59489;
  assign n59491 = pi18 ? n20563 : n59490;
  assign n59492 = pi17 ? n41169 : n59491;
  assign n59493 = pi16 ? n32 : n59492;
  assign n59494 = pi19 ? n56687 : n40791;
  assign n59495 = pi18 ? n32 : n59494;
  assign n59496 = pi20 ? n43010 : n55475;
  assign n59497 = pi23 ? n8319 : n204;
  assign n59498 = pi22 ? n59497 : n13481;
  assign n59499 = pi21 ? n36659 : n59498;
  assign n59500 = pi20 ? n59499 : n32;
  assign n59501 = pi19 ? n59496 : n59500;
  assign n59502 = pi18 ? n20563 : n59501;
  assign n59503 = pi17 ? n59495 : n59502;
  assign n59504 = pi16 ? n32 : n59503;
  assign n59505 = pi15 ? n59493 : n59504;
  assign n59506 = pi14 ? n59486 : n59505;
  assign n59507 = pi13 ? n59473 : n59506;
  assign n59508 = pi21 ? n39394 : n37768;
  assign n59509 = pi20 ? n32 : n59508;
  assign n59510 = pi20 ? n53326 : n54468;
  assign n59511 = pi19 ? n59509 : n59510;
  assign n59512 = pi18 ? n32 : n59511;
  assign n59513 = pi20 ? n33792 : n56539;
  assign n59514 = pi22 ? n58553 : n58452;
  assign n59515 = pi21 ? n36781 : n59514;
  assign n59516 = pi20 ? n59515 : n32;
  assign n59517 = pi19 ? n59513 : n59516;
  assign n59518 = pi18 ? n20563 : n59517;
  assign n59519 = pi17 ? n59512 : n59518;
  assign n59520 = pi16 ? n32 : n59519;
  assign n59521 = pi19 ? n59509 : n20563;
  assign n59522 = pi18 ? n32 : n59521;
  assign n59523 = pi20 ? n47280 : n20563;
  assign n59524 = pi22 ? n30868 : n36798;
  assign n59525 = pi23 ? n35938 : n233;
  assign n59526 = pi22 ? n59525 : n317;
  assign n59527 = pi21 ? n59524 : n59526;
  assign n59528 = pi20 ? n59527 : n32;
  assign n59529 = pi19 ? n59523 : n59528;
  assign n59530 = pi18 ? n20563 : n59529;
  assign n59531 = pi17 ? n59522 : n59530;
  assign n59532 = pi16 ? n32 : n59531;
  assign n59533 = pi15 ? n59520 : n59532;
  assign n59534 = pi21 ? n39394 : n37784;
  assign n59535 = pi20 ? n32 : n59534;
  assign n59536 = pi19 ? n59535 : n20563;
  assign n59537 = pi18 ? n32 : n59536;
  assign n59538 = pi20 ? n47280 : n38754;
  assign n59539 = pi22 ? n14626 : n53982;
  assign n59540 = pi21 ? n36798 : n59539;
  assign n59541 = pi20 ? n59540 : n32;
  assign n59542 = pi19 ? n59538 : n59541;
  assign n59543 = pi18 ? n20563 : n59542;
  assign n59544 = pi17 ? n59537 : n59543;
  assign n59545 = pi16 ? n32 : n59544;
  assign n59546 = pi21 ? n45620 : n20563;
  assign n59547 = pi20 ? n32 : n59546;
  assign n59548 = pi19 ? n59547 : n20563;
  assign n59549 = pi18 ? n32 : n59548;
  assign n59550 = pi21 ? n45049 : n39801;
  assign n59551 = pi20 ? n59550 : n51188;
  assign n59552 = pi19 ? n59551 : n42915;
  assign n59553 = pi21 ? n46116 : n36489;
  assign n59554 = pi20 ? n20563 : n59553;
  assign n59555 = pi22 ? n33792 : n204;
  assign n59556 = pi21 ? n59555 : n57563;
  assign n59557 = pi20 ? n59556 : n32;
  assign n59558 = pi19 ? n59554 : n59557;
  assign n59559 = pi18 ? n59552 : n59558;
  assign n59560 = pi17 ? n59549 : n59559;
  assign n59561 = pi16 ? n32 : n59560;
  assign n59562 = pi15 ? n59545 : n59561;
  assign n59563 = pi14 ? n59533 : n59562;
  assign n59564 = pi21 ? n43198 : n2320;
  assign n59565 = pi20 ? n59564 : n32;
  assign n59566 = pi19 ? n42915 : n59565;
  assign n59567 = pi18 ? n20563 : n59566;
  assign n59568 = pi17 ? n47057 : n59567;
  assign n59569 = pi16 ? n32 : n59568;
  assign n59570 = pi21 ? n14626 : n2320;
  assign n59571 = pi20 ? n59570 : n32;
  assign n59572 = pi19 ? n47159 : n59571;
  assign n59573 = pi18 ? n20563 : n59572;
  assign n59574 = pi17 ? n40024 : n59573;
  assign n59575 = pi16 ? n32 : n59574;
  assign n59576 = pi15 ? n59569 : n59575;
  assign n59577 = pi21 ? n14626 : n2700;
  assign n59578 = pi20 ? n59577 : n32;
  assign n59579 = pi19 ? n47159 : n59578;
  assign n59580 = pi18 ? n20563 : n59579;
  assign n59581 = pi17 ? n40024 : n59580;
  assign n59582 = pi16 ? n32 : n59581;
  assign n59583 = pi21 ? n51564 : n53983;
  assign n59584 = pi20 ? n59583 : n32;
  assign n59585 = pi19 ? n55476 : n59584;
  assign n59586 = pi18 ? n20563 : n59585;
  assign n59587 = pi17 ? n41182 : n59586;
  assign n59588 = pi16 ? n32 : n59587;
  assign n59589 = pi15 ? n59582 : n59588;
  assign n59590 = pi14 ? n59576 : n59589;
  assign n59591 = pi13 ? n59563 : n59590;
  assign n59592 = pi12 ? n59507 : n59591;
  assign n59593 = pi21 ? n20563 : n55685;
  assign n59594 = pi20 ? n20563 : n59593;
  assign n59595 = pi22 ? n14626 : n51564;
  assign n59596 = pi21 ? n59595 : n1009;
  assign n59597 = pi20 ? n59596 : n32;
  assign n59598 = pi19 ? n59594 : n59597;
  assign n59599 = pi18 ? n20563 : n59598;
  assign n59600 = pi17 ? n41182 : n59599;
  assign n59601 = pi16 ? n32 : n59600;
  assign n59602 = pi21 ? n20563 : n39952;
  assign n59603 = pi20 ? n20563 : n59602;
  assign n59604 = pi21 ? n13481 : n32;
  assign n59605 = pi20 ? n59604 : n32;
  assign n59606 = pi19 ? n59603 : n59605;
  assign n59607 = pi18 ? n20563 : n59606;
  assign n59608 = pi17 ? n41182 : n59607;
  assign n59609 = pi16 ? n32 : n59608;
  assign n59610 = pi15 ? n59601 : n59609;
  assign n59611 = pi21 ? n28156 : n45049;
  assign n59612 = pi20 ? n32 : n59611;
  assign n59613 = pi19 ? n59612 : n40791;
  assign n59614 = pi18 ? n32 : n59613;
  assign n59615 = pi20 ? n36489 : n42006;
  assign n59616 = pi20 ? n40915 : n43010;
  assign n59617 = pi19 ? n59615 : n59616;
  assign n59618 = pi22 ? n33792 : n40004;
  assign n59619 = pi21 ? n36489 : n59618;
  assign n59620 = pi20 ? n40915 : n59619;
  assign n59621 = pi22 ? n51564 : n58452;
  assign n59622 = pi21 ? n59621 : n32;
  assign n59623 = pi20 ? n59622 : n32;
  assign n59624 = pi19 ? n59620 : n59623;
  assign n59625 = pi18 ? n59617 : n59624;
  assign n59626 = pi17 ? n59614 : n59625;
  assign n59627 = pi16 ? n32 : n59626;
  assign n59628 = pi21 ? n58125 : n30868;
  assign n59629 = pi20 ? n32 : n59628;
  assign n59630 = pi19 ? n59629 : n30868;
  assign n59631 = pi18 ? n32 : n59630;
  assign n59632 = pi21 ? n30868 : n46260;
  assign n59633 = pi20 ? n30868 : n59632;
  assign n59634 = pi22 ? n13481 : n317;
  assign n59635 = pi21 ? n59634 : n32;
  assign n59636 = pi20 ? n59635 : n32;
  assign n59637 = pi19 ? n59633 : n59636;
  assign n59638 = pi18 ? n30868 : n59637;
  assign n59639 = pi17 ? n59631 : n59638;
  assign n59640 = pi16 ? n32 : n59639;
  assign n59641 = pi15 ? n59627 : n59640;
  assign n59642 = pi14 ? n59610 : n59641;
  assign n59643 = pi20 ? n32 : n58144;
  assign n59644 = pi19 ? n59643 : n30868;
  assign n59645 = pi18 ? n32 : n59644;
  assign n59646 = pi21 ? n30868 : n50795;
  assign n59647 = pi20 ? n30868 : n59646;
  assign n59648 = pi22 ? n13481 : n21502;
  assign n59649 = pi21 ? n59648 : n32;
  assign n59650 = pi20 ? n59649 : n32;
  assign n59651 = pi19 ? n59647 : n59650;
  assign n59652 = pi18 ? n30868 : n59651;
  assign n59653 = pi17 ? n59645 : n59652;
  assign n59654 = pi16 ? n32 : n59653;
  assign n59655 = pi21 ? n59524 : n57774;
  assign n59656 = pi20 ? n30868 : n59655;
  assign n59657 = pi22 ? n59395 : n32;
  assign n59658 = pi21 ? n59657 : n32;
  assign n59659 = pi20 ? n59658 : n32;
  assign n59660 = pi19 ? n59656 : n59659;
  assign n59661 = pi18 ? n30868 : n59660;
  assign n59662 = pi17 ? n59645 : n59661;
  assign n59663 = pi16 ? n32 : n59662;
  assign n59664 = pi15 ? n59654 : n59663;
  assign n59665 = pi21 ? n37332 : n36489;
  assign n59666 = pi20 ? n32 : n59665;
  assign n59667 = pi20 ? n40791 : n30868;
  assign n59668 = pi19 ? n59666 : n59667;
  assign n59669 = pi18 ? n32 : n59668;
  assign n59670 = pi21 ? n36659 : n55708;
  assign n59671 = pi20 ? n30868 : n59670;
  assign n59672 = pi23 ? n51564 : n51565;
  assign n59673 = pi22 ? n59672 : n32;
  assign n59674 = pi21 ? n59673 : n32;
  assign n59675 = pi20 ? n59674 : n32;
  assign n59676 = pi19 ? n59671 : n59675;
  assign n59677 = pi18 ? n30868 : n59676;
  assign n59678 = pi17 ? n59669 : n59677;
  assign n59679 = pi16 ? n32 : n59678;
  assign n59680 = pi18 ? n32 : n53953;
  assign n59681 = pi22 ? n36798 : n51564;
  assign n59682 = pi21 ? n50338 : n59681;
  assign n59683 = pi20 ? n30868 : n59682;
  assign n59684 = pi19 ? n59683 : n54566;
  assign n59685 = pi18 ? n30868 : n59684;
  assign n59686 = pi17 ? n59680 : n59685;
  assign n59687 = pi16 ? n32 : n59686;
  assign n59688 = pi15 ? n59679 : n59687;
  assign n59689 = pi14 ? n59664 : n59688;
  assign n59690 = pi13 ? n59642 : n59689;
  assign n59691 = pi22 ? n43198 : n13481;
  assign n59692 = pi21 ? n43198 : n59691;
  assign n59693 = pi20 ? n30868 : n59692;
  assign n59694 = pi19 ? n59693 : n37641;
  assign n59695 = pi18 ? n30868 : n59694;
  assign n59696 = pi17 ? n59680 : n59695;
  assign n59697 = pi16 ? n32 : n59696;
  assign n59698 = pi21 ? n46276 : n55715;
  assign n59699 = pi20 ? n32 : n59698;
  assign n59700 = pi20 ? n49401 : n43198;
  assign n59701 = pi19 ? n59699 : n59700;
  assign n59702 = pi18 ? n32 : n59701;
  assign n59703 = pi21 ? n46280 : n43198;
  assign n59704 = pi20 ? n59703 : n54655;
  assign n59705 = pi21 ? n47396 : n53471;
  assign n59706 = pi21 ? n36659 : n43198;
  assign n59707 = pi20 ? n59705 : n59706;
  assign n59708 = pi19 ? n59704 : n59707;
  assign n59709 = pi20 ? n54591 : n59692;
  assign n59710 = pi19 ? n59709 : n32;
  assign n59711 = pi18 ? n59708 : n59710;
  assign n59712 = pi17 ? n59702 : n59711;
  assign n59713 = pi16 ? n32 : n59712;
  assign n59714 = pi15 ? n59697 : n59713;
  assign n59715 = pi21 ? n55516 : n33792;
  assign n59716 = pi20 ? n32 : n59715;
  assign n59717 = pi19 ? n59716 : n33792;
  assign n59718 = pi18 ? n32 : n59717;
  assign n59719 = pi23 ? n204 : n43198;
  assign n59720 = pi22 ? n59719 : n13481;
  assign n59721 = pi21 ? n43198 : n59720;
  assign n59722 = pi20 ? n33792 : n59721;
  assign n59723 = pi19 ? n59722 : n32;
  assign n59724 = pi18 ? n33792 : n59723;
  assign n59725 = pi17 ? n59718 : n59724;
  assign n59726 = pi16 ? n32 : n59725;
  assign n59727 = pi21 ? n32 : n50338;
  assign n59728 = pi20 ? n32 : n59727;
  assign n59729 = pi20 ? n46284 : n43198;
  assign n59730 = pi19 ? n59728 : n59729;
  assign n59731 = pi18 ? n32 : n59730;
  assign n59732 = pi20 ? n43198 : n55701;
  assign n59733 = pi19 ? n43198 : n59732;
  assign n59734 = pi21 ? n43198 : n59415;
  assign n59735 = pi20 ? n43198 : n59734;
  assign n59736 = pi19 ? n59735 : n32;
  assign n59737 = pi18 ? n59733 : n59736;
  assign n59738 = pi17 ? n59731 : n59737;
  assign n59739 = pi16 ? n32 : n59738;
  assign n59740 = pi15 ? n59726 : n59739;
  assign n59741 = pi14 ? n59714 : n59740;
  assign n59742 = pi20 ? n54009 : n43198;
  assign n59743 = pi19 ? n59728 : n59742;
  assign n59744 = pi18 ? n32 : n59743;
  assign n59745 = pi21 ? n55717 : n57433;
  assign n59746 = pi20 ? n43198 : n59745;
  assign n59747 = pi19 ? n59746 : n32;
  assign n59748 = pi18 ? n43198 : n59747;
  assign n59749 = pi17 ? n59744 : n59748;
  assign n59750 = pi16 ? n32 : n59749;
  assign n59751 = pi22 ? n45634 : n36781;
  assign n59752 = pi21 ? n32 : n59751;
  assign n59753 = pi20 ? n32 : n59752;
  assign n59754 = pi19 ? n59753 : n43198;
  assign n59755 = pi18 ? n32 : n59754;
  assign n59756 = pi21 ? n56760 : n58778;
  assign n59757 = pi20 ? n43198 : n59756;
  assign n59758 = pi19 ? n59757 : n32;
  assign n59759 = pi18 ? n43198 : n59758;
  assign n59760 = pi17 ? n59755 : n59759;
  assign n59761 = pi16 ? n32 : n59760;
  assign n59762 = pi15 ? n59750 : n59761;
  assign n59763 = pi22 ? n53550 : n36781;
  assign n59764 = pi21 ? n59763 : n36781;
  assign n59765 = pi22 ? n58221 : n36798;
  assign n59766 = pi21 ? n46283 : n59765;
  assign n59767 = pi20 ? n59764 : n59766;
  assign n59768 = pi19 ? n45664 : n59767;
  assign n59769 = pi18 ? n32 : n59768;
  assign n59770 = pi20 ? n46289 : n38901;
  assign n59771 = pi20 ? n38901 : n45140;
  assign n59772 = pi19 ? n59770 : n59771;
  assign n59773 = pi21 ? n39972 : n38901;
  assign n59774 = pi22 ? n36798 : n13481;
  assign n59775 = pi21 ? n59774 : n55560;
  assign n59776 = pi20 ? n59773 : n59775;
  assign n59777 = pi19 ? n59776 : n32;
  assign n59778 = pi18 ? n59772 : n59777;
  assign n59779 = pi17 ? n59769 : n59778;
  assign n59780 = pi16 ? n32 : n59779;
  assign n59781 = pi20 ? n47398 : n49401;
  assign n59782 = pi19 ? n45671 : n59781;
  assign n59783 = pi18 ? n32 : n59782;
  assign n59784 = pi23 ? n316 : n13481;
  assign n59785 = pi22 ? n59784 : n32;
  assign n59786 = pi21 ? n59691 : n59785;
  assign n59787 = pi20 ? n55701 : n59786;
  assign n59788 = pi19 ? n59787 : n32;
  assign n59789 = pi18 ? n54659 : n59788;
  assign n59790 = pi17 ? n59783 : n59789;
  assign n59791 = pi16 ? n32 : n59790;
  assign n59792 = pi15 ? n59780 : n59791;
  assign n59793 = pi14 ? n59762 : n59792;
  assign n59794 = pi13 ? n59741 : n59793;
  assign n59795 = pi12 ? n59690 : n59794;
  assign n59796 = pi11 ? n59592 : n59795;
  assign n59797 = pi10 ? n59442 : n59796;
  assign n59798 = pi09 ? n59225 : n59797;
  assign n59799 = pi18 ? n45392 : n59205;
  assign n59800 = pi17 ? n32 : n59799;
  assign n59801 = pi16 ? n32 : n59800;
  assign n59802 = pi15 ? n32 : n59801;
  assign n59803 = pi18 ? n45392 : n59210;
  assign n59804 = pi17 ? n32 : n59803;
  assign n59805 = pi16 ? n32 : n59804;
  assign n59806 = pi18 ? n45392 : n59216;
  assign n59807 = pi17 ? n32 : n59806;
  assign n59808 = pi16 ? n32 : n59807;
  assign n59809 = pi15 ? n59805 : n59808;
  assign n59810 = pi14 ? n59802 : n59809;
  assign n59811 = pi13 ? n32 : n59810;
  assign n59812 = pi12 ? n32 : n59811;
  assign n59813 = pi11 ? n32 : n59812;
  assign n59814 = pi10 ? n32 : n59813;
  assign n59815 = pi18 ? n45413 : n59229;
  assign n59816 = pi17 ? n32 : n59815;
  assign n59817 = pi16 ? n32 : n59816;
  assign n59818 = pi15 ? n59817 : n59239;
  assign n59819 = pi22 ? n335 : n47;
  assign n59820 = pi21 ? n4938 : n59819;
  assign n59821 = pi20 ? n20563 : n59820;
  assign n59822 = pi19 ? n20563 : n59821;
  assign n59823 = pi18 ? n20563 : n59822;
  assign n59824 = pi17 ? n45739 : n59823;
  assign n59825 = pi16 ? n32 : n59824;
  assign n59826 = pi22 ? n335 : n103;
  assign n59827 = pi21 ? n59247 : n59826;
  assign n59828 = pi20 ? n20563 : n59827;
  assign n59829 = pi19 ? n20563 : n59828;
  assign n59830 = pi18 ? n20563 : n59829;
  assign n59831 = pi17 ? n46884 : n59830;
  assign n59832 = pi16 ? n32 : n59831;
  assign n59833 = pi15 ? n59825 : n59832;
  assign n59834 = pi14 ? n59818 : n59833;
  assign n59835 = pi22 ? n52290 : n335;
  assign n59836 = pi21 ? n59835 : n59826;
  assign n59837 = pi20 ? n31220 : n59836;
  assign n59838 = pi19 ? n20563 : n59837;
  assign n59839 = pi18 ? n20563 : n59838;
  assign n59840 = pi17 ? n46884 : n59839;
  assign n59841 = pi16 ? n32 : n59840;
  assign n59842 = pi22 ? n55429 : n335;
  assign n59843 = pi22 ? n335 : n261;
  assign n59844 = pi21 ? n59842 : n59843;
  assign n59845 = pi20 ? n31220 : n59844;
  assign n59846 = pi19 ? n20563 : n59845;
  assign n59847 = pi18 ? n20563 : n59846;
  assign n59848 = pi17 ? n44643 : n59847;
  assign n59849 = pi16 ? n32 : n59848;
  assign n59850 = pi15 ? n59841 : n59849;
  assign n59851 = pi17 ? n44652 : n59847;
  assign n59852 = pi16 ? n32 : n59851;
  assign n59853 = pi17 ? n44222 : n59260;
  assign n59854 = pi16 ? n32 : n59853;
  assign n59855 = pi15 ? n59852 : n59854;
  assign n59856 = pi14 ? n59850 : n59855;
  assign n59857 = pi13 ? n59834 : n59856;
  assign n59858 = pi17 ? n43674 : n59278;
  assign n59859 = pi16 ? n32 : n59858;
  assign n59860 = pi17 ? n43674 : n59286;
  assign n59861 = pi16 ? n32 : n59860;
  assign n59862 = pi17 ? n44687 : n59286;
  assign n59863 = pi16 ? n32 : n59862;
  assign n59864 = pi15 ? n59861 : n59863;
  assign n59865 = pi14 ? n59859 : n59864;
  assign n59866 = pi17 ? n44247 : n59297;
  assign n59867 = pi16 ? n32 : n59866;
  assign n59868 = pi17 ? n43223 : n59297;
  assign n59869 = pi16 ? n32 : n59868;
  assign n59870 = pi15 ? n59867 : n59869;
  assign n59871 = pi17 ? n43223 : n59308;
  assign n59872 = pi16 ? n32 : n59871;
  assign n59873 = pi17 ? n43223 : n58894;
  assign n59874 = pi16 ? n32 : n59873;
  assign n59875 = pi15 ? n59872 : n59874;
  assign n59876 = pi14 ? n59870 : n59875;
  assign n59877 = pi13 ? n59865 : n59876;
  assign n59878 = pi12 ? n59857 : n59877;
  assign n59879 = pi21 ? n59324 : n37547;
  assign n59880 = pi20 ? n54354 : n59879;
  assign n59881 = pi19 ? n20563 : n59880;
  assign n59882 = pi18 ? n20563 : n59881;
  assign n59883 = pi17 ? n43223 : n59882;
  assign n59884 = pi16 ? n32 : n59883;
  assign n59885 = pi24 ? n157 : n51564;
  assign n59886 = pi23 ? n59885 : n316;
  assign n59887 = pi22 ? n59886 : n316;
  assign n59888 = pi21 ? n59887 : n2320;
  assign n59889 = pi20 ? n54354 : n59888;
  assign n59890 = pi19 ? n20563 : n59889;
  assign n59891 = pi18 ? n20563 : n59890;
  assign n59892 = pi17 ? n43227 : n59891;
  assign n59893 = pi16 ? n32 : n59892;
  assign n59894 = pi15 ? n59884 : n59893;
  assign n59895 = pi17 ? n43248 : n58925;
  assign n59896 = pi16 ? n32 : n59895;
  assign n59897 = pi17 ? n44274 : n59346;
  assign n59898 = pi16 ? n32 : n59897;
  assign n59899 = pi15 ? n59896 : n59898;
  assign n59900 = pi14 ? n59894 : n59899;
  assign n59901 = pi17 ? n44274 : n59354;
  assign n59902 = pi16 ? n32 : n59901;
  assign n59903 = pi17 ? n44274 : n59361;
  assign n59904 = pi16 ? n32 : n59903;
  assign n59905 = pi15 ? n59902 : n59904;
  assign n59906 = pi17 ? n48624 : n59370;
  assign n59907 = pi16 ? n32 : n59906;
  assign n59908 = pi17 ? n42645 : n59376;
  assign n59909 = pi16 ? n32 : n59908;
  assign n59910 = pi15 ? n59907 : n59909;
  assign n59911 = pi14 ? n59905 : n59910;
  assign n59912 = pi13 ? n59900 : n59911;
  assign n59913 = pi17 ? n42655 : n59385;
  assign n59914 = pi16 ? n32 : n59913;
  assign n59915 = pi17 ? n43255 : n59391;
  assign n59916 = pi16 ? n32 : n59915;
  assign n59917 = pi15 ? n59914 : n59916;
  assign n59918 = pi17 ? n43255 : n59400;
  assign n59919 = pi16 ? n32 : n59918;
  assign n59920 = pi17 ? n43255 : n56406;
  assign n59921 = pi16 ? n32 : n59920;
  assign n59922 = pi15 ? n59919 : n59921;
  assign n59923 = pi14 ? n59917 : n59922;
  assign n59924 = pi17 ? n43255 : n59409;
  assign n59925 = pi16 ? n32 : n59924;
  assign n59926 = pi17 ? n43262 : n59419;
  assign n59927 = pi16 ? n32 : n59926;
  assign n59928 = pi15 ? n59925 : n59927;
  assign n59929 = pi17 ? n43262 : n59428;
  assign n59930 = pi16 ? n32 : n59929;
  assign n59931 = pi17 ? n48121 : n59435;
  assign n59932 = pi16 ? n32 : n59931;
  assign n59933 = pi15 ? n59930 : n59932;
  assign n59934 = pi14 ? n59928 : n59933;
  assign n59935 = pi13 ? n59923 : n59934;
  assign n59936 = pi12 ? n59912 : n59935;
  assign n59937 = pi11 ? n59878 : n59936;
  assign n59938 = pi17 ? n48121 : n59445;
  assign n59939 = pi16 ? n32 : n59938;
  assign n59940 = pi17 ? n48121 : n59454;
  assign n59941 = pi16 ? n32 : n59940;
  assign n59942 = pi15 ? n59939 : n59941;
  assign n59943 = pi17 ? n48121 : n59462;
  assign n59944 = pi16 ? n32 : n59943;
  assign n59945 = pi17 ? n42207 : n59469;
  assign n59946 = pi16 ? n32 : n59945;
  assign n59947 = pi15 ? n59944 : n59946;
  assign n59948 = pi14 ? n59942 : n59947;
  assign n59949 = pi17 ? n42207 : n59477;
  assign n59950 = pi16 ? n32 : n59949;
  assign n59951 = pi20 ? n59480 : n53984;
  assign n59952 = pi19 ? n47159 : n59951;
  assign n59953 = pi18 ? n20563 : n59952;
  assign n59954 = pi17 ? n41642 : n59953;
  assign n59955 = pi16 ? n32 : n59954;
  assign n59956 = pi15 ? n59950 : n59955;
  assign n59957 = pi24 ? n36659 : n157;
  assign n59958 = pi23 ? n59957 : n157;
  assign n59959 = pi22 ? n59958 : n316;
  assign n59960 = pi21 ? n36659 : n59959;
  assign n59961 = pi20 ? n59960 : n1822;
  assign n59962 = pi19 ? n56631 : n59961;
  assign n59963 = pi18 ? n20563 : n59962;
  assign n59964 = pi17 ? n42688 : n59963;
  assign n59965 = pi16 ? n32 : n59964;
  assign n59966 = pi19 ? n51234 : n40791;
  assign n59967 = pi18 ? n32 : n59966;
  assign n59968 = pi17 ? n59967 : n59502;
  assign n59969 = pi16 ? n32 : n59968;
  assign n59970 = pi15 ? n59965 : n59969;
  assign n59971 = pi14 ? n59956 : n59970;
  assign n59972 = pi13 ? n59948 : n59971;
  assign n59973 = pi22 ? n49720 : n20563;
  assign n59974 = pi21 ? n32 : n59973;
  assign n59975 = pi20 ? n32 : n59974;
  assign n59976 = pi19 ? n59975 : n59510;
  assign n59977 = pi18 ? n32 : n59976;
  assign n59978 = pi23 ? n15293 : n204;
  assign n59979 = pi22 ? n59978 : n58452;
  assign n59980 = pi21 ? n36781 : n59979;
  assign n59981 = pi20 ? n59980 : n32;
  assign n59982 = pi19 ? n59513 : n59981;
  assign n59983 = pi18 ? n20563 : n59982;
  assign n59984 = pi17 ? n59977 : n59983;
  assign n59985 = pi16 ? n32 : n59984;
  assign n59986 = pi19 ? n59975 : n20563;
  assign n59987 = pi18 ? n32 : n59986;
  assign n59988 = pi17 ? n59987 : n59530;
  assign n59989 = pi16 ? n32 : n59988;
  assign n59990 = pi15 ? n59985 : n59989;
  assign n59991 = pi22 ? n51754 : n20563;
  assign n59992 = pi21 ? n32 : n59991;
  assign n59993 = pi20 ? n32 : n59992;
  assign n59994 = pi19 ? n59993 : n20563;
  assign n59995 = pi18 ? n32 : n59994;
  assign n59996 = pi17 ? n59995 : n59543;
  assign n59997 = pi16 ? n32 : n59996;
  assign n59998 = pi20 ? n20563 : n51188;
  assign n59999 = pi19 ? n59551 : n59998;
  assign n60000 = pi18 ? n59999 : n59558;
  assign n60001 = pi17 ? n46998 : n60000;
  assign n60002 = pi16 ? n32 : n60001;
  assign n60003 = pi15 ? n59997 : n60002;
  assign n60004 = pi14 ? n59990 : n60003;
  assign n60005 = pi17 ? n46998 : n59567;
  assign n60006 = pi16 ? n32 : n60005;
  assign n60007 = pi17 ? n46998 : n59573;
  assign n60008 = pi16 ? n32 : n60007;
  assign n60009 = pi15 ? n60006 : n60008;
  assign n60010 = pi17 ? n46998 : n59580;
  assign n60011 = pi16 ? n32 : n60010;
  assign n60012 = pi17 ? n40486 : n59586;
  assign n60013 = pi16 ? n32 : n60012;
  assign n60014 = pi15 ? n60011 : n60013;
  assign n60015 = pi14 ? n60009 : n60014;
  assign n60016 = pi13 ? n60004 : n60015;
  assign n60017 = pi12 ? n59972 : n60016;
  assign n60018 = pi17 ? n46998 : n59599;
  assign n60019 = pi16 ? n32 : n60018;
  assign n60020 = pi17 ? n46998 : n59607;
  assign n60021 = pi16 ? n32 : n60020;
  assign n60022 = pi15 ? n60019 : n60021;
  assign n60023 = pi21 ? n32 : n39801;
  assign n60024 = pi20 ? n32 : n60023;
  assign n60025 = pi19 ? n60024 : n40791;
  assign n60026 = pi18 ? n32 : n60025;
  assign n60027 = pi21 ? n36489 : n39191;
  assign n60028 = pi20 ? n36489 : n60027;
  assign n60029 = pi21 ? n30868 : n39191;
  assign n60030 = pi20 ? n40915 : n60029;
  assign n60031 = pi19 ? n60028 : n60030;
  assign n60032 = pi22 ? n33792 : n3944;
  assign n60033 = pi21 ? n36489 : n60032;
  assign n60034 = pi20 ? n40915 : n60033;
  assign n60035 = pi19 ? n60034 : n59623;
  assign n60036 = pi18 ? n60031 : n60035;
  assign n60037 = pi17 ? n60026 : n60036;
  assign n60038 = pi16 ? n32 : n60037;
  assign n60039 = pi19 ? n48790 : n30868;
  assign n60040 = pi18 ? n32 : n60039;
  assign n60041 = pi17 ? n60040 : n59638;
  assign n60042 = pi16 ? n32 : n60041;
  assign n60043 = pi15 ? n60038 : n60042;
  assign n60044 = pi14 ? n60022 : n60043;
  assign n60045 = pi21 ? n55560 : n32;
  assign n60046 = pi20 ? n60045 : n32;
  assign n60047 = pi19 ? n59647 : n60046;
  assign n60048 = pi18 ? n30868 : n60047;
  assign n60049 = pi17 ? n48799 : n60048;
  assign n60050 = pi16 ? n32 : n60049;
  assign n60051 = pi17 ? n48799 : n59661;
  assign n60052 = pi16 ? n32 : n60051;
  assign n60053 = pi15 ? n60050 : n60052;
  assign n60054 = pi22 ? n30115 : n30868;
  assign n60055 = pi21 ? n32 : n60054;
  assign n60056 = pi20 ? n32 : n60055;
  assign n60057 = pi19 ? n60056 : n59667;
  assign n60058 = pi18 ? n32 : n60057;
  assign n60059 = pi17 ? n60058 : n59677;
  assign n60060 = pi16 ? n32 : n60059;
  assign n60061 = pi17 ? n48806 : n59685;
  assign n60062 = pi16 ? n32 : n60061;
  assign n60063 = pi15 ? n60060 : n60062;
  assign n60064 = pi14 ? n60053 : n60063;
  assign n60065 = pi13 ? n60044 : n60064;
  assign n60066 = pi17 ? n48806 : n59695;
  assign n60067 = pi16 ? n32 : n60066;
  assign n60068 = pi19 ? n48858 : n59700;
  assign n60069 = pi18 ? n32 : n60068;
  assign n60070 = pi17 ? n60069 : n59711;
  assign n60071 = pi16 ? n32 : n60070;
  assign n60072 = pi15 ? n60067 : n60071;
  assign n60073 = pi19 ? n46078 : n33792;
  assign n60074 = pi18 ? n32 : n60073;
  assign n60075 = pi24 ? n43198 : n14626;
  assign n60076 = pi23 ? n204 : n60075;
  assign n60077 = pi22 ? n60076 : n13481;
  assign n60078 = pi21 ? n43198 : n60077;
  assign n60079 = pi20 ? n33792 : n60078;
  assign n60080 = pi19 ? n60079 : n32;
  assign n60081 = pi18 ? n33792 : n60080;
  assign n60082 = pi17 ? n60074 : n60081;
  assign n60083 = pi16 ? n32 : n60082;
  assign n60084 = pi19 ? n46202 : n59729;
  assign n60085 = pi18 ? n32 : n60084;
  assign n60086 = pi17 ? n60085 : n59737;
  assign n60087 = pi16 ? n32 : n60086;
  assign n60088 = pi15 ? n60083 : n60087;
  assign n60089 = pi14 ? n60072 : n60088;
  assign n60090 = pi19 ? n46226 : n59742;
  assign n60091 = pi18 ? n32 : n60090;
  assign n60092 = pi23 ? n36781 : n13481;
  assign n60093 = pi22 ? n43198 : n60092;
  assign n60094 = pi21 ? n60093 : n58966;
  assign n60095 = pi20 ? n43198 : n60094;
  assign n60096 = pi19 ? n60095 : n32;
  assign n60097 = pi18 ? n43198 : n60096;
  assign n60098 = pi17 ? n60091 : n60097;
  assign n60099 = pi16 ? n32 : n60098;
  assign n60100 = pi18 ? n32 : n54588;
  assign n60101 = pi17 ? n60100 : n59759;
  assign n60102 = pi16 ? n32 : n60101;
  assign n60103 = pi15 ? n60099 : n60102;
  assign n60104 = pi21 ? n57185 : n39972;
  assign n60105 = pi20 ? n59764 : n60104;
  assign n60106 = pi19 ? n46226 : n60105;
  assign n60107 = pi18 ? n32 : n60106;
  assign n60108 = pi17 ? n60107 : n59778;
  assign n60109 = pi16 ? n32 : n60108;
  assign n60110 = pi19 ? n46278 : n59781;
  assign n60111 = pi18 ? n32 : n60110;
  assign n60112 = pi21 ? n59691 : n928;
  assign n60113 = pi20 ? n55701 : n60112;
  assign n60114 = pi19 ? n60113 : n32;
  assign n60115 = pi18 ? n54659 : n60114;
  assign n60116 = pi17 ? n60111 : n60115;
  assign n60117 = pi16 ? n32 : n60116;
  assign n60118 = pi15 ? n60109 : n60117;
  assign n60119 = pi14 ? n60103 : n60118;
  assign n60120 = pi13 ? n60089 : n60119;
  assign n60121 = pi12 ? n60065 : n60120;
  assign n60122 = pi11 ? n60017 : n60121;
  assign n60123 = pi10 ? n59937 : n60122;
  assign n60124 = pi09 ? n59814 : n60123;
  assign n60125 = pi08 ? n59798 : n60124;
  assign n60126 = pi22 ? n139 : n119;
  assign n60127 = pi21 ? n297 : n60126;
  assign n60128 = pi20 ? n31220 : n60127;
  assign n60129 = pi19 ? n38478 : n60128;
  assign n60130 = pi18 ? n38957 : n60129;
  assign n60131 = pi17 ? n32 : n60130;
  assign n60132 = pi16 ? n32 : n60131;
  assign n60133 = pi15 ? n32 : n60132;
  assign n60134 = pi22 ? n139 : n1617;
  assign n60135 = pi21 ? n297 : n60134;
  assign n60136 = pi20 ? n31220 : n60135;
  assign n60137 = pi19 ? n20563 : n60136;
  assign n60138 = pi18 ? n38957 : n60137;
  assign n60139 = pi17 ? n32 : n60138;
  assign n60140 = pi16 ? n32 : n60139;
  assign n60141 = pi20 ? n33821 : n60135;
  assign n60142 = pi19 ? n38478 : n60141;
  assign n60143 = pi18 ? n40045 : n60142;
  assign n60144 = pi17 ? n32 : n60143;
  assign n60145 = pi16 ? n32 : n60144;
  assign n60146 = pi15 ? n60140 : n60145;
  assign n60147 = pi14 ? n60133 : n60146;
  assign n60148 = pi13 ? n32 : n60147;
  assign n60149 = pi12 ? n32 : n60148;
  assign n60150 = pi11 ? n32 : n60149;
  assign n60151 = pi10 ? n32 : n60150;
  assign n60152 = pi22 ? n335 : n1617;
  assign n60153 = pi21 ? n569 : n60152;
  assign n60154 = pi20 ? n31220 : n60153;
  assign n60155 = pi19 ? n20563 : n60154;
  assign n60156 = pi18 ? n40045 : n60155;
  assign n60157 = pi17 ? n32 : n60156;
  assign n60158 = pi16 ? n32 : n60157;
  assign n60159 = pi18 ? n38316 : n60155;
  assign n60160 = pi17 ? n32 : n60159;
  assign n60161 = pi16 ? n32 : n60160;
  assign n60162 = pi15 ? n60158 : n60161;
  assign n60163 = pi20 ? n20563 : n60153;
  assign n60164 = pi19 ? n20563 : n60163;
  assign n60165 = pi18 ? n20563 : n60164;
  assign n60166 = pi17 ? n32 : n60165;
  assign n60167 = pi16 ? n32 : n60166;
  assign n60168 = pi19 ? n53012 : n60163;
  assign n60169 = pi18 ? n20563 : n60168;
  assign n60170 = pi17 ? n32 : n60169;
  assign n60171 = pi16 ? n32 : n60170;
  assign n60172 = pi15 ? n60167 : n60171;
  assign n60173 = pi14 ? n60162 : n60172;
  assign n60174 = pi18 ? n20563 : n60155;
  assign n60175 = pi17 ? n45232 : n60174;
  assign n60176 = pi16 ? n32 : n60175;
  assign n60177 = pi17 ? n44634 : n60174;
  assign n60178 = pi16 ? n32 : n60177;
  assign n60179 = pi17 ? n45739 : n60174;
  assign n60180 = pi16 ? n32 : n60179;
  assign n60181 = pi15 ? n60178 : n60180;
  assign n60182 = pi14 ? n60176 : n60181;
  assign n60183 = pi13 ? n60173 : n60182;
  assign n60184 = pi22 ? n363 : n1617;
  assign n60185 = pi21 ? n3392 : n60184;
  assign n60186 = pi20 ? n20563 : n60185;
  assign n60187 = pi19 ? n20563 : n60186;
  assign n60188 = pi18 ? n20563 : n60187;
  assign n60189 = pi17 ? n44222 : n60188;
  assign n60190 = pi16 ? n32 : n60189;
  assign n60191 = pi22 ? n157 : n1617;
  assign n60192 = pi21 ? n244 : n60191;
  assign n60193 = pi20 ? n31220 : n60192;
  assign n60194 = pi19 ? n20563 : n60193;
  assign n60195 = pi18 ? n20563 : n60194;
  assign n60196 = pi17 ? n45242 : n60195;
  assign n60197 = pi16 ? n32 : n60196;
  assign n60198 = pi17 ? n46348 : n60195;
  assign n60199 = pi16 ? n32 : n60198;
  assign n60200 = pi15 ? n60197 : n60199;
  assign n60201 = pi14 ? n60190 : n60200;
  assign n60202 = pi17 ? n44670 : n59297;
  assign n60203 = pi16 ? n32 : n60202;
  assign n60204 = pi17 ? n43674 : n59297;
  assign n60205 = pi16 ? n32 : n60204;
  assign n60206 = pi15 ? n60203 : n60205;
  assign n60207 = pi17 ? n43674 : n59308;
  assign n60208 = pi16 ? n32 : n60207;
  assign n60209 = pi24 ? n37 : n14626;
  assign n60210 = pi23 ? n60209 : n14626;
  assign n60211 = pi22 ? n60210 : n685;
  assign n60212 = pi21 ? n60211 : n696;
  assign n60213 = pi20 ? n20563 : n60212;
  assign n60214 = pi19 ? n20563 : n60213;
  assign n60215 = pi18 ? n20563 : n60214;
  assign n60216 = pi17 ? n43674 : n60215;
  assign n60217 = pi16 ? n32 : n60216;
  assign n60218 = pi15 ? n60208 : n60217;
  assign n60219 = pi14 ? n60206 : n60218;
  assign n60220 = pi13 ? n60201 : n60219;
  assign n60221 = pi12 ? n60183 : n60220;
  assign n60222 = pi17 ? n43674 : n59882;
  assign n60223 = pi16 ? n32 : n60222;
  assign n60224 = pi17 ? n44687 : n59333;
  assign n60225 = pi16 ? n32 : n60224;
  assign n60226 = pi15 ? n60223 : n60225;
  assign n60227 = pi17 ? n44247 : n58925;
  assign n60228 = pi16 ? n32 : n60227;
  assign n60229 = pi17 ? n44247 : n59346;
  assign n60230 = pi16 ? n32 : n60229;
  assign n60231 = pi15 ? n60228 : n60230;
  assign n60232 = pi14 ? n60226 : n60231;
  assign n60233 = pi20 ? n59340 : n59351;
  assign n60234 = pi19 ? n20563 : n60233;
  assign n60235 = pi18 ? n20563 : n60234;
  assign n60236 = pi17 ? n44247 : n60235;
  assign n60237 = pi16 ? n32 : n60236;
  assign n60238 = pi21 ? n14626 : n928;
  assign n60239 = pi20 ? n56361 : n60238;
  assign n60240 = pi19 ? n20563 : n60239;
  assign n60241 = pi18 ? n20563 : n60240;
  assign n60242 = pi17 ? n44247 : n60241;
  assign n60243 = pi16 ? n32 : n60242;
  assign n60244 = pi15 ? n60237 : n60243;
  assign n60245 = pi20 ? n56374 : n59367;
  assign n60246 = pi19 ? n20563 : n60245;
  assign n60247 = pi18 ? n20563 : n60246;
  assign n60248 = pi17 ? n44247 : n60247;
  assign n60249 = pi16 ? n32 : n60248;
  assign n60250 = pi21 ? n51564 : n2700;
  assign n60251 = pi20 ? n56374 : n60250;
  assign n60252 = pi19 ? n20563 : n60251;
  assign n60253 = pi18 ? n20563 : n60252;
  assign n60254 = pi17 ? n43223 : n60253;
  assign n60255 = pi16 ? n32 : n60254;
  assign n60256 = pi15 ? n60249 : n60255;
  assign n60257 = pi14 ? n60244 : n60256;
  assign n60258 = pi13 ? n60232 : n60257;
  assign n60259 = pi20 ? n55343 : n59388;
  assign n60260 = pi19 ? n20563 : n60259;
  assign n60261 = pi18 ? n20563 : n60260;
  assign n60262 = pi17 ? n43227 : n60261;
  assign n60263 = pi16 ? n32 : n60262;
  assign n60264 = pi23 ? n30868 : n157;
  assign n60265 = pi22 ? n37 : n60264;
  assign n60266 = pi21 ? n20563 : n60265;
  assign n60267 = pi20 ? n60266 : n59388;
  assign n60268 = pi19 ? n20563 : n60267;
  assign n60269 = pi18 ? n20563 : n60268;
  assign n60270 = pi17 ? n43248 : n60269;
  assign n60271 = pi16 ? n32 : n60270;
  assign n60272 = pi15 ? n60263 : n60271;
  assign n60273 = pi17 ? n43248 : n59400;
  assign n60274 = pi16 ? n32 : n60273;
  assign n60275 = pi23 ? n33792 : n204;
  assign n60276 = pi22 ? n37 : n60275;
  assign n60277 = pi21 ? n20563 : n60276;
  assign n60278 = pi20 ? n60277 : n15407;
  assign n60279 = pi19 ? n20563 : n60278;
  assign n60280 = pi18 ? n20563 : n60279;
  assign n60281 = pi17 ? n43248 : n60280;
  assign n60282 = pi16 ? n32 : n60281;
  assign n60283 = pi15 ? n60274 : n60282;
  assign n60284 = pi14 ? n60272 : n60283;
  assign n60285 = pi21 ? n20563 : n2084;
  assign n60286 = pi20 ? n60285 : n8917;
  assign n60287 = pi19 ? n20563 : n60286;
  assign n60288 = pi18 ? n20563 : n60287;
  assign n60289 = pi17 ? n44274 : n60288;
  assign n60290 = pi16 ? n32 : n60289;
  assign n60291 = pi23 ? n363 : n14626;
  assign n60292 = pi22 ? n20563 : n60291;
  assign n60293 = pi21 ? n20563 : n60292;
  assign n60294 = pi20 ? n60293 : n59416;
  assign n60295 = pi19 ? n20563 : n60294;
  assign n60296 = pi18 ? n20563 : n60295;
  assign n60297 = pi17 ? n48624 : n60296;
  assign n60298 = pi16 ? n32 : n60297;
  assign n60299 = pi15 ? n60290 : n60298;
  assign n60300 = pi23 ? n157 : n51564;
  assign n60301 = pi22 ? n99 : n60300;
  assign n60302 = pi21 ? n20563 : n60301;
  assign n60303 = pi20 ? n60302 : n57434;
  assign n60304 = pi19 ? n20563 : n60303;
  assign n60305 = pi18 ? n20563 : n60304;
  assign n60306 = pi17 ? n48624 : n60305;
  assign n60307 = pi16 ? n32 : n60306;
  assign n60308 = pi22 ? n30868 : n1484;
  assign n60309 = pi21 ? n20563 : n60308;
  assign n60310 = pi20 ? n60309 : n4008;
  assign n60311 = pi19 ? n20563 : n60310;
  assign n60312 = pi18 ? n20563 : n60311;
  assign n60313 = pi17 ? n42681 : n60312;
  assign n60314 = pi16 ? n32 : n60313;
  assign n60315 = pi15 ? n60307 : n60314;
  assign n60316 = pi14 ? n60299 : n60315;
  assign n60317 = pi13 ? n60284 : n60316;
  assign n60318 = pi12 ? n60258 : n60317;
  assign n60319 = pi11 ? n60221 : n60318;
  assign n60320 = pi17 ? n42681 : n59445;
  assign n60321 = pi16 ? n32 : n60320;
  assign n60322 = pi20 ? n59448 : n57459;
  assign n60323 = pi19 ? n40792 : n60322;
  assign n60324 = pi18 ? n20563 : n60323;
  assign n60325 = pi17 ? n42681 : n60324;
  assign n60326 = pi16 ? n32 : n60325;
  assign n60327 = pi15 ? n60321 : n60326;
  assign n60328 = pi21 ? n52632 : n14626;
  assign n60329 = pi20 ? n60328 : n5830;
  assign n60330 = pi19 ? n59458 : n60329;
  assign n60331 = pi18 ? n20563 : n60330;
  assign n60332 = pi17 ? n42681 : n60331;
  assign n60333 = pi16 ? n32 : n60332;
  assign n60334 = pi22 ? n37 : n39190;
  assign n60335 = pi21 ? n60334 : n14626;
  assign n60336 = pi20 ? n60335 : n2653;
  assign n60337 = pi19 ? n20563 : n60336;
  assign n60338 = pi18 ? n20563 : n60337;
  assign n60339 = pi17 ? n43255 : n60338;
  assign n60340 = pi16 ? n32 : n60339;
  assign n60341 = pi15 ? n60333 : n60340;
  assign n60342 = pi14 ? n60327 : n60341;
  assign n60343 = pi21 ? n47664 : n685;
  assign n60344 = pi20 ? n60343 : n37640;
  assign n60345 = pi19 ? n20563 : n60344;
  assign n60346 = pi18 ? n20563 : n60345;
  assign n60347 = pi17 ? n43255 : n60346;
  assign n60348 = pi16 ? n32 : n60347;
  assign n60349 = pi20 ? n59480 : n1822;
  assign n60350 = pi19 ? n47159 : n60349;
  assign n60351 = pi18 ? n20563 : n60350;
  assign n60352 = pi17 ? n42201 : n60351;
  assign n60353 = pi16 ? n32 : n60352;
  assign n60354 = pi15 ? n60348 : n60353;
  assign n60355 = pi23 ? n59957 : n36798;
  assign n60356 = pi22 ? n60355 : n316;
  assign n60357 = pi21 ? n36659 : n60356;
  assign n60358 = pi20 ? n60357 : n1822;
  assign n60359 = pi19 ? n56631 : n60358;
  assign n60360 = pi18 ? n20563 : n60359;
  assign n60361 = pi17 ? n42201 : n60360;
  assign n60362 = pi16 ? n32 : n60361;
  assign n60363 = pi20 ? n59020 : n40791;
  assign n60364 = pi19 ? n32 : n60363;
  assign n60365 = pi18 ? n32 : n60364;
  assign n60366 = pi20 ? n43010 : n59593;
  assign n60367 = pi22 ? n59497 : n1407;
  assign n60368 = pi21 ? n36659 : n60367;
  assign n60369 = pi20 ? n60368 : n32;
  assign n60370 = pi19 ? n60366 : n60369;
  assign n60371 = pi18 ? n20563 : n60370;
  assign n60372 = pi17 ? n60365 : n60371;
  assign n60373 = pi16 ? n32 : n60372;
  assign n60374 = pi15 ? n60362 : n60373;
  assign n60375 = pi14 ? n60354 : n60374;
  assign n60376 = pi13 ? n60342 : n60375;
  assign n60377 = pi21 ? n30866 : n33792;
  assign n60378 = pi20 ? n60377 : n53326;
  assign n60379 = pi19 ? n32 : n60378;
  assign n60380 = pi18 ? n32 : n60379;
  assign n60381 = pi20 ? n33792 : n59602;
  assign n60382 = pi23 ? n15293 : n43198;
  assign n60383 = pi22 ? n60382 : n317;
  assign n60384 = pi21 ? n36781 : n60383;
  assign n60385 = pi20 ? n60384 : n32;
  assign n60386 = pi19 ? n60381 : n60385;
  assign n60387 = pi18 ? n20563 : n60386;
  assign n60388 = pi17 ? n60380 : n60387;
  assign n60389 = pi16 ? n32 : n60388;
  assign n60390 = pi22 ? n36617 : n55535;
  assign n60391 = pi21 ? n20563 : n60390;
  assign n60392 = pi20 ? n55014 : n60391;
  assign n60393 = pi19 ? n32 : n60392;
  assign n60394 = pi18 ? n32 : n60393;
  assign n60395 = pi20 ? n20563 : n54468;
  assign n60396 = pi23 ? n36659 : n157;
  assign n60397 = pi22 ? n30868 : n60396;
  assign n60398 = pi23 ? n35938 : n14626;
  assign n60399 = pi22 ? n60398 : n317;
  assign n60400 = pi21 ? n60397 : n60399;
  assign n60401 = pi20 ? n60400 : n32;
  assign n60402 = pi19 ? n60395 : n60401;
  assign n60403 = pi18 ? n20563 : n60402;
  assign n60404 = pi17 ? n60394 : n60403;
  assign n60405 = pi16 ? n32 : n60404;
  assign n60406 = pi15 ? n60389 : n60405;
  assign n60407 = pi21 ? n20563 : n45092;
  assign n60408 = pi24 ? n36659 : n20563;
  assign n60409 = pi23 ? n36659 : n60408;
  assign n60410 = pi22 ? n59056 : n60409;
  assign n60411 = pi21 ? n20563 : n60410;
  assign n60412 = pi20 ? n60407 : n60411;
  assign n60413 = pi19 ? n32 : n60412;
  assign n60414 = pi18 ? n32 : n60413;
  assign n60415 = pi21 ? n40986 : n20563;
  assign n60416 = pi20 ? n60415 : n38754;
  assign n60417 = pi19 ? n60416 : n59541;
  assign n60418 = pi18 ? n20563 : n60417;
  assign n60419 = pi17 ? n60414 : n60418;
  assign n60420 = pi16 ? n32 : n60419;
  assign n60421 = pi22 ? n51564 : n32;
  assign n60422 = pi21 ? n59555 : n60421;
  assign n60423 = pi20 ? n60422 : n32;
  assign n60424 = pi19 ? n39193 : n60423;
  assign n60425 = pi18 ? n20563 : n60424;
  assign n60426 = pi17 ? n41631 : n60425;
  assign n60427 = pi16 ? n32 : n60426;
  assign n60428 = pi15 ? n60420 : n60427;
  assign n60429 = pi14 ? n60406 : n60428;
  assign n60430 = pi19 ? n56605 : n59565;
  assign n60431 = pi18 ? n20563 : n60430;
  assign n60432 = pi17 ? n41631 : n60431;
  assign n60433 = pi16 ? n32 : n60432;
  assign n60434 = pi21 ? n14626 : n59785;
  assign n60435 = pi20 ? n60434 : n32;
  assign n60436 = pi19 ? n56605 : n60435;
  assign n60437 = pi18 ? n20563 : n60436;
  assign n60438 = pi17 ? n42207 : n60437;
  assign n60439 = pi16 ? n32 : n60438;
  assign n60440 = pi15 ? n60433 : n60439;
  assign n60441 = pi22 ? n20563 : n58710;
  assign n60442 = pi21 ? n20563 : n60441;
  assign n60443 = pi20 ? n20563 : n60442;
  assign n60444 = pi19 ? n60443 : n59578;
  assign n60445 = pi18 ? n20563 : n60444;
  assign n60446 = pi17 ? n42207 : n60445;
  assign n60447 = pi16 ? n32 : n60446;
  assign n60448 = pi23 ? n37 : n56976;
  assign n60449 = pi22 ? n60448 : n36659;
  assign n60450 = pi21 ? n20563 : n60449;
  assign n60451 = pi20 ? n20563 : n60450;
  assign n60452 = pi19 ? n60451 : n59584;
  assign n60453 = pi18 ? n20563 : n60452;
  assign n60454 = pi17 ? n47593 : n60453;
  assign n60455 = pi16 ? n32 : n60454;
  assign n60456 = pi15 ? n60447 : n60455;
  assign n60457 = pi14 ? n60440 : n60456;
  assign n60458 = pi13 ? n60429 : n60457;
  assign n60459 = pi12 ? n60376 : n60458;
  assign n60460 = pi22 ? n30868 : n38284;
  assign n60461 = pi21 ? n20563 : n60460;
  assign n60462 = pi20 ? n20563 : n60461;
  assign n60463 = pi22 ? n14626 : n56678;
  assign n60464 = pi21 ? n60463 : n1009;
  assign n60465 = pi20 ? n60464 : n32;
  assign n60466 = pi19 ? n60462 : n60465;
  assign n60467 = pi18 ? n20563 : n60466;
  assign n60468 = pi17 ? n48121 : n60467;
  assign n60469 = pi16 ? n32 : n60468;
  assign n60470 = pi22 ? n33792 : n37276;
  assign n60471 = pi21 ? n20563 : n60470;
  assign n60472 = pi20 ? n20563 : n60471;
  assign n60473 = pi19 ? n60472 : n59605;
  assign n60474 = pi18 ? n20563 : n60473;
  assign n60475 = pi17 ? n48121 : n60474;
  assign n60476 = pi16 ? n32 : n60475;
  assign n60477 = pi15 ? n60469 : n60476;
  assign n60478 = pi20 ? n48184 : n42005;
  assign n60479 = pi19 ? n37927 : n60478;
  assign n60480 = pi18 ? n32 : n60479;
  assign n60481 = pi20 ? n39805 : n36489;
  assign n60482 = pi19 ? n60481 : n40915;
  assign n60483 = pi22 ? n33792 : n46796;
  assign n60484 = pi21 ? n36489 : n60483;
  assign n60485 = pi20 ? n40915 : n60484;
  assign n60486 = pi19 ? n60485 : n55658;
  assign n60487 = pi18 ? n60482 : n60486;
  assign n60488 = pi17 ? n60480 : n60487;
  assign n60489 = pi16 ? n32 : n60488;
  assign n60490 = pi20 ? n48184 : n30868;
  assign n60491 = pi19 ? n37927 : n60490;
  assign n60492 = pi18 ? n32 : n60491;
  assign n60493 = pi22 ? n36659 : n52451;
  assign n60494 = pi21 ? n30868 : n60493;
  assign n60495 = pi20 ? n30868 : n60494;
  assign n60496 = pi19 ? n60495 : n59650;
  assign n60497 = pi18 ? n30868 : n60496;
  assign n60498 = pi17 ? n60492 : n60497;
  assign n60499 = pi16 ? n32 : n60498;
  assign n60500 = pi15 ? n60489 : n60499;
  assign n60501 = pi14 ? n60477 : n60500;
  assign n60502 = pi21 ? n48173 : n30868;
  assign n60503 = pi20 ? n60502 : n30868;
  assign n60504 = pi19 ? n49331 : n60503;
  assign n60505 = pi18 ? n32 : n60504;
  assign n60506 = pi17 ? n60505 : n60048;
  assign n60507 = pi16 ? n32 : n60506;
  assign n60508 = pi19 ? n59656 : n59675;
  assign n60509 = pi18 ? n30868 : n60508;
  assign n60510 = pi17 ? n60505 : n60509;
  assign n60511 = pi16 ? n32 : n60510;
  assign n60512 = pi15 ? n60507 : n60511;
  assign n60513 = pi21 ? n45049 : n30868;
  assign n60514 = pi20 ? n60513 : n30868;
  assign n60515 = pi19 ? n32 : n60514;
  assign n60516 = pi18 ? n32 : n60515;
  assign n60517 = pi17 ? n60516 : n59677;
  assign n60518 = pi16 ? n32 : n60517;
  assign n60519 = pi21 ? n43198 : n59681;
  assign n60520 = pi20 ? n30868 : n60519;
  assign n60521 = pi19 ? n60520 : n55691;
  assign n60522 = pi18 ? n30868 : n60521;
  assign n60523 = pi17 ? n49323 : n60522;
  assign n60524 = pi16 ? n32 : n60523;
  assign n60525 = pi15 ? n60518 : n60524;
  assign n60526 = pi14 ? n60512 : n60525;
  assign n60527 = pi13 ? n60501 : n60526;
  assign n60528 = pi18 ? n32 : n55004;
  assign n60529 = pi19 ? n59693 : n1823;
  assign n60530 = pi18 ? n30868 : n60529;
  assign n60531 = pi17 ? n60528 : n60530;
  assign n60532 = pi16 ? n32 : n60531;
  assign n60533 = pi22 ? n45652 : n37276;
  assign n60534 = pi21 ? n60533 : n52879;
  assign n60535 = pi21 ? n53480 : n43198;
  assign n60536 = pi20 ? n60534 : n60535;
  assign n60537 = pi19 ? n32 : n60536;
  assign n60538 = pi18 ? n32 : n60537;
  assign n60539 = pi22 ? n55799 : n33792;
  assign n60540 = pi21 ? n60539 : n43198;
  assign n60541 = pi23 ? n36659 : n139;
  assign n60542 = pi22 ? n60541 : n36798;
  assign n60543 = pi22 ? n58710 : n43198;
  assign n60544 = pi21 ? n60542 : n60543;
  assign n60545 = pi20 ? n60540 : n60544;
  assign n60546 = pi22 ? n54574 : n33792;
  assign n60547 = pi21 ? n53463 : n60546;
  assign n60548 = pi21 ? n36659 : n53484;
  assign n60549 = pi20 ? n60547 : n60548;
  assign n60550 = pi19 ? n60545 : n60549;
  assign n60551 = pi22 ? n54574 : n58736;
  assign n60552 = pi21 ? n43198 : n60551;
  assign n60553 = pi20 ? n60552 : n59692;
  assign n60554 = pi19 ? n60553 : n32;
  assign n60555 = pi18 ? n60550 : n60554;
  assign n60556 = pi17 ? n60538 : n60555;
  assign n60557 = pi16 ? n32 : n60556;
  assign n60558 = pi15 ? n60532 : n60557;
  assign n60559 = pi21 ? n52742 : n33792;
  assign n60560 = pi20 ? n60559 : n33792;
  assign n60561 = pi19 ? n32 : n60560;
  assign n60562 = pi18 ? n32 : n60561;
  assign n60563 = pi20 ? n33792 : n59734;
  assign n60564 = pi19 ? n60563 : n32;
  assign n60565 = pi18 ? n33792 : n60564;
  assign n60566 = pi17 ? n60562 : n60565;
  assign n60567 = pi16 ? n32 : n60566;
  assign n60568 = pi21 ? n57755 : n43198;
  assign n60569 = pi20 ? n60568 : n43198;
  assign n60570 = pi19 ? n32 : n60569;
  assign n60571 = pi18 ? n32 : n60570;
  assign n60572 = pi17 ? n60571 : n59737;
  assign n60573 = pi16 ? n32 : n60572;
  assign n60574 = pi15 ? n60567 : n60573;
  assign n60575 = pi14 ? n60558 : n60574;
  assign n60576 = pi22 ? n57197 : n53982;
  assign n60577 = pi21 ? n58777 : n60576;
  assign n60578 = pi20 ? n43198 : n60577;
  assign n60579 = pi19 ? n60578 : n32;
  assign n60580 = pi18 ? n43198 : n60579;
  assign n60581 = pi17 ? n60571 : n60580;
  assign n60582 = pi16 ? n32 : n60581;
  assign n60583 = pi21 ? n48856 : n46283;
  assign n60584 = pi20 ? n60583 : n43198;
  assign n60585 = pi19 ? n32 : n60584;
  assign n60586 = pi18 ? n32 : n60585;
  assign n60587 = pi17 ? n60586 : n59759;
  assign n60588 = pi16 ? n32 : n60587;
  assign n60589 = pi15 ? n60582 : n60588;
  assign n60590 = pi21 ? n58708 : n53551;
  assign n60591 = pi22 ? n36798 : n55799;
  assign n60592 = pi21 ? n60591 : n55800;
  assign n60593 = pi20 ? n60590 : n60592;
  assign n60594 = pi19 ? n32 : n60593;
  assign n60595 = pi18 ? n32 : n60594;
  assign n60596 = pi21 ? n53551 : n56212;
  assign n60597 = pi21 ? n60591 : n53551;
  assign n60598 = pi20 ? n60596 : n60597;
  assign n60599 = pi21 ? n56212 : n36798;
  assign n60600 = pi20 ? n36798 : n60599;
  assign n60601 = pi19 ? n60598 : n60600;
  assign n60602 = pi22 ? n51907 : n36798;
  assign n60603 = pi21 ? n60602 : n60591;
  assign n60604 = pi21 ? n59691 : n55560;
  assign n60605 = pi20 ? n60603 : n60604;
  assign n60606 = pi19 ? n60605 : n32;
  assign n60607 = pi18 ? n60601 : n60606;
  assign n60608 = pi17 ? n60595 : n60607;
  assign n60609 = pi16 ? n32 : n60608;
  assign n60610 = pi21 ? n46772 : n47397;
  assign n60611 = pi20 ? n60610 : n49401;
  assign n60612 = pi19 ? n32 : n60611;
  assign n60613 = pi18 ? n32 : n60612;
  assign n60614 = pi21 ? n59691 : n37639;
  assign n60615 = pi20 ? n55701 : n60614;
  assign n60616 = pi19 ? n60615 : n32;
  assign n60617 = pi18 ? n54659 : n60616;
  assign n60618 = pi17 ? n60613 : n60617;
  assign n60619 = pi16 ? n32 : n60618;
  assign n60620 = pi15 ? n60609 : n60619;
  assign n60621 = pi14 ? n60589 : n60620;
  assign n60622 = pi13 ? n60575 : n60621;
  assign n60623 = pi12 ? n60527 : n60622;
  assign n60624 = pi11 ? n60459 : n60623;
  assign n60625 = pi10 ? n60319 : n60624;
  assign n60626 = pi09 ? n60151 : n60625;
  assign n60627 = pi18 ? n40497 : n60129;
  assign n60628 = pi17 ? n32 : n60627;
  assign n60629 = pi16 ? n32 : n60628;
  assign n60630 = pi15 ? n32 : n60629;
  assign n60631 = pi18 ? n41682 : n60137;
  assign n60632 = pi17 ? n32 : n60631;
  assign n60633 = pi16 ? n32 : n60632;
  assign n60634 = pi18 ? n41682 : n60142;
  assign n60635 = pi17 ? n32 : n60634;
  assign n60636 = pi16 ? n32 : n60635;
  assign n60637 = pi15 ? n60633 : n60636;
  assign n60638 = pi14 ? n60630 : n60637;
  assign n60639 = pi13 ? n32 : n60638;
  assign n60640 = pi12 ? n32 : n60639;
  assign n60641 = pi11 ? n32 : n60640;
  assign n60642 = pi10 ? n32 : n60641;
  assign n60643 = pi18 ? n40510 : n60155;
  assign n60644 = pi17 ? n32 : n60643;
  assign n60645 = pi16 ? n32 : n60644;
  assign n60646 = pi18 ? n39397 : n60155;
  assign n60647 = pi17 ? n32 : n60646;
  assign n60648 = pi16 ? n32 : n60647;
  assign n60649 = pi15 ? n60645 : n60648;
  assign n60650 = pi18 ? n40550 : n60164;
  assign n60651 = pi17 ? n32 : n60650;
  assign n60652 = pi16 ? n32 : n60651;
  assign n60653 = pi18 ? n45413 : n60168;
  assign n60654 = pi17 ? n32 : n60653;
  assign n60655 = pi16 ? n32 : n60654;
  assign n60656 = pi15 ? n60652 : n60655;
  assign n60657 = pi14 ? n60649 : n60656;
  assign n60658 = pi18 ? n45413 : n60155;
  assign n60659 = pi17 ? n32 : n60658;
  assign n60660 = pi16 ? n32 : n60659;
  assign n60661 = pi15 ? n60161 : n60180;
  assign n60662 = pi14 ? n60660 : n60661;
  assign n60663 = pi13 ? n60657 : n60662;
  assign n60664 = pi17 ? n45739 : n60188;
  assign n60665 = pi16 ? n32 : n60664;
  assign n60666 = pi17 ? n46884 : n60188;
  assign n60667 = pi16 ? n32 : n60666;
  assign n60668 = pi15 ? n60665 : n60667;
  assign n60669 = pi17 ? n46884 : n60195;
  assign n60670 = pi16 ? n32 : n60669;
  assign n60671 = pi17 ? n44643 : n60195;
  assign n60672 = pi16 ? n32 : n60671;
  assign n60673 = pi15 ? n60670 : n60672;
  assign n60674 = pi14 ? n60668 : n60673;
  assign n60675 = pi17 ? n44652 : n59297;
  assign n60676 = pi16 ? n32 : n60675;
  assign n60677 = pi17 ? n44222 : n59297;
  assign n60678 = pi16 ? n32 : n60677;
  assign n60679 = pi15 ? n60676 : n60678;
  assign n60680 = pi17 ? n44222 : n59308;
  assign n60681 = pi16 ? n32 : n60680;
  assign n60682 = pi21 ? n60211 : n58086;
  assign n60683 = pi20 ? n20563 : n60682;
  assign n60684 = pi19 ? n20563 : n60683;
  assign n60685 = pi18 ? n20563 : n60684;
  assign n60686 = pi17 ? n44222 : n60685;
  assign n60687 = pi16 ? n32 : n60686;
  assign n60688 = pi15 ? n60681 : n60687;
  assign n60689 = pi14 ? n60679 : n60688;
  assign n60690 = pi13 ? n60674 : n60689;
  assign n60691 = pi12 ? n60663 : n60690;
  assign n60692 = pi17 ? n45242 : n59882;
  assign n60693 = pi16 ? n32 : n60692;
  assign n60694 = pi17 ? n46348 : n59333;
  assign n60695 = pi16 ? n32 : n60694;
  assign n60696 = pi15 ? n60693 : n60695;
  assign n60697 = pi17 ? n44670 : n58925;
  assign n60698 = pi16 ? n32 : n60697;
  assign n60699 = pi17 ? n44670 : n59346;
  assign n60700 = pi16 ? n32 : n60699;
  assign n60701 = pi15 ? n60698 : n60700;
  assign n60702 = pi14 ? n60696 : n60701;
  assign n60703 = pi17 ? n44670 : n60235;
  assign n60704 = pi16 ? n32 : n60703;
  assign n60705 = pi17 ? n44670 : n60241;
  assign n60706 = pi16 ? n32 : n60705;
  assign n60707 = pi15 ? n60704 : n60706;
  assign n60708 = pi17 ? n44670 : n60247;
  assign n60709 = pi16 ? n32 : n60708;
  assign n60710 = pi17 ? n43684 : n60253;
  assign n60711 = pi16 ? n32 : n60710;
  assign n60712 = pi15 ? n60709 : n60711;
  assign n60713 = pi14 ? n60707 : n60712;
  assign n60714 = pi13 ? n60702 : n60713;
  assign n60715 = pi17 ? n43218 : n60261;
  assign n60716 = pi16 ? n32 : n60715;
  assign n60717 = pi17 ? n43218 : n60269;
  assign n60718 = pi16 ? n32 : n60717;
  assign n60719 = pi15 ? n60716 : n60718;
  assign n60720 = pi17 ? n43218 : n59400;
  assign n60721 = pi16 ? n32 : n60720;
  assign n60722 = pi17 ? n43218 : n60280;
  assign n60723 = pi16 ? n32 : n60722;
  assign n60724 = pi15 ? n60721 : n60723;
  assign n60725 = pi14 ? n60719 : n60724;
  assign n60726 = pi17 ? n43218 : n60288;
  assign n60727 = pi16 ? n32 : n60726;
  assign n60728 = pi17 ? n44247 : n60296;
  assign n60729 = pi16 ? n32 : n60728;
  assign n60730 = pi15 ? n60727 : n60729;
  assign n60731 = pi20 ? n60302 : n58967;
  assign n60732 = pi19 ? n20563 : n60731;
  assign n60733 = pi18 ? n20563 : n60732;
  assign n60734 = pi17 ? n44247 : n60733;
  assign n60735 = pi16 ? n32 : n60734;
  assign n60736 = pi17 ? n43223 : n60312;
  assign n60737 = pi16 ? n32 : n60736;
  assign n60738 = pi15 ? n60735 : n60737;
  assign n60739 = pi14 ? n60730 : n60738;
  assign n60740 = pi13 ? n60725 : n60739;
  assign n60741 = pi12 ? n60714 : n60740;
  assign n60742 = pi11 ? n60691 : n60741;
  assign n60743 = pi19 ? n40792 : n58490;
  assign n60744 = pi18 ? n20563 : n60743;
  assign n60745 = pi17 ? n43223 : n60744;
  assign n60746 = pi16 ? n32 : n60745;
  assign n60747 = pi17 ? n43223 : n60324;
  assign n60748 = pi16 ? n32 : n60747;
  assign n60749 = pi15 ? n60746 : n60748;
  assign n60750 = pi22 ? n20563 : n112;
  assign n60751 = pi21 ? n60750 : n14626;
  assign n60752 = pi20 ? n60751 : n5830;
  assign n60753 = pi19 ? n59458 : n60752;
  assign n60754 = pi18 ? n20563 : n60753;
  assign n60755 = pi17 ? n43227 : n60754;
  assign n60756 = pi16 ? n32 : n60755;
  assign n60757 = pi17 ? n43248 : n60338;
  assign n60758 = pi16 ? n32 : n60757;
  assign n60759 = pi15 ? n60756 : n60758;
  assign n60760 = pi14 ? n60749 : n60759;
  assign n60761 = pi17 ? n43248 : n60346;
  assign n60762 = pi16 ? n32 : n60761;
  assign n60763 = pi17 ? n42645 : n60351;
  assign n60764 = pi16 ? n32 : n60763;
  assign n60765 = pi15 ? n60762 : n60764;
  assign n60766 = pi17 ? n42645 : n60360;
  assign n60767 = pi16 ? n32 : n60766;
  assign n60768 = pi21 ? n38375 : n30868;
  assign n60769 = pi20 ? n60768 : n40791;
  assign n60770 = pi19 ? n32 : n60769;
  assign n60771 = pi18 ? n32 : n60770;
  assign n60772 = pi17 ? n60771 : n60371;
  assign n60773 = pi16 ? n32 : n60772;
  assign n60774 = pi15 ? n60767 : n60773;
  assign n60775 = pi14 ? n60765 : n60774;
  assign n60776 = pi13 ? n60760 : n60775;
  assign n60777 = pi21 ? n38375 : n33792;
  assign n60778 = pi20 ? n60777 : n53326;
  assign n60779 = pi19 ? n32 : n60778;
  assign n60780 = pi18 ? n32 : n60779;
  assign n60781 = pi17 ? n60780 : n60387;
  assign n60782 = pi16 ? n32 : n60781;
  assign n60783 = pi21 ? n20563 : n36618;
  assign n60784 = pi20 ? n39395 : n60783;
  assign n60785 = pi19 ? n32 : n60784;
  assign n60786 = pi18 ? n32 : n60785;
  assign n60787 = pi17 ? n60786 : n60403;
  assign n60788 = pi16 ? n32 : n60787;
  assign n60789 = pi15 ? n60782 : n60788;
  assign n60790 = pi22 ? n59056 : n37;
  assign n60791 = pi21 ? n20563 : n60790;
  assign n60792 = pi20 ? n39395 : n60791;
  assign n60793 = pi19 ? n32 : n60792;
  assign n60794 = pi18 ? n32 : n60793;
  assign n60795 = pi22 ? n14626 : n706;
  assign n60796 = pi21 ? n36798 : n60795;
  assign n60797 = pi20 ? n60796 : n32;
  assign n60798 = pi19 ? n60416 : n60797;
  assign n60799 = pi18 ? n20563 : n60798;
  assign n60800 = pi17 ? n60794 : n60799;
  assign n60801 = pi16 ? n32 : n60800;
  assign n60802 = pi17 ? n42201 : n60425;
  assign n60803 = pi16 ? n32 : n60802;
  assign n60804 = pi15 ? n60801 : n60803;
  assign n60805 = pi14 ? n60789 : n60804;
  assign n60806 = pi23 ? n56976 : n33792;
  assign n60807 = pi22 ? n20563 : n60806;
  assign n60808 = pi21 ? n20563 : n60807;
  assign n60809 = pi20 ? n20563 : n60808;
  assign n60810 = pi19 ? n60809 : n59565;
  assign n60811 = pi18 ? n20563 : n60810;
  assign n60812 = pi17 ? n42201 : n60811;
  assign n60813 = pi16 ? n32 : n60812;
  assign n60814 = pi20 ? n60238 : n32;
  assign n60815 = pi19 ? n60809 : n60814;
  assign n60816 = pi18 ? n20563 : n60815;
  assign n60817 = pi17 ? n42681 : n60816;
  assign n60818 = pi16 ? n32 : n60817;
  assign n60819 = pi15 ? n60813 : n60818;
  assign n60820 = pi23 ? n56467 : n36659;
  assign n60821 = pi22 ? n20563 : n60820;
  assign n60822 = pi21 ? n20563 : n60821;
  assign n60823 = pi20 ? n20563 : n60822;
  assign n60824 = pi19 ? n60823 : n59578;
  assign n60825 = pi18 ? n20563 : n60824;
  assign n60826 = pi17 ? n42681 : n60825;
  assign n60827 = pi16 ? n32 : n60826;
  assign n60828 = pi22 ? n112 : n36659;
  assign n60829 = pi21 ? n20563 : n60828;
  assign n60830 = pi20 ? n20563 : n60829;
  assign n60831 = pi21 ? n51564 : n1009;
  assign n60832 = pi20 ? n60831 : n32;
  assign n60833 = pi19 ? n60830 : n60832;
  assign n60834 = pi18 ? n20563 : n60833;
  assign n60835 = pi17 ? n42194 : n60834;
  assign n60836 = pi16 ? n32 : n60835;
  assign n60837 = pi15 ? n60827 : n60836;
  assign n60838 = pi14 ? n60819 : n60837;
  assign n60839 = pi13 ? n60805 : n60838;
  assign n60840 = pi12 ? n60776 : n60839;
  assign n60841 = pi23 ? n56478 : n36781;
  assign n60842 = pi22 ? n30868 : n60841;
  assign n60843 = pi21 ? n20563 : n60842;
  assign n60844 = pi20 ? n20563 : n60843;
  assign n60845 = pi19 ? n60844 : n60465;
  assign n60846 = pi18 ? n20563 : n60845;
  assign n60847 = pi17 ? n42194 : n60846;
  assign n60848 = pi16 ? n32 : n60847;
  assign n60849 = pi17 ? n42194 : n60474;
  assign n60850 = pi16 ? n32 : n60849;
  assign n60851 = pi15 ? n60848 : n60850;
  assign n60852 = pi20 ? n46699 : n42005;
  assign n60853 = pi19 ? n32 : n60852;
  assign n60854 = pi18 ? n32 : n60853;
  assign n60855 = pi17 ? n60854 : n60487;
  assign n60856 = pi16 ? n32 : n60855;
  assign n60857 = pi18 ? n32 : n55089;
  assign n60858 = pi23 ? n157 : n13481;
  assign n60859 = pi22 ? n36659 : n60858;
  assign n60860 = pi21 ? n30868 : n60859;
  assign n60861 = pi20 ? n30868 : n60860;
  assign n60862 = pi19 ? n60861 : n59650;
  assign n60863 = pi18 ? n30868 : n60862;
  assign n60864 = pi17 ? n60857 : n60863;
  assign n60865 = pi16 ? n32 : n60864;
  assign n60866 = pi15 ? n60856 : n60865;
  assign n60867 = pi14 ? n60851 : n60866;
  assign n60868 = pi19 ? n32 : n52230;
  assign n60869 = pi18 ? n32 : n60868;
  assign n60870 = pi17 ? n60869 : n60048;
  assign n60871 = pi16 ? n32 : n60870;
  assign n60872 = pi17 ? n60869 : n60509;
  assign n60873 = pi16 ? n32 : n60872;
  assign n60874 = pi15 ? n60871 : n60873;
  assign n60875 = pi20 ? n45502 : n30868;
  assign n60876 = pi19 ? n32 : n60875;
  assign n60877 = pi18 ? n32 : n60876;
  assign n60878 = pi19 ? n59671 : n52867;
  assign n60879 = pi18 ? n30868 : n60878;
  assign n60880 = pi17 ? n60877 : n60879;
  assign n60881 = pi16 ? n32 : n60880;
  assign n60882 = pi19 ? n60520 : n57717;
  assign n60883 = pi18 ? n30868 : n60882;
  assign n60884 = pi17 ? n49798 : n60883;
  assign n60885 = pi16 ? n32 : n60884;
  assign n60886 = pi15 ? n60881 : n60885;
  assign n60887 = pi14 ? n60874 : n60886;
  assign n60888 = pi13 ? n60867 : n60887;
  assign n60889 = pi17 ? n49798 : n60530;
  assign n60890 = pi16 ? n32 : n60889;
  assign n60891 = pi21 ? n55516 : n54597;
  assign n60892 = pi20 ? n60891 : n55729;
  assign n60893 = pi19 ? n32 : n60892;
  assign n60894 = pi18 ? n32 : n60893;
  assign n60895 = pi22 ? n36762 : n36798;
  assign n60896 = pi21 ? n60895 : n53471;
  assign n60897 = pi20 ? n55729 : n60896;
  assign n60898 = pi19 ? n60897 : n60549;
  assign n60899 = pi18 ? n60898 : n60554;
  assign n60900 = pi17 ? n60894 : n60899;
  assign n60901 = pi16 ? n32 : n60900;
  assign n60902 = pi15 ? n60890 : n60901;
  assign n60903 = pi20 ? n59715 : n33792;
  assign n60904 = pi19 ? n32 : n60903;
  assign n60905 = pi18 ? n32 : n60904;
  assign n60906 = pi17 ? n60905 : n60565;
  assign n60907 = pi16 ? n32 : n60906;
  assign n60908 = pi19 ? n32 : n52446;
  assign n60909 = pi18 ? n32 : n60908;
  assign n60910 = pi22 ? n57197 : n317;
  assign n60911 = pi21 ? n43198 : n60910;
  assign n60912 = pi20 ? n43198 : n60911;
  assign n60913 = pi19 ? n60912 : n32;
  assign n60914 = pi18 ? n59733 : n60913;
  assign n60915 = pi17 ? n60909 : n60914;
  assign n60916 = pi16 ? n32 : n60915;
  assign n60917 = pi15 ? n60907 : n60916;
  assign n60918 = pi14 ? n60902 : n60917;
  assign n60919 = pi22 ? n56622 : n706;
  assign n60920 = pi21 ? n58777 : n60919;
  assign n60921 = pi20 ? n43198 : n60920;
  assign n60922 = pi19 ? n60921 : n32;
  assign n60923 = pi18 ? n43198 : n60922;
  assign n60924 = pi17 ? n60909 : n60923;
  assign n60925 = pi16 ? n32 : n60924;
  assign n60926 = pi21 ? n56760 : n56698;
  assign n60927 = pi20 ? n43198 : n60926;
  assign n60928 = pi19 ? n60927 : n32;
  assign n60929 = pi18 ? n43198 : n60928;
  assign n60930 = pi17 ? n49869 : n60929;
  assign n60931 = pi16 ? n32 : n60930;
  assign n60932 = pi15 ? n60925 : n60931;
  assign n60933 = pi21 ? n32 : n57755;
  assign n60934 = pi22 ? n53550 : n55799;
  assign n60935 = pi21 ? n60934 : n55800;
  assign n60936 = pi20 ? n60933 : n60935;
  assign n60937 = pi19 ? n32 : n60936;
  assign n60938 = pi18 ? n32 : n60937;
  assign n60939 = pi21 ? n47397 : n47396;
  assign n60940 = pi20 ? n60939 : n60597;
  assign n60941 = pi20 ? n60591 : n60599;
  assign n60942 = pi19 ? n60940 : n60941;
  assign n60943 = pi22 ? n157 : n36798;
  assign n60944 = pi21 ? n60943 : n60591;
  assign n60945 = pi20 ? n60944 : n60614;
  assign n60946 = pi19 ? n60945 : n32;
  assign n60947 = pi18 ? n60942 : n60946;
  assign n60948 = pi17 ? n60938 : n60947;
  assign n60949 = pi16 ? n32 : n60948;
  assign n60950 = pi22 ? n45652 : n43198;
  assign n60951 = pi21 ? n32 : n60950;
  assign n60952 = pi20 ? n60951 : n49401;
  assign n60953 = pi19 ? n32 : n60952;
  assign n60954 = pi18 ? n32 : n60953;
  assign n60955 = pi17 ? n60954 : n60617;
  assign n60956 = pi16 ? n32 : n60955;
  assign n60957 = pi15 ? n60949 : n60956;
  assign n60958 = pi14 ? n60932 : n60957;
  assign n60959 = pi13 ? n60918 : n60958;
  assign n60960 = pi12 ? n60888 : n60959;
  assign n60961 = pi11 ? n60840 : n60960;
  assign n60962 = pi10 ? n60742 : n60961;
  assign n60963 = pi09 ? n60642 : n60962;
  assign n60964 = pi08 ? n60626 : n60963;
  assign n60965 = pi07 ? n60125 : n60964;
  assign n60966 = pi20 ? n36250 : n12225;
  assign n60967 = pi19 ? n32294 : n60966;
  assign n60968 = pi18 ? n42239 : n60967;
  assign n60969 = pi17 ? n32 : n60968;
  assign n60970 = pi16 ? n32 : n60969;
  assign n60971 = pi15 ? n32 : n60970;
  assign n60972 = pi20 ? n20563 : n54701;
  assign n60973 = pi23 ? n20563 : n54737;
  assign n60974 = pi22 ? n37 : n60973;
  assign n60975 = pi21 ? n60974 : n37;
  assign n60976 = pi20 ? n60975 : n1619;
  assign n60977 = pi19 ? n60972 : n60976;
  assign n60978 = pi18 ? n42239 : n60977;
  assign n60979 = pi17 ? n32 : n60978;
  assign n60980 = pi16 ? n32 : n60979;
  assign n60981 = pi19 ? n31264 : n34246;
  assign n60982 = pi20 ? n47433 : n39118;
  assign n60983 = pi19 ? n60982 : n60976;
  assign n60984 = pi18 ? n60981 : n60983;
  assign n60985 = pi17 ? n32 : n60984;
  assign n60986 = pi16 ? n32 : n60985;
  assign n60987 = pi15 ? n60980 : n60986;
  assign n60988 = pi14 ? n60971 : n60987;
  assign n60989 = pi13 ? n32 : n60988;
  assign n60990 = pi12 ? n32 : n60989;
  assign n60991 = pi11 ? n32 : n60990;
  assign n60992 = pi10 ? n32 : n60991;
  assign n60993 = pi21 ? n31924 : n35230;
  assign n60994 = pi20 ? n38340 : n60993;
  assign n60995 = pi19 ? n31314 : n60994;
  assign n60996 = pi20 ? n38028 : n37;
  assign n60997 = pi20 ? n33821 : n1619;
  assign n60998 = pi19 ? n60996 : n60997;
  assign n60999 = pi18 ? n60995 : n60998;
  assign n61000 = pi17 ? n32 : n60999;
  assign n61001 = pi16 ? n32 : n61000;
  assign n61002 = pi20 ? n31220 : n1619;
  assign n61003 = pi19 ? n32898 : n61002;
  assign n61004 = pi18 ? n38957 : n61003;
  assign n61005 = pi17 ? n32 : n61004;
  assign n61006 = pi16 ? n32 : n61005;
  assign n61007 = pi15 ? n61001 : n61006;
  assign n61008 = pi21 ? n20563 : n1618;
  assign n61009 = pi20 ? n31220 : n61008;
  assign n61010 = pi19 ? n38478 : n61009;
  assign n61011 = pi18 ? n40045 : n61010;
  assign n61012 = pi17 ? n32 : n61011;
  assign n61013 = pi16 ? n32 : n61012;
  assign n61014 = pi20 ? n20563 : n46815;
  assign n61015 = pi19 ? n61014 : n61009;
  assign n61016 = pi18 ? n40045 : n61015;
  assign n61017 = pi17 ? n32 : n61016;
  assign n61018 = pi16 ? n32 : n61017;
  assign n61019 = pi15 ? n61013 : n61018;
  assign n61020 = pi14 ? n61007 : n61019;
  assign n61021 = pi20 ? n30096 : n1619;
  assign n61022 = pi19 ? n32348 : n61021;
  assign n61023 = pi18 ? n40045 : n61022;
  assign n61024 = pi17 ? n32 : n61023;
  assign n61025 = pi16 ? n32 : n61024;
  assign n61026 = pi20 ? n20563 : n54233;
  assign n61027 = pi19 ? n61026 : n61021;
  assign n61028 = pi18 ? n39397 : n61027;
  assign n61029 = pi17 ? n32 : n61028;
  assign n61030 = pi16 ? n32 : n61029;
  assign n61031 = pi15 ? n61025 : n61030;
  assign n61032 = pi19 ? n61014 : n61021;
  assign n61033 = pi18 ? n39397 : n61032;
  assign n61034 = pi17 ? n32 : n61033;
  assign n61035 = pi16 ? n32 : n61034;
  assign n61036 = pi19 ? n38478 : n61002;
  assign n61037 = pi18 ? n20563 : n61036;
  assign n61038 = pi17 ? n32 : n61037;
  assign n61039 = pi16 ? n32 : n61038;
  assign n61040 = pi15 ? n61035 : n61039;
  assign n61041 = pi14 ? n61031 : n61040;
  assign n61042 = pi13 ? n61020 : n61041;
  assign n61043 = pi19 ? n53012 : n61009;
  assign n61044 = pi18 ? n20563 : n61043;
  assign n61045 = pi17 ? n32 : n61044;
  assign n61046 = pi16 ? n32 : n61045;
  assign n61047 = pi19 ? n53012 : n61021;
  assign n61048 = pi18 ? n20563 : n61047;
  assign n61049 = pi17 ? n45232 : n61048;
  assign n61050 = pi16 ? n32 : n61049;
  assign n61051 = pi20 ? n31903 : n1619;
  assign n61052 = pi19 ? n53012 : n61051;
  assign n61053 = pi18 ? n20563 : n61052;
  assign n61054 = pi17 ? n45232 : n61053;
  assign n61055 = pi16 ? n32 : n61054;
  assign n61056 = pi15 ? n61050 : n61055;
  assign n61057 = pi14 ? n61046 : n61056;
  assign n61058 = pi17 ? n44634 : n59297;
  assign n61059 = pi16 ? n32 : n61058;
  assign n61060 = pi24 ? n37 : n43198;
  assign n61061 = pi23 ? n61060 : n43198;
  assign n61062 = pi22 ? n61061 : n43198;
  assign n61063 = pi24 ? n43198 : n32;
  assign n61064 = pi23 ? n61063 : n32;
  assign n61065 = pi22 ? n43198 : n61064;
  assign n61066 = pi21 ? n61062 : n61065;
  assign n61067 = pi20 ? n20563 : n61066;
  assign n61068 = pi19 ? n20563 : n61067;
  assign n61069 = pi18 ? n20563 : n61068;
  assign n61070 = pi17 ? n45739 : n61069;
  assign n61071 = pi16 ? n32 : n61070;
  assign n61072 = pi15 ? n61059 : n61071;
  assign n61073 = pi20 ? n20563 : n52962;
  assign n61074 = pi20 ? n31220 : n59305;
  assign n61075 = pi19 ? n61073 : n61074;
  assign n61076 = pi18 ? n20563 : n61075;
  assign n61077 = pi17 ? n45739 : n61076;
  assign n61078 = pi16 ? n32 : n61077;
  assign n61079 = pi19 ? n38478 : n20563;
  assign n61080 = pi23 ? n60209 : n685;
  assign n61081 = pi22 ? n61080 : n685;
  assign n61082 = pi21 ? n61081 : n58086;
  assign n61083 = pi20 ? n31220 : n61082;
  assign n61084 = pi19 ? n53012 : n61083;
  assign n61085 = pi18 ? n61079 : n61084;
  assign n61086 = pi17 ? n46884 : n61085;
  assign n61087 = pi16 ? n32 : n61086;
  assign n61088 = pi15 ? n61078 : n61087;
  assign n61089 = pi14 ? n61072 : n61088;
  assign n61090 = pi13 ? n61057 : n61089;
  assign n61091 = pi12 ? n61042 : n61090;
  assign n61092 = pi17 ? n46884 : n59882;
  assign n61093 = pi16 ? n32 : n61092;
  assign n61094 = pi20 ? n45947 : n58922;
  assign n61095 = pi19 ? n20563 : n61094;
  assign n61096 = pi18 ? n20563 : n61095;
  assign n61097 = pi17 ? n44643 : n61096;
  assign n61098 = pi16 ? n32 : n61097;
  assign n61099 = pi15 ? n61093 : n61098;
  assign n61100 = pi22 ? n22383 : n13481;
  assign n61101 = pi21 ? n61100 : n55560;
  assign n61102 = pi20 ? n57578 : n61101;
  assign n61103 = pi19 ? n20563 : n61102;
  assign n61104 = pi18 ? n20563 : n61103;
  assign n61105 = pi17 ? n44652 : n61104;
  assign n61106 = pi16 ? n32 : n61105;
  assign n61107 = pi21 ? n20563 : n569;
  assign n61108 = pi21 ? n43198 : n2637;
  assign n61109 = pi20 ? n61107 : n61108;
  assign n61110 = pi19 ? n20563 : n61109;
  assign n61111 = pi18 ? n20563 : n61110;
  assign n61112 = pi17 ? n44652 : n61111;
  assign n61113 = pi16 ? n32 : n61112;
  assign n61114 = pi15 ? n61106 : n61113;
  assign n61115 = pi14 ? n61099 : n61114;
  assign n61116 = pi21 ? n20563 : n57491;
  assign n61117 = pi20 ? n61116 : n59351;
  assign n61118 = pi19 ? n20563 : n61117;
  assign n61119 = pi18 ? n20563 : n61118;
  assign n61120 = pi17 ? n44652 : n61119;
  assign n61121 = pi16 ? n32 : n61120;
  assign n61122 = pi22 ? n37 : n37783;
  assign n61123 = pi21 ? n20563 : n61122;
  assign n61124 = pi20 ? n61123 : n60238;
  assign n61125 = pi19 ? n20563 : n61124;
  assign n61126 = pi18 ? n20563 : n61125;
  assign n61127 = pi17 ? n44652 : n61126;
  assign n61128 = pi16 ? n32 : n61127;
  assign n61129 = pi15 ? n61121 : n61128;
  assign n61130 = pi17 ? n44222 : n60247;
  assign n61131 = pi16 ? n32 : n61130;
  assign n61132 = pi23 ? n37 : n36781;
  assign n61133 = pi22 ? n37 : n61132;
  assign n61134 = pi21 ? n20563 : n61133;
  assign n61135 = pi20 ? n61134 : n60250;
  assign n61136 = pi19 ? n20563 : n61135;
  assign n61137 = pi18 ? n20563 : n61136;
  assign n61138 = pi17 ? n45242 : n61137;
  assign n61139 = pi16 ? n32 : n61138;
  assign n61140 = pi15 ? n61131 : n61139;
  assign n61141 = pi14 ? n61129 : n61140;
  assign n61142 = pi13 ? n61115 : n61141;
  assign n61143 = pi17 ? n43663 : n60261;
  assign n61144 = pi16 ? n32 : n61143;
  assign n61145 = pi23 ? n37 : n36798;
  assign n61146 = pi22 ? n37 : n61145;
  assign n61147 = pi21 ? n20563 : n61146;
  assign n61148 = pi20 ? n61147 : n59388;
  assign n61149 = pi19 ? n20563 : n61148;
  assign n61150 = pi18 ? n20563 : n61149;
  assign n61151 = pi17 ? n43663 : n61150;
  assign n61152 = pi16 ? n32 : n61151;
  assign n61153 = pi15 ? n61144 : n61152;
  assign n61154 = pi22 ? n37 : n52875;
  assign n61155 = pi21 ? n20563 : n61154;
  assign n61156 = pi22 ? n43198 : n759;
  assign n61157 = pi21 ? n61156 : n32;
  assign n61158 = pi20 ? n61155 : n61157;
  assign n61159 = pi19 ? n20563 : n61158;
  assign n61160 = pi18 ? n20563 : n61159;
  assign n61161 = pi17 ? n43663 : n61160;
  assign n61162 = pi16 ? n32 : n61161;
  assign n61163 = pi23 ? n335 : n43198;
  assign n61164 = pi22 ? n37 : n61163;
  assign n61165 = pi21 ? n20563 : n61164;
  assign n61166 = pi20 ? n61165 : n16944;
  assign n61167 = pi19 ? n20563 : n61166;
  assign n61168 = pi18 ? n20563 : n61167;
  assign n61169 = pi17 ? n43663 : n61168;
  assign n61170 = pi16 ? n32 : n61169;
  assign n61171 = pi15 ? n61162 : n61170;
  assign n61172 = pi14 ? n61153 : n61171;
  assign n61173 = pi20 ? n60293 : n9963;
  assign n61174 = pi19 ? n50863 : n61173;
  assign n61175 = pi18 ? n20563 : n61174;
  assign n61176 = pi17 ? n43663 : n61175;
  assign n61177 = pi16 ? n32 : n61176;
  assign n61178 = pi20 ? n59425 : n55657;
  assign n61179 = pi19 ? n20563 : n61178;
  assign n61180 = pi18 ? n20563 : n61179;
  assign n61181 = pi17 ? n43674 : n61180;
  assign n61182 = pi16 ? n32 : n61181;
  assign n61183 = pi15 ? n61177 : n61182;
  assign n61184 = pi22 ? n13481 : n53982;
  assign n61185 = pi21 ? n61184 : n32;
  assign n61186 = pi20 ? n60309 : n61185;
  assign n61187 = pi19 ? n20563 : n61186;
  assign n61188 = pi18 ? n20563 : n61187;
  assign n61189 = pi17 ? n43684 : n61188;
  assign n61190 = pi16 ? n32 : n61189;
  assign n61191 = pi23 ? n36798 : n316;
  assign n61192 = pi22 ? n33792 : n61191;
  assign n61193 = pi21 ? n20563 : n61192;
  assign n61194 = pi20 ? n61193 : n55668;
  assign n61195 = pi19 ? n20563 : n61194;
  assign n61196 = pi18 ? n20563 : n61195;
  assign n61197 = pi17 ? n43684 : n61196;
  assign n61198 = pi16 ? n32 : n61197;
  assign n61199 = pi15 ? n61190 : n61198;
  assign n61200 = pi14 ? n61183 : n61199;
  assign n61201 = pi13 ? n61172 : n61200;
  assign n61202 = pi12 ? n61142 : n61201;
  assign n61203 = pi11 ? n61091 : n61202;
  assign n61204 = pi22 ? n335 : n13481;
  assign n61205 = pi21 ? n20563 : n61204;
  assign n61206 = pi20 ? n61205 : n56130;
  assign n61207 = pi19 ? n40792 : n61206;
  assign n61208 = pi18 ? n20563 : n61207;
  assign n61209 = pi17 ? n43684 : n61208;
  assign n61210 = pi16 ? n32 : n61209;
  assign n61211 = pi22 ? n36659 : n233;
  assign n61212 = pi21 ? n31294 : n61211;
  assign n61213 = pi20 ? n61212 : n5830;
  assign n61214 = pi19 ? n40792 : n61213;
  assign n61215 = pi18 ? n53297 : n61214;
  assign n61216 = pi17 ? n43684 : n61215;
  assign n61217 = pi16 ? n32 : n61216;
  assign n61218 = pi15 ? n61210 : n61217;
  assign n61219 = pi21 ? n36489 : n2721;
  assign n61220 = pi20 ? n61219 : n10011;
  assign n61221 = pi19 ? n20563 : n61220;
  assign n61222 = pi18 ? n53297 : n61221;
  assign n61223 = pi17 ? n43684 : n61222;
  assign n61224 = pi16 ? n32 : n61223;
  assign n61225 = pi21 ? n39191 : n6461;
  assign n61226 = pi20 ? n61225 : n2653;
  assign n61227 = pi19 ? n20563 : n61226;
  assign n61228 = pi18 ? n55016 : n61227;
  assign n61229 = pi17 ? n44687 : n61228;
  assign n61230 = pi16 ? n32 : n61229;
  assign n61231 = pi15 ? n61224 : n61230;
  assign n61232 = pi14 ? n61218 : n61231;
  assign n61233 = pi22 ? n20563 : n53450;
  assign n61234 = pi22 ? n157 : n13481;
  assign n61235 = pi21 ? n61233 : n61234;
  assign n61236 = pi20 ? n61235 : n37640;
  assign n61237 = pi19 ? n40792 : n61236;
  assign n61238 = pi18 ? n55016 : n61237;
  assign n61239 = pi17 ? n44687 : n61238;
  assign n61240 = pi16 ? n32 : n61239;
  assign n61241 = pi21 ? n20563 : n40912;
  assign n61242 = pi20 ? n40054 : n61241;
  assign n61243 = pi19 ? n32 : n61242;
  assign n61244 = pi18 ? n32 : n61243;
  assign n61245 = pi20 ? n39192 : n42005;
  assign n61246 = pi21 ? n40917 : n39801;
  assign n61247 = pi20 ? n61246 : n42005;
  assign n61248 = pi19 ? n61245 : n61247;
  assign n61249 = pi20 ? n42006 : n53326;
  assign n61250 = pi22 ? n20563 : n40428;
  assign n61251 = pi22 ? n204 : n13481;
  assign n61252 = pi21 ? n61250 : n61251;
  assign n61253 = pi20 ? n61252 : n1822;
  assign n61254 = pi19 ? n61249 : n61253;
  assign n61255 = pi18 ? n61248 : n61254;
  assign n61256 = pi17 ? n61244 : n61255;
  assign n61257 = pi16 ? n32 : n61256;
  assign n61258 = pi15 ? n61240 : n61257;
  assign n61259 = pi20 ? n57040 : n48184;
  assign n61260 = pi19 ? n32 : n61259;
  assign n61261 = pi18 ? n32 : n61260;
  assign n61262 = pi21 ? n36489 : n36659;
  assign n61263 = pi20 ? n20563 : n61262;
  assign n61264 = pi22 ? n30868 : n58710;
  assign n61265 = pi21 ? n61264 : n59691;
  assign n61266 = pi20 ? n61265 : n20953;
  assign n61267 = pi19 ? n61263 : n61266;
  assign n61268 = pi18 ? n30868 : n61267;
  assign n61269 = pi17 ? n61261 : n61268;
  assign n61270 = pi16 ? n32 : n61269;
  assign n61271 = pi21 ? n20563 : n45008;
  assign n61272 = pi20 ? n40054 : n61271;
  assign n61273 = pi19 ? n32 : n61272;
  assign n61274 = pi18 ? n32 : n61273;
  assign n61275 = pi21 ? n30868 : n41489;
  assign n61276 = pi20 ? n61275 : n53307;
  assign n61277 = pi21 ? n40960 : n40957;
  assign n61278 = pi20 ? n61277 : n53307;
  assign n61279 = pi19 ? n61276 : n61278;
  assign n61280 = pi21 ? n45016 : n20563;
  assign n61281 = pi20 ? n61280 : n61262;
  assign n61282 = pi22 ? n30868 : n10400;
  assign n61283 = pi23 ? n8319 : n43198;
  assign n61284 = pi22 ? n61283 : n1407;
  assign n61285 = pi21 ? n61282 : n61284;
  assign n61286 = pi20 ? n61285 : n32;
  assign n61287 = pi19 ? n61281 : n61286;
  assign n61288 = pi18 ? n61279 : n61287;
  assign n61289 = pi17 ? n61274 : n61288;
  assign n61290 = pi16 ? n32 : n61289;
  assign n61291 = pi15 ? n61270 : n61290;
  assign n61292 = pi14 ? n61258 : n61291;
  assign n61293 = pi13 ? n61232 : n61292;
  assign n61294 = pi22 ? n49720 : n36615;
  assign n61295 = pi21 ? n32 : n61294;
  assign n61296 = pi21 ? n45016 : n33792;
  assign n61297 = pi20 ? n61295 : n61296;
  assign n61298 = pi19 ? n32 : n61297;
  assign n61299 = pi18 ? n32 : n61298;
  assign n61300 = pi20 ? n53326 : n40958;
  assign n61301 = pi21 ? n45016 : n40957;
  assign n61302 = pi20 ? n61301 : n40957;
  assign n61303 = pi19 ? n61300 : n61302;
  assign n61304 = pi21 ? n47220 : n36781;
  assign n61305 = pi20 ? n20563 : n61304;
  assign n61306 = pi22 ? n33792 : n56776;
  assign n61307 = pi23 ? n15293 : n14626;
  assign n61308 = pi22 ? n61307 : n317;
  assign n61309 = pi21 ? n61306 : n61308;
  assign n61310 = pi20 ? n61309 : n32;
  assign n61311 = pi19 ? n61305 : n61310;
  assign n61312 = pi18 ? n61303 : n61311;
  assign n61313 = pi17 ? n61299 : n61312;
  assign n61314 = pi16 ? n32 : n61313;
  assign n61315 = pi22 ? n39190 : n37173;
  assign n61316 = pi21 ? n61315 : n36781;
  assign n61317 = pi20 ? n20563 : n61316;
  assign n61318 = pi23 ? n35938 : n685;
  assign n61319 = pi22 ? n61318 : n317;
  assign n61320 = pi21 ? n60483 : n61319;
  assign n61321 = pi20 ? n61320 : n32;
  assign n61322 = pi19 ? n61317 : n61321;
  assign n61323 = pi18 ? n20563 : n61322;
  assign n61324 = pi17 ? n44247 : n61323;
  assign n61325 = pi16 ? n32 : n61324;
  assign n61326 = pi15 ? n61314 : n61325;
  assign n61327 = pi22 ? n42109 : n37783;
  assign n61328 = pi21 ? n61327 : n51270;
  assign n61329 = pi20 ? n20563 : n61328;
  assign n61330 = pi22 ? n36659 : n56026;
  assign n61331 = pi21 ? n61330 : n37547;
  assign n61332 = pi20 ? n61331 : n32;
  assign n61333 = pi19 ? n61329 : n61332;
  assign n61334 = pi18 ? n20563 : n61333;
  assign n61335 = pi17 ? n44247 : n61334;
  assign n61336 = pi16 ? n32 : n61335;
  assign n61337 = pi21 ? n46283 : n55560;
  assign n61338 = pi20 ? n61337 : n32;
  assign n61339 = pi19 ? n56540 : n61338;
  assign n61340 = pi18 ? n20563 : n61339;
  assign n61341 = pi17 ? n44274 : n61340;
  assign n61342 = pi16 ? n32 : n61341;
  assign n61343 = pi15 ? n61336 : n61342;
  assign n61344 = pi14 ? n61326 : n61343;
  assign n61345 = pi22 ? n36781 : n55641;
  assign n61346 = pi21 ? n61345 : n55560;
  assign n61347 = pi20 ? n61346 : n32;
  assign n61348 = pi19 ? n56540 : n61347;
  assign n61349 = pi18 ? n20563 : n61348;
  assign n61350 = pi17 ? n44274 : n61349;
  assign n61351 = pi16 ? n32 : n61350;
  assign n61352 = pi22 ? n20563 : n36798;
  assign n61353 = pi21 ? n20563 : n61352;
  assign n61354 = pi20 ? n20563 : n61353;
  assign n61355 = pi22 ? n36781 : n54664;
  assign n61356 = pi21 ? n61355 : n928;
  assign n61357 = pi20 ? n61356 : n32;
  assign n61358 = pi19 ? n61354 : n61357;
  assign n61359 = pi18 ? n20563 : n61358;
  assign n61360 = pi17 ? n43248 : n61359;
  assign n61361 = pi16 ? n32 : n61360;
  assign n61362 = pi15 ? n61351 : n61361;
  assign n61363 = pi22 ? n30868 : n60820;
  assign n61364 = pi21 ? n20563 : n61363;
  assign n61365 = pi20 ? n20563 : n61364;
  assign n61366 = pi22 ? n36798 : n57197;
  assign n61367 = pi21 ? n61366 : n2700;
  assign n61368 = pi20 ? n61367 : n32;
  assign n61369 = pi19 ? n61365 : n61368;
  assign n61370 = pi18 ? n20563 : n61369;
  assign n61371 = pi17 ? n43248 : n61370;
  assign n61372 = pi16 ? n32 : n61371;
  assign n61373 = pi22 ? n39190 : n36798;
  assign n61374 = pi21 ? n20563 : n61373;
  assign n61375 = pi20 ? n20563 : n61374;
  assign n61376 = pi22 ? n43198 : n56678;
  assign n61377 = pi21 ? n61376 : n1009;
  assign n61378 = pi20 ? n61377 : n32;
  assign n61379 = pi19 ? n61375 : n61378;
  assign n61380 = pi18 ? n20563 : n61379;
  assign n61381 = pi17 ? n44274 : n61380;
  assign n61382 = pi16 ? n32 : n61381;
  assign n61383 = pi15 ? n61372 : n61382;
  assign n61384 = pi14 ? n61362 : n61383;
  assign n61385 = pi13 ? n61344 : n61384;
  assign n61386 = pi12 ? n61293 : n61385;
  assign n61387 = pi22 ? n42109 : n36798;
  assign n61388 = pi21 ? n20563 : n61387;
  assign n61389 = pi20 ? n20563 : n61388;
  assign n61390 = pi22 ? n14626 : n56186;
  assign n61391 = pi21 ? n61390 : n1009;
  assign n61392 = pi20 ? n61391 : n32;
  assign n61393 = pi19 ? n61389 : n61392;
  assign n61394 = pi18 ? n20563 : n61393;
  assign n61395 = pi17 ? n44274 : n61394;
  assign n61396 = pi16 ? n32 : n61395;
  assign n61397 = pi23 ? n55053 : n36798;
  assign n61398 = pi22 ? n33792 : n61397;
  assign n61399 = pi21 ? n20563 : n61398;
  assign n61400 = pi20 ? n20563 : n61399;
  assign n61401 = pi22 ? n51564 : n396;
  assign n61402 = pi21 ? n61401 : n32;
  assign n61403 = pi20 ? n61402 : n32;
  assign n61404 = pi19 ? n61400 : n61403;
  assign n61405 = pi18 ? n44911 : n61404;
  assign n61406 = pi17 ? n44274 : n61405;
  assign n61407 = pi16 ? n32 : n61406;
  assign n61408 = pi15 ? n61396 : n61407;
  assign n61409 = pi20 ? n60023 : n30868;
  assign n61410 = pi19 ? n32 : n61409;
  assign n61411 = pi18 ? n32 : n61410;
  assign n61412 = pi22 ? n36659 : n49412;
  assign n61413 = pi21 ? n30868 : n61412;
  assign n61414 = pi20 ? n30868 : n61413;
  assign n61415 = pi20 ? n58471 : n32;
  assign n61416 = pi19 ? n61414 : n61415;
  assign n61417 = pi18 ? n30868 : n61416;
  assign n61418 = pi17 ? n61411 : n61417;
  assign n61419 = pi16 ? n32 : n61418;
  assign n61420 = pi19 ? n56697 : n60046;
  assign n61421 = pi18 ? n30868 : n61420;
  assign n61422 = pi17 ? n61411 : n61421;
  assign n61423 = pi16 ? n32 : n61422;
  assign n61424 = pi15 ? n61419 : n61423;
  assign n61425 = pi14 ? n61408 : n61424;
  assign n61426 = pi21 ? n32 : n58125;
  assign n61427 = pi20 ? n61426 : n30868;
  assign n61428 = pi19 ? n32 : n61427;
  assign n61429 = pi18 ? n32 : n61428;
  assign n61430 = pi21 ? n30868 : n53551;
  assign n61431 = pi20 ? n30868 : n61430;
  assign n61432 = pi19 ? n61431 : n60046;
  assign n61433 = pi18 ? n30868 : n61432;
  assign n61434 = pi17 ? n61429 : n61433;
  assign n61435 = pi16 ? n32 : n61434;
  assign n61436 = pi21 ? n51313 : n55708;
  assign n61437 = pi20 ? n30868 : n61436;
  assign n61438 = pi19 ? n61437 : n52867;
  assign n61439 = pi18 ? n30868 : n61438;
  assign n61440 = pi17 ? n61429 : n61439;
  assign n61441 = pi16 ? n32 : n61440;
  assign n61442 = pi15 ? n61435 : n61441;
  assign n61443 = pi20 ? n37933 : n41912;
  assign n61444 = pi19 ? n32 : n61443;
  assign n61445 = pi18 ? n32 : n61444;
  assign n61446 = pi22 ? n30868 : n43198;
  assign n61447 = pi21 ? n61446 : n56760;
  assign n61448 = pi20 ? n30868 : n61447;
  assign n61449 = pi19 ? n61448 : n55691;
  assign n61450 = pi18 ? n30868 : n61449;
  assign n61451 = pi17 ? n61445 : n61450;
  assign n61452 = pi16 ? n32 : n61451;
  assign n61453 = pi20 ? n46061 : n30868;
  assign n61454 = pi19 ? n32 : n61453;
  assign n61455 = pi18 ? n32 : n61454;
  assign n61456 = pi21 ? n36798 : n59691;
  assign n61457 = pi20 ? n30868 : n61456;
  assign n61458 = pi19 ? n61457 : n57717;
  assign n61459 = pi18 ? n30868 : n61458;
  assign n61460 = pi17 ? n61455 : n61459;
  assign n61461 = pi16 ? n32 : n61460;
  assign n61462 = pi15 ? n61452 : n61461;
  assign n61463 = pi14 ? n61442 : n61462;
  assign n61464 = pi13 ? n61425 : n61463;
  assign n61465 = pi17 ? n61455 : n60530;
  assign n61466 = pi16 ? n32 : n61465;
  assign n61467 = pi20 ? n54444 : n33792;
  assign n61468 = pi19 ? n32 : n61467;
  assign n61469 = pi18 ? n32 : n61468;
  assign n61470 = pi22 ? n56607 : n56186;
  assign n61471 = pi21 ? n43198 : n61470;
  assign n61472 = pi20 ? n33792 : n61471;
  assign n61473 = pi19 ? n61472 : n32;
  assign n61474 = pi18 ? n33792 : n61473;
  assign n61475 = pi17 ? n61469 : n61474;
  assign n61476 = pi16 ? n32 : n61475;
  assign n61477 = pi15 ? n61466 : n61476;
  assign n61478 = pi21 ? n53463 : n33792;
  assign n61479 = pi20 ? n58727 : n61478;
  assign n61480 = pi21 ? n33792 : n53471;
  assign n61481 = pi20 ? n53485 : n61480;
  assign n61482 = pi19 ? n61479 : n61481;
  assign n61483 = pi21 ? n43198 : n39952;
  assign n61484 = pi23 ? n43198 : n13481;
  assign n61485 = pi22 ? n61484 : n21502;
  assign n61486 = pi21 ? n43198 : n61485;
  assign n61487 = pi20 ? n61483 : n61486;
  assign n61488 = pi19 ? n61487 : n32;
  assign n61489 = pi18 ? n61482 : n61488;
  assign n61490 = pi17 ? n61469 : n61489;
  assign n61491 = pi16 ? n32 : n61490;
  assign n61492 = pi20 ? n46277 : n55716;
  assign n61493 = pi19 ? n32 : n61492;
  assign n61494 = pi18 ? n32 : n61493;
  assign n61495 = pi22 ? n43198 : n61484;
  assign n61496 = pi21 ? n61495 : n59648;
  assign n61497 = pi20 ? n49401 : n61496;
  assign n61498 = pi19 ? n61497 : n32;
  assign n61499 = pi18 ? n43198 : n61498;
  assign n61500 = pi17 ? n61494 : n61499;
  assign n61501 = pi16 ? n32 : n61500;
  assign n61502 = pi15 ? n61491 : n61501;
  assign n61503 = pi14 ? n61477 : n61502;
  assign n61504 = pi21 ? n55792 : n43198;
  assign n61505 = pi20 ? n46277 : n61504;
  assign n61506 = pi19 ? n32 : n61505;
  assign n61507 = pi18 ? n32 : n61506;
  assign n61508 = pi24 ? n43198 : n51564;
  assign n61509 = pi23 ? n36798 : n61508;
  assign n61510 = pi22 ? n43198 : n61509;
  assign n61511 = pi21 ? n61510 : n56129;
  assign n61512 = pi20 ? n43198 : n61511;
  assign n61513 = pi19 ? n61512 : n32;
  assign n61514 = pi18 ? n43198 : n61513;
  assign n61515 = pi17 ? n61507 : n61514;
  assign n61516 = pi16 ? n32 : n61515;
  assign n61517 = pi20 ? n32 : n47397;
  assign n61518 = pi19 ? n32 : n61517;
  assign n61519 = pi18 ? n32 : n61518;
  assign n61520 = pi24 ? n43198 : n13481;
  assign n61521 = pi23 ? n43198 : n61520;
  assign n61522 = pi22 ? n43198 : n61521;
  assign n61523 = pi21 ? n61522 : n56129;
  assign n61524 = pi20 ? n43198 : n61523;
  assign n61525 = pi19 ? n61524 : n32;
  assign n61526 = pi18 ? n43198 : n61525;
  assign n61527 = pi17 ? n61519 : n61526;
  assign n61528 = pi16 ? n32 : n61527;
  assign n61529 = pi15 ? n61516 : n61528;
  assign n61530 = pi20 ? n32 : n54655;
  assign n61531 = pi19 ? n32 : n61530;
  assign n61532 = pi18 ? n32 : n61531;
  assign n61533 = pi21 ? n43198 : n60602;
  assign n61534 = pi20 ? n61533 : n43198;
  assign n61535 = pi19 ? n61534 : n43198;
  assign n61536 = pi21 ? n52452 : n43198;
  assign n61537 = pi21 ? n13481 : n37639;
  assign n61538 = pi20 ? n61536 : n61537;
  assign n61539 = pi19 ? n61538 : n32;
  assign n61540 = pi18 ? n61535 : n61539;
  assign n61541 = pi17 ? n61532 : n61540;
  assign n61542 = pi16 ? n32 : n61541;
  assign n61543 = pi23 ? n14626 : n43198;
  assign n61544 = pi22 ? n55799 : n61543;
  assign n61545 = pi22 ? n43198 : n55799;
  assign n61546 = pi21 ? n61544 : n61545;
  assign n61547 = pi20 ? n46277 : n61546;
  assign n61548 = pi19 ? n32 : n61547;
  assign n61549 = pi18 ? n32 : n61548;
  assign n61550 = pi21 ? n55800 : n43198;
  assign n61551 = pi20 ? n43198 : n61550;
  assign n61552 = pi19 ? n61551 : n43198;
  assign n61553 = pi18 ? n61552 : n60616;
  assign n61554 = pi17 ? n61549 : n61553;
  assign n61555 = pi16 ? n32 : n61554;
  assign n61556 = pi15 ? n61542 : n61555;
  assign n61557 = pi14 ? n61529 : n61556;
  assign n61558 = pi13 ? n61503 : n61557;
  assign n61559 = pi12 ? n61464 : n61558;
  assign n61560 = pi11 ? n61386 : n61559;
  assign n61561 = pi10 ? n61203 : n61560;
  assign n61562 = pi09 ? n60992 : n61561;
  assign n61563 = pi18 ? n41157 : n60967;
  assign n61564 = pi17 ? n32 : n61563;
  assign n61565 = pi16 ? n32 : n61564;
  assign n61566 = pi15 ? n32 : n61565;
  assign n61567 = pi20 ? n20563 : n54155;
  assign n61568 = pi19 ? n38377 : n61567;
  assign n61569 = pi20 ? n36250 : n1619;
  assign n61570 = pi19 ? n60972 : n61569;
  assign n61571 = pi18 ? n61568 : n61570;
  assign n61572 = pi17 ? n32 : n61571;
  assign n61573 = pi16 ? n32 : n61572;
  assign n61574 = pi21 ? n38375 : n31877;
  assign n61575 = pi20 ? n32 : n61574;
  assign n61576 = pi21 ? n31885 : n30867;
  assign n61577 = pi21 ? n31877 : n30843;
  assign n61578 = pi20 ? n61576 : n61577;
  assign n61579 = pi19 ? n61575 : n61578;
  assign n61580 = pi21 ? n29133 : n35230;
  assign n61581 = pi20 ? n61580 : n36250;
  assign n61582 = pi19 ? n61581 : n1620;
  assign n61583 = pi18 ? n61579 : n61582;
  assign n61584 = pi17 ? n32 : n61583;
  assign n61585 = pi16 ? n32 : n61584;
  assign n61586 = pi15 ? n61573 : n61585;
  assign n61587 = pi14 ? n61566 : n61586;
  assign n61588 = pi13 ? n32 : n61587;
  assign n61589 = pi12 ? n32 : n61588;
  assign n61590 = pi11 ? n32 : n61589;
  assign n61591 = pi10 ? n32 : n61590;
  assign n61592 = pi20 ? n46815 : n33821;
  assign n61593 = pi19 ? n28158 : n61592;
  assign n61594 = pi18 ? n61593 : n60998;
  assign n61595 = pi17 ? n32 : n61594;
  assign n61596 = pi16 ? n32 : n61595;
  assign n61597 = pi18 ? n41682 : n61003;
  assign n61598 = pi17 ? n32 : n61597;
  assign n61599 = pi16 ? n32 : n61598;
  assign n61600 = pi15 ? n61596 : n61599;
  assign n61601 = pi18 ? n41682 : n61010;
  assign n61602 = pi17 ? n32 : n61601;
  assign n61603 = pi16 ? n32 : n61602;
  assign n61604 = pi21 ? n31924 : n36249;
  assign n61605 = pi20 ? n20563 : n61604;
  assign n61606 = pi19 ? n61605 : n61009;
  assign n61607 = pi18 ? n41682 : n61606;
  assign n61608 = pi17 ? n32 : n61607;
  assign n61609 = pi16 ? n32 : n61608;
  assign n61610 = pi15 ? n61603 : n61609;
  assign n61611 = pi14 ? n61600 : n61610;
  assign n61612 = pi18 ? n40510 : n61022;
  assign n61613 = pi17 ? n32 : n61612;
  assign n61614 = pi16 ? n32 : n61613;
  assign n61615 = pi18 ? n40510 : n61027;
  assign n61616 = pi17 ? n32 : n61615;
  assign n61617 = pi16 ? n32 : n61616;
  assign n61618 = pi15 ? n61614 : n61617;
  assign n61619 = pi18 ? n39373 : n61032;
  assign n61620 = pi17 ? n32 : n61619;
  assign n61621 = pi16 ? n32 : n61620;
  assign n61622 = pi18 ? n40550 : n61036;
  assign n61623 = pi17 ? n32 : n61622;
  assign n61624 = pi16 ? n32 : n61623;
  assign n61625 = pi15 ? n61621 : n61624;
  assign n61626 = pi14 ? n61618 : n61625;
  assign n61627 = pi13 ? n61611 : n61626;
  assign n61628 = pi18 ? n40550 : n61043;
  assign n61629 = pi17 ? n32 : n61628;
  assign n61630 = pi16 ? n32 : n61629;
  assign n61631 = pi18 ? n45413 : n61043;
  assign n61632 = pi17 ? n32 : n61631;
  assign n61633 = pi16 ? n32 : n61632;
  assign n61634 = pi15 ? n61630 : n61633;
  assign n61635 = pi18 ? n45413 : n61047;
  assign n61636 = pi17 ? n32 : n61635;
  assign n61637 = pi16 ? n32 : n61636;
  assign n61638 = pi18 ? n45413 : n61052;
  assign n61639 = pi17 ? n32 : n61638;
  assign n61640 = pi16 ? n32 : n61639;
  assign n61641 = pi15 ? n61637 : n61640;
  assign n61642 = pi14 ? n61634 : n61641;
  assign n61643 = pi18 ? n38316 : n59296;
  assign n61644 = pi17 ? n32 : n61643;
  assign n61645 = pi16 ? n32 : n61644;
  assign n61646 = pi17 ? n32 : n61069;
  assign n61647 = pi16 ? n32 : n61646;
  assign n61648 = pi15 ? n61645 : n61647;
  assign n61649 = pi17 ? n32 : n61076;
  assign n61650 = pi16 ? n32 : n61649;
  assign n61651 = pi21 ? n58878 : n58086;
  assign n61652 = pi20 ? n31220 : n61651;
  assign n61653 = pi19 ? n53012 : n61652;
  assign n61654 = pi18 ? n61079 : n61653;
  assign n61655 = pi17 ? n32 : n61654;
  assign n61656 = pi16 ? n32 : n61655;
  assign n61657 = pi15 ? n61650 : n61656;
  assign n61658 = pi14 ? n61648 : n61657;
  assign n61659 = pi13 ? n61642 : n61658;
  assign n61660 = pi12 ? n61627 : n61659;
  assign n61661 = pi17 ? n45232 : n59328;
  assign n61662 = pi16 ? n32 : n61661;
  assign n61663 = pi17 ? n45232 : n61096;
  assign n61664 = pi16 ? n32 : n61663;
  assign n61665 = pi15 ? n61662 : n61664;
  assign n61666 = pi17 ? n44634 : n61104;
  assign n61667 = pi16 ? n32 : n61666;
  assign n61668 = pi17 ? n44634 : n61111;
  assign n61669 = pi16 ? n32 : n61668;
  assign n61670 = pi15 ? n61667 : n61669;
  assign n61671 = pi14 ? n61665 : n61670;
  assign n61672 = pi17 ? n44634 : n61119;
  assign n61673 = pi16 ? n32 : n61672;
  assign n61674 = pi17 ? n45739 : n61126;
  assign n61675 = pi16 ? n32 : n61674;
  assign n61676 = pi15 ? n61673 : n61675;
  assign n61677 = pi17 ? n45739 : n60247;
  assign n61678 = pi16 ? n32 : n61677;
  assign n61679 = pi17 ? n50066 : n61137;
  assign n61680 = pi16 ? n32 : n61679;
  assign n61681 = pi15 ? n61678 : n61680;
  assign n61682 = pi14 ? n61676 : n61681;
  assign n61683 = pi13 ? n61671 : n61682;
  assign n61684 = pi17 ? n44643 : n60261;
  assign n61685 = pi16 ? n32 : n61684;
  assign n61686 = pi17 ? n44643 : n61150;
  assign n61687 = pi16 ? n32 : n61686;
  assign n61688 = pi15 ? n61685 : n61687;
  assign n61689 = pi17 ? n44643 : n61160;
  assign n61690 = pi16 ? n32 : n61689;
  assign n61691 = pi17 ? n44643 : n61168;
  assign n61692 = pi16 ? n32 : n61691;
  assign n61693 = pi15 ? n61690 : n61692;
  assign n61694 = pi14 ? n61688 : n61693;
  assign n61695 = pi17 ? n44652 : n61175;
  assign n61696 = pi16 ? n32 : n61695;
  assign n61697 = pi17 ? n44222 : n61180;
  assign n61698 = pi16 ? n32 : n61697;
  assign n61699 = pi15 ? n61696 : n61698;
  assign n61700 = pi20 ? n60309 : n55668;
  assign n61701 = pi19 ? n20563 : n61700;
  assign n61702 = pi18 ? n20563 : n61701;
  assign n61703 = pi17 ? n49594 : n61702;
  assign n61704 = pi16 ? n32 : n61703;
  assign n61705 = pi17 ? n49594 : n61196;
  assign n61706 = pi16 ? n32 : n61705;
  assign n61707 = pi15 ? n61704 : n61706;
  assign n61708 = pi14 ? n61699 : n61707;
  assign n61709 = pi13 ? n61694 : n61708;
  assign n61710 = pi12 ? n61683 : n61709;
  assign n61711 = pi11 ? n61660 : n61710;
  assign n61712 = pi23 ? n13481 : n687;
  assign n61713 = pi22 ? n61712 : n32;
  assign n61714 = pi21 ? n61713 : n32;
  assign n61715 = pi20 ? n61205 : n61714;
  assign n61716 = pi19 ? n40792 : n61715;
  assign n61717 = pi18 ? n20563 : n61716;
  assign n61718 = pi17 ? n49594 : n61717;
  assign n61719 = pi16 ? n32 : n61718;
  assign n61720 = pi22 ? n20563 : n60448;
  assign n61721 = pi21 ? n61720 : n61211;
  assign n61722 = pi20 ? n61721 : n5830;
  assign n61723 = pi19 ? n40792 : n61722;
  assign n61724 = pi18 ? n53297 : n61723;
  assign n61725 = pi17 ? n49594 : n61724;
  assign n61726 = pi16 ? n32 : n61725;
  assign n61727 = pi15 ? n61719 : n61726;
  assign n61728 = pi18 ? n55000 : n61221;
  assign n61729 = pi17 ? n49594 : n61728;
  assign n61730 = pi16 ? n32 : n61729;
  assign n61731 = pi22 ? n20563 : n3492;
  assign n61732 = pi21 ? n61731 : n6461;
  assign n61733 = pi20 ? n61732 : n2653;
  assign n61734 = pi19 ? n20563 : n61733;
  assign n61735 = pi18 ? n55016 : n61734;
  assign n61736 = pi17 ? n43663 : n61735;
  assign n61737 = pi16 ? n32 : n61736;
  assign n61738 = pi15 ? n61730 : n61737;
  assign n61739 = pi14 ? n61727 : n61738;
  assign n61740 = pi20 ? n61235 : n53984;
  assign n61741 = pi19 ? n40792 : n61740;
  assign n61742 = pi18 ? n55016 : n61741;
  assign n61743 = pi17 ? n44670 : n61742;
  assign n61744 = pi16 ? n32 : n61743;
  assign n61745 = pi22 ? n41458 : n40386;
  assign n61746 = pi21 ? n61745 : n30868;
  assign n61747 = pi20 ? n32 : n61746;
  assign n61748 = pi19 ? n32 : n61747;
  assign n61749 = pi18 ? n32 : n61748;
  assign n61750 = pi20 ? n48174 : n42005;
  assign n61751 = pi19 ? n61750 : n61247;
  assign n61752 = pi22 ? n20563 : n49452;
  assign n61753 = pi21 ? n61752 : n61251;
  assign n61754 = pi20 ? n61753 : n1822;
  assign n61755 = pi19 ? n61249 : n61754;
  assign n61756 = pi18 ? n61751 : n61755;
  assign n61757 = pi17 ? n61749 : n61756;
  assign n61758 = pi16 ? n32 : n61757;
  assign n61759 = pi15 ? n61744 : n61758;
  assign n61760 = pi18 ? n32 : n41462;
  assign n61761 = pi23 ? n33792 : n55053;
  assign n61762 = pi22 ? n30868 : n61761;
  assign n61763 = pi21 ? n61762 : n59691;
  assign n61764 = pi20 ? n61763 : n20953;
  assign n61765 = pi19 ? n61263 : n61764;
  assign n61766 = pi18 ? n30868 : n61765;
  assign n61767 = pi17 ? n61760 : n61766;
  assign n61768 = pi16 ? n32 : n61767;
  assign n61769 = pi22 ? n41481 : n36615;
  assign n61770 = pi21 ? n61769 : n33792;
  assign n61771 = pi20 ? n32 : n61770;
  assign n61772 = pi19 ? n32 : n61771;
  assign n61773 = pi18 ? n32 : n61772;
  assign n61774 = pi21 ? n30868 : n54446;
  assign n61775 = pi20 ? n61774 : n53307;
  assign n61776 = pi19 ? n61775 : n61278;
  assign n61777 = pi18 ? n61776 : n61287;
  assign n61778 = pi17 ? n61773 : n61777;
  assign n61779 = pi16 ? n32 : n61778;
  assign n61780 = pi15 ? n61768 : n61779;
  assign n61781 = pi14 ? n61759 : n61780;
  assign n61782 = pi13 ? n61739 : n61781;
  assign n61783 = pi18 ? n32 : n41485;
  assign n61784 = pi24 ? n157 : n43198;
  assign n61785 = pi23 ? n61784 : n14626;
  assign n61786 = pi22 ? n61785 : n317;
  assign n61787 = pi21 ? n61306 : n61786;
  assign n61788 = pi20 ? n61787 : n32;
  assign n61789 = pi19 ? n61305 : n61788;
  assign n61790 = pi18 ? n61303 : n61789;
  assign n61791 = pi17 ? n61783 : n61790;
  assign n61792 = pi16 ? n32 : n61791;
  assign n61793 = pi22 ? n37783 : n43571;
  assign n61794 = pi21 ? n20563 : n61793;
  assign n61795 = pi20 ? n61794 : n20563;
  assign n61796 = pi19 ? n61795 : n20563;
  assign n61797 = pi23 ? n57029 : n685;
  assign n61798 = pi22 ? n61797 : n317;
  assign n61799 = pi21 ? n60483 : n61798;
  assign n61800 = pi20 ? n61799 : n32;
  assign n61801 = pi19 ? n61317 : n61800;
  assign n61802 = pi18 ? n61796 : n61801;
  assign n61803 = pi17 ? n44670 : n61802;
  assign n61804 = pi16 ? n32 : n61803;
  assign n61805 = pi15 ? n61792 : n61804;
  assign n61806 = pi23 ? n685 : n51564;
  assign n61807 = pi22 ? n61806 : n14363;
  assign n61808 = pi21 ? n61330 : n61807;
  assign n61809 = pi20 ? n61808 : n32;
  assign n61810 = pi19 ? n61329 : n61809;
  assign n61811 = pi18 ? n20563 : n61810;
  assign n61812 = pi17 ? n44670 : n61811;
  assign n61813 = pi16 ? n32 : n61812;
  assign n61814 = pi17 ? n43218 : n61340;
  assign n61815 = pi16 ? n32 : n61814;
  assign n61816 = pi15 ? n61813 : n61815;
  assign n61817 = pi14 ? n61805 : n61816;
  assign n61818 = pi17 ? n43218 : n61349;
  assign n61819 = pi16 ? n32 : n61818;
  assign n61820 = pi17 ? n43218 : n61359;
  assign n61821 = pi16 ? n32 : n61820;
  assign n61822 = pi15 ? n61819 : n61821;
  assign n61823 = pi21 ? n20563 : n61264;
  assign n61824 = pi20 ? n20563 : n61823;
  assign n61825 = pi21 ? n61366 : n53983;
  assign n61826 = pi20 ? n61825 : n32;
  assign n61827 = pi19 ? n61824 : n61826;
  assign n61828 = pi18 ? n20563 : n61827;
  assign n61829 = pi17 ? n43674 : n61828;
  assign n61830 = pi16 ? n32 : n61829;
  assign n61831 = pi17 ? n43684 : n61380;
  assign n61832 = pi16 ? n32 : n61831;
  assign n61833 = pi15 ? n61830 : n61832;
  assign n61834 = pi14 ? n61822 : n61833;
  assign n61835 = pi13 ? n61817 : n61834;
  assign n61836 = pi12 ? n61782 : n61835;
  assign n61837 = pi21 ? n61390 : n20952;
  assign n61838 = pi20 ? n61837 : n32;
  assign n61839 = pi19 ? n61389 : n61838;
  assign n61840 = pi18 ? n20563 : n61839;
  assign n61841 = pi17 ? n43684 : n61840;
  assign n61842 = pi16 ? n32 : n61841;
  assign n61843 = pi24 ? n33792 : n36781;
  assign n61844 = pi23 ? n61843 : n36798;
  assign n61845 = pi22 ? n33792 : n61844;
  assign n61846 = pi21 ? n20563 : n61845;
  assign n61847 = pi20 ? n20563 : n61846;
  assign n61848 = pi19 ? n61847 : n61403;
  assign n61849 = pi18 ? n44911 : n61848;
  assign n61850 = pi17 ? n43684 : n61849;
  assign n61851 = pi16 ? n32 : n61850;
  assign n61852 = pi15 ? n61842 : n61851;
  assign n61853 = pi18 ? n32 : n56127;
  assign n61854 = pi17 ? n61853 : n61417;
  assign n61855 = pi16 ? n32 : n61854;
  assign n61856 = pi17 ? n61853 : n61421;
  assign n61857 = pi16 ? n32 : n61856;
  assign n61858 = pi15 ? n61855 : n61857;
  assign n61859 = pi14 ? n61852 : n61858;
  assign n61860 = pi19 ? n32 : n53290;
  assign n61861 = pi18 ? n32 : n61860;
  assign n61862 = pi22 ? n36798 : n55622;
  assign n61863 = pi21 ? n30868 : n61862;
  assign n61864 = pi20 ? n30868 : n61863;
  assign n61865 = pi19 ? n61864 : n60046;
  assign n61866 = pi18 ? n30868 : n61865;
  assign n61867 = pi17 ? n61861 : n61866;
  assign n61868 = pi16 ? n32 : n61867;
  assign n61869 = pi19 ? n61437 : n10012;
  assign n61870 = pi18 ? n30868 : n61869;
  assign n61871 = pi17 ? n61861 : n61870;
  assign n61872 = pi16 ? n32 : n61871;
  assign n61873 = pi15 ? n61868 : n61872;
  assign n61874 = pi20 ? n32 : n41912;
  assign n61875 = pi19 ? n32 : n61874;
  assign n61876 = pi18 ? n32 : n61875;
  assign n61877 = pi17 ? n61876 : n61450;
  assign n61878 = pi16 ? n32 : n61877;
  assign n61879 = pi19 ? n32 : n48328;
  assign n61880 = pi18 ? n32 : n61879;
  assign n61881 = pi19 ? n61457 : n1823;
  assign n61882 = pi18 ? n30868 : n61881;
  assign n61883 = pi17 ? n61880 : n61882;
  assign n61884 = pi16 ? n32 : n61883;
  assign n61885 = pi15 ? n61878 : n61884;
  assign n61886 = pi14 ? n61873 : n61885;
  assign n61887 = pi13 ? n61859 : n61886;
  assign n61888 = pi19 ? n59693 : n35482;
  assign n61889 = pi18 ? n30868 : n61888;
  assign n61890 = pi17 ? n61880 : n61889;
  assign n61891 = pi16 ? n32 : n61890;
  assign n61892 = pi18 ? n32 : n45520;
  assign n61893 = pi22 ? n56607 : n58452;
  assign n61894 = pi21 ? n43198 : n61893;
  assign n61895 = pi20 ? n33792 : n61894;
  assign n61896 = pi19 ? n61895 : n32;
  assign n61897 = pi18 ? n33792 : n61896;
  assign n61898 = pi17 ? n61892 : n61897;
  assign n61899 = pi16 ? n32 : n61898;
  assign n61900 = pi15 ? n61891 : n61899;
  assign n61901 = pi17 ? n61892 : n61489;
  assign n61902 = pi16 ? n32 : n61901;
  assign n61903 = pi19 ? n32 : n53549;
  assign n61904 = pi18 ? n32 : n61903;
  assign n61905 = pi17 ? n61904 : n61499;
  assign n61906 = pi16 ? n32 : n61905;
  assign n61907 = pi15 ? n61902 : n61906;
  assign n61908 = pi14 ? n61900 : n61907;
  assign n61909 = pi22 ? n43198 : n55622;
  assign n61910 = pi21 ? n61909 : n56129;
  assign n61911 = pi20 ? n43198 : n61910;
  assign n61912 = pi19 ? n61911 : n32;
  assign n61913 = pi18 ? n43198 : n61912;
  assign n61914 = pi17 ? n61904 : n61913;
  assign n61915 = pi16 ? n32 : n61914;
  assign n61916 = pi21 ? n48856 : n47397;
  assign n61917 = pi20 ? n32 : n61916;
  assign n61918 = pi19 ? n32 : n61917;
  assign n61919 = pi18 ? n32 : n61918;
  assign n61920 = pi21 ? n55732 : n56129;
  assign n61921 = pi20 ? n43198 : n61920;
  assign n61922 = pi19 ? n61921 : n32;
  assign n61923 = pi18 ? n43198 : n61922;
  assign n61924 = pi17 ? n61919 : n61923;
  assign n61925 = pi16 ? n32 : n61924;
  assign n61926 = pi15 ? n61915 : n61925;
  assign n61927 = pi17 ? n50836 : n61540;
  assign n61928 = pi16 ? n32 : n61927;
  assign n61929 = pi22 ? n32 : n61543;
  assign n61930 = pi22 ? n43198 : n55641;
  assign n61931 = pi21 ? n61929 : n61930;
  assign n61932 = pi20 ? n32 : n61931;
  assign n61933 = pi19 ? n32 : n61932;
  assign n61934 = pi18 ? n32 : n61933;
  assign n61935 = pi24 ? n14626 : n43198;
  assign n61936 = pi23 ? n61935 : n36798;
  assign n61937 = pi22 ? n55641 : n61936;
  assign n61938 = pi21 ? n61937 : n43198;
  assign n61939 = pi20 ? n43198 : n61938;
  assign n61940 = pi19 ? n61939 : n43198;
  assign n61941 = pi21 ? n59691 : n32;
  assign n61942 = pi20 ? n55701 : n61941;
  assign n61943 = pi19 ? n61942 : n32;
  assign n61944 = pi18 ? n61940 : n61943;
  assign n61945 = pi17 ? n61934 : n61944;
  assign n61946 = pi16 ? n32 : n61945;
  assign n61947 = pi15 ? n61928 : n61946;
  assign n61948 = pi14 ? n61926 : n61947;
  assign n61949 = pi13 ? n61908 : n61948;
  assign n61950 = pi12 ? n61887 : n61949;
  assign n61951 = pi11 ? n61836 : n61950;
  assign n61952 = pi10 ? n61711 : n61951;
  assign n61953 = pi09 ? n61591 : n61952;
  assign n61954 = pi08 ? n61562 : n61953;
  assign n61955 = pi20 ? n37439 : n12225;
  assign n61956 = pi19 ? n20563 : n61955;
  assign n61957 = pi18 ? n42206 : n61956;
  assign n61958 = pi17 ? n32 : n61957;
  assign n61959 = pi16 ? n32 : n61958;
  assign n61960 = pi15 ? n32 : n61959;
  assign n61961 = pi20 ? n37439 : n1619;
  assign n61962 = pi19 ? n20563 : n61961;
  assign n61963 = pi18 ? n42206 : n61962;
  assign n61964 = pi17 ? n32 : n61963;
  assign n61965 = pi16 ? n32 : n61964;
  assign n61966 = pi19 ? n32294 : n61569;
  assign n61967 = pi18 ? n40023 : n61966;
  assign n61968 = pi17 ? n32 : n61967;
  assign n61969 = pi16 ? n32 : n61968;
  assign n61970 = pi15 ? n61965 : n61969;
  assign n61971 = pi14 ? n61960 : n61970;
  assign n61972 = pi13 ? n32 : n61971;
  assign n61973 = pi12 ? n32 : n61972;
  assign n61974 = pi11 ? n32 : n61973;
  assign n61975 = pi10 ? n32 : n61974;
  assign n61976 = pi20 ? n31266 : n1619;
  assign n61977 = pi19 ? n60972 : n61976;
  assign n61978 = pi18 ? n41181 : n61977;
  assign n61979 = pi17 ? n32 : n61978;
  assign n61980 = pi16 ? n32 : n61979;
  assign n61981 = pi19 ? n32294 : n61002;
  assign n61982 = pi18 ? n42239 : n61981;
  assign n61983 = pi17 ? n32 : n61982;
  assign n61984 = pi16 ? n32 : n61983;
  assign n61985 = pi15 ? n61980 : n61984;
  assign n61986 = pi19 ? n20563 : n61009;
  assign n61987 = pi18 ? n42239 : n61986;
  assign n61988 = pi17 ? n32 : n61987;
  assign n61989 = pi16 ? n32 : n61988;
  assign n61990 = pi20 ? n33821 : n61008;
  assign n61991 = pi19 ? n37309 : n61990;
  assign n61992 = pi18 ? n47056 : n61991;
  assign n61993 = pi17 ? n32 : n61992;
  assign n61994 = pi16 ? n32 : n61993;
  assign n61995 = pi15 ? n61989 : n61994;
  assign n61996 = pi14 ? n61985 : n61995;
  assign n61997 = pi19 ? n33822 : n60997;
  assign n61998 = pi18 ? n47056 : n61997;
  assign n61999 = pi17 ? n32 : n61998;
  assign n62000 = pi16 ? n32 : n61999;
  assign n62001 = pi20 ? n38961 : n61604;
  assign n62002 = pi19 ? n31314 : n62001;
  assign n62003 = pi19 ? n20563 : n61002;
  assign n62004 = pi18 ? n62002 : n62003;
  assign n62005 = pi17 ? n32 : n62004;
  assign n62006 = pi16 ? n32 : n62005;
  assign n62007 = pi15 ? n62000 : n62006;
  assign n62008 = pi22 ? n60973 : n30195;
  assign n62009 = pi23 ? n54737 : n20563;
  assign n62010 = pi22 ? n30867 : n62009;
  assign n62011 = pi21 ? n62008 : n62010;
  assign n62012 = pi20 ? n32 : n62011;
  assign n62013 = pi21 ? n30195 : n31294;
  assign n62014 = pi20 ? n62013 : n61580;
  assign n62015 = pi19 ? n62012 : n62014;
  assign n62016 = pi21 ? n31885 : n31200;
  assign n62017 = pi20 ? n62016 : n30096;
  assign n62018 = pi19 ? n62017 : n1620;
  assign n62019 = pi18 ? n62015 : n62018;
  assign n62020 = pi17 ? n32 : n62019;
  assign n62021 = pi16 ? n32 : n62020;
  assign n62022 = pi19 ? n38956 : n52963;
  assign n62023 = pi18 ? n62022 : n61003;
  assign n62024 = pi17 ? n32 : n62023;
  assign n62025 = pi16 ? n32 : n62024;
  assign n62026 = pi15 ? n62021 : n62025;
  assign n62027 = pi14 ? n62007 : n62026;
  assign n62028 = pi13 ? n61996 : n62027;
  assign n62029 = pi18 ? n40045 : n61986;
  assign n62030 = pi17 ? n32 : n62029;
  assign n62031 = pi16 ? n32 : n62030;
  assign n62032 = pi15 ? n61013 : n62031;
  assign n62033 = pi20 ? n54155 : n20563;
  assign n62034 = pi19 ? n40044 : n62033;
  assign n62035 = pi19 ? n31904 : n61021;
  assign n62036 = pi18 ? n62034 : n62035;
  assign n62037 = pi17 ? n32 : n62036;
  assign n62038 = pi16 ? n32 : n62037;
  assign n62039 = pi15 ? n62038 : n61030;
  assign n62040 = pi14 ? n62032 : n62039;
  assign n62041 = pi19 ? n39396 : n62033;
  assign n62042 = pi18 ? n62041 : n59296;
  assign n62043 = pi17 ? n32 : n62042;
  assign n62044 = pi16 ? n32 : n62043;
  assign n62045 = pi18 ? n40550 : n61068;
  assign n62046 = pi17 ? n32 : n62045;
  assign n62047 = pi16 ? n32 : n62046;
  assign n62048 = pi15 ? n62044 : n62047;
  assign n62049 = pi20 ? n28157 : n31266;
  assign n62050 = pi19 ? n62049 : n53601;
  assign n62051 = pi20 ? n38966 : n49916;
  assign n62052 = pi19 ? n62051 : n61074;
  assign n62053 = pi18 ? n62050 : n62052;
  assign n62054 = pi17 ? n32 : n62053;
  assign n62055 = pi16 ? n32 : n62054;
  assign n62056 = pi18 ? n45413 : n61653;
  assign n62057 = pi17 ? n32 : n62056;
  assign n62058 = pi16 ? n32 : n62057;
  assign n62059 = pi15 ? n62055 : n62058;
  assign n62060 = pi14 ? n62048 : n62059;
  assign n62061 = pi13 ? n62040 : n62060;
  assign n62062 = pi12 ? n62028 : n62061;
  assign n62063 = pi18 ? n45413 : n59327;
  assign n62064 = pi17 ? n32 : n62063;
  assign n62065 = pi16 ? n32 : n62064;
  assign n62066 = pi20 ? n31263 : n31913;
  assign n62067 = pi20 ? n54701 : n20563;
  assign n62068 = pi19 ? n62066 : n62067;
  assign n62069 = pi21 ? n30843 : n36249;
  assign n62070 = pi20 ? n20563 : n62069;
  assign n62071 = pi21 ? n30843 : n181;
  assign n62072 = pi20 ? n62071 : n58922;
  assign n62073 = pi19 ? n62070 : n62072;
  assign n62074 = pi18 ? n62068 : n62073;
  assign n62075 = pi17 ? n32 : n62074;
  assign n62076 = pi16 ? n32 : n62075;
  assign n62077 = pi15 ? n62065 : n62076;
  assign n62078 = pi23 ? n842 : n13481;
  assign n62079 = pi22 ? n62078 : n13481;
  assign n62080 = pi21 ? n62079 : n55560;
  assign n62081 = pi20 ? n57578 : n62080;
  assign n62082 = pi19 ? n20563 : n62081;
  assign n62083 = pi18 ? n38316 : n62082;
  assign n62084 = pi17 ? n32 : n62083;
  assign n62085 = pi16 ? n32 : n62084;
  assign n62086 = pi20 ? n31313 : n31913;
  assign n62087 = pi19 ? n62086 : n20563;
  assign n62088 = pi18 ? n62087 : n61110;
  assign n62089 = pi17 ? n32 : n62088;
  assign n62090 = pi16 ? n32 : n62089;
  assign n62091 = pi15 ? n62085 : n62090;
  assign n62092 = pi14 ? n62077 : n62091;
  assign n62093 = pi20 ? n61107 : n59351;
  assign n62094 = pi19 ? n20563 : n62093;
  assign n62095 = pi18 ? n38316 : n62094;
  assign n62096 = pi17 ? n32 : n62095;
  assign n62097 = pi16 ? n32 : n62096;
  assign n62098 = pi20 ? n31313 : n47428;
  assign n62099 = pi20 ? n37308 : n54068;
  assign n62100 = pi19 ? n62098 : n62099;
  assign n62101 = pi20 ? n56374 : n60238;
  assign n62102 = pi19 ? n62070 : n62101;
  assign n62103 = pi18 ? n62100 : n62102;
  assign n62104 = pi17 ? n32 : n62103;
  assign n62105 = pi16 ? n32 : n62104;
  assign n62106 = pi15 ? n62097 : n62105;
  assign n62107 = pi17 ? n46325 : n59376;
  assign n62108 = pi16 ? n32 : n62107;
  assign n62109 = pi20 ? n55343 : n59583;
  assign n62110 = pi19 ? n20563 : n62109;
  assign n62111 = pi18 ? n20563 : n62110;
  assign n62112 = pi17 ? n46325 : n62111;
  assign n62113 = pi16 ? n32 : n62112;
  assign n62114 = pi15 ? n62108 : n62113;
  assign n62115 = pi14 ? n62106 : n62114;
  assign n62116 = pi13 ? n62092 : n62115;
  assign n62117 = pi17 ? n45232 : n61150;
  assign n62118 = pi16 ? n32 : n62117;
  assign n62119 = pi21 ? n20563 : n1313;
  assign n62120 = pi20 ? n62119 : n58439;
  assign n62121 = pi19 ? n20563 : n62120;
  assign n62122 = pi18 ? n20563 : n62121;
  assign n62123 = pi17 ? n45232 : n62122;
  assign n62124 = pi16 ? n32 : n62123;
  assign n62125 = pi15 ? n62118 : n62124;
  assign n62126 = pi19 ? n38962 : n20563;
  assign n62127 = pi23 ? n20563 : n43198;
  assign n62128 = pi22 ? n37 : n62127;
  assign n62129 = pi21 ? n20563 : n62128;
  assign n62130 = pi20 ? n62129 : n61157;
  assign n62131 = pi19 ? n20563 : n62130;
  assign n62132 = pi18 ? n62126 : n62131;
  assign n62133 = pi17 ? n45232 : n62132;
  assign n62134 = pi16 ? n32 : n62133;
  assign n62135 = pi23 ? n36659 : n233;
  assign n62136 = pi22 ? n37 : n62135;
  assign n62137 = pi21 ? n20563 : n62136;
  assign n62138 = pi22 ? n233 : n54563;
  assign n62139 = pi21 ? n62138 : n32;
  assign n62140 = pi20 ? n62137 : n62139;
  assign n62141 = pi19 ? n20563 : n62140;
  assign n62142 = pi18 ? n20563 : n62141;
  assign n62143 = pi17 ? n44634 : n62142;
  assign n62144 = pi16 ? n32 : n62143;
  assign n62145 = pi15 ? n62134 : n62144;
  assign n62146 = pi14 ? n62125 : n62145;
  assign n62147 = pi20 ? n20563 : n38340;
  assign n62148 = pi20 ? n38966 : n54155;
  assign n62149 = pi19 ? n62147 : n62148;
  assign n62150 = pi20 ? n31925 : n48905;
  assign n62151 = pi21 ? n36249 : n58463;
  assign n62152 = pi20 ? n62151 : n57425;
  assign n62153 = pi19 ? n62150 : n62152;
  assign n62154 = pi18 ? n62149 : n62153;
  assign n62155 = pi17 ? n44634 : n62154;
  assign n62156 = pi16 ? n32 : n62155;
  assign n62157 = pi20 ? n60302 : n58471;
  assign n62158 = pi19 ? n20563 : n62157;
  assign n62159 = pi18 ? n20563 : n62158;
  assign n62160 = pi17 ? n46884 : n62159;
  assign n62161 = pi16 ? n32 : n62160;
  assign n62162 = pi15 ? n62156 : n62161;
  assign n62163 = pi22 ? n30868 : n60858;
  assign n62164 = pi21 ? n20563 : n62163;
  assign n62165 = pi20 ? n62164 : n55668;
  assign n62166 = pi19 ? n20563 : n62165;
  assign n62167 = pi18 ? n20563 : n62166;
  assign n62168 = pi17 ? n46884 : n62167;
  assign n62169 = pi16 ? n32 : n62168;
  assign n62170 = pi22 ? n33792 : n56936;
  assign n62171 = pi21 ? n20563 : n62170;
  assign n62172 = pi20 ? n62171 : n55668;
  assign n62173 = pi19 ? n20563 : n62172;
  assign n62174 = pi18 ? n20563 : n62173;
  assign n62175 = pi17 ? n46884 : n62174;
  assign n62176 = pi16 ? n32 : n62175;
  assign n62177 = pi15 ? n62169 : n62176;
  assign n62178 = pi14 ? n62162 : n62177;
  assign n62179 = pi13 ? n62146 : n62178;
  assign n62180 = pi12 ? n62116 : n62179;
  assign n62181 = pi11 ? n62062 : n62180;
  assign n62182 = pi20 ? n61205 : n4116;
  assign n62183 = pi19 ? n40792 : n62182;
  assign n62184 = pi18 ? n20563 : n62183;
  assign n62185 = pi17 ? n46884 : n62184;
  assign n62186 = pi16 ? n32 : n62185;
  assign n62187 = pi20 ? n20563 : n54068;
  assign n62188 = pi19 ? n62187 : n20563;
  assign n62189 = pi20 ? n31913 : n40791;
  assign n62190 = pi22 ? n20563 : n20628;
  assign n62191 = pi21 ? n62190 : n61211;
  assign n62192 = pi20 ? n62191 : n5830;
  assign n62193 = pi19 ? n62189 : n62192;
  assign n62194 = pi18 ? n62188 : n62193;
  assign n62195 = pi17 ? n46884 : n62194;
  assign n62196 = pi16 ? n32 : n62195;
  assign n62197 = pi15 ? n62186 : n62196;
  assign n62198 = pi21 ? n39191 : n2721;
  assign n62199 = pi20 ? n62198 : n55690;
  assign n62200 = pi19 ? n20563 : n62199;
  assign n62201 = pi18 ? n20563 : n62200;
  assign n62202 = pi17 ? n50066 : n62201;
  assign n62203 = pi16 ? n32 : n62202;
  assign n62204 = pi23 ? n99 : n54954;
  assign n62205 = pi22 ? n20563 : n62204;
  assign n62206 = pi21 ? n62205 : n6461;
  assign n62207 = pi20 ? n62206 : n37640;
  assign n62208 = pi19 ? n20563 : n62207;
  assign n62209 = pi18 ? n20563 : n62208;
  assign n62210 = pi17 ? n44643 : n62209;
  assign n62211 = pi16 ? n32 : n62210;
  assign n62212 = pi15 ? n62203 : n62211;
  assign n62213 = pi14 ? n62197 : n62212;
  assign n62214 = pi21 ? n56603 : n61234;
  assign n62215 = pi20 ? n62214 : n1822;
  assign n62216 = pi19 ? n40792 : n62215;
  assign n62217 = pi18 ? n20563 : n62216;
  assign n62218 = pi17 ? n45242 : n62217;
  assign n62219 = pi16 ? n32 : n62218;
  assign n62220 = pi21 ? n38375 : n48173;
  assign n62221 = pi20 ? n32 : n62220;
  assign n62222 = pi19 ? n32 : n62221;
  assign n62223 = pi18 ? n32 : n62222;
  assign n62224 = pi20 ? n20563 : n42005;
  assign n62225 = pi19 ? n62224 : n60478;
  assign n62226 = pi20 ? n43010 : n53326;
  assign n62227 = pi23 ? n33792 : n55580;
  assign n62228 = pi22 ? n20563 : n62227;
  assign n62229 = pi21 ? n62228 : n61251;
  assign n62230 = pi20 ? n62229 : n1822;
  assign n62231 = pi19 ? n62226 : n62230;
  assign n62232 = pi18 ? n62225 : n62231;
  assign n62233 = pi17 ? n62223 : n62232;
  assign n62234 = pi16 ? n32 : n62233;
  assign n62235 = pi15 ? n62219 : n62234;
  assign n62236 = pi23 ? n36659 : n55053;
  assign n62237 = pi22 ? n30868 : n62236;
  assign n62238 = pi22 ? n43198 : n2192;
  assign n62239 = pi21 ? n62237 : n62238;
  assign n62240 = pi20 ? n62239 : n32;
  assign n62241 = pi19 ? n61263 : n62240;
  assign n62242 = pi18 ? n30868 : n62241;
  assign n62243 = pi17 ? n45242 : n62242;
  assign n62244 = pi16 ? n32 : n62243;
  assign n62245 = pi20 ? n43010 : n53307;
  assign n62246 = pi20 ? n53326 : n53307;
  assign n62247 = pi19 ? n62245 : n62246;
  assign n62248 = pi23 ? n58538 : n233;
  assign n62249 = pi22 ? n62248 : n1407;
  assign n62250 = pi21 ? n60460 : n62249;
  assign n62251 = pi20 ? n62250 : n32;
  assign n62252 = pi19 ? n61281 : n62251;
  assign n62253 = pi18 ? n62247 : n62252;
  assign n62254 = pi17 ? n45242 : n62253;
  assign n62255 = pi16 ? n32 : n62254;
  assign n62256 = pi15 ? n62244 : n62255;
  assign n62257 = pi14 ? n62235 : n62256;
  assign n62258 = pi13 ? n62213 : n62257;
  assign n62259 = pi22 ? n33792 : n30867;
  assign n62260 = pi21 ? n40917 : n62259;
  assign n62261 = pi23 ? n30868 : n54737;
  assign n62262 = pi22 ? n62261 : n30195;
  assign n62263 = pi21 ? n31877 : n62262;
  assign n62264 = pi20 ? n62260 : n62263;
  assign n62265 = pi22 ? n30867 : n39291;
  assign n62266 = pi21 ? n20563 : n62265;
  assign n62267 = pi20 ? n62266 : n38966;
  assign n62268 = pi19 ? n62264 : n62267;
  assign n62269 = pi21 ? n30195 : n36249;
  assign n62270 = pi20 ? n62269 : n61304;
  assign n62271 = pi23 ? n61784 : n685;
  assign n62272 = pi22 ? n62271 : n21502;
  assign n62273 = pi21 ? n60032 : n62272;
  assign n62274 = pi20 ? n62273 : n32;
  assign n62275 = pi19 ? n62270 : n62274;
  assign n62276 = pi18 ? n62268 : n62275;
  assign n62277 = pi17 ? n45242 : n62276;
  assign n62278 = pi16 ? n32 : n62277;
  assign n62279 = pi20 ? n20563 : n55014;
  assign n62280 = pi19 ? n62279 : n20563;
  assign n62281 = pi21 ? n45016 : n36781;
  assign n62282 = pi20 ? n20563 : n62281;
  assign n62283 = pi23 ? n36781 : n204;
  assign n62284 = pi22 ? n33792 : n62283;
  assign n62285 = pi22 ? n61797 : n21502;
  assign n62286 = pi21 ? n62284 : n62285;
  assign n62287 = pi20 ? n62286 : n32;
  assign n62288 = pi19 ? n62282 : n62287;
  assign n62289 = pi18 ? n62280 : n62288;
  assign n62290 = pi17 ? n46348 : n62289;
  assign n62291 = pi16 ? n32 : n62290;
  assign n62292 = pi15 ? n62278 : n62291;
  assign n62293 = pi22 ? n36659 : n53550;
  assign n62294 = pi21 ? n62293 : n7048;
  assign n62295 = pi20 ? n62294 : n32;
  assign n62296 = pi19 ? n56540 : n62295;
  assign n62297 = pi18 ? n20563 : n62296;
  assign n62298 = pi17 ? n44670 : n62297;
  assign n62299 = pi16 ? n32 : n62298;
  assign n62300 = pi23 ? n36798 : n233;
  assign n62301 = pi22 ? n36781 : n62300;
  assign n62302 = pi21 ? n62301 : n55560;
  assign n62303 = pi20 ? n62302 : n32;
  assign n62304 = pi19 ? n56540 : n62303;
  assign n62305 = pi18 ? n20563 : n62304;
  assign n62306 = pi17 ? n44670 : n62305;
  assign n62307 = pi16 ? n32 : n62306;
  assign n62308 = pi15 ? n62299 : n62307;
  assign n62309 = pi14 ? n62292 : n62308;
  assign n62310 = pi19 ? n56540 : n61357;
  assign n62311 = pi18 ? n20563 : n62310;
  assign n62312 = pi17 ? n49594 : n62311;
  assign n62313 = pi16 ? n32 : n62312;
  assign n62314 = pi21 ? n61355 : n37639;
  assign n62315 = pi20 ? n62314 : n32;
  assign n62316 = pi19 ? n61354 : n62315;
  assign n62317 = pi18 ? n20563 : n62316;
  assign n62318 = pi17 ? n49594 : n62317;
  assign n62319 = pi16 ? n32 : n62318;
  assign n62320 = pi15 ? n62313 : n62319;
  assign n62321 = pi23 ? n20563 : n36798;
  assign n62322 = pi22 ? n62321 : n36798;
  assign n62323 = pi21 ? n20563 : n62322;
  assign n62324 = pi20 ? n20563 : n62323;
  assign n62325 = pi22 ? n36798 : n56678;
  assign n62326 = pi21 ? n62325 : n53983;
  assign n62327 = pi20 ? n62326 : n32;
  assign n62328 = pi19 ? n62324 : n62327;
  assign n62329 = pi18 ? n20563 : n62328;
  assign n62330 = pi17 ? n46348 : n62329;
  assign n62331 = pi16 ? n32 : n62330;
  assign n62332 = pi24 ? n20563 : n33792;
  assign n62333 = pi23 ? n20563 : n62332;
  assign n62334 = pi22 ? n62333 : n36798;
  assign n62335 = pi21 ? n20563 : n62334;
  assign n62336 = pi20 ? n20563 : n62335;
  assign n62337 = pi21 ? n59691 : n1009;
  assign n62338 = pi20 ? n62337 : n32;
  assign n62339 = pi19 ? n62336 : n62338;
  assign n62340 = pi18 ? n20563 : n62339;
  assign n62341 = pi17 ? n49594 : n62340;
  assign n62342 = pi16 ? n32 : n62341;
  assign n62343 = pi15 ? n62331 : n62342;
  assign n62344 = pi14 ? n62320 : n62343;
  assign n62345 = pi13 ? n62309 : n62344;
  assign n62346 = pi12 ? n62258 : n62345;
  assign n62347 = pi22 ? n46172 : n36798;
  assign n62348 = pi21 ? n20563 : n62347;
  assign n62349 = pi20 ? n20563 : n62348;
  assign n62350 = pi19 ? n62349 : n61838;
  assign n62351 = pi18 ? n20563 : n62350;
  assign n62352 = pi17 ? n49594 : n62351;
  assign n62353 = pi16 ? n32 : n62352;
  assign n62354 = pi21 ? n28156 : n39801;
  assign n62355 = pi20 ? n32 : n62354;
  assign n62356 = pi19 ? n32 : n62355;
  assign n62357 = pi18 ? n32 : n62356;
  assign n62358 = pi20 ? n42006 : n38754;
  assign n62359 = pi19 ? n20563 : n62358;
  assign n62360 = pi23 ? n36659 : n56064;
  assign n62361 = pi23 ? n56079 : n51564;
  assign n62362 = pi22 ? n62360 : n62361;
  assign n62363 = pi21 ? n36489 : n62362;
  assign n62364 = pi20 ? n20563 : n62363;
  assign n62365 = pi22 ? n51564 : n55688;
  assign n62366 = pi21 ? n62365 : n32;
  assign n62367 = pi20 ? n62366 : n32;
  assign n62368 = pi19 ? n62364 : n62367;
  assign n62369 = pi18 ? n62359 : n62368;
  assign n62370 = pi17 ? n62357 : n62369;
  assign n62371 = pi16 ? n32 : n62370;
  assign n62372 = pi15 ? n62353 : n62371;
  assign n62373 = pi21 ? n28156 : n30868;
  assign n62374 = pi20 ? n32 : n62373;
  assign n62375 = pi19 ? n32 : n62374;
  assign n62376 = pi18 ? n32 : n62375;
  assign n62377 = pi23 ? n36781 : n51564;
  assign n62378 = pi22 ? n38284 : n62377;
  assign n62379 = pi21 ? n30868 : n62378;
  assign n62380 = pi20 ? n30868 : n62379;
  assign n62381 = pi19 ? n62380 : n61415;
  assign n62382 = pi18 ? n30868 : n62381;
  assign n62383 = pi17 ? n62376 : n62382;
  assign n62384 = pi16 ? n32 : n62383;
  assign n62385 = pi21 ? n46060 : n36489;
  assign n62386 = pi20 ? n32 : n62385;
  assign n62387 = pi19 ? n32 : n62386;
  assign n62388 = pi18 ? n32 : n62387;
  assign n62389 = pi23 ? n36798 : n13481;
  assign n62390 = pi22 ? n49412 : n62389;
  assign n62391 = pi21 ? n55685 : n62390;
  assign n62392 = pi20 ? n30868 : n62391;
  assign n62393 = pi19 ? n62392 : n60046;
  assign n62394 = pi18 ? n30868 : n62393;
  assign n62395 = pi17 ? n62388 : n62394;
  assign n62396 = pi16 ? n32 : n62395;
  assign n62397 = pi15 ? n62384 : n62396;
  assign n62398 = pi14 ? n62372 : n62397;
  assign n62399 = pi22 ? n36798 : n62389;
  assign n62400 = pi21 ? n55685 : n62399;
  assign n62401 = pi20 ? n30868 : n62400;
  assign n62402 = pi19 ? n62401 : n60046;
  assign n62403 = pi18 ? n30868 : n62402;
  assign n62404 = pi17 ? n62388 : n62403;
  assign n62405 = pi16 ? n32 : n62404;
  assign n62406 = pi21 ? n47321 : n48173;
  assign n62407 = pi20 ? n32 : n62406;
  assign n62408 = pi19 ? n32 : n62407;
  assign n62409 = pi18 ? n32 : n62408;
  assign n62410 = pi24 ? n36798 : n13481;
  assign n62411 = pi23 ? n62410 : n13481;
  assign n62412 = pi22 ? n36798 : n62411;
  assign n62413 = pi21 ? n51313 : n62412;
  assign n62414 = pi20 ? n30868 : n62413;
  assign n62415 = pi19 ? n62414 : n55691;
  assign n62416 = pi18 ? n30868 : n62415;
  assign n62417 = pi17 ? n62409 : n62416;
  assign n62418 = pi16 ? n32 : n62417;
  assign n62419 = pi15 ? n62405 : n62418;
  assign n62420 = pi22 ? n43198 : n56607;
  assign n62421 = pi21 ? n51313 : n62420;
  assign n62422 = pi20 ? n30868 : n62421;
  assign n62423 = pi19 ? n62422 : n57717;
  assign n62424 = pi18 ? n30868 : n62423;
  assign n62425 = pi17 ? n62409 : n62424;
  assign n62426 = pi16 ? n32 : n62425;
  assign n62427 = pi23 ? n61520 : n13481;
  assign n62428 = pi22 ? n43198 : n62427;
  assign n62429 = pi21 ? n36798 : n62428;
  assign n62430 = pi20 ? n30868 : n62429;
  assign n62431 = pi19 ? n62430 : n35482;
  assign n62432 = pi18 ? n30868 : n62431;
  assign n62433 = pi17 ? n51290 : n62432;
  assign n62434 = pi16 ? n32 : n62433;
  assign n62435 = pi15 ? n62426 : n62434;
  assign n62436 = pi14 ? n62419 : n62435;
  assign n62437 = pi13 ? n62398 : n62436;
  assign n62438 = pi22 ? n55641 : n56186;
  assign n62439 = pi21 ? n43198 : n62438;
  assign n62440 = pi20 ? n30868 : n62439;
  assign n62441 = pi19 ? n62440 : n35482;
  assign n62442 = pi18 ? n30868 : n62441;
  assign n62443 = pi17 ? n51290 : n62442;
  assign n62444 = pi16 ? n32 : n62443;
  assign n62445 = pi21 ? n32 : n33792;
  assign n62446 = pi20 ? n32 : n62445;
  assign n62447 = pi19 ? n32 : n62446;
  assign n62448 = pi18 ? n32 : n62447;
  assign n62449 = pi22 ? n54664 : n58452;
  assign n62450 = pi21 ? n43198 : n62449;
  assign n62451 = pi20 ? n33792 : n62450;
  assign n62452 = pi19 ? n62451 : n32;
  assign n62453 = pi18 ? n33792 : n62452;
  assign n62454 = pi17 ? n62448 : n62453;
  assign n62455 = pi16 ? n32 : n62454;
  assign n62456 = pi15 ? n62444 : n62455;
  assign n62457 = pi21 ? n46260 : n43198;
  assign n62458 = pi20 ? n43198 : n62457;
  assign n62459 = pi21 ? n50795 : n56148;
  assign n62460 = pi20 ? n62459 : n54655;
  assign n62461 = pi19 ? n62458 : n62460;
  assign n62462 = pi21 ? n43198 : n37878;
  assign n62463 = pi20 ? n62462 : n59156;
  assign n62464 = pi19 ? n62463 : n32;
  assign n62465 = pi18 ? n62461 : n62464;
  assign n62466 = pi17 ? n62448 : n62465;
  assign n62467 = pi16 ? n32 : n62466;
  assign n62468 = pi22 ? n43198 : n37276;
  assign n62469 = pi21 ? n32 : n62468;
  assign n62470 = pi20 ? n32 : n62469;
  assign n62471 = pi19 ? n32 : n62470;
  assign n62472 = pi18 ? n32 : n62471;
  assign n62473 = pi23 ? n51564 : n316;
  assign n62474 = pi22 ? n62473 : n21502;
  assign n62475 = pi21 ? n58777 : n62474;
  assign n62476 = pi20 ? n49401 : n62475;
  assign n62477 = pi19 ? n62476 : n32;
  assign n62478 = pi18 ? n43198 : n62477;
  assign n62479 = pi17 ? n62472 : n62478;
  assign n62480 = pi16 ? n32 : n62479;
  assign n62481 = pi15 ? n62467 : n62480;
  assign n62482 = pi14 ? n62456 : n62481;
  assign n62483 = pi22 ? n46275 : n43199;
  assign n62484 = pi21 ? n32 : n62483;
  assign n62485 = pi20 ? n32 : n62484;
  assign n62486 = pi19 ? n32 : n62485;
  assign n62487 = pi18 ? n32 : n62486;
  assign n62488 = pi21 ? n56760 : n56129;
  assign n62489 = pi20 ? n43198 : n62488;
  assign n62490 = pi19 ? n62489 : n32;
  assign n62491 = pi18 ? n43198 : n62490;
  assign n62492 = pi17 ? n62487 : n62491;
  assign n62493 = pi16 ? n32 : n62492;
  assign n62494 = pi21 ? n56760 : n57097;
  assign n62495 = pi20 ? n43198 : n62494;
  assign n62496 = pi19 ? n62495 : n32;
  assign n62497 = pi18 ? n43198 : n62496;
  assign n62498 = pi17 ? n62487 : n62497;
  assign n62499 = pi16 ? n32 : n62498;
  assign n62500 = pi15 ? n62493 : n62499;
  assign n62501 = pi19 ? n59700 : n43198;
  assign n62502 = pi20 ? n54009 : n59604;
  assign n62503 = pi19 ? n62502 : n32;
  assign n62504 = pi18 ? n62501 : n62503;
  assign n62505 = pi17 ? n51333 : n62504;
  assign n62506 = pi16 ? n32 : n62505;
  assign n62507 = pi20 ? n32 : n47342;
  assign n62508 = pi19 ? n32 : n62507;
  assign n62509 = pi18 ? n32 : n62508;
  assign n62510 = pi23 ? n14626 : n36798;
  assign n62511 = pi22 ? n62510 : n43198;
  assign n62512 = pi21 ? n62511 : n43198;
  assign n62513 = pi20 ? n62512 : n55701;
  assign n62514 = pi19 ? n62513 : n43198;
  assign n62515 = pi22 ? n56607 : n13481;
  assign n62516 = pi21 ? n62515 : n32;
  assign n62517 = pi20 ? n55701 : n62516;
  assign n62518 = pi19 ? n62517 : n32;
  assign n62519 = pi18 ? n62514 : n62518;
  assign n62520 = pi17 ? n62509 : n62519;
  assign n62521 = pi16 ? n32 : n62520;
  assign n62522 = pi15 ? n62506 : n62521;
  assign n62523 = pi14 ? n62500 : n62522;
  assign n62524 = pi13 ? n62482 : n62523;
  assign n62525 = pi12 ? n62437 : n62524;
  assign n62526 = pi11 ? n62346 : n62525;
  assign n62527 = pi10 ? n62181 : n62526;
  assign n62528 = pi09 ? n61975 : n62527;
  assign n62529 = pi18 ? n43254 : n61956;
  assign n62530 = pi17 ? n32 : n62529;
  assign n62531 = pi16 ? n32 : n62530;
  assign n62532 = pi15 ? n32 : n62531;
  assign n62533 = pi18 ? n42200 : n61962;
  assign n62534 = pi17 ? n32 : n62533;
  assign n62535 = pi16 ? n32 : n62534;
  assign n62536 = pi20 ? n51988 : n1619;
  assign n62537 = pi19 ? n32294 : n62536;
  assign n62538 = pi18 ? n46997 : n62537;
  assign n62539 = pi17 ? n32 : n62538;
  assign n62540 = pi16 ? n32 : n62539;
  assign n62541 = pi15 ? n62535 : n62540;
  assign n62542 = pi14 ? n62532 : n62541;
  assign n62543 = pi13 ? n32 : n62542;
  assign n62544 = pi12 ? n32 : n62543;
  assign n62545 = pi11 ? n32 : n62544;
  assign n62546 = pi10 ? n32 : n62545;
  assign n62547 = pi19 ? n20563 : n61976;
  assign n62548 = pi18 ? n40485 : n62547;
  assign n62549 = pi17 ? n32 : n62548;
  assign n62550 = pi16 ? n32 : n62549;
  assign n62551 = pi18 ? n41157 : n61981;
  assign n62552 = pi17 ? n32 : n62551;
  assign n62553 = pi16 ? n32 : n62552;
  assign n62554 = pi15 ? n62550 : n62553;
  assign n62555 = pi18 ? n41157 : n61986;
  assign n62556 = pi17 ? n32 : n62555;
  assign n62557 = pi16 ? n32 : n62556;
  assign n62558 = pi19 ? n60972 : n61009;
  assign n62559 = pi18 ? n41168 : n62558;
  assign n62560 = pi17 ? n32 : n62559;
  assign n62561 = pi16 ? n32 : n62560;
  assign n62562 = pi15 ? n62557 : n62561;
  assign n62563 = pi14 ? n62554 : n62562;
  assign n62564 = pi19 ? n31221 : n60997;
  assign n62565 = pi18 ? n41168 : n62564;
  assign n62566 = pi17 ? n32 : n62565;
  assign n62567 = pi16 ? n32 : n62566;
  assign n62568 = pi19 ? n39454 : n38962;
  assign n62569 = pi18 ? n62568 : n62003;
  assign n62570 = pi17 ? n32 : n62569;
  assign n62571 = pi16 ? n32 : n62570;
  assign n62572 = pi15 ? n62567 : n62571;
  assign n62573 = pi20 ? n38966 : n61604;
  assign n62574 = pi19 ? n30118 : n62573;
  assign n62575 = pi20 ? n38028 : n33821;
  assign n62576 = pi20 ? n35231 : n1619;
  assign n62577 = pi19 ? n62575 : n62576;
  assign n62578 = pi18 ? n62574 : n62577;
  assign n62579 = pi17 ? n32 : n62578;
  assign n62580 = pi16 ? n32 : n62579;
  assign n62581 = pi19 ? n41681 : n62033;
  assign n62582 = pi19 ? n33822 : n61002;
  assign n62583 = pi18 ? n62581 : n62582;
  assign n62584 = pi17 ? n32 : n62583;
  assign n62585 = pi16 ? n32 : n62584;
  assign n62586 = pi15 ? n62580 : n62585;
  assign n62587 = pi14 ? n62572 : n62586;
  assign n62588 = pi13 ? n62563 : n62587;
  assign n62589 = pi19 ? n54080 : n61009;
  assign n62590 = pi18 ? n41682 : n62589;
  assign n62591 = pi17 ? n32 : n62590;
  assign n62592 = pi16 ? n32 : n62591;
  assign n62593 = pi18 ? n41682 : n61986;
  assign n62594 = pi17 ? n32 : n62593;
  assign n62595 = pi16 ? n32 : n62594;
  assign n62596 = pi15 ? n62592 : n62595;
  assign n62597 = pi19 ? n32898 : n60997;
  assign n62598 = pi18 ? n40510 : n62597;
  assign n62599 = pi17 ? n32 : n62598;
  assign n62600 = pi16 ? n32 : n62599;
  assign n62601 = pi19 ? n38478 : n60997;
  assign n62602 = pi18 ? n40510 : n62601;
  assign n62603 = pi17 ? n32 : n62602;
  assign n62604 = pi16 ? n32 : n62603;
  assign n62605 = pi15 ? n62600 : n62604;
  assign n62606 = pi14 ? n62596 : n62605;
  assign n62607 = pi18 ? n39373 : n59296;
  assign n62608 = pi17 ? n32 : n62607;
  assign n62609 = pi16 ? n32 : n62608;
  assign n62610 = pi18 ? n38957 : n61068;
  assign n62611 = pi17 ? n32 : n62610;
  assign n62612 = pi16 ? n32 : n62611;
  assign n62613 = pi15 ? n62609 : n62612;
  assign n62614 = pi20 ? n38376 : n31913;
  assign n62615 = pi19 ? n62614 : n20563;
  assign n62616 = pi19 ? n62070 : n61074;
  assign n62617 = pi18 ? n62615 : n62616;
  assign n62618 = pi17 ? n32 : n62617;
  assign n62619 = pi16 ? n32 : n62618;
  assign n62620 = pi19 ? n61026 : n61652;
  assign n62621 = pi18 ? n40045 : n62620;
  assign n62622 = pi17 ? n32 : n62621;
  assign n62623 = pi16 ? n32 : n62622;
  assign n62624 = pi15 ? n62619 : n62623;
  assign n62625 = pi14 ? n62613 : n62624;
  assign n62626 = pi13 ? n62606 : n62625;
  assign n62627 = pi12 ? n62588 : n62626;
  assign n62628 = pi24 ? n36781 : n685;
  assign n62629 = pi23 ? n62628 : n685;
  assign n62630 = pi22 ? n62629 : n685;
  assign n62631 = pi21 ? n62630 : n7723;
  assign n62632 = pi20 ? n54354 : n62631;
  assign n62633 = pi19 ? n20563 : n62632;
  assign n62634 = pi18 ? n40045 : n62633;
  assign n62635 = pi17 ? n32 : n62634;
  assign n62636 = pi16 ? n32 : n62635;
  assign n62637 = pi24 ? n36798 : n316;
  assign n62638 = pi23 ? n62637 : n316;
  assign n62639 = pi22 ? n62638 : n316;
  assign n62640 = pi21 ? n62639 : n2320;
  assign n62641 = pi20 ? n45947 : n62640;
  assign n62642 = pi19 ? n62070 : n62641;
  assign n62643 = pi18 ? n39397 : n62642;
  assign n62644 = pi17 ? n32 : n62643;
  assign n62645 = pi16 ? n32 : n62644;
  assign n62646 = pi15 ? n62636 : n62645;
  assign n62647 = pi22 ? n62411 : n13481;
  assign n62648 = pi21 ? n62647 : n55560;
  assign n62649 = pi20 ? n57578 : n62648;
  assign n62650 = pi19 ? n20563 : n62649;
  assign n62651 = pi18 ? n39397 : n62650;
  assign n62652 = pi17 ? n32 : n62651;
  assign n62653 = pi16 ? n32 : n62652;
  assign n62654 = pi18 ? n39397 : n61110;
  assign n62655 = pi17 ? n32 : n62654;
  assign n62656 = pi16 ? n32 : n62655;
  assign n62657 = pi15 ? n62653 : n62656;
  assign n62658 = pi14 ? n62646 : n62657;
  assign n62659 = pi18 ? n39397 : n62094;
  assign n62660 = pi17 ? n32 : n62659;
  assign n62661 = pi16 ? n32 : n62660;
  assign n62662 = pi19 ? n42192 : n62067;
  assign n62663 = pi18 ? n62662 : n62102;
  assign n62664 = pi17 ? n32 : n62663;
  assign n62665 = pi16 ? n32 : n62664;
  assign n62666 = pi15 ? n62661 : n62665;
  assign n62667 = pi18 ? n45392 : n59375;
  assign n62668 = pi17 ? n32 : n62667;
  assign n62669 = pi16 ? n32 : n62668;
  assign n62670 = pi18 ? n45392 : n62110;
  assign n62671 = pi17 ? n32 : n62670;
  assign n62672 = pi16 ? n32 : n62671;
  assign n62673 = pi15 ? n62669 : n62672;
  assign n62674 = pi14 ? n62666 : n62673;
  assign n62675 = pi13 ? n62658 : n62674;
  assign n62676 = pi20 ? n61147 : n58439;
  assign n62677 = pi19 ? n20563 : n62676;
  assign n62678 = pi18 ? n45413 : n62677;
  assign n62679 = pi17 ? n32 : n62678;
  assign n62680 = pi16 ? n32 : n62679;
  assign n62681 = pi18 ? n45413 : n62121;
  assign n62682 = pi17 ? n32 : n62681;
  assign n62683 = pi16 ? n32 : n62682;
  assign n62684 = pi15 ? n62680 : n62683;
  assign n62685 = pi18 ? n45413 : n62131;
  assign n62686 = pi17 ? n32 : n62685;
  assign n62687 = pi16 ? n32 : n62686;
  assign n62688 = pi18 ? n45413 : n62141;
  assign n62689 = pi17 ? n32 : n62688;
  assign n62690 = pi16 ? n32 : n62689;
  assign n62691 = pi15 ? n62687 : n62690;
  assign n62692 = pi14 ? n62684 : n62691;
  assign n62693 = pi21 ? n31924 : n31877;
  assign n62694 = pi20 ? n20563 : n62693;
  assign n62695 = pi19 ? n62694 : n20563;
  assign n62696 = pi21 ? n31885 : n58463;
  assign n62697 = pi20 ? n62696 : n57425;
  assign n62698 = pi19 ? n53012 : n62697;
  assign n62699 = pi18 ? n62695 : n62698;
  assign n62700 = pi17 ? n32 : n62699;
  assign n62701 = pi16 ? n32 : n62700;
  assign n62702 = pi17 ? n32 : n62159;
  assign n62703 = pi16 ? n32 : n62702;
  assign n62704 = pi15 ? n62701 : n62703;
  assign n62705 = pi20 ? n62164 : n56130;
  assign n62706 = pi19 ? n20563 : n62705;
  assign n62707 = pi18 ? n20563 : n62706;
  assign n62708 = pi17 ? n32 : n62707;
  assign n62709 = pi16 ? n32 : n62708;
  assign n62710 = pi20 ? n62171 : n56130;
  assign n62711 = pi19 ? n20563 : n62710;
  assign n62712 = pi18 ? n20563 : n62711;
  assign n62713 = pi17 ? n32 : n62712;
  assign n62714 = pi16 ? n32 : n62713;
  assign n62715 = pi15 ? n62709 : n62714;
  assign n62716 = pi14 ? n62704 : n62715;
  assign n62717 = pi13 ? n62692 : n62716;
  assign n62718 = pi12 ? n62675 : n62717;
  assign n62719 = pi11 ? n62627 : n62718;
  assign n62720 = pi17 ? n32 : n62184;
  assign n62721 = pi16 ? n32 : n62720;
  assign n62722 = pi18 ? n20563 : n61723;
  assign n62723 = pi17 ? n46325 : n62722;
  assign n62724 = pi16 ? n32 : n62723;
  assign n62725 = pi15 ? n62721 : n62724;
  assign n62726 = pi21 ? n57086 : n2721;
  assign n62727 = pi20 ? n62726 : n57716;
  assign n62728 = pi19 ? n20563 : n62727;
  assign n62729 = pi18 ? n20563 : n62728;
  assign n62730 = pi17 ? n46325 : n62729;
  assign n62731 = pi16 ? n32 : n62730;
  assign n62732 = pi23 ? n99 : n55567;
  assign n62733 = pi22 ? n20563 : n62732;
  assign n62734 = pi21 ? n62733 : n6461;
  assign n62735 = pi20 ? n62734 : n37640;
  assign n62736 = pi19 ? n20563 : n62735;
  assign n62737 = pi18 ? n20563 : n62736;
  assign n62738 = pi17 ? n50066 : n62737;
  assign n62739 = pi16 ? n32 : n62738;
  assign n62740 = pi15 ? n62731 : n62739;
  assign n62741 = pi14 ? n62725 : n62740;
  assign n62742 = pi23 ? n30868 : n56478;
  assign n62743 = pi22 ? n20563 : n62742;
  assign n62744 = pi21 ? n62743 : n61234;
  assign n62745 = pi20 ? n62744 : n20953;
  assign n62746 = pi19 ? n40792 : n62745;
  assign n62747 = pi18 ? n20563 : n62746;
  assign n62748 = pi17 ? n44634 : n62747;
  assign n62749 = pi16 ? n32 : n62748;
  assign n62750 = pi20 ? n62229 : n20953;
  assign n62751 = pi19 ? n62226 : n62750;
  assign n62752 = pi18 ? n62225 : n62751;
  assign n62753 = pi17 ? n51210 : n62752;
  assign n62754 = pi16 ? n32 : n62753;
  assign n62755 = pi15 ? n62749 : n62754;
  assign n62756 = pi23 ? n36659 : n19714;
  assign n62757 = pi22 ? n30868 : n62756;
  assign n62758 = pi21 ? n62757 : n62238;
  assign n62759 = pi20 ? n62758 : n32;
  assign n62760 = pi19 ? n61263 : n62759;
  assign n62761 = pi18 ? n30868 : n62760;
  assign n62762 = pi17 ? n44634 : n62761;
  assign n62763 = pi16 ? n32 : n62762;
  assign n62764 = pi17 ? n44634 : n62253;
  assign n62765 = pi16 ? n32 : n62764;
  assign n62766 = pi15 ? n62763 : n62765;
  assign n62767 = pi14 ? n62755 : n62766;
  assign n62768 = pi13 ? n62741 : n62767;
  assign n62769 = pi21 ? n40917 : n40957;
  assign n62770 = pi22 ? n55502 : n20563;
  assign n62771 = pi21 ? n31877 : n62770;
  assign n62772 = pi20 ? n62769 : n62771;
  assign n62773 = pi19 ? n62772 : n50863;
  assign n62774 = pi20 ? n37308 : n61304;
  assign n62775 = pi19 ? n62774 : n62274;
  assign n62776 = pi18 ? n62773 : n62775;
  assign n62777 = pi17 ? n45739 : n62776;
  assign n62778 = pi16 ? n32 : n62777;
  assign n62779 = pi21 ? n20563 : n58594;
  assign n62780 = pi20 ? n40961 : n62779;
  assign n62781 = pi19 ? n62780 : n20563;
  assign n62782 = pi22 ? n34132 : n21502;
  assign n62783 = pi21 ? n62284 : n62782;
  assign n62784 = pi20 ? n62783 : n32;
  assign n62785 = pi19 ? n62282 : n62784;
  assign n62786 = pi18 ? n62781 : n62785;
  assign n62787 = pi17 ? n45739 : n62786;
  assign n62788 = pi16 ? n32 : n62787;
  assign n62789 = pi15 ? n62778 : n62788;
  assign n62790 = pi17 ? n44652 : n62297;
  assign n62791 = pi16 ? n32 : n62790;
  assign n62792 = pi22 ? n36781 : n55766;
  assign n62793 = pi21 ? n62792 : n55560;
  assign n62794 = pi20 ? n62793 : n32;
  assign n62795 = pi19 ? n56540 : n62794;
  assign n62796 = pi18 ? n20563 : n62795;
  assign n62797 = pi17 ? n44652 : n62796;
  assign n62798 = pi16 ? n32 : n62797;
  assign n62799 = pi15 ? n62791 : n62798;
  assign n62800 = pi14 ? n62789 : n62799;
  assign n62801 = pi17 ? n44643 : n62311;
  assign n62802 = pi16 ? n32 : n62801;
  assign n62803 = pi23 ? n14626 : n685;
  assign n62804 = pi22 ? n36781 : n62803;
  assign n62805 = pi21 ? n62804 : n37639;
  assign n62806 = pi20 ? n62805 : n32;
  assign n62807 = pi19 ? n61354 : n62806;
  assign n62808 = pi18 ? n20563 : n62807;
  assign n62809 = pi17 ? n44643 : n62808;
  assign n62810 = pi16 ? n32 : n62809;
  assign n62811 = pi15 ? n62802 : n62810;
  assign n62812 = pi22 ? n36798 : n1475;
  assign n62813 = pi21 ? n62812 : n1009;
  assign n62814 = pi20 ? n62813 : n32;
  assign n62815 = pi19 ? n62324 : n62814;
  assign n62816 = pi18 ? n20563 : n62815;
  assign n62817 = pi17 ? n44643 : n62816;
  assign n62818 = pi16 ? n32 : n62817;
  assign n62819 = pi22 ? n53450 : n36798;
  assign n62820 = pi21 ? n20563 : n62819;
  assign n62821 = pi20 ? n20563 : n62820;
  assign n62822 = pi21 ? n59691 : n20952;
  assign n62823 = pi20 ? n62822 : n32;
  assign n62824 = pi19 ? n62821 : n62823;
  assign n62825 = pi18 ? n20563 : n62824;
  assign n62826 = pi17 ? n44652 : n62825;
  assign n62827 = pi16 ? n32 : n62826;
  assign n62828 = pi15 ? n62818 : n62827;
  assign n62829 = pi14 ? n62811 : n62828;
  assign n62830 = pi13 ? n62800 : n62829;
  assign n62831 = pi12 ? n62768 : n62830;
  assign n62832 = pi24 ? n33792 : n335;
  assign n62833 = pi23 ? n33792 : n62832;
  assign n62834 = pi22 ? n62833 : n36798;
  assign n62835 = pi21 ? n20563 : n62834;
  assign n62836 = pi20 ? n20563 : n62835;
  assign n62837 = pi22 ? n14626 : n56665;
  assign n62838 = pi21 ? n62837 : n32;
  assign n62839 = pi20 ? n62838 : n32;
  assign n62840 = pi19 ? n62836 : n62839;
  assign n62841 = pi18 ? n20563 : n62840;
  assign n62842 = pi17 ? n44652 : n62841;
  assign n62843 = pi16 ? n32 : n62842;
  assign n62844 = pi19 ? n32 : n60024;
  assign n62845 = pi18 ? n32 : n62844;
  assign n62846 = pi22 ? n36659 : n62361;
  assign n62847 = pi21 ? n36489 : n62846;
  assign n62848 = pi20 ? n20563 : n62847;
  assign n62849 = pi22 ? n51564 : n56665;
  assign n62850 = pi21 ? n62849 : n32;
  assign n62851 = pi20 ? n62850 : n32;
  assign n62852 = pi19 ? n62848 : n62851;
  assign n62853 = pi18 ? n62359 : n62852;
  assign n62854 = pi17 ? n62845 : n62853;
  assign n62855 = pi16 ? n32 : n62854;
  assign n62856 = pi15 ? n62843 : n62855;
  assign n62857 = pi21 ? n60421 : n32;
  assign n62858 = pi20 ? n62857 : n32;
  assign n62859 = pi19 ? n62380 : n62858;
  assign n62860 = pi18 ? n30868 : n62859;
  assign n62861 = pi17 ? n51290 : n62860;
  assign n62862 = pi16 ? n32 : n62861;
  assign n62863 = pi18 ? n32 : n46169;
  assign n62864 = pi17 ? n62863 : n62394;
  assign n62865 = pi16 ? n32 : n62864;
  assign n62866 = pi15 ? n62862 : n62865;
  assign n62867 = pi14 ? n62856 : n62866;
  assign n62868 = pi17 ? n62863 : n62403;
  assign n62869 = pi16 ? n32 : n62868;
  assign n62870 = pi18 ? n32 : n46063;
  assign n62871 = pi23 ? n55783 : n13481;
  assign n62872 = pi22 ? n36798 : n62871;
  assign n62873 = pi21 ? n51313 : n62872;
  assign n62874 = pi20 ? n30868 : n62873;
  assign n62875 = pi19 ? n62874 : n57717;
  assign n62876 = pi18 ? n30868 : n62875;
  assign n62877 = pi17 ? n62870 : n62876;
  assign n62878 = pi16 ? n32 : n62877;
  assign n62879 = pi15 ? n62869 : n62878;
  assign n62880 = pi23 ? n43198 : n316;
  assign n62881 = pi22 ? n43198 : n62880;
  assign n62882 = pi21 ? n51313 : n62881;
  assign n62883 = pi20 ? n30868 : n62882;
  assign n62884 = pi19 ? n62883 : n57717;
  assign n62885 = pi18 ? n30868 : n62884;
  assign n62886 = pi17 ? n62870 : n62885;
  assign n62887 = pi16 ? n32 : n62886;
  assign n62888 = pi23 ? n60075 : n13481;
  assign n62889 = pi22 ? n43198 : n62888;
  assign n62890 = pi21 ? n36798 : n62889;
  assign n62891 = pi20 ? n30868 : n62890;
  assign n62892 = pi19 ? n62891 : n35482;
  assign n62893 = pi18 ? n30868 : n62892;
  assign n62894 = pi17 ? n62870 : n62893;
  assign n62895 = pi16 ? n32 : n62894;
  assign n62896 = pi15 ? n62887 : n62895;
  assign n62897 = pi14 ? n62879 : n62896;
  assign n62898 = pi13 ? n62867 : n62897;
  assign n62899 = pi22 ? n55641 : n54563;
  assign n62900 = pi21 ? n43198 : n62899;
  assign n62901 = pi20 ? n30868 : n62900;
  assign n62902 = pi19 ? n62901 : n32;
  assign n62903 = pi18 ? n30868 : n62902;
  assign n62904 = pi17 ? n62870 : n62903;
  assign n62905 = pi16 ? n32 : n62904;
  assign n62906 = pi19 ? n32 : n54445;
  assign n62907 = pi18 ? n32 : n62906;
  assign n62908 = pi22 ? n62803 : n58452;
  assign n62909 = pi21 ? n43198 : n62908;
  assign n62910 = pi20 ? n33792 : n62909;
  assign n62911 = pi19 ? n62910 : n32;
  assign n62912 = pi18 ? n33792 : n62911;
  assign n62913 = pi17 ? n62907 : n62912;
  assign n62914 = pi16 ? n32 : n62913;
  assign n62915 = pi15 ? n62905 : n62914;
  assign n62916 = pi18 ? n32 : n46279;
  assign n62917 = pi22 ? n43198 : n36801;
  assign n62918 = pi21 ? n50795 : n62917;
  assign n62919 = pi20 ? n62918 : n54655;
  assign n62920 = pi19 ? n62458 : n62919;
  assign n62921 = pi18 ? n62920 : n62464;
  assign n62922 = pi17 ? n62916 : n62921;
  assign n62923 = pi16 ? n32 : n62922;
  assign n62924 = pi17 ? n62916 : n62478;
  assign n62925 = pi16 ? n32 : n62924;
  assign n62926 = pi15 ? n62923 : n62925;
  assign n62927 = pi14 ? n62915 : n62926;
  assign n62928 = pi17 ? n32 : n62491;
  assign n62929 = pi16 ? n32 : n62928;
  assign n62930 = pi17 ? n32 : n62497;
  assign n62931 = pi16 ? n32 : n62930;
  assign n62932 = pi15 ? n62929 : n62931;
  assign n62933 = pi17 ? n32 : n62504;
  assign n62934 = pi16 ? n32 : n62933;
  assign n62935 = pi17 ? n32 : n62519;
  assign n62936 = pi16 ? n32 : n62935;
  assign n62937 = pi15 ? n62934 : n62936;
  assign n62938 = pi14 ? n62932 : n62937;
  assign n62939 = pi13 ? n62927 : n62938;
  assign n62940 = pi12 ? n62898 : n62939;
  assign n62941 = pi11 ? n62831 : n62940;
  assign n62942 = pi10 ? n62719 : n62941;
  assign n62943 = pi09 ? n62546 : n62942;
  assign n62944 = pi08 ? n62528 : n62943;
  assign n62945 = pi07 ? n61954 : n62944;
  assign n62946 = pi06 ? n60965 : n62945;
  assign n62947 = pi05 ? n59202 : n62946;
  assign n62948 = pi20 ? n20563 : n12225;
  assign n62949 = pi19 ? n20563 : n62948;
  assign n62950 = pi18 ? n42644 : n62949;
  assign n62951 = pi17 ? n32 : n62950;
  assign n62952 = pi16 ? n32 : n62951;
  assign n62953 = pi15 ? n32 : n62952;
  assign n62954 = pi20 ? n20563 : n61008;
  assign n62955 = pi19 ? n20563 : n62954;
  assign n62956 = pi18 ? n42654 : n62955;
  assign n62957 = pi17 ? n32 : n62956;
  assign n62958 = pi16 ? n32 : n62957;
  assign n62959 = pi18 ? n43261 : n62955;
  assign n62960 = pi17 ? n32 : n62959;
  assign n62961 = pi16 ? n32 : n62960;
  assign n62962 = pi15 ? n62958 : n62961;
  assign n62963 = pi14 ? n62953 : n62962;
  assign n62964 = pi13 ? n32 : n62963;
  assign n62965 = pi12 ? n32 : n62964;
  assign n62966 = pi11 ? n32 : n62965;
  assign n62967 = pi10 ? n32 : n62966;
  assign n62968 = pi18 ? n48120 : n62955;
  assign n62969 = pi17 ? n32 : n62968;
  assign n62970 = pi16 ? n32 : n62969;
  assign n62971 = pi18 ? n47592 : n62955;
  assign n62972 = pi17 ? n32 : n62971;
  assign n62973 = pi16 ? n32 : n62972;
  assign n62974 = pi15 ? n62970 : n62973;
  assign n62975 = pi20 ? n20563 : n1619;
  assign n62976 = pi19 ? n20563 : n62975;
  assign n62977 = pi18 ? n47592 : n62976;
  assign n62978 = pi17 ? n32 : n62977;
  assign n62979 = pi16 ? n32 : n62978;
  assign n62980 = pi18 ? n42206 : n62976;
  assign n62981 = pi17 ? n32 : n62980;
  assign n62982 = pi16 ? n32 : n62981;
  assign n62983 = pi15 ? n62979 : n62982;
  assign n62984 = pi14 ? n62974 : n62983;
  assign n62985 = pi18 ? n41630 : n62976;
  assign n62986 = pi17 ? n32 : n62985;
  assign n62987 = pi16 ? n32 : n62986;
  assign n62988 = pi18 ? n41181 : n62976;
  assign n62989 = pi17 ? n32 : n62988;
  assign n62990 = pi16 ? n32 : n62989;
  assign n62991 = pi18 ? n42239 : n62976;
  assign n62992 = pi17 ? n32 : n62991;
  assign n62993 = pi16 ? n32 : n62992;
  assign n62994 = pi15 ? n62990 : n62993;
  assign n62995 = pi14 ? n62987 : n62994;
  assign n62996 = pi13 ? n62984 : n62995;
  assign n62997 = pi18 ? n47056 : n62955;
  assign n62998 = pi17 ? n32 : n62997;
  assign n62999 = pi16 ? n32 : n62998;
  assign n63000 = pi14 ? n62993 : n62999;
  assign n63001 = pi18 ? n46446 : n59296;
  assign n63002 = pi17 ? n32 : n63001;
  assign n63003 = pi16 ? n32 : n63002;
  assign n63004 = pi18 ? n40497 : n59307;
  assign n63005 = pi17 ? n32 : n63004;
  assign n63006 = pi16 ? n32 : n63005;
  assign n63007 = pi15 ? n63003 : n63006;
  assign n63008 = pi24 ? n14626 : n32;
  assign n63009 = pi23 ? n63008 : n32;
  assign n63010 = pi22 ? n233 : n63009;
  assign n63011 = pi21 ? n59304 : n63010;
  assign n63012 = pi20 ? n20563 : n63011;
  assign n63013 = pi19 ? n20563 : n63012;
  assign n63014 = pi18 ? n41682 : n63013;
  assign n63015 = pi17 ? n32 : n63014;
  assign n63016 = pi16 ? n32 : n63015;
  assign n63017 = pi20 ? n53343 : n61651;
  assign n63018 = pi19 ? n20563 : n63017;
  assign n63019 = pi18 ? n41682 : n63018;
  assign n63020 = pi17 ? n32 : n63019;
  assign n63021 = pi16 ? n32 : n63020;
  assign n63022 = pi15 ? n63016 : n63021;
  assign n63023 = pi14 ? n63007 : n63022;
  assign n63024 = pi13 ? n63000 : n63023;
  assign n63025 = pi12 ? n62996 : n63024;
  assign n63026 = pi22 ? n62629 : n51564;
  assign n63027 = pi21 ? n63026 : n60421;
  assign n63028 = pi20 ? n53356 : n63027;
  assign n63029 = pi19 ? n20563 : n63028;
  assign n63030 = pi18 ? n41682 : n63029;
  assign n63031 = pi17 ? n32 : n63030;
  assign n63032 = pi16 ? n32 : n63031;
  assign n63033 = pi20 ? n53356 : n62640;
  assign n63034 = pi19 ? n20563 : n63033;
  assign n63035 = pi18 ? n40510 : n63034;
  assign n63036 = pi17 ? n32 : n63035;
  assign n63037 = pi16 ? n32 : n63036;
  assign n63038 = pi15 ? n63032 : n63037;
  assign n63039 = pi20 ? n53367 : n62648;
  assign n63040 = pi19 ? n20563 : n63039;
  assign n63041 = pi18 ? n40510 : n63040;
  assign n63042 = pi17 ? n32 : n63041;
  assign n63043 = pi16 ? n32 : n63042;
  assign n63044 = pi20 ? n53367 : n23203;
  assign n63045 = pi19 ? n20563 : n63044;
  assign n63046 = pi18 ? n39373 : n63045;
  assign n63047 = pi17 ? n32 : n63046;
  assign n63048 = pi16 ? n32 : n63047;
  assign n63049 = pi15 ? n63043 : n63048;
  assign n63050 = pi14 ? n63038 : n63049;
  assign n63051 = pi20 ? n53386 : n27076;
  assign n63052 = pi19 ? n20563 : n63051;
  assign n63053 = pi18 ? n38948 : n63052;
  assign n63054 = pi17 ? n32 : n63053;
  assign n63055 = pi16 ? n32 : n63054;
  assign n63056 = pi22 ? n20563 : n5011;
  assign n63057 = pi21 ? n20563 : n63056;
  assign n63058 = pi20 ? n63057 : n14723;
  assign n63059 = pi19 ? n20563 : n63058;
  assign n63060 = pi18 ? n38957 : n63059;
  assign n63061 = pi17 ? n32 : n63060;
  assign n63062 = pi16 ? n32 : n63061;
  assign n63063 = pi15 ? n63055 : n63062;
  assign n63064 = pi22 ? n20563 : n61132;
  assign n63065 = pi21 ? n20563 : n63064;
  assign n63066 = pi21 ? n316 : n37639;
  assign n63067 = pi20 ? n63065 : n63066;
  assign n63068 = pi19 ? n20563 : n63067;
  assign n63069 = pi18 ? n38957 : n63068;
  assign n63070 = pi17 ? n32 : n63069;
  assign n63071 = pi16 ? n32 : n63070;
  assign n63072 = pi22 ? n20563 : n61145;
  assign n63073 = pi21 ? n20563 : n63072;
  assign n63074 = pi20 ? n63073 : n1010;
  assign n63075 = pi19 ? n20563 : n63074;
  assign n63076 = pi18 ? n38957 : n63075;
  assign n63077 = pi17 ? n32 : n63076;
  assign n63078 = pi16 ? n32 : n63077;
  assign n63079 = pi15 ? n63071 : n63078;
  assign n63080 = pi14 ? n63063 : n63079;
  assign n63081 = pi13 ? n63050 : n63080;
  assign n63082 = pi18 ? n40045 : n62677;
  assign n63083 = pi17 ? n32 : n63082;
  assign n63084 = pi16 ? n32 : n63083;
  assign n63085 = pi20 ? n62129 : n17510;
  assign n63086 = pi19 ? n20563 : n63085;
  assign n63087 = pi18 ? n40045 : n63086;
  assign n63088 = pi17 ? n32 : n63087;
  assign n63089 = pi16 ? n32 : n63088;
  assign n63090 = pi15 ? n63084 : n63089;
  assign n63091 = pi23 ? n30868 : n233;
  assign n63092 = pi22 ? n20563 : n63091;
  assign n63093 = pi21 ? n45016 : n63092;
  assign n63094 = pi20 ? n63093 : n19727;
  assign n63095 = pi19 ? n20563 : n63094;
  assign n63096 = pi18 ? n40045 : n63095;
  assign n63097 = pi17 ? n32 : n63096;
  assign n63098 = pi16 ? n32 : n63097;
  assign n63099 = pi23 ? n30868 : n14626;
  assign n63100 = pi22 ? n30868 : n63099;
  assign n63101 = pi21 ? n20563 : n63100;
  assign n63102 = pi20 ? n63101 : n10326;
  assign n63103 = pi19 ? n20563 : n63102;
  assign n63104 = pi18 ? n40045 : n63103;
  assign n63105 = pi17 ? n32 : n63104;
  assign n63106 = pi16 ? n32 : n63105;
  assign n63107 = pi15 ? n63098 : n63106;
  assign n63108 = pi14 ? n63090 : n63107;
  assign n63109 = pi22 ? n139 : n59423;
  assign n63110 = pi21 ? n40986 : n63109;
  assign n63111 = pi20 ? n63110 : n58471;
  assign n63112 = pi19 ? n20563 : n63111;
  assign n63113 = pi18 ? n40550 : n63112;
  assign n63114 = pi17 ? n32 : n63113;
  assign n63115 = pi16 ? n32 : n63114;
  assign n63116 = pi21 ? n36489 : n61192;
  assign n63117 = pi20 ? n63116 : n54547;
  assign n63118 = pi19 ? n20563 : n63117;
  assign n63119 = pi18 ? n40550 : n63118;
  assign n63120 = pi17 ? n32 : n63119;
  assign n63121 = pi16 ? n32 : n63120;
  assign n63122 = pi15 ? n63115 : n63121;
  assign n63123 = pi22 ? n335 : n62389;
  assign n63124 = pi21 ? n45016 : n63123;
  assign n63125 = pi20 ? n63124 : n56130;
  assign n63126 = pi19 ? n40792 : n63125;
  assign n63127 = pi18 ? n40550 : n63126;
  assign n63128 = pi17 ? n32 : n63127;
  assign n63129 = pi16 ? n32 : n63128;
  assign n63130 = pi22 ? n36659 : n61484;
  assign n63131 = pi21 ? n39801 : n63130;
  assign n63132 = pi20 ? n63131 : n56130;
  assign n63133 = pi19 ? n40792 : n63132;
  assign n63134 = pi18 ? n40550 : n63133;
  assign n63135 = pi17 ? n32 : n63134;
  assign n63136 = pi16 ? n32 : n63135;
  assign n63137 = pi15 ? n63129 : n63136;
  assign n63138 = pi14 ? n63122 : n63137;
  assign n63139 = pi13 ? n63108 : n63138;
  assign n63140 = pi12 ? n63081 : n63139;
  assign n63141 = pi11 ? n63025 : n63140;
  assign n63142 = pi21 ? n40249 : n57671;
  assign n63143 = pi20 ? n63142 : n4116;
  assign n63144 = pi19 ? n59458 : n63143;
  assign n63145 = pi18 ? n40550 : n63144;
  assign n63146 = pi17 ? n32 : n63145;
  assign n63147 = pi16 ? n32 : n63146;
  assign n63148 = pi22 ? n33792 : n57085;
  assign n63149 = pi21 ? n63148 : n58999;
  assign n63150 = pi20 ? n63149 : n10011;
  assign n63151 = pi19 ? n59458 : n63150;
  assign n63152 = pi18 ? n40550 : n63151;
  assign n63153 = pi17 ? n32 : n63152;
  assign n63154 = pi16 ? n32 : n63153;
  assign n63155 = pi15 ? n63147 : n63154;
  assign n63156 = pi22 ? n36659 : n42109;
  assign n63157 = pi21 ? n63156 : n59681;
  assign n63158 = pi20 ? n63157 : n57716;
  assign n63159 = pi19 ? n50091 : n63158;
  assign n63160 = pi18 ? n40550 : n63159;
  assign n63161 = pi17 ? n32 : n63160;
  assign n63162 = pi16 ? n32 : n63161;
  assign n63163 = pi21 ? n62743 : n57733;
  assign n63164 = pi20 ? n63163 : n37640;
  assign n63165 = pi19 ? n20563 : n63164;
  assign n63166 = pi18 ? n45413 : n63165;
  assign n63167 = pi17 ? n32 : n63166;
  assign n63168 = pi16 ? n32 : n63167;
  assign n63169 = pi15 ? n63162 : n63168;
  assign n63170 = pi14 ? n63155 : n63169;
  assign n63171 = pi20 ? n31263 : n40791;
  assign n63172 = pi19 ? n63171 : n20563;
  assign n63173 = pi21 ? n60441 : n59691;
  assign n63174 = pi20 ? n63173 : n20953;
  assign n63175 = pi19 ? n40792 : n63174;
  assign n63176 = pi18 ? n63172 : n63175;
  assign n63177 = pi17 ? n32 : n63176;
  assign n63178 = pi16 ? n32 : n63177;
  assign n63179 = pi22 ? n30154 : n40386;
  assign n63180 = pi21 ? n63179 : n30868;
  assign n63181 = pi20 ? n63180 : n40791;
  assign n63182 = pi19 ? n63181 : n50101;
  assign n63183 = pi21 ? n56645 : n57746;
  assign n63184 = pi20 ? n63183 : n20953;
  assign n63185 = pi19 ? n40792 : n63184;
  assign n63186 = pi18 ? n63182 : n63185;
  assign n63187 = pi17 ? n32 : n63186;
  assign n63188 = pi16 ? n32 : n63187;
  assign n63189 = pi15 ? n63178 : n63188;
  assign n63190 = pi20 ? n20563 : n61280;
  assign n63191 = pi19 ? n43253 : n63190;
  assign n63192 = pi21 ? n36489 : n33792;
  assign n63193 = pi20 ? n20563 : n63192;
  assign n63194 = pi24 ? n36659 : n363;
  assign n63195 = pi23 ? n36659 : n63194;
  assign n63196 = pi22 ? n30868 : n63195;
  assign n63197 = pi22 ? n14626 : n2192;
  assign n63198 = pi21 ? n63196 : n63197;
  assign n63199 = pi20 ? n63198 : n32;
  assign n63200 = pi19 ? n63193 : n63199;
  assign n63201 = pi18 ? n63191 : n63200;
  assign n63202 = pi17 ? n32 : n63201;
  assign n63203 = pi16 ? n32 : n63202;
  assign n63204 = pi20 ? n20563 : n51280;
  assign n63205 = pi19 ? n43253 : n63204;
  assign n63206 = pi21 ? n29133 : n33792;
  assign n63207 = pi20 ? n20563 : n63206;
  assign n63208 = pi22 ? n33792 : n57501;
  assign n63209 = pi21 ? n63208 : n59621;
  assign n63210 = pi20 ? n63209 : n32;
  assign n63211 = pi19 ? n63207 : n63210;
  assign n63212 = pi18 ? n63205 : n63211;
  assign n63213 = pi17 ? n32 : n63212;
  assign n63214 = pi16 ? n32 : n63213;
  assign n63215 = pi15 ? n63203 : n63214;
  assign n63216 = pi14 ? n63189 : n63215;
  assign n63217 = pi13 ? n63170 : n63216;
  assign n63218 = pi20 ? n31313 : n37308;
  assign n63219 = pi19 ? n63218 : n20563;
  assign n63220 = pi21 ? n29133 : n36659;
  assign n63221 = pi20 ? n20563 : n63220;
  assign n63222 = pi21 ? n53463 : n62285;
  assign n63223 = pi20 ? n63222 : n32;
  assign n63224 = pi19 ? n63221 : n63223;
  assign n63225 = pi18 ? n63219 : n63224;
  assign n63226 = pi17 ? n32 : n63225;
  assign n63227 = pi16 ? n32 : n63226;
  assign n63228 = pi20 ? n53428 : n20563;
  assign n63229 = pi19 ? n63228 : n20563;
  assign n63230 = pi23 ? n58566 : n51564;
  assign n63231 = pi22 ? n63230 : n21502;
  assign n63232 = pi21 ? n50795 : n63231;
  assign n63233 = pi20 ? n63232 : n32;
  assign n63234 = pi19 ? n56631 : n63233;
  assign n63235 = pi18 ? n63229 : n63234;
  assign n63236 = pi17 ? n32 : n63235;
  assign n63237 = pi16 ? n32 : n63236;
  assign n63238 = pi15 ? n63227 : n63237;
  assign n63239 = pi20 ? n20563 : n57630;
  assign n63240 = pi22 ? n57674 : n32;
  assign n63241 = pi21 ? n57774 : n63240;
  assign n63242 = pi20 ? n63241 : n32;
  assign n63243 = pi19 ? n63239 : n63242;
  assign n63244 = pi18 ? n20563 : n63243;
  assign n63245 = pi17 ? n44634 : n63244;
  assign n63246 = pi16 ? n32 : n63245;
  assign n63247 = pi19 ? n56540 : n63242;
  assign n63248 = pi18 ? n20563 : n63247;
  assign n63249 = pi17 ? n44634 : n63248;
  assign n63250 = pi16 ? n32 : n63249;
  assign n63251 = pi15 ? n63246 : n63250;
  assign n63252 = pi14 ? n63238 : n63251;
  assign n63253 = pi22 ? n36781 : n51564;
  assign n63254 = pi21 ? n63253 : n928;
  assign n63255 = pi20 ? n63254 : n32;
  assign n63256 = pi19 ? n56540 : n63255;
  assign n63257 = pi18 ? n20563 : n63256;
  assign n63258 = pi17 ? n44634 : n63257;
  assign n63259 = pi16 ? n32 : n63258;
  assign n63260 = pi23 ? n20563 : n56976;
  assign n63261 = pi22 ? n63260 : n36798;
  assign n63262 = pi21 ? n20563 : n63261;
  assign n63263 = pi20 ? n20563 : n63262;
  assign n63264 = pi21 ? n59681 : n37639;
  assign n63265 = pi20 ? n63264 : n32;
  assign n63266 = pi19 ? n63263 : n63265;
  assign n63267 = pi18 ? n20563 : n63266;
  assign n63268 = pi17 ? n32 : n63267;
  assign n63269 = pi16 ? n32 : n63268;
  assign n63270 = pi15 ? n63259 : n63269;
  assign n63271 = pi22 ? n42106 : n36798;
  assign n63272 = pi21 ? n20563 : n63271;
  assign n63273 = pi20 ? n20563 : n63272;
  assign n63274 = pi21 ? n59774 : n20952;
  assign n63275 = pi20 ? n63274 : n32;
  assign n63276 = pi19 ? n63273 : n63275;
  assign n63277 = pi18 ? n20563 : n63276;
  assign n63278 = pi17 ? n32 : n63277;
  assign n63279 = pi16 ? n32 : n63278;
  assign n63280 = pi23 ? n335 : n55567;
  assign n63281 = pi22 ? n63280 : n36798;
  assign n63282 = pi21 ? n20563 : n63281;
  assign n63283 = pi20 ? n20563 : n63282;
  assign n63284 = pi21 ? n55606 : n20952;
  assign n63285 = pi20 ? n63284 : n32;
  assign n63286 = pi19 ? n63283 : n63285;
  assign n63287 = pi18 ? n20563 : n63286;
  assign n63288 = pi17 ? n46325 : n63287;
  assign n63289 = pi16 ? n32 : n63288;
  assign n63290 = pi15 ? n63279 : n63289;
  assign n63291 = pi14 ? n63270 : n63290;
  assign n63292 = pi13 ? n63252 : n63291;
  assign n63293 = pi12 ? n63217 : n63292;
  assign n63294 = pi23 ? n36659 : n62832;
  assign n63295 = pi22 ? n63294 : n233;
  assign n63296 = pi21 ? n36489 : n63295;
  assign n63297 = pi20 ? n20563 : n63296;
  assign n63298 = pi19 ? n63297 : n62839;
  assign n63299 = pi18 ? n20563 : n63298;
  assign n63300 = pi17 ? n46325 : n63299;
  assign n63301 = pi16 ? n32 : n63300;
  assign n63302 = pi19 ? n60503 : n59667;
  assign n63303 = pi22 ? n52421 : n51564;
  assign n63304 = pi21 ? n30868 : n63303;
  assign n63305 = pi20 ? n30868 : n63304;
  assign n63306 = pi24 ? n14626 : n51564;
  assign n63307 = pi23 ? n14626 : n63306;
  assign n63308 = pi22 ? n63307 : n56665;
  assign n63309 = pi21 ? n63308 : n32;
  assign n63310 = pi20 ? n63309 : n32;
  assign n63311 = pi19 ? n63305 : n63310;
  assign n63312 = pi18 ? n63302 : n63311;
  assign n63313 = pi17 ? n51824 : n63312;
  assign n63314 = pi16 ? n32 : n63313;
  assign n63315 = pi15 ? n63301 : n63314;
  assign n63316 = pi19 ? n60503 : n30868;
  assign n63317 = pi23 ? n36781 : n14626;
  assign n63318 = pi22 ? n38284 : n63317;
  assign n63319 = pi21 ? n36489 : n63318;
  assign n63320 = pi20 ? n30868 : n63319;
  assign n63321 = pi19 ? n63320 : n62858;
  assign n63322 = pi18 ? n63316 : n63321;
  assign n63323 = pi17 ? n51824 : n63322;
  assign n63324 = pi16 ? n32 : n63323;
  assign n63325 = pi20 ? n36489 : n30868;
  assign n63326 = pi19 ? n63325 : n30868;
  assign n63327 = pi22 ? n36659 : n30868;
  assign n63328 = pi23 ? n36798 : n51564;
  assign n63329 = pi22 ? n36798 : n63328;
  assign n63330 = pi21 ? n63327 : n63329;
  assign n63331 = pi20 ? n30868 : n63330;
  assign n63332 = pi19 ? n63331 : n60046;
  assign n63333 = pi18 ? n63326 : n63332;
  assign n63334 = pi17 ? n32 : n63333;
  assign n63335 = pi16 ? n32 : n63334;
  assign n63336 = pi15 ? n63324 : n63335;
  assign n63337 = pi14 ? n63315 : n63336;
  assign n63338 = pi20 ? n42005 : n43010;
  assign n63339 = pi19 ? n63338 : n30868;
  assign n63340 = pi21 ? n42146 : n57104;
  assign n63341 = pi20 ? n30868 : n63340;
  assign n63342 = pi19 ? n63341 : n60046;
  assign n63343 = pi18 ? n63339 : n63342;
  assign n63344 = pi17 ? n32 : n63343;
  assign n63345 = pi16 ? n32 : n63344;
  assign n63346 = pi21 ? n36781 : n57112;
  assign n63347 = pi20 ? n30868 : n63346;
  assign n63348 = pi19 ? n63347 : n57717;
  assign n63349 = pi18 ? n63339 : n63348;
  assign n63350 = pi17 ? n32 : n63349;
  assign n63351 = pi16 ? n32 : n63350;
  assign n63352 = pi15 ? n63345 : n63351;
  assign n63353 = pi21 ? n30116 : n30868;
  assign n63354 = pi20 ? n63353 : n30868;
  assign n63355 = pi19 ? n63354 : n30868;
  assign n63356 = pi22 ? n55622 : n56622;
  assign n63357 = pi21 ? n38901 : n63356;
  assign n63358 = pi20 ? n30868 : n63357;
  assign n63359 = pi19 ? n63358 : n35482;
  assign n63360 = pi18 ? n63355 : n63359;
  assign n63361 = pi17 ? n32 : n63360;
  assign n63362 = pi16 ? n32 : n63361;
  assign n63363 = pi21 ? n30868 : n59524;
  assign n63364 = pi21 ? n36798 : n62899;
  assign n63365 = pi20 ? n63363 : n63364;
  assign n63366 = pi19 ? n63365 : n32;
  assign n63367 = pi18 ? n46701 : n63366;
  assign n63368 = pi17 ? n32 : n63367;
  assign n63369 = pi16 ? n32 : n63368;
  assign n63370 = pi15 ? n63362 : n63369;
  assign n63371 = pi14 ? n63352 : n63370;
  assign n63372 = pi13 ? n63337 : n63371;
  assign n63373 = pi21 ? n46166 : n33792;
  assign n63374 = pi20 ? n63373 : n33792;
  assign n63375 = pi19 ? n63374 : n33792;
  assign n63376 = pi22 ? n56607 : n57647;
  assign n63377 = pi21 ? n47396 : n63376;
  assign n63378 = pi20 ? n33792 : n63377;
  assign n63379 = pi19 ? n63378 : n32;
  assign n63380 = pi18 ? n63375 : n63379;
  assign n63381 = pi17 ? n32 : n63380;
  assign n63382 = pi16 ? n32 : n63381;
  assign n63383 = pi20 ? n45518 : n33792;
  assign n63384 = pi19 ? n63383 : n33792;
  assign n63385 = pi21 ? n36798 : n59648;
  assign n63386 = pi20 ? n61480 : n63385;
  assign n63387 = pi19 ? n63386 : n32;
  assign n63388 = pi18 ? n63384 : n63387;
  assign n63389 = pi17 ? n32 : n63388;
  assign n63390 = pi16 ? n32 : n63389;
  assign n63391 = pi15 ? n63382 : n63390;
  assign n63392 = pi21 ? n46727 : n47396;
  assign n63393 = pi20 ? n63392 : n54009;
  assign n63394 = pi19 ? n63393 : n43198;
  assign n63395 = pi21 ? n47397 : n59648;
  assign n63396 = pi20 ? n43198 : n63395;
  assign n63397 = pi19 ? n63396 : n32;
  assign n63398 = pi18 ? n63394 : n63397;
  assign n63399 = pi17 ? n32 : n63398;
  assign n63400 = pi16 ? n32 : n63399;
  assign n63401 = pi22 ? n37276 : n36798;
  assign n63402 = pi21 ? n48856 : n63401;
  assign n63403 = pi20 ? n63402 : n43198;
  assign n63404 = pi19 ? n63403 : n43198;
  assign n63405 = pi21 ? n58777 : n55560;
  assign n63406 = pi20 ? n43198 : n63405;
  assign n63407 = pi19 ? n63406 : n32;
  assign n63408 = pi18 ? n63404 : n63407;
  assign n63409 = pi17 ? n32 : n63408;
  assign n63410 = pi16 ? n32 : n63409;
  assign n63411 = pi15 ? n63400 : n63410;
  assign n63412 = pi14 ? n63391 : n63411;
  assign n63413 = pi21 ? n48856 : n58755;
  assign n63414 = pi20 ? n63413 : n43198;
  assign n63415 = pi19 ? n63414 : n43198;
  assign n63416 = pi20 ? n43198 : n60250;
  assign n63417 = pi19 ? n63416 : n32;
  assign n63418 = pi18 ? n63415 : n63417;
  assign n63419 = pi17 ? n32 : n63418;
  assign n63420 = pi16 ? n32 : n63419;
  assign n63421 = pi20 ? n59698 : n43198;
  assign n63422 = pi19 ? n63421 : n43198;
  assign n63423 = pi22 ? n13481 : n51564;
  assign n63424 = pi21 ? n63423 : n1009;
  assign n63425 = pi20 ? n59703 : n63424;
  assign n63426 = pi19 ? n63425 : n32;
  assign n63427 = pi18 ? n63422 : n63426;
  assign n63428 = pi17 ? n32 : n63427;
  assign n63429 = pi16 ? n32 : n63428;
  assign n63430 = pi15 ? n63420 : n63429;
  assign n63431 = pi24 ? n32 : n14626;
  assign n63432 = pi23 ? n32 : n63431;
  assign n63433 = pi22 ? n32 : n63432;
  assign n63434 = pi22 ? n53550 : n14626;
  assign n63435 = pi21 ? n63433 : n63434;
  assign n63436 = pi20 ? n63435 : n14626;
  assign n63437 = pi19 ? n63436 : n14626;
  assign n63438 = pi20 ? n14626 : n59604;
  assign n63439 = pi19 ? n63438 : n32;
  assign n63440 = pi18 ? n63437 : n63439;
  assign n63441 = pi17 ? n32 : n63440;
  assign n63442 = pi16 ? n32 : n63441;
  assign n63443 = pi22 ? n14626 : n36798;
  assign n63444 = pi21 ? n63443 : n36798;
  assign n63445 = pi20 ? n63444 : n36798;
  assign n63446 = pi19 ? n52381 : n63445;
  assign n63447 = pi20 ? n36798 : n59604;
  assign n63448 = pi19 ? n63447 : n32;
  assign n63449 = pi18 ? n63446 : n63448;
  assign n63450 = pi17 ? n32 : n63449;
  assign n63451 = pi16 ? n32 : n63450;
  assign n63452 = pi15 ? n63442 : n63451;
  assign n63453 = pi14 ? n63430 : n63452;
  assign n63454 = pi13 ? n63412 : n63453;
  assign n63455 = pi12 ? n63372 : n63454;
  assign n63456 = pi11 ? n63293 : n63455;
  assign n63457 = pi10 ? n63141 : n63456;
  assign n63458 = pi09 ? n62967 : n63457;
  assign n63459 = pi18 ? n43226 : n62949;
  assign n63460 = pi17 ? n32 : n63459;
  assign n63461 = pi16 ? n32 : n63460;
  assign n63462 = pi15 ? n32 : n63461;
  assign n63463 = pi18 ? n43247 : n62955;
  assign n63464 = pi17 ? n32 : n63463;
  assign n63465 = pi16 ? n32 : n63464;
  assign n63466 = pi18 ? n42680 : n62955;
  assign n63467 = pi17 ? n32 : n63466;
  assign n63468 = pi16 ? n32 : n63467;
  assign n63469 = pi15 ? n63465 : n63468;
  assign n63470 = pi14 ? n63462 : n63469;
  assign n63471 = pi13 ? n32 : n63470;
  assign n63472 = pi12 ? n32 : n63471;
  assign n63473 = pi11 ? n32 : n63472;
  assign n63474 = pi10 ? n32 : n63473;
  assign n63475 = pi18 ? n42193 : n62955;
  assign n63476 = pi17 ? n32 : n63475;
  assign n63477 = pi16 ? n32 : n63476;
  assign n63478 = pi18 ? n43254 : n62955;
  assign n63479 = pi17 ? n32 : n63478;
  assign n63480 = pi16 ? n32 : n63479;
  assign n63481 = pi15 ? n63477 : n63480;
  assign n63482 = pi18 ? n43254 : n62976;
  assign n63483 = pi17 ? n32 : n63482;
  assign n63484 = pi16 ? n32 : n63483;
  assign n63485 = pi18 ? n42200 : n62976;
  assign n63486 = pi17 ? n32 : n63485;
  assign n63487 = pi16 ? n32 : n63486;
  assign n63488 = pi15 ? n63484 : n63487;
  assign n63489 = pi14 ? n63481 : n63488;
  assign n63490 = pi18 ? n43261 : n62976;
  assign n63491 = pi17 ? n32 : n63490;
  assign n63492 = pi16 ? n32 : n63491;
  assign n63493 = pi15 ? n63487 : n63492;
  assign n63494 = pi18 ? n40485 : n62976;
  assign n63495 = pi17 ? n32 : n63494;
  assign n63496 = pi16 ? n32 : n63495;
  assign n63497 = pi18 ? n41157 : n62976;
  assign n63498 = pi17 ? n32 : n63497;
  assign n63499 = pi16 ? n32 : n63498;
  assign n63500 = pi15 ? n63496 : n63499;
  assign n63501 = pi14 ? n63493 : n63500;
  assign n63502 = pi13 ? n63489 : n63501;
  assign n63503 = pi18 ? n41168 : n62955;
  assign n63504 = pi17 ? n32 : n63503;
  assign n63505 = pi16 ? n32 : n63504;
  assign n63506 = pi14 ? n63499 : n63505;
  assign n63507 = pi18 ? n41168 : n59296;
  assign n63508 = pi17 ? n32 : n63507;
  assign n63509 = pi16 ? n32 : n63508;
  assign n63510 = pi18 ? n41181 : n59307;
  assign n63511 = pi17 ? n32 : n63510;
  assign n63512 = pi16 ? n32 : n63511;
  assign n63513 = pi15 ? n63509 : n63512;
  assign n63514 = pi18 ? n42239 : n63013;
  assign n63515 = pi17 ? n32 : n63514;
  assign n63516 = pi16 ? n32 : n63515;
  assign n63517 = pi24 ? n20563 : n685;
  assign n63518 = pi23 ? n63517 : n685;
  assign n63519 = pi22 ? n63518 : n685;
  assign n63520 = pi21 ? n63519 : n8486;
  assign n63521 = pi20 ? n53343 : n63520;
  assign n63522 = pi19 ? n20563 : n63521;
  assign n63523 = pi18 ? n42239 : n63522;
  assign n63524 = pi17 ? n32 : n63523;
  assign n63525 = pi16 ? n32 : n63524;
  assign n63526 = pi15 ? n63516 : n63525;
  assign n63527 = pi14 ? n63513 : n63526;
  assign n63528 = pi13 ? n63506 : n63527;
  assign n63529 = pi12 ? n63502 : n63528;
  assign n63530 = pi24 ? n30868 : n685;
  assign n63531 = pi23 ? n63530 : n685;
  assign n63532 = pi22 ? n63531 : n51564;
  assign n63533 = pi21 ? n63532 : n60421;
  assign n63534 = pi20 ? n53356 : n63533;
  assign n63535 = pi19 ? n20563 : n63534;
  assign n63536 = pi18 ? n42239 : n63535;
  assign n63537 = pi17 ? n32 : n63536;
  assign n63538 = pi16 ? n32 : n63537;
  assign n63539 = pi18 ? n47056 : n63034;
  assign n63540 = pi17 ? n32 : n63539;
  assign n63541 = pi16 ? n32 : n63540;
  assign n63542 = pi15 ? n63538 : n63541;
  assign n63543 = pi23 ? n32126 : n13481;
  assign n63544 = pi22 ? n63543 : n13481;
  assign n63545 = pi21 ? n63544 : n55560;
  assign n63546 = pi20 ? n53367 : n63545;
  assign n63547 = pi19 ? n20563 : n63546;
  assign n63548 = pi18 ? n47056 : n63547;
  assign n63549 = pi17 ? n32 : n63548;
  assign n63550 = pi16 ? n32 : n63549;
  assign n63551 = pi18 ? n46446 : n63045;
  assign n63552 = pi17 ? n32 : n63551;
  assign n63553 = pi16 ? n32 : n63552;
  assign n63554 = pi15 ? n63550 : n63553;
  assign n63555 = pi14 ? n63542 : n63554;
  assign n63556 = pi18 ? n46446 : n63052;
  assign n63557 = pi17 ? n32 : n63556;
  assign n63558 = pi16 ? n32 : n63557;
  assign n63559 = pi18 ? n40497 : n63059;
  assign n63560 = pi17 ? n32 : n63559;
  assign n63561 = pi16 ? n32 : n63560;
  assign n63562 = pi15 ? n63558 : n63561;
  assign n63563 = pi18 ? n40497 : n63068;
  assign n63564 = pi17 ? n32 : n63563;
  assign n63565 = pi16 ? n32 : n63564;
  assign n63566 = pi18 ? n40497 : n63075;
  assign n63567 = pi17 ? n32 : n63566;
  assign n63568 = pi16 ? n32 : n63567;
  assign n63569 = pi15 ? n63565 : n63568;
  assign n63570 = pi14 ? n63562 : n63569;
  assign n63571 = pi13 ? n63555 : n63570;
  assign n63572 = pi18 ? n41682 : n62677;
  assign n63573 = pi17 ? n32 : n63572;
  assign n63574 = pi16 ? n32 : n63573;
  assign n63575 = pi18 ? n41682 : n63086;
  assign n63576 = pi17 ? n32 : n63575;
  assign n63577 = pi16 ? n32 : n63576;
  assign n63578 = pi15 ? n63574 : n63577;
  assign n63579 = pi18 ? n40510 : n63095;
  assign n63580 = pi17 ? n32 : n63579;
  assign n63581 = pi16 ? n32 : n63580;
  assign n63582 = pi18 ? n45366 : n63103;
  assign n63583 = pi17 ? n32 : n63582;
  assign n63584 = pi16 ? n32 : n63583;
  assign n63585 = pi15 ? n63581 : n63584;
  assign n63586 = pi14 ? n63578 : n63585;
  assign n63587 = pi18 ? n38948 : n63112;
  assign n63588 = pi17 ? n32 : n63587;
  assign n63589 = pi16 ? n32 : n63588;
  assign n63590 = pi20 ? n63116 : n4008;
  assign n63591 = pi19 ? n20563 : n63590;
  assign n63592 = pi18 ? n38948 : n63591;
  assign n63593 = pi17 ? n32 : n63592;
  assign n63594 = pi16 ? n32 : n63593;
  assign n63595 = pi15 ? n63589 : n63594;
  assign n63596 = pi18 ? n38948 : n63126;
  assign n63597 = pi17 ? n32 : n63596;
  assign n63598 = pi16 ? n32 : n63597;
  assign n63599 = pi20 ? n63131 : n61714;
  assign n63600 = pi19 ? n40792 : n63599;
  assign n63601 = pi18 ? n38948 : n63600;
  assign n63602 = pi17 ? n32 : n63601;
  assign n63603 = pi16 ? n32 : n63602;
  assign n63604 = pi15 ? n63598 : n63603;
  assign n63605 = pi14 ? n63595 : n63604;
  assign n63606 = pi13 ? n63586 : n63605;
  assign n63607 = pi12 ? n63571 : n63606;
  assign n63608 = pi11 ? n63529 : n63607;
  assign n63609 = pi18 ? n38948 : n63144;
  assign n63610 = pi17 ? n32 : n63609;
  assign n63611 = pi16 ? n32 : n63610;
  assign n63612 = pi22 ? n33792 : n39190;
  assign n63613 = pi21 ? n63612 : n58999;
  assign n63614 = pi20 ? n63613 : n10011;
  assign n63615 = pi19 ? n59458 : n63614;
  assign n63616 = pi18 ? n38948 : n63615;
  assign n63617 = pi17 ? n32 : n63616;
  assign n63618 = pi16 ? n32 : n63617;
  assign n63619 = pi15 ? n63611 : n63618;
  assign n63620 = pi18 ? n38948 : n63159;
  assign n63621 = pi17 ? n32 : n63620;
  assign n63622 = pi16 ? n32 : n63621;
  assign n63623 = pi23 ? n30868 : n335;
  assign n63624 = pi22 ? n20563 : n63623;
  assign n63625 = pi21 ? n63624 : n57733;
  assign n63626 = pi20 ? n63625 : n1822;
  assign n63627 = pi19 ? n20563 : n63626;
  assign n63628 = pi18 ? n40045 : n63627;
  assign n63629 = pi17 ? n32 : n63628;
  assign n63630 = pi16 ? n32 : n63629;
  assign n63631 = pi15 ? n63622 : n63630;
  assign n63632 = pi14 ? n63619 : n63631;
  assign n63633 = pi20 ? n38376 : n40791;
  assign n63634 = pi19 ? n63633 : n20563;
  assign n63635 = pi18 ? n63634 : n63175;
  assign n63636 = pi17 ? n32 : n63635;
  assign n63637 = pi16 ? n32 : n63636;
  assign n63638 = pi19 ? n60769 : n50101;
  assign n63639 = pi22 ? n30868 : n56065;
  assign n63640 = pi22 ? n14626 : n61712;
  assign n63641 = pi21 ? n63639 : n63640;
  assign n63642 = pi20 ? n63641 : n32;
  assign n63643 = pi19 ? n40792 : n63642;
  assign n63644 = pi18 ? n63638 : n63643;
  assign n63645 = pi17 ? n32 : n63644;
  assign n63646 = pi16 ? n32 : n63645;
  assign n63647 = pi15 ? n63637 : n63646;
  assign n63648 = pi19 ? n40044 : n63190;
  assign n63649 = pi23 ? n36659 : n56079;
  assign n63650 = pi22 ? n30868 : n63649;
  assign n63651 = pi21 ? n63650 : n63197;
  assign n63652 = pi20 ? n63651 : n32;
  assign n63653 = pi19 ? n63193 : n63652;
  assign n63654 = pi18 ? n63648 : n63653;
  assign n63655 = pi17 ? n32 : n63654;
  assign n63656 = pi16 ? n32 : n63655;
  assign n63657 = pi19 ? n40044 : n63204;
  assign n63658 = pi22 ? n33792 : n58044;
  assign n63659 = pi21 ? n63658 : n59621;
  assign n63660 = pi20 ? n63659 : n32;
  assign n63661 = pi19 ? n63207 : n63660;
  assign n63662 = pi18 ? n63657 : n63661;
  assign n63663 = pi17 ? n32 : n63662;
  assign n63664 = pi16 ? n32 : n63663;
  assign n63665 = pi15 ? n63656 : n63664;
  assign n63666 = pi14 ? n63647 : n63665;
  assign n63667 = pi13 ? n63632 : n63666;
  assign n63668 = pi20 ? n39395 : n37308;
  assign n63669 = pi19 ? n63668 : n20563;
  assign n63670 = pi18 ? n63669 : n63224;
  assign n63671 = pi17 ? n32 : n63670;
  assign n63672 = pi16 ? n32 : n63671;
  assign n63673 = pi20 ? n53943 : n20563;
  assign n63674 = pi19 ? n63673 : n20563;
  assign n63675 = pi22 ? n63230 : n32;
  assign n63676 = pi21 ? n50795 : n63675;
  assign n63677 = pi20 ? n63676 : n32;
  assign n63678 = pi19 ? n56631 : n63677;
  assign n63679 = pi18 ? n63674 : n63678;
  assign n63680 = pi17 ? n32 : n63679;
  assign n63681 = pi16 ? n32 : n63680;
  assign n63682 = pi15 ? n63672 : n63681;
  assign n63683 = pi18 ? n38316 : n63243;
  assign n63684 = pi17 ? n32 : n63683;
  assign n63685 = pi16 ? n32 : n63684;
  assign n63686 = pi21 ? n57774 : n2637;
  assign n63687 = pi20 ? n63686 : n32;
  assign n63688 = pi19 ? n56540 : n63687;
  assign n63689 = pi18 ? n40550 : n63688;
  assign n63690 = pi17 ? n32 : n63689;
  assign n63691 = pi16 ? n32 : n63690;
  assign n63692 = pi15 ? n63685 : n63691;
  assign n63693 = pi14 ? n63682 : n63692;
  assign n63694 = pi22 ? n56712 : n51564;
  assign n63695 = pi21 ? n63694 : n928;
  assign n63696 = pi20 ? n63695 : n32;
  assign n63697 = pi19 ? n56540 : n63696;
  assign n63698 = pi18 ? n39397 : n63697;
  assign n63699 = pi17 ? n32 : n63698;
  assign n63700 = pi16 ? n32 : n63699;
  assign n63701 = pi22 ? n57085 : n36798;
  assign n63702 = pi21 ? n20563 : n63701;
  assign n63703 = pi20 ? n20563 : n63702;
  assign n63704 = pi19 ? n63703 : n63265;
  assign n63705 = pi18 ? n39397 : n63704;
  assign n63706 = pi17 ? n32 : n63705;
  assign n63707 = pi16 ? n32 : n63706;
  assign n63708 = pi15 ? n63700 : n63707;
  assign n63709 = pi21 ? n20563 : n53463;
  assign n63710 = pi20 ? n20563 : n63709;
  assign n63711 = pi19 ? n63710 : n63275;
  assign n63712 = pi18 ? n39397 : n63711;
  assign n63713 = pi17 ? n32 : n63712;
  assign n63714 = pi16 ? n32 : n63713;
  assign n63715 = pi21 ? n20563 : n57562;
  assign n63716 = pi20 ? n20563 : n63715;
  assign n63717 = pi23 ? n55783 : n43198;
  assign n63718 = pi22 ? n63717 : n13481;
  assign n63719 = pi21 ? n63718 : n20952;
  assign n63720 = pi20 ? n63719 : n32;
  assign n63721 = pi19 ? n63716 : n63720;
  assign n63722 = pi18 ? n40550 : n63721;
  assign n63723 = pi17 ? n32 : n63722;
  assign n63724 = pi16 ? n32 : n63723;
  assign n63725 = pi15 ? n63714 : n63724;
  assign n63726 = pi14 ? n63708 : n63725;
  assign n63727 = pi13 ? n63693 : n63726;
  assign n63728 = pi12 ? n63667 : n63727;
  assign n63729 = pi21 ? n36489 : n61211;
  assign n63730 = pi20 ? n20563 : n63729;
  assign n63731 = pi19 ? n63730 : n62839;
  assign n63732 = pi18 ? n40550 : n63731;
  assign n63733 = pi17 ? n32 : n63732;
  assign n63734 = pi16 ? n32 : n63733;
  assign n63735 = pi19 ? n52230 : n59667;
  assign n63736 = pi22 ? n363 : n51564;
  assign n63737 = pi21 ? n30868 : n63736;
  assign n63738 = pi20 ? n30868 : n63737;
  assign n63739 = pi22 ? n62803 : n53982;
  assign n63740 = pi21 ? n63739 : n32;
  assign n63741 = pi20 ? n63740 : n32;
  assign n63742 = pi19 ? n63738 : n63741;
  assign n63743 = pi18 ? n63735 : n63742;
  assign n63744 = pi17 ? n32 : n63743;
  assign n63745 = pi16 ? n32 : n63744;
  assign n63746 = pi15 ? n63734 : n63745;
  assign n63747 = pi19 ? n52230 : n30868;
  assign n63748 = pi21 ? n36489 : n58794;
  assign n63749 = pi20 ? n30868 : n63748;
  assign n63750 = pi19 ? n63749 : n62858;
  assign n63751 = pi18 ? n63747 : n63750;
  assign n63752 = pi17 ? n32 : n63751;
  assign n63753 = pi16 ? n32 : n63752;
  assign n63754 = pi20 ? n62385 : n30868;
  assign n63755 = pi19 ? n63754 : n30868;
  assign n63756 = pi18 ? n63755 : n63332;
  assign n63757 = pi17 ? n32 : n63756;
  assign n63758 = pi16 ? n32 : n63757;
  assign n63759 = pi15 ? n63753 : n63758;
  assign n63760 = pi14 ? n63746 : n63759;
  assign n63761 = pi20 ? n47322 : n43010;
  assign n63762 = pi19 ? n63761 : n30868;
  assign n63763 = pi21 ? n42146 : n58804;
  assign n63764 = pi20 ? n30868 : n63763;
  assign n63765 = pi19 ? n63764 : n60046;
  assign n63766 = pi18 ? n63762 : n63765;
  assign n63767 = pi17 ? n32 : n63766;
  assign n63768 = pi16 ? n32 : n63767;
  assign n63769 = pi20 ? n47192 : n43010;
  assign n63770 = pi19 ? n63769 : n30868;
  assign n63771 = pi22 ? n43198 : n56622;
  assign n63772 = pi21 ? n36781 : n63771;
  assign n63773 = pi20 ? n30868 : n63772;
  assign n63774 = pi19 ? n63773 : n57717;
  assign n63775 = pi18 ? n63770 : n63774;
  assign n63776 = pi17 ? n32 : n63775;
  assign n63777 = pi16 ? n32 : n63776;
  assign n63778 = pi15 ? n63768 : n63777;
  assign n63779 = pi22 ? n14626 : n56622;
  assign n63780 = pi21 ? n38901 : n63779;
  assign n63781 = pi20 ? n30868 : n63780;
  assign n63782 = pi19 ? n63781 : n35482;
  assign n63783 = pi18 ? n47194 : n63782;
  assign n63784 = pi17 ? n32 : n63783;
  assign n63785 = pi16 ? n32 : n63784;
  assign n63786 = pi22 ? n14626 : n54563;
  assign n63787 = pi21 ? n36798 : n63786;
  assign n63788 = pi20 ? n63363 : n63787;
  assign n63789 = pi19 ? n63788 : n32;
  assign n63790 = pi18 ? n47194 : n63789;
  assign n63791 = pi17 ? n32 : n63790;
  assign n63792 = pi16 ? n32 : n63791;
  assign n63793 = pi15 ? n63785 : n63792;
  assign n63794 = pi14 ? n63778 : n63793;
  assign n63795 = pi13 ? n63760 : n63794;
  assign n63796 = pi20 ? n62445 : n33792;
  assign n63797 = pi19 ? n63796 : n33792;
  assign n63798 = pi21 ? n47396 : n58665;
  assign n63799 = pi20 ? n33792 : n63798;
  assign n63800 = pi19 ? n63799 : n32;
  assign n63801 = pi18 ? n63797 : n63800;
  assign n63802 = pi17 ? n32 : n63801;
  assign n63803 = pi16 ? n32 : n63802;
  assign n63804 = pi18 ? n63797 : n63387;
  assign n63805 = pi17 ? n32 : n63804;
  assign n63806 = pi16 ? n32 : n63805;
  assign n63807 = pi15 ? n63803 : n63806;
  assign n63808 = pi18 ? n58194 : n63397;
  assign n63809 = pi17 ? n32 : n63808;
  assign n63810 = pi16 ? n32 : n63809;
  assign n63811 = pi22 ? n46275 : n36798;
  assign n63812 = pi21 ? n32 : n63811;
  assign n63813 = pi20 ? n63812 : n43198;
  assign n63814 = pi19 ? n63813 : n43198;
  assign n63815 = pi18 ? n63814 : n63407;
  assign n63816 = pi17 ? n32 : n63815;
  assign n63817 = pi16 ? n32 : n63816;
  assign n63818 = pi15 ? n63810 : n63817;
  assign n63819 = pi14 ? n63807 : n63818;
  assign n63820 = pi20 ? n48857 : n43198;
  assign n63821 = pi19 ? n63820 : n43198;
  assign n63822 = pi18 ? n63821 : n63417;
  assign n63823 = pi17 ? n32 : n63822;
  assign n63824 = pi16 ? n32 : n63823;
  assign n63825 = pi18 ? n63821 : n63426;
  assign n63826 = pi17 ? n32 : n63825;
  assign n63827 = pi16 ? n32 : n63826;
  assign n63828 = pi15 ? n63824 : n63827;
  assign n63829 = pi22 ? n32 : n14626;
  assign n63830 = pi21 ? n32 : n63829;
  assign n63831 = pi20 ? n63830 : n14626;
  assign n63832 = pi19 ? n63831 : n14626;
  assign n63833 = pi18 ? n63832 : n63439;
  assign n63834 = pi17 ? n32 : n63833;
  assign n63835 = pi16 ? n32 : n63834;
  assign n63836 = pi22 ? n62510 : n36798;
  assign n63837 = pi21 ? n63836 : n36798;
  assign n63838 = pi20 ? n63837 : n36798;
  assign n63839 = pi19 ? n47343 : n63838;
  assign n63840 = pi21 ? n36798 : n42622;
  assign n63841 = pi20 ? n63840 : n59604;
  assign n63842 = pi19 ? n63841 : n32;
  assign n63843 = pi18 ? n63839 : n63842;
  assign n63844 = pi17 ? n32 : n63843;
  assign n63845 = pi16 ? n32 : n63844;
  assign n63846 = pi15 ? n63835 : n63845;
  assign n63847 = pi14 ? n63828 : n63846;
  assign n63848 = pi13 ? n63819 : n63847;
  assign n63849 = pi12 ? n63795 : n63848;
  assign n63850 = pi11 ? n63728 : n63849;
  assign n63851 = pi10 ? n63608 : n63850;
  assign n63852 = pi09 ? n63474 : n63851;
  assign n63853 = pi08 ? n63458 : n63852;
  assign n63854 = pi18 ? n31265 : n62949;
  assign n63855 = pi17 ? n32 : n63854;
  assign n63856 = pi16 ? n32 : n63855;
  assign n63857 = pi15 ? n32 : n63856;
  assign n63858 = pi18 ? n43217 : n62955;
  assign n63859 = pi17 ? n32 : n63858;
  assign n63860 = pi16 ? n32 : n63859;
  assign n63861 = pi18 ? n44273 : n62955;
  assign n63862 = pi17 ? n32 : n63861;
  assign n63863 = pi16 ? n32 : n63862;
  assign n63864 = pi15 ? n63860 : n63863;
  assign n63865 = pi14 ? n63857 : n63864;
  assign n63866 = pi13 ? n32 : n63865;
  assign n63867 = pi12 ? n32 : n63866;
  assign n63868 = pi11 ? n32 : n63867;
  assign n63869 = pi10 ? n32 : n63868;
  assign n63870 = pi18 ? n48623 : n62955;
  assign n63871 = pi17 ? n32 : n63870;
  assign n63872 = pi16 ? n32 : n63871;
  assign n63873 = pi18 ? n42644 : n62955;
  assign n63874 = pi17 ? n32 : n63873;
  assign n63875 = pi16 ? n32 : n63874;
  assign n63876 = pi15 ? n63872 : n63875;
  assign n63877 = pi18 ? n42644 : n62976;
  assign n63878 = pi17 ? n32 : n63877;
  assign n63879 = pi16 ? n32 : n63878;
  assign n63880 = pi18 ? n42654 : n62976;
  assign n63881 = pi17 ? n32 : n63880;
  assign n63882 = pi16 ? n32 : n63881;
  assign n63883 = pi15 ? n63879 : n63882;
  assign n63884 = pi14 ? n63876 : n63883;
  assign n63885 = pi18 ? n42680 : n62976;
  assign n63886 = pi17 ? n32 : n63885;
  assign n63887 = pi16 ? n32 : n63886;
  assign n63888 = pi15 ? n63882 : n63887;
  assign n63889 = pi18 ? n48120 : n62976;
  assign n63890 = pi17 ? n32 : n63889;
  assign n63891 = pi16 ? n32 : n63890;
  assign n63892 = pi15 ? n63891 : n62979;
  assign n63893 = pi14 ? n63888 : n63892;
  assign n63894 = pi13 ? n63884 : n63893;
  assign n63895 = pi18 ? n42206 : n62955;
  assign n63896 = pi17 ? n32 : n63895;
  assign n63897 = pi16 ? n32 : n63896;
  assign n63898 = pi18 ? n41630 : n62955;
  assign n63899 = pi17 ? n32 : n63898;
  assign n63900 = pi16 ? n32 : n63899;
  assign n63901 = pi15 ? n63897 : n63900;
  assign n63902 = pi14 ? n62979 : n63901;
  assign n63903 = pi18 ? n41630 : n59296;
  assign n63904 = pi17 ? n32 : n63903;
  assign n63905 = pi16 ? n32 : n63904;
  assign n63906 = pi18 ? n40485 : n59307;
  assign n63907 = pi17 ? n32 : n63906;
  assign n63908 = pi16 ? n32 : n63907;
  assign n63909 = pi15 ? n63905 : n63908;
  assign n63910 = pi18 ? n41157 : n63013;
  assign n63911 = pi17 ? n32 : n63910;
  assign n63912 = pi16 ? n32 : n63911;
  assign n63913 = pi18 ? n41157 : n63522;
  assign n63914 = pi17 ? n32 : n63913;
  assign n63915 = pi16 ? n32 : n63914;
  assign n63916 = pi15 ? n63912 : n63915;
  assign n63917 = pi14 ? n63909 : n63916;
  assign n63918 = pi13 ? n63902 : n63917;
  assign n63919 = pi12 ? n63894 : n63918;
  assign n63920 = pi24 ? n30868 : n51564;
  assign n63921 = pi23 ? n63920 : n51564;
  assign n63922 = pi22 ? n63921 : n51564;
  assign n63923 = pi21 ? n63922 : n60421;
  assign n63924 = pi20 ? n53356 : n63923;
  assign n63925 = pi19 ? n20563 : n63924;
  assign n63926 = pi18 ? n41157 : n63925;
  assign n63927 = pi17 ? n32 : n63926;
  assign n63928 = pi16 ? n32 : n63927;
  assign n63929 = pi18 ? n41168 : n63034;
  assign n63930 = pi17 ? n32 : n63929;
  assign n63931 = pi16 ? n32 : n63930;
  assign n63932 = pi15 ? n63928 : n63931;
  assign n63933 = pi18 ? n41168 : n63547;
  assign n63934 = pi17 ? n32 : n63933;
  assign n63935 = pi16 ? n32 : n63934;
  assign n63936 = pi18 ? n41168 : n63045;
  assign n63937 = pi17 ? n32 : n63936;
  assign n63938 = pi16 ? n32 : n63937;
  assign n63939 = pi15 ? n63935 : n63938;
  assign n63940 = pi14 ? n63932 : n63939;
  assign n63941 = pi21 ? n685 : n59357;
  assign n63942 = pi20 ? n53386 : n63941;
  assign n63943 = pi19 ? n20563 : n63942;
  assign n63944 = pi18 ? n40023 : n63943;
  assign n63945 = pi17 ? n32 : n63944;
  assign n63946 = pi16 ? n32 : n63945;
  assign n63947 = pi20 ? n63065 : n14723;
  assign n63948 = pi19 ? n20563 : n63947;
  assign n63949 = pi18 ? n41181 : n63948;
  assign n63950 = pi17 ? n32 : n63949;
  assign n63951 = pi16 ? n32 : n63950;
  assign n63952 = pi15 ? n63946 : n63951;
  assign n63953 = pi22 ? n20563 : n893;
  assign n63954 = pi21 ? n20563 : n63953;
  assign n63955 = pi20 ? n63954 : n63066;
  assign n63956 = pi19 ? n20563 : n63955;
  assign n63957 = pi18 ? n41181 : n63956;
  assign n63958 = pi17 ? n32 : n63957;
  assign n63959 = pi16 ? n32 : n63958;
  assign n63960 = pi22 ? n20563 : n456;
  assign n63961 = pi21 ? n20563 : n63960;
  assign n63962 = pi20 ? n63961 : n1010;
  assign n63963 = pi19 ? n20563 : n63962;
  assign n63964 = pi18 ? n41181 : n63963;
  assign n63965 = pi17 ? n32 : n63964;
  assign n63966 = pi16 ? n32 : n63965;
  assign n63967 = pi15 ? n63959 : n63966;
  assign n63968 = pi14 ? n63952 : n63967;
  assign n63969 = pi13 ? n63940 : n63968;
  assign n63970 = pi18 ? n42239 : n62121;
  assign n63971 = pi17 ? n32 : n63970;
  assign n63972 = pi16 ? n32 : n63971;
  assign n63973 = pi21 ? n20563 : n11146;
  assign n63974 = pi20 ? n63973 : n17510;
  assign n63975 = pi19 ? n20563 : n63974;
  assign n63976 = pi18 ? n42239 : n63975;
  assign n63977 = pi17 ? n32 : n63976;
  assign n63978 = pi16 ? n32 : n63977;
  assign n63979 = pi15 ? n63972 : n63978;
  assign n63980 = pi22 ? n20563 : n6833;
  assign n63981 = pi21 ? n45016 : n63980;
  assign n63982 = pi22 ? n233 : n54520;
  assign n63983 = pi21 ? n63982 : n32;
  assign n63984 = pi20 ? n63981 : n63983;
  assign n63985 = pi19 ? n20563 : n63984;
  assign n63986 = pi18 ? n47056 : n63985;
  assign n63987 = pi17 ? n32 : n63986;
  assign n63988 = pi16 ? n32 : n63987;
  assign n63989 = pi22 ? n30868 : n3472;
  assign n63990 = pi21 ? n20563 : n63989;
  assign n63991 = pi20 ? n63990 : n10326;
  assign n63992 = pi19 ? n20563 : n63991;
  assign n63993 = pi18 ? n47056 : n63992;
  assign n63994 = pi17 ? n32 : n63993;
  assign n63995 = pi16 ? n32 : n63994;
  assign n63996 = pi15 ? n63988 : n63995;
  assign n63997 = pi14 ? n63979 : n63996;
  assign n63998 = pi22 ? n139 : n60300;
  assign n63999 = pi21 ? n40986 : n63998;
  assign n64000 = pi20 ? n63999 : n58471;
  assign n64001 = pi19 ? n20563 : n64000;
  assign n64002 = pi18 ? n46446 : n64001;
  assign n64003 = pi17 ? n32 : n64002;
  assign n64004 = pi16 ? n32 : n64003;
  assign n64005 = pi22 ? n33792 : n2299;
  assign n64006 = pi21 ? n36489 : n64005;
  assign n64007 = pi20 ? n64006 : n4008;
  assign n64008 = pi19 ? n20563 : n64007;
  assign n64009 = pi18 ? n46446 : n64008;
  assign n64010 = pi17 ? n32 : n64009;
  assign n64011 = pi16 ? n32 : n64010;
  assign n64012 = pi15 ? n64004 : n64011;
  assign n64013 = pi22 ? n335 : n56936;
  assign n64014 = pi21 ? n45016 : n64013;
  assign n64015 = pi20 ? n64014 : n56130;
  assign n64016 = pi19 ? n40792 : n64015;
  assign n64017 = pi18 ? n46446 : n64016;
  assign n64018 = pi17 ? n32 : n64017;
  assign n64019 = pi16 ? n32 : n64018;
  assign n64020 = pi21 ? n47220 : n61211;
  assign n64021 = pi20 ? n64020 : n4116;
  assign n64022 = pi19 ? n40792 : n64021;
  assign n64023 = pi18 ? n46446 : n64022;
  assign n64024 = pi17 ? n32 : n64023;
  assign n64025 = pi16 ? n32 : n64024;
  assign n64026 = pi15 ? n64019 : n64025;
  assign n64027 = pi14 ? n64012 : n64026;
  assign n64028 = pi13 ? n63997 : n64027;
  assign n64029 = pi12 ? n63969 : n64028;
  assign n64030 = pi11 ? n63919 : n64029;
  assign n64031 = pi21 ? n55685 : n57671;
  assign n64032 = pi20 ? n64031 : n59674;
  assign n64033 = pi19 ? n59458 : n64032;
  assign n64034 = pi18 ? n46446 : n64033;
  assign n64035 = pi17 ? n32 : n64034;
  assign n64036 = pi16 ? n32 : n64035;
  assign n64037 = pi21 ? n47360 : n58999;
  assign n64038 = pi20 ? n64037 : n10011;
  assign n64039 = pi19 ? n59458 : n64038;
  assign n64040 = pi18 ? n40497 : n64039;
  assign n64041 = pi17 ? n32 : n64040;
  assign n64042 = pi16 ? n32 : n64041;
  assign n64043 = pi15 ? n64036 : n64042;
  assign n64044 = pi23 ? n62332 : n36659;
  assign n64045 = pi22 ? n36659 : n64044;
  assign n64046 = pi21 ? n64045 : n59681;
  assign n64047 = pi20 ? n64046 : n57716;
  assign n64048 = pi19 ? n50091 : n64047;
  assign n64049 = pi18 ? n40532 : n64048;
  assign n64050 = pi17 ? n32 : n64049;
  assign n64051 = pi16 ? n32 : n64050;
  assign n64052 = pi22 ? n20563 : n64044;
  assign n64053 = pi21 ? n64052 : n57733;
  assign n64054 = pi20 ? n64053 : n1822;
  assign n64055 = pi19 ? n20563 : n64054;
  assign n64056 = pi18 ? n41708 : n64055;
  assign n64057 = pi17 ? n32 : n64056;
  assign n64058 = pi16 ? n32 : n64057;
  assign n64059 = pi15 ? n64051 : n64058;
  assign n64060 = pi14 ? n64043 : n64059;
  assign n64061 = pi20 ? n37955 : n40791;
  assign n64062 = pi19 ? n64061 : n20563;
  assign n64063 = pi24 ? n20563 : n36659;
  assign n64064 = pi23 ? n64063 : n36781;
  assign n64065 = pi22 ? n30868 : n64064;
  assign n64066 = pi21 ? n64065 : n59691;
  assign n64067 = pi20 ? n64066 : n20953;
  assign n64068 = pi19 ? n40792 : n64067;
  assign n64069 = pi18 ? n64062 : n64068;
  assign n64070 = pi17 ? n32 : n64069;
  assign n64071 = pi16 ? n32 : n64070;
  assign n64072 = pi20 ? n57040 : n40791;
  assign n64073 = pi19 ? n64072 : n50101;
  assign n64074 = pi23 ? n56064 : n36781;
  assign n64075 = pi22 ? n40387 : n64074;
  assign n64076 = pi22 ? n14626 : n759;
  assign n64077 = pi21 ? n64075 : n64076;
  assign n64078 = pi20 ? n64077 : n32;
  assign n64079 = pi19 ? n40792 : n64078;
  assign n64080 = pi18 ? n64073 : n64079;
  assign n64081 = pi17 ? n32 : n64080;
  assign n64082 = pi16 ? n32 : n64081;
  assign n64083 = pi15 ? n64071 : n64082;
  assign n64084 = pi20 ? n61295 : n20563;
  assign n64085 = pi19 ? n64084 : n63190;
  assign n64086 = pi22 ? n37783 : n30868;
  assign n64087 = pi21 ? n64086 : n33792;
  assign n64088 = pi20 ? n20563 : n64087;
  assign n64089 = pi23 ? n61843 : n14626;
  assign n64090 = pi22 ? n33792 : n64089;
  assign n64091 = pi21 ? n64090 : n63786;
  assign n64092 = pi20 ? n64091 : n32;
  assign n64093 = pi19 ? n64088 : n64092;
  assign n64094 = pi18 ? n64085 : n64093;
  assign n64095 = pi17 ? n32 : n64094;
  assign n64096 = pi16 ? n32 : n64095;
  assign n64097 = pi19 ? n64084 : n63204;
  assign n64098 = pi22 ? n40428 : n58044;
  assign n64099 = pi21 ? n64098 : n53559;
  assign n64100 = pi20 ? n64099 : n32;
  assign n64101 = pi19 ? n59458 : n64100;
  assign n64102 = pi18 ? n64097 : n64101;
  assign n64103 = pi17 ? n32 : n64102;
  assign n64104 = pi16 ? n32 : n64103;
  assign n64105 = pi15 ? n64096 : n64104;
  assign n64106 = pi14 ? n64083 : n64105;
  assign n64107 = pi13 ? n64060 : n64106;
  assign n64108 = pi20 ? n59992 : n20563;
  assign n64109 = pi19 ? n64108 : n58562;
  assign n64110 = pi24 ? n36659 : n36798;
  assign n64111 = pi23 ? n64110 : n55783;
  assign n64112 = pi22 ? n335 : n64111;
  assign n64113 = pi21 ? n64112 : n58470;
  assign n64114 = pi20 ? n64113 : n32;
  assign n64115 = pi19 ? n56631 : n64114;
  assign n64116 = pi18 ? n64109 : n64115;
  assign n64117 = pi17 ? n32 : n64116;
  assign n64118 = pi16 ? n32 : n64117;
  assign n64119 = pi23 ? n60408 : n20563;
  assign n64120 = pi22 ? n51754 : n64119;
  assign n64121 = pi21 ? n32 : n64120;
  assign n64122 = pi22 ? n20563 : n55502;
  assign n64123 = pi21 ? n64122 : n20563;
  assign n64124 = pi20 ? n64121 : n64123;
  assign n64125 = pi22 ? n20563 : n59056;
  assign n64126 = pi21 ? n64125 : n20563;
  assign n64127 = pi20 ? n43935 : n64126;
  assign n64128 = pi19 ? n64124 : n64127;
  assign n64129 = pi24 ? n36659 : n43198;
  assign n64130 = pi23 ? n64129 : n60075;
  assign n64131 = pi22 ? n36781 : n64130;
  assign n64132 = pi21 ? n64131 : n55560;
  assign n64133 = pi20 ? n64132 : n32;
  assign n64134 = pi19 ? n56631 : n64133;
  assign n64135 = pi18 ? n64128 : n64134;
  assign n64136 = pi17 ? n32 : n64135;
  assign n64137 = pi16 ? n32 : n64136;
  assign n64138 = pi15 ? n64118 : n64137;
  assign n64139 = pi24 ? n36781 : n14626;
  assign n64140 = pi23 ? n64139 : n14626;
  assign n64141 = pi22 ? n36781 : n64140;
  assign n64142 = pi21 ? n64141 : n63240;
  assign n64143 = pi20 ? n64142 : n32;
  assign n64144 = pi19 ? n63239 : n64143;
  assign n64145 = pi18 ? n45366 : n64144;
  assign n64146 = pi17 ? n32 : n64145;
  assign n64147 = pi16 ? n32 : n64146;
  assign n64148 = pi24 ? n36781 : n51564;
  assign n64149 = pi23 ? n64148 : n51564;
  assign n64150 = pi22 ? n36781 : n64149;
  assign n64151 = pi21 ? n64150 : n59357;
  assign n64152 = pi20 ? n64151 : n32;
  assign n64153 = pi19 ? n56540 : n64152;
  assign n64154 = pi18 ? n45366 : n64153;
  assign n64155 = pi17 ? n32 : n64154;
  assign n64156 = pi16 ? n32 : n64155;
  assign n64157 = pi15 ? n64147 : n64156;
  assign n64158 = pi14 ? n64138 : n64157;
  assign n64159 = pi23 ? n157 : n36781;
  assign n64160 = pi24 ? n36798 : n51564;
  assign n64161 = pi23 ? n64160 : n51564;
  assign n64162 = pi22 ? n64159 : n64161;
  assign n64163 = pi21 ? n64162 : n37639;
  assign n64164 = pi20 ? n64163 : n32;
  assign n64165 = pi19 ? n59603 : n64164;
  assign n64166 = pi18 ? n45366 : n64165;
  assign n64167 = pi17 ? n32 : n64166;
  assign n64168 = pi16 ? n32 : n64167;
  assign n64169 = pi23 ? n204 : n36798;
  assign n64170 = pi22 ? n64169 : n62411;
  assign n64171 = pi21 ? n64170 : n37639;
  assign n64172 = pi20 ? n64171 : n32;
  assign n64173 = pi19 ? n63710 : n64172;
  assign n64174 = pi18 ? n45366 : n64173;
  assign n64175 = pi17 ? n32 : n64174;
  assign n64176 = pi16 ? n32 : n64175;
  assign n64177 = pi15 ? n64168 : n64176;
  assign n64178 = pi21 ? n20563 : n46260;
  assign n64179 = pi20 ? n20563 : n64178;
  assign n64180 = pi22 ? n55799 : n13481;
  assign n64181 = pi21 ? n64180 : n20952;
  assign n64182 = pi20 ? n64181 : n32;
  assign n64183 = pi19 ? n64179 : n64182;
  assign n64184 = pi18 ? n45366 : n64183;
  assign n64185 = pi17 ? n32 : n64184;
  assign n64186 = pi16 ? n32 : n64185;
  assign n64187 = pi21 ? n20563 : n53432;
  assign n64188 = pi20 ? n20563 : n64187;
  assign n64189 = pi22 ? n233 : n56665;
  assign n64190 = pi21 ? n64189 : n32;
  assign n64191 = pi20 ? n64190 : n32;
  assign n64192 = pi19 ? n64188 : n64191;
  assign n64193 = pi18 ? n38948 : n64192;
  assign n64194 = pi17 ? n32 : n64193;
  assign n64195 = pi16 ? n32 : n64194;
  assign n64196 = pi15 ? n64186 : n64195;
  assign n64197 = pi14 ? n64177 : n64196;
  assign n64198 = pi13 ? n64158 : n64197;
  assign n64199 = pi12 ? n64107 : n64198;
  assign n64200 = pi21 ? n36489 : n57671;
  assign n64201 = pi20 ? n20563 : n64200;
  assign n64202 = pi19 ? n64201 : n8296;
  assign n64203 = pi18 ? n38948 : n64202;
  assign n64204 = pi17 ? n32 : n64203;
  assign n64205 = pi16 ? n32 : n64204;
  assign n64206 = pi19 ? n61409 : n59667;
  assign n64207 = pi21 ? n30868 : n63253;
  assign n64208 = pi20 ? n30868 : n64207;
  assign n64209 = pi20 ? n58967 : n32;
  assign n64210 = pi19 ? n64208 : n64209;
  assign n64211 = pi18 ? n64206 : n64210;
  assign n64212 = pi17 ? n32 : n64211;
  assign n64213 = pi16 ? n32 : n64212;
  assign n64214 = pi15 ? n64205 : n64213;
  assign n64215 = pi20 ? n54401 : n30868;
  assign n64216 = pi19 ? n64215 : n30868;
  assign n64217 = pi22 ? n39190 : n33792;
  assign n64218 = pi21 ? n64217 : n63694;
  assign n64219 = pi20 ? n30868 : n64218;
  assign n64220 = pi19 ? n64219 : n60046;
  assign n64221 = pi18 ? n64216 : n64220;
  assign n64222 = pi17 ? n32 : n64221;
  assign n64223 = pi16 ? n32 : n64222;
  assign n64224 = pi22 ? n32 : n39190;
  assign n64225 = pi21 ? n32 : n64224;
  assign n64226 = pi20 ? n64225 : n30868;
  assign n64227 = pi19 ? n64226 : n30868;
  assign n64228 = pi22 ? n36659 : n62227;
  assign n64229 = pi23 ? n51564 : n36798;
  assign n64230 = pi22 ? n64229 : n62389;
  assign n64231 = pi21 ? n64228 : n64230;
  assign n64232 = pi20 ? n30868 : n64231;
  assign n64233 = pi19 ? n64232 : n60046;
  assign n64234 = pi18 ? n64227 : n64233;
  assign n64235 = pi17 ? n32 : n64234;
  assign n64236 = pi16 ? n32 : n64235;
  assign n64237 = pi15 ? n64223 : n64236;
  assign n64238 = pi14 ? n64214 : n64237;
  assign n64239 = pi20 ? n37933 : n43010;
  assign n64240 = pi19 ? n64239 : n30868;
  assign n64241 = pi22 ? n64229 : n13481;
  assign n64242 = pi21 ? n42146 : n64241;
  assign n64243 = pi20 ? n30868 : n64242;
  assign n64244 = pi19 ? n64243 : n37641;
  assign n64245 = pi18 ? n64240 : n64244;
  assign n64246 = pi17 ? n32 : n64245;
  assign n64247 = pi16 ? n32 : n64246;
  assign n64248 = pi22 ? n14626 : n59395;
  assign n64249 = pi21 ? n36781 : n64248;
  assign n64250 = pi20 ? n30868 : n64249;
  assign n64251 = pi19 ? n64250 : n32;
  assign n64252 = pi18 ? n64240 : n64251;
  assign n64253 = pi17 ? n32 : n64252;
  assign n64254 = pi16 ? n32 : n64253;
  assign n64255 = pi15 ? n64247 : n64254;
  assign n64256 = pi20 ? n37933 : n30868;
  assign n64257 = pi19 ? n64256 : n30868;
  assign n64258 = pi23 ? n51564 : n687;
  assign n64259 = pi22 ? n51564 : n64258;
  assign n64260 = pi21 ? n38901 : n64259;
  assign n64261 = pi20 ? n30868 : n64260;
  assign n64262 = pi19 ? n64261 : n32;
  assign n64263 = pi18 ? n64257 : n64262;
  assign n64264 = pi17 ? n32 : n64263;
  assign n64265 = pi16 ? n32 : n64264;
  assign n64266 = pi19 ? n61453 : n30868;
  assign n64267 = pi21 ? n36798 : n61401;
  assign n64268 = pi20 ? n63363 : n64267;
  assign n64269 = pi19 ? n64268 : n32;
  assign n64270 = pi18 ? n64266 : n64269;
  assign n64271 = pi17 ? n32 : n64270;
  assign n64272 = pi16 ? n32 : n64271;
  assign n64273 = pi15 ? n64265 : n64272;
  assign n64274 = pi14 ? n64255 : n64273;
  assign n64275 = pi13 ? n64238 : n64274;
  assign n64276 = pi20 ? n46061 : n33792;
  assign n64277 = pi19 ? n64276 : n33792;
  assign n64278 = pi22 ? n13481 : n56665;
  assign n64279 = pi21 ? n47396 : n64278;
  assign n64280 = pi20 ? n33792 : n64279;
  assign n64281 = pi19 ? n64280 : n32;
  assign n64282 = pi18 ? n64277 : n64281;
  assign n64283 = pi17 ? n32 : n64282;
  assign n64284 = pi16 ? n32 : n64283;
  assign n64285 = pi19 ? n61467 : n33792;
  assign n64286 = pi21 ? n55792 : n59648;
  assign n64287 = pi20 ? n61480 : n64286;
  assign n64288 = pi19 ? n64287 : n32;
  assign n64289 = pi18 ? n64285 : n64288;
  assign n64290 = pi17 ? n32 : n64289;
  assign n64291 = pi16 ? n32 : n64290;
  assign n64292 = pi15 ? n64284 : n64291;
  assign n64293 = pi22 ? n37276 : n43198;
  assign n64294 = pi21 ? n64293 : n43198;
  assign n64295 = pi20 ? n46277 : n64294;
  assign n64296 = pi19 ? n64295 : n43198;
  assign n64297 = pi23 ? n43198 : n60075;
  assign n64298 = pi22 ? n55766 : n64297;
  assign n64299 = pi21 ? n64298 : n55560;
  assign n64300 = pi20 ? n43198 : n64299;
  assign n64301 = pi19 ? n64300 : n32;
  assign n64302 = pi18 ? n64296 : n64301;
  assign n64303 = pi17 ? n32 : n64302;
  assign n64304 = pi16 ? n32 : n64303;
  assign n64305 = pi20 ? n32 : n55716;
  assign n64306 = pi19 ? n64305 : n43198;
  assign n64307 = pi22 ? n51564 : n57197;
  assign n64308 = pi21 ? n64307 : n53983;
  assign n64309 = pi20 ? n43198 : n64308;
  assign n64310 = pi19 ? n64309 : n32;
  assign n64311 = pi18 ? n64306 : n64310;
  assign n64312 = pi17 ? n32 : n64311;
  assign n64313 = pi16 ? n32 : n64312;
  assign n64314 = pi15 ? n64304 : n64313;
  assign n64315 = pi14 ? n64292 : n64314;
  assign n64316 = pi20 ? n32 : n46284;
  assign n64317 = pi19 ? n64316 : n43198;
  assign n64318 = pi22 ? n51564 : n61806;
  assign n64319 = pi21 ? n64318 : n2700;
  assign n64320 = pi20 ? n43198 : n64319;
  assign n64321 = pi19 ? n64320 : n32;
  assign n64322 = pi18 ? n64317 : n64321;
  assign n64323 = pi17 ? n32 : n64322;
  assign n64324 = pi16 ? n32 : n64323;
  assign n64325 = pi23 ? n14626 : n36781;
  assign n64326 = pi22 ? n36798 : n64325;
  assign n64327 = pi21 ? n64326 : n43198;
  assign n64328 = pi20 ? n32 : n64327;
  assign n64329 = pi21 ? n58777 : n43198;
  assign n64330 = pi20 ? n64329 : n43198;
  assign n64331 = pi19 ? n64328 : n64330;
  assign n64332 = pi22 ? n14626 : n36781;
  assign n64333 = pi22 ? n14626 : n43198;
  assign n64334 = pi21 ? n64332 : n64333;
  assign n64335 = pi22 ? n13481 : n56186;
  assign n64336 = pi21 ? n64335 : n20952;
  assign n64337 = pi20 ? n64334 : n64336;
  assign n64338 = pi19 ? n64337 : n32;
  assign n64339 = pi18 ? n64331 : n64338;
  assign n64340 = pi17 ? n32 : n64339;
  assign n64341 = pi16 ? n32 : n64340;
  assign n64342 = pi15 ? n64324 : n64341;
  assign n64343 = pi21 ? n55708 : n14626;
  assign n64344 = pi20 ? n32 : n64343;
  assign n64345 = pi19 ? n64344 : n14626;
  assign n64346 = pi18 ? n64345 : n63439;
  assign n64347 = pi17 ? n32 : n64346;
  assign n64348 = pi16 ? n32 : n64347;
  assign n64349 = pi21 ? n55800 : n36798;
  assign n64350 = pi20 ? n32 : n64349;
  assign n64351 = pi19 ? n64350 : n60600;
  assign n64352 = pi21 ? n36798 : n53551;
  assign n64353 = pi22 ? n56622 : n21502;
  assign n64354 = pi21 ? n64353 : n32;
  assign n64355 = pi20 ? n64352 : n64354;
  assign n64356 = pi19 ? n64355 : n32;
  assign n64357 = pi18 ? n64351 : n64356;
  assign n64358 = pi17 ? n32 : n64357;
  assign n64359 = pi16 ? n32 : n64358;
  assign n64360 = pi15 ? n64348 : n64359;
  assign n64361 = pi14 ? n64342 : n64360;
  assign n64362 = pi13 ? n64315 : n64361;
  assign n64363 = pi12 ? n64275 : n64362;
  assign n64364 = pi11 ? n64199 : n64363;
  assign n64365 = pi10 ? n64030 : n64364;
  assign n64366 = pi09 ? n63869 : n64365;
  assign n64367 = pi18 ? n38378 : n62949;
  assign n64368 = pi17 ? n32 : n64367;
  assign n64369 = pi16 ? n32 : n64368;
  assign n64370 = pi15 ? n32 : n64369;
  assign n64371 = pi18 ? n44246 : n62955;
  assign n64372 = pi17 ? n32 : n64371;
  assign n64373 = pi16 ? n32 : n64372;
  assign n64374 = pi15 ? n63860 : n64373;
  assign n64375 = pi14 ? n64370 : n64374;
  assign n64376 = pi13 ? n32 : n64375;
  assign n64377 = pi12 ? n32 : n64376;
  assign n64378 = pi11 ? n32 : n64377;
  assign n64379 = pi10 ? n32 : n64378;
  assign n64380 = pi18 ? n43222 : n62955;
  assign n64381 = pi17 ? n32 : n64380;
  assign n64382 = pi16 ? n32 : n64381;
  assign n64383 = pi18 ? n43226 : n62955;
  assign n64384 = pi17 ? n32 : n64383;
  assign n64385 = pi16 ? n32 : n64384;
  assign n64386 = pi15 ? n64382 : n64385;
  assign n64387 = pi18 ? n43226 : n62976;
  assign n64388 = pi17 ? n32 : n64387;
  assign n64389 = pi16 ? n32 : n64388;
  assign n64390 = pi18 ? n43247 : n62976;
  assign n64391 = pi17 ? n32 : n64390;
  assign n64392 = pi16 ? n32 : n64391;
  assign n64393 = pi15 ? n64389 : n64392;
  assign n64394 = pi14 ? n64386 : n64393;
  assign n64395 = pi18 ? n44273 : n62976;
  assign n64396 = pi17 ? n32 : n64395;
  assign n64397 = pi16 ? n32 : n64396;
  assign n64398 = pi15 ? n64392 : n64397;
  assign n64399 = pi18 ? n42193 : n62976;
  assign n64400 = pi17 ? n32 : n64399;
  assign n64401 = pi16 ? n32 : n64400;
  assign n64402 = pi15 ? n64401 : n63484;
  assign n64403 = pi14 ? n64398 : n64402;
  assign n64404 = pi13 ? n64394 : n64403;
  assign n64405 = pi18 ? n42200 : n62955;
  assign n64406 = pi17 ? n32 : n64405;
  assign n64407 = pi16 ? n32 : n64406;
  assign n64408 = pi14 ? n63484 : n64407;
  assign n64409 = pi18 ? n43261 : n59296;
  assign n64410 = pi17 ? n32 : n64409;
  assign n64411 = pi16 ? n32 : n64410;
  assign n64412 = pi18 ? n48120 : n59307;
  assign n64413 = pi17 ? n32 : n64412;
  assign n64414 = pi16 ? n32 : n64413;
  assign n64415 = pi15 ? n64411 : n64414;
  assign n64416 = pi18 ? n47592 : n63013;
  assign n64417 = pi17 ? n32 : n64416;
  assign n64418 = pi16 ? n32 : n64417;
  assign n64419 = pi24 ? n99 : n685;
  assign n64420 = pi23 ? n64419 : n685;
  assign n64421 = pi22 ? n64420 : n685;
  assign n64422 = pi21 ? n64421 : n8486;
  assign n64423 = pi20 ? n53343 : n64422;
  assign n64424 = pi19 ? n20563 : n64423;
  assign n64425 = pi18 ? n47592 : n64424;
  assign n64426 = pi17 ? n32 : n64425;
  assign n64427 = pi16 ? n32 : n64426;
  assign n64428 = pi15 ? n64418 : n64427;
  assign n64429 = pi14 ? n64415 : n64428;
  assign n64430 = pi13 ? n64408 : n64429;
  assign n64431 = pi12 ? n64404 : n64430;
  assign n64432 = pi24 ? n139 : n51564;
  assign n64433 = pi23 ? n64432 : n51564;
  assign n64434 = pi22 ? n64433 : n51564;
  assign n64435 = pi21 ? n64434 : n60421;
  assign n64436 = pi20 ? n53356 : n64435;
  assign n64437 = pi19 ? n20563 : n64436;
  assign n64438 = pi18 ? n47592 : n64437;
  assign n64439 = pi17 ? n32 : n64438;
  assign n64440 = pi16 ? n32 : n64439;
  assign n64441 = pi21 ? n57350 : n2320;
  assign n64442 = pi20 ? n53356 : n64441;
  assign n64443 = pi19 ? n20563 : n64442;
  assign n64444 = pi18 ? n42206 : n64443;
  assign n64445 = pi17 ? n32 : n64444;
  assign n64446 = pi16 ? n32 : n64445;
  assign n64447 = pi15 ? n64440 : n64446;
  assign n64448 = pi22 ? n56936 : n13481;
  assign n64449 = pi21 ? n64448 : n37639;
  assign n64450 = pi20 ? n53367 : n64449;
  assign n64451 = pi19 ? n20563 : n64450;
  assign n64452 = pi18 ? n41630 : n64451;
  assign n64453 = pi17 ? n32 : n64452;
  assign n64454 = pi16 ? n32 : n64453;
  assign n64455 = pi18 ? n41630 : n63045;
  assign n64456 = pi17 ? n32 : n64455;
  assign n64457 = pi16 ? n32 : n64456;
  assign n64458 = pi15 ? n64454 : n64457;
  assign n64459 = pi14 ? n64447 : n64458;
  assign n64460 = pi18 ? n46997 : n63943;
  assign n64461 = pi17 ? n32 : n64460;
  assign n64462 = pi16 ? n32 : n64461;
  assign n64463 = pi18 ? n40485 : n63948;
  assign n64464 = pi17 ? n32 : n64463;
  assign n64465 = pi16 ? n32 : n64464;
  assign n64466 = pi15 ? n64462 : n64465;
  assign n64467 = pi20 ? n63954 : n58944;
  assign n64468 = pi19 ? n20563 : n64467;
  assign n64469 = pi18 ? n40485 : n64468;
  assign n64470 = pi17 ? n32 : n64469;
  assign n64471 = pi16 ? n32 : n64470;
  assign n64472 = pi18 ? n40485 : n63963;
  assign n64473 = pi17 ? n32 : n64472;
  assign n64474 = pi16 ? n32 : n64473;
  assign n64475 = pi15 ? n64471 : n64474;
  assign n64476 = pi14 ? n64466 : n64475;
  assign n64477 = pi13 ? n64459 : n64476;
  assign n64478 = pi18 ? n41157 : n62121;
  assign n64479 = pi17 ? n32 : n64478;
  assign n64480 = pi16 ? n32 : n64479;
  assign n64481 = pi18 ? n41157 : n63975;
  assign n64482 = pi17 ? n32 : n64481;
  assign n64483 = pi16 ? n32 : n64482;
  assign n64484 = pi15 ? n64480 : n64483;
  assign n64485 = pi18 ? n41157 : n63985;
  assign n64486 = pi17 ? n32 : n64485;
  assign n64487 = pi16 ? n32 : n64486;
  assign n64488 = pi18 ? n41168 : n63992;
  assign n64489 = pi17 ? n32 : n64488;
  assign n64490 = pi16 ? n32 : n64489;
  assign n64491 = pi15 ? n64487 : n64490;
  assign n64492 = pi14 ? n64484 : n64491;
  assign n64493 = pi18 ? n40023 : n64001;
  assign n64494 = pi17 ? n32 : n64493;
  assign n64495 = pi16 ? n32 : n64494;
  assign n64496 = pi18 ? n40023 : n64008;
  assign n64497 = pi17 ? n32 : n64496;
  assign n64498 = pi16 ? n32 : n64497;
  assign n64499 = pi15 ? n64495 : n64498;
  assign n64500 = pi18 ? n40023 : n64016;
  assign n64501 = pi17 ? n32 : n64500;
  assign n64502 = pi16 ? n32 : n64501;
  assign n64503 = pi18 ? n40023 : n64022;
  assign n64504 = pi17 ? n32 : n64503;
  assign n64505 = pi16 ? n32 : n64504;
  assign n64506 = pi15 ? n64502 : n64505;
  assign n64507 = pi14 ? n64499 : n64506;
  assign n64508 = pi13 ? n64492 : n64507;
  assign n64509 = pi12 ? n64477 : n64508;
  assign n64510 = pi11 ? n64431 : n64509;
  assign n64511 = pi18 ? n40023 : n64033;
  assign n64512 = pi17 ? n32 : n64511;
  assign n64513 = pi16 ? n32 : n64512;
  assign n64514 = pi18 ? n41181 : n64039;
  assign n64515 = pi17 ? n32 : n64514;
  assign n64516 = pi16 ? n32 : n64515;
  assign n64517 = pi15 ? n64513 : n64516;
  assign n64518 = pi22 ? n36659 : n58710;
  assign n64519 = pi21 ? n64518 : n59681;
  assign n64520 = pi20 ? n64519 : n57716;
  assign n64521 = pi19 ? n50091 : n64520;
  assign n64522 = pi18 ? n41181 : n64521;
  assign n64523 = pi17 ? n32 : n64522;
  assign n64524 = pi16 ? n32 : n64523;
  assign n64525 = pi23 ? n1342 : n36659;
  assign n64526 = pi22 ? n20563 : n64525;
  assign n64527 = pi21 ? n64526 : n57733;
  assign n64528 = pi20 ? n64527 : n1822;
  assign n64529 = pi19 ? n20563 : n64528;
  assign n64530 = pi18 ? n42239 : n64529;
  assign n64531 = pi17 ? n32 : n64530;
  assign n64532 = pi16 ? n32 : n64531;
  assign n64533 = pi15 ? n64524 : n64532;
  assign n64534 = pi14 ? n64517 : n64533;
  assign n64535 = pi21 ? n30155 : n30868;
  assign n64536 = pi20 ? n32 : n64535;
  assign n64537 = pi19 ? n64536 : n20563;
  assign n64538 = pi24 ? n99 : n36659;
  assign n64539 = pi23 ? n64538 : n36781;
  assign n64540 = pi22 ? n30868 : n64539;
  assign n64541 = pi21 ? n64540 : n59691;
  assign n64542 = pi20 ? n64541 : n20953;
  assign n64543 = pi19 ? n40792 : n64542;
  assign n64544 = pi18 ? n64537 : n64543;
  assign n64545 = pi17 ? n32 : n64544;
  assign n64546 = pi16 ? n32 : n64545;
  assign n64547 = pi19 ? n64536 : n50101;
  assign n64548 = pi24 ? n139 : n36781;
  assign n64549 = pi23 ? n64548 : n36781;
  assign n64550 = pi22 ? n745 : n64549;
  assign n64551 = pi21 ? n64550 : n64076;
  assign n64552 = pi20 ? n64551 : n32;
  assign n64553 = pi19 ? n40792 : n64552;
  assign n64554 = pi18 ? n64547 : n64553;
  assign n64555 = pi17 ? n32 : n64554;
  assign n64556 = pi16 ? n32 : n64555;
  assign n64557 = pi15 ? n64546 : n64556;
  assign n64558 = pi19 ? n31264 : n63190;
  assign n64559 = pi23 ? n64548 : n14626;
  assign n64560 = pi22 ? n33792 : n64559;
  assign n64561 = pi21 ? n64560 : n63786;
  assign n64562 = pi20 ? n64561 : n32;
  assign n64563 = pi19 ? n64088 : n64562;
  assign n64564 = pi18 ? n64558 : n64563;
  assign n64565 = pi17 ? n32 : n64564;
  assign n64566 = pi16 ? n32 : n64565;
  assign n64567 = pi19 ? n31264 : n63204;
  assign n64568 = pi21 ? n40960 : n33792;
  assign n64569 = pi20 ? n20563 : n64568;
  assign n64570 = pi24 ? n335 : n36798;
  assign n64571 = pi23 ? n64570 : n14626;
  assign n64572 = pi22 ? n9827 : n64571;
  assign n64573 = pi21 ? n64572 : n53559;
  assign n64574 = pi20 ? n64573 : n32;
  assign n64575 = pi19 ? n64569 : n64574;
  assign n64576 = pi18 ? n64567 : n64575;
  assign n64577 = pi17 ? n32 : n64576;
  assign n64578 = pi16 ? n32 : n64577;
  assign n64579 = pi15 ? n64566 : n64578;
  assign n64580 = pi14 ? n64557 : n64579;
  assign n64581 = pi13 ? n64534 : n64580;
  assign n64582 = pi21 ? n30866 : n62770;
  assign n64583 = pi20 ? n32 : n64582;
  assign n64584 = pi19 ? n64583 : n59029;
  assign n64585 = pi21 ? n40960 : n36659;
  assign n64586 = pi20 ? n20563 : n64585;
  assign n64587 = pi24 ? n335 : n204;
  assign n64588 = pi23 ? n64587 : n51564;
  assign n64589 = pi22 ? n335 : n64588;
  assign n64590 = pi21 ? n64589 : n58470;
  assign n64591 = pi20 ? n64590 : n32;
  assign n64592 = pi19 ? n64586 : n64591;
  assign n64593 = pi18 ? n64584 : n64592;
  assign n64594 = pi17 ? n32 : n64593;
  assign n64595 = pi16 ? n32 : n64594;
  assign n64596 = pi19 ? n40509 : n38478;
  assign n64597 = pi23 ? n43198 : n61508;
  assign n64598 = pi22 ? n36781 : n64597;
  assign n64599 = pi21 ? n64598 : n55560;
  assign n64600 = pi20 ? n64599 : n32;
  assign n64601 = pi19 ? n56631 : n64600;
  assign n64602 = pi18 ? n64596 : n64601;
  assign n64603 = pi17 ? n32 : n64602;
  assign n64604 = pi16 ? n32 : n64603;
  assign n64605 = pi15 ? n64595 : n64604;
  assign n64606 = pi23 ? n233 : n14626;
  assign n64607 = pi22 ? n36781 : n64606;
  assign n64608 = pi23 ? n63306 : n32;
  assign n64609 = pi22 ? n64608 : n32;
  assign n64610 = pi21 ? n64607 : n64609;
  assign n64611 = pi20 ? n64610 : n32;
  assign n64612 = pi19 ? n63239 : n64611;
  assign n64613 = pi18 ? n40510 : n64612;
  assign n64614 = pi17 ? n32 : n64613;
  assign n64615 = pi16 ? n32 : n64614;
  assign n64616 = pi22 ? n56776 : n57197;
  assign n64617 = pi21 ? n64616 : n59357;
  assign n64618 = pi20 ? n64617 : n32;
  assign n64619 = pi19 ? n56540 : n64618;
  assign n64620 = pi18 ? n40510 : n64619;
  assign n64621 = pi17 ? n32 : n64620;
  assign n64622 = pi16 ? n32 : n64621;
  assign n64623 = pi15 ? n64615 : n64622;
  assign n64624 = pi14 ? n64605 : n64623;
  assign n64625 = pi22 ? n18448 : n51564;
  assign n64626 = pi21 ? n64625 : n37639;
  assign n64627 = pi20 ? n64626 : n32;
  assign n64628 = pi19 ? n59603 : n64627;
  assign n64629 = pi18 ? n40510 : n64628;
  assign n64630 = pi17 ? n32 : n64629;
  assign n64631 = pi16 ? n32 : n64630;
  assign n64632 = pi22 ? n204 : n56186;
  assign n64633 = pi21 ? n64632 : n37639;
  assign n64634 = pi20 ? n64633 : n32;
  assign n64635 = pi19 ? n63710 : n64634;
  assign n64636 = pi18 ? n40510 : n64635;
  assign n64637 = pi17 ? n32 : n64636;
  assign n64638 = pi16 ? n32 : n64637;
  assign n64639 = pi15 ? n64631 : n64638;
  assign n64640 = pi21 ? n55767 : n20952;
  assign n64641 = pi20 ? n64640 : n32;
  assign n64642 = pi19 ? n64179 : n64641;
  assign n64643 = pi18 ? n46446 : n64642;
  assign n64644 = pi17 ? n32 : n64643;
  assign n64645 = pi16 ? n32 : n64644;
  assign n64646 = pi18 ? n40497 : n64192;
  assign n64647 = pi17 ? n32 : n64646;
  assign n64648 = pi16 ? n32 : n64647;
  assign n64649 = pi15 ? n64645 : n64648;
  assign n64650 = pi14 ? n64639 : n64649;
  assign n64651 = pi13 ? n64624 : n64650;
  assign n64652 = pi12 ? n64581 : n64651;
  assign n64653 = pi21 ? n48173 : n57671;
  assign n64654 = pi20 ? n20563 : n64653;
  assign n64655 = pi21 ? n58086 : n32;
  assign n64656 = pi20 ? n64655 : n32;
  assign n64657 = pi19 ? n64654 : n64656;
  assign n64658 = pi18 ? n40497 : n64657;
  assign n64659 = pi17 ? n32 : n64658;
  assign n64660 = pi16 ? n32 : n64659;
  assign n64661 = pi19 ? n47836 : n59667;
  assign n64662 = pi23 ? n30868 : n55567;
  assign n64663 = pi22 ? n30868 : n64662;
  assign n64664 = pi21 ? n64663 : n63253;
  assign n64665 = pi20 ? n30868 : n64664;
  assign n64666 = pi19 ? n64665 : n64209;
  assign n64667 = pi18 ? n64661 : n64666;
  assign n64668 = pi17 ? n32 : n64667;
  assign n64669 = pi16 ? n32 : n64668;
  assign n64670 = pi15 ? n64660 : n64669;
  assign n64671 = pi22 ? n37218 : n58710;
  assign n64672 = pi21 ? n64671 : n59681;
  assign n64673 = pi20 ? n30868 : n64672;
  assign n64674 = pi19 ? n64673 : n60046;
  assign n64675 = pi18 ? n59115 : n64674;
  assign n64676 = pi17 ? n32 : n64675;
  assign n64677 = pi16 ? n32 : n64676;
  assign n64678 = pi23 ? n51564 : n43198;
  assign n64679 = pi22 ? n64678 : n56622;
  assign n64680 = pi21 ? n50801 : n64679;
  assign n64681 = pi20 ? n30868 : n64680;
  assign n64682 = pi19 ? n64681 : n60046;
  assign n64683 = pi18 ? n59115 : n64682;
  assign n64684 = pi17 ? n32 : n64683;
  assign n64685 = pi16 ? n32 : n64684;
  assign n64686 = pi15 ? n64677 : n64685;
  assign n64687 = pi14 ? n64670 : n64686;
  assign n64688 = pi19 ? n59109 : n30868;
  assign n64689 = pi23 ? n51564 : n14626;
  assign n64690 = pi22 ? n64689 : n13481;
  assign n64691 = pi21 ? n40002 : n64690;
  assign n64692 = pi20 ? n30868 : n64691;
  assign n64693 = pi19 ? n64692 : n37641;
  assign n64694 = pi18 ? n64688 : n64693;
  assign n64695 = pi17 ? n32 : n64694;
  assign n64696 = pi16 ? n32 : n64695;
  assign n64697 = pi22 ? n14626 : n64258;
  assign n64698 = pi21 ? n36781 : n64697;
  assign n64699 = pi20 ? n30868 : n64698;
  assign n64700 = pi19 ? n64699 : n32;
  assign n64701 = pi18 ? n64688 : n64700;
  assign n64702 = pi17 ? n32 : n64701;
  assign n64703 = pi16 ? n32 : n64702;
  assign n64704 = pi15 ? n64696 : n64703;
  assign n64705 = pi22 ? n36798 : n49412;
  assign n64706 = pi22 ? n51564 : n59672;
  assign n64707 = pi21 ? n64705 : n64706;
  assign n64708 = pi20 ? n30868 : n64707;
  assign n64709 = pi19 ? n64708 : n32;
  assign n64710 = pi18 ? n59115 : n64709;
  assign n64711 = pi17 ? n32 : n64710;
  assign n64712 = pi16 ? n32 : n64711;
  assign n64713 = pi18 ? n48361 : n64269;
  assign n64714 = pi17 ? n32 : n64713;
  assign n64715 = pi16 ? n32 : n64714;
  assign n64716 = pi15 ? n64712 : n64715;
  assign n64717 = pi14 ? n64704 : n64716;
  assign n64718 = pi13 ? n64687 : n64717;
  assign n64719 = pi21 ? n56207 : n64278;
  assign n64720 = pi20 ? n33792 : n64719;
  assign n64721 = pi19 ? n64720 : n32;
  assign n64722 = pi18 ? n53321 : n64721;
  assign n64723 = pi17 ? n32 : n64722;
  assign n64724 = pi16 ? n32 : n64723;
  assign n64725 = pi19 ? n45519 : n33792;
  assign n64726 = pi22 ? n61543 : n55766;
  assign n64727 = pi21 ? n64726 : n56129;
  assign n64728 = pi20 ? n61480 : n64727;
  assign n64729 = pi19 ? n64728 : n32;
  assign n64730 = pi18 ? n64725 : n64729;
  assign n64731 = pi17 ? n32 : n64730;
  assign n64732 = pi16 ? n32 : n64731;
  assign n64733 = pi15 ? n64724 : n64732;
  assign n64734 = pi19 ? n53549 : n43198;
  assign n64735 = pi23 ? n14626 : n233;
  assign n64736 = pi22 ? n64735 : n233;
  assign n64737 = pi21 ? n64736 : n2678;
  assign n64738 = pi20 ? n43198 : n64737;
  assign n64739 = pi19 ? n64738 : n32;
  assign n64740 = pi18 ? n64734 : n64739;
  assign n64741 = pi17 ? n32 : n64740;
  assign n64742 = pi16 ? n32 : n64741;
  assign n64743 = pi18 ? n64734 : n64310;
  assign n64744 = pi17 ? n32 : n64743;
  assign n64745 = pi16 ? n32 : n64744;
  assign n64746 = pi15 ? n64742 : n64745;
  assign n64747 = pi14 ? n64733 : n64746;
  assign n64748 = pi20 ? n43198 : n59583;
  assign n64749 = pi19 ? n64748 : n32;
  assign n64750 = pi18 ? n64734 : n64749;
  assign n64751 = pi17 ? n32 : n64750;
  assign n64752 = pi16 ? n32 : n64751;
  assign n64753 = pi21 ? n63829 : n43198;
  assign n64754 = pi20 ? n32 : n64753;
  assign n64755 = pi19 ? n64754 : n64330;
  assign n64756 = pi18 ? n64755 : n64338;
  assign n64757 = pi17 ? n32 : n64756;
  assign n64758 = pi16 ? n32 : n64757;
  assign n64759 = pi15 ? n64752 : n64758;
  assign n64760 = pi21 ? n63829 : n14626;
  assign n64761 = pi20 ? n32 : n64760;
  assign n64762 = pi19 ? n64761 : n14626;
  assign n64763 = pi18 ? n64762 : n63439;
  assign n64764 = pi17 ? n32 : n64763;
  assign n64765 = pi16 ? n32 : n64764;
  assign n64766 = pi21 ? n45653 : n53551;
  assign n64767 = pi20 ? n32 : n64766;
  assign n64768 = pi24 ? n43198 : n36798;
  assign n64769 = pi23 ? n64768 : n36798;
  assign n64770 = pi22 ? n64769 : n36798;
  assign n64771 = pi21 ? n64770 : n36798;
  assign n64772 = pi21 ? n60934 : n36798;
  assign n64773 = pi20 ? n64771 : n64772;
  assign n64774 = pi19 ? n64767 : n64773;
  assign n64775 = pi18 ? n64774 : n64356;
  assign n64776 = pi17 ? n32 : n64775;
  assign n64777 = pi16 ? n32 : n64776;
  assign n64778 = pi15 ? n64765 : n64777;
  assign n64779 = pi14 ? n64759 : n64778;
  assign n64780 = pi13 ? n64747 : n64779;
  assign n64781 = pi12 ? n64718 : n64780;
  assign n64782 = pi11 ? n64652 : n64781;
  assign n64783 = pi10 ? n64510 : n64782;
  assign n64784 = pi09 ? n64379 : n64783;
  assign n64785 = pi08 ? n64366 : n64784;
  assign n64786 = pi07 ? n63853 : n64785;
  assign n64787 = pi21 ? n20563 : n12224;
  assign n64788 = pi20 ? n20563 : n64787;
  assign n64789 = pi19 ? n20563 : n64788;
  assign n64790 = pi18 ? n37957 : n64789;
  assign n64791 = pi17 ? n32 : n64790;
  assign n64792 = pi16 ? n32 : n64791;
  assign n64793 = pi15 ? n32 : n64792;
  assign n64794 = pi18 ? n39455 : n62955;
  assign n64795 = pi17 ? n32 : n64794;
  assign n64796 = pi16 ? n32 : n64795;
  assign n64797 = pi18 ? n28159 : n62955;
  assign n64798 = pi17 ? n32 : n64797;
  assign n64799 = pi16 ? n32 : n64798;
  assign n64800 = pi15 ? n64796 : n64799;
  assign n64801 = pi14 ? n64793 : n64800;
  assign n64802 = pi13 ? n32 : n64801;
  assign n64803 = pi12 ? n32 : n64802;
  assign n64804 = pi11 ? n32 : n64803;
  assign n64805 = pi10 ? n32 : n64804;
  assign n64806 = pi18 ? n30119 : n62955;
  assign n64807 = pi17 ? n32 : n64806;
  assign n64808 = pi16 ? n32 : n64807;
  assign n64809 = pi18 ? n31265 : n62955;
  assign n64810 = pi17 ? n32 : n64809;
  assign n64811 = pi16 ? n32 : n64810;
  assign n64812 = pi15 ? n64808 : n64811;
  assign n64813 = pi18 ? n31265 : n62976;
  assign n64814 = pi17 ? n32 : n64813;
  assign n64815 = pi16 ? n32 : n64814;
  assign n64816 = pi18 ? n31315 : n62976;
  assign n64817 = pi17 ? n32 : n64816;
  assign n64818 = pi16 ? n32 : n64817;
  assign n64819 = pi15 ? n64815 : n64818;
  assign n64820 = pi14 ? n64812 : n64819;
  assign n64821 = pi18 ? n44246 : n62976;
  assign n64822 = pi17 ? n32 : n64821;
  assign n64823 = pi16 ? n32 : n64822;
  assign n64824 = pi15 ? n64818 : n64823;
  assign n64825 = pi18 ? n48623 : n62976;
  assign n64826 = pi17 ? n32 : n64825;
  assign n64827 = pi16 ? n32 : n64826;
  assign n64828 = pi15 ? n64827 : n63879;
  assign n64829 = pi14 ? n64824 : n64828;
  assign n64830 = pi13 ? n64820 : n64829;
  assign n64831 = pi14 ? n63879 : n62958;
  assign n64832 = pi18 ? n42680 : n59296;
  assign n64833 = pi17 ? n32 : n64832;
  assign n64834 = pi16 ? n32 : n64833;
  assign n64835 = pi18 ? n42193 : n59307;
  assign n64836 = pi17 ? n32 : n64835;
  assign n64837 = pi16 ? n32 : n64836;
  assign n64838 = pi15 ? n64834 : n64837;
  assign n64839 = pi24 ? n20563 : n233;
  assign n64840 = pi23 ? n64839 : n14626;
  assign n64841 = pi22 ? n64840 : n14626;
  assign n64842 = pi22 ? n14626 : n63009;
  assign n64843 = pi21 ? n64841 : n64842;
  assign n64844 = pi20 ? n38754 : n64843;
  assign n64845 = pi19 ? n20563 : n64844;
  assign n64846 = pi18 ? n43254 : n64845;
  assign n64847 = pi17 ? n32 : n64846;
  assign n64848 = pi16 ? n32 : n64847;
  assign n64849 = pi20 ? n38754 : n64422;
  assign n64850 = pi19 ? n20563 : n64849;
  assign n64851 = pi18 ? n43254 : n64850;
  assign n64852 = pi17 ? n32 : n64851;
  assign n64853 = pi16 ? n32 : n64852;
  assign n64854 = pi15 ? n64848 : n64853;
  assign n64855 = pi14 ? n64838 : n64854;
  assign n64856 = pi13 ? n64831 : n64855;
  assign n64857 = pi12 ? n64830 : n64856;
  assign n64858 = pi22 ? n64433 : n316;
  assign n64859 = pi21 ? n64858 : n2320;
  assign n64860 = pi20 ? n47158 : n64859;
  assign n64861 = pi19 ? n20563 : n64860;
  assign n64862 = pi18 ? n43254 : n64861;
  assign n64863 = pi17 ? n32 : n64862;
  assign n64864 = pi16 ? n32 : n64863;
  assign n64865 = pi18 ? n42200 : n64443;
  assign n64866 = pi17 ? n32 : n64865;
  assign n64867 = pi16 ? n32 : n64866;
  assign n64868 = pi15 ? n64864 : n64867;
  assign n64869 = pi20 ? n55475 : n59343;
  assign n64870 = pi19 ? n20563 : n64869;
  assign n64871 = pi18 ? n42200 : n64870;
  assign n64872 = pi17 ? n32 : n64871;
  assign n64873 = pi16 ? n32 : n64872;
  assign n64874 = pi20 ? n55475 : n23203;
  assign n64875 = pi19 ? n20563 : n64874;
  assign n64876 = pi18 ? n43261 : n64875;
  assign n64877 = pi17 ? n32 : n64876;
  assign n64878 = pi16 ? n32 : n64877;
  assign n64879 = pi15 ? n64873 : n64878;
  assign n64880 = pi14 ? n64868 : n64879;
  assign n64881 = pi21 ? n20563 : n51313;
  assign n64882 = pi20 ? n64881 : n63941;
  assign n64883 = pi19 ? n20563 : n64882;
  assign n64884 = pi18 ? n43261 : n64883;
  assign n64885 = pi17 ? n32 : n64884;
  assign n64886 = pi16 ? n32 : n64885;
  assign n64887 = pi22 ? n30868 : n58428;
  assign n64888 = pi21 ? n20563 : n64887;
  assign n64889 = pi20 ? n64888 : n14723;
  assign n64890 = pi19 ? n20563 : n64889;
  assign n64891 = pi18 ? n48120 : n64890;
  assign n64892 = pi17 ? n32 : n64891;
  assign n64893 = pi16 ? n32 : n64892;
  assign n64894 = pi15 ? n64886 : n64893;
  assign n64895 = pi22 ? n33792 : n893;
  assign n64896 = pi21 ? n30868 : n64895;
  assign n64897 = pi20 ? n64896 : n58944;
  assign n64898 = pi19 ? n20563 : n64897;
  assign n64899 = pi18 ? n48120 : n64898;
  assign n64900 = pi17 ? n32 : n64899;
  assign n64901 = pi16 ? n32 : n64900;
  assign n64902 = pi22 ? n33792 : n456;
  assign n64903 = pi21 ? n45016 : n64902;
  assign n64904 = pi20 ? n64903 : n1010;
  assign n64905 = pi19 ? n20563 : n64904;
  assign n64906 = pi18 ? n48120 : n64905;
  assign n64907 = pi17 ? n32 : n64906;
  assign n64908 = pi16 ? n32 : n64907;
  assign n64909 = pi15 ? n64901 : n64908;
  assign n64910 = pi14 ? n64894 : n64909;
  assign n64911 = pi13 ? n64880 : n64910;
  assign n64912 = pi22 ? n20563 : n3961;
  assign n64913 = pi21 ? n20563 : n64912;
  assign n64914 = pi20 ? n64913 : n21338;
  assign n64915 = pi19 ? n20563 : n64914;
  assign n64916 = pi18 ? n47592 : n64915;
  assign n64917 = pi17 ? n32 : n64916;
  assign n64918 = pi16 ? n32 : n64917;
  assign n64919 = pi22 ? n30868 : n11047;
  assign n64920 = pi21 ? n20563 : n64919;
  assign n64921 = pi20 ? n64920 : n17510;
  assign n64922 = pi19 ? n20563 : n64921;
  assign n64923 = pi18 ? n42206 : n64922;
  assign n64924 = pi17 ? n32 : n64923;
  assign n64925 = pi16 ? n32 : n64924;
  assign n64926 = pi15 ? n64918 : n64925;
  assign n64927 = pi23 ? n139 : n14626;
  assign n64928 = pi22 ? n30868 : n64927;
  assign n64929 = pi21 ? n20563 : n64928;
  assign n64930 = pi22 ? n14626 : n54520;
  assign n64931 = pi21 ? n64930 : n32;
  assign n64932 = pi20 ? n64929 : n64931;
  assign n64933 = pi19 ? n20563 : n64932;
  assign n64934 = pi18 ? n42206 : n64933;
  assign n64935 = pi17 ? n32 : n64934;
  assign n64936 = pi16 ? n32 : n64935;
  assign n64937 = pi22 ? n33792 : n3472;
  assign n64938 = pi21 ? n20563 : n64937;
  assign n64939 = pi20 ? n64938 : n61402;
  assign n64940 = pi19 ? n20563 : n64939;
  assign n64941 = pi18 ? n42699 : n64940;
  assign n64942 = pi17 ? n32 : n64941;
  assign n64943 = pi16 ? n32 : n64942;
  assign n64944 = pi15 ? n64936 : n64943;
  assign n64945 = pi14 ? n64926 : n64944;
  assign n64946 = pi22 ? n33792 : n60300;
  assign n64947 = pi21 ? n30868 : n64946;
  assign n64948 = pi20 ? n64947 : n54547;
  assign n64949 = pi19 ? n20563 : n64948;
  assign n64950 = pi18 ? n46997 : n64949;
  assign n64951 = pi17 ? n32 : n64950;
  assign n64952 = pi16 ? n32 : n64951;
  assign n64953 = pi22 ? n36659 : n2299;
  assign n64954 = pi21 ? n45016 : n64953;
  assign n64955 = pi20 ? n64954 : n55668;
  assign n64956 = pi19 ? n20563 : n64955;
  assign n64957 = pi18 ? n46997 : n64956;
  assign n64958 = pi17 ? n32 : n64957;
  assign n64959 = pi16 ? n32 : n64958;
  assign n64960 = pi15 ? n64952 : n64959;
  assign n64961 = pi22 ? n36659 : n14626;
  assign n64962 = pi21 ? n45016 : n64961;
  assign n64963 = pi23 ? n14626 : n624;
  assign n64964 = pi22 ? n64963 : n32;
  assign n64965 = pi21 ? n64964 : n32;
  assign n64966 = pi20 ? n64962 : n64965;
  assign n64967 = pi19 ? n20563 : n64966;
  assign n64968 = pi18 ? n46997 : n64967;
  assign n64969 = pi17 ? n32 : n64968;
  assign n64970 = pi16 ? n32 : n64969;
  assign n64971 = pi22 ? n52395 : n14626;
  assign n64972 = pi21 ? n40986 : n64971;
  assign n64973 = pi20 ? n64972 : n4116;
  assign n64974 = pi19 ? n20563 : n64973;
  assign n64975 = pi18 ? n46997 : n64974;
  assign n64976 = pi17 ? n32 : n64975;
  assign n64977 = pi16 ? n32 : n64976;
  assign n64978 = pi15 ? n64970 : n64977;
  assign n64979 = pi14 ? n64960 : n64978;
  assign n64980 = pi13 ? n64945 : n64979;
  assign n64981 = pi12 ? n64911 : n64980;
  assign n64982 = pi11 ? n64857 : n64981;
  assign n64983 = pi20 ? n64972 : n59674;
  assign n64984 = pi19 ? n40792 : n64983;
  assign n64985 = pi18 ? n46997 : n64984;
  assign n64986 = pi17 ? n32 : n64985;
  assign n64987 = pi16 ? n32 : n64986;
  assign n64988 = pi22 ? n37276 : n51564;
  assign n64989 = pi21 ? n45016 : n64988;
  assign n64990 = pi20 ? n64989 : n10011;
  assign n64991 = pi19 ? n40792 : n64990;
  assign n64992 = pi18 ? n46997 : n64991;
  assign n64993 = pi17 ? n32 : n64992;
  assign n64994 = pi16 ? n32 : n64993;
  assign n64995 = pi15 ? n64987 : n64994;
  assign n64996 = pi22 ? n50339 : n51564;
  assign n64997 = pi21 ? n40986 : n64996;
  assign n64998 = pi20 ? n64997 : n53984;
  assign n64999 = pi19 ? n59458 : n64998;
  assign n65000 = pi18 ? n40485 : n64999;
  assign n65001 = pi17 ? n32 : n65000;
  assign n65002 = pi16 ? n32 : n65001;
  assign n65003 = pi24 ? n20563 : n335;
  assign n65004 = pi23 ? n65003 : n335;
  assign n65005 = pi22 ? n20563 : n65004;
  assign n65006 = pi21 ? n65005 : n55597;
  assign n65007 = pi20 ? n65006 : n20953;
  assign n65008 = pi19 ? n20563 : n65007;
  assign n65009 = pi18 ? n41157 : n65008;
  assign n65010 = pi17 ? n32 : n65009;
  assign n65011 = pi16 ? n32 : n65010;
  assign n65012 = pi15 ? n65002 : n65011;
  assign n65013 = pi14 ? n64995 : n65012;
  assign n65014 = pi20 ? n42006 : n48184;
  assign n65015 = pi22 ? n63317 : n1388;
  assign n65016 = pi21 ? n63639 : n65015;
  assign n65017 = pi20 ? n65016 : n32;
  assign n65018 = pi19 ? n65014 : n65017;
  assign n65019 = pi18 ? n41157 : n65018;
  assign n65020 = pi17 ? n32 : n65019;
  assign n65021 = pi16 ? n32 : n65020;
  assign n65022 = pi21 ? n47220 : n30868;
  assign n65023 = pi20 ? n20563 : n65022;
  assign n65024 = pi22 ? n33792 : n64549;
  assign n65025 = pi22 ? n51564 : n759;
  assign n65026 = pi21 ? n65024 : n65025;
  assign n65027 = pi20 ? n65026 : n32;
  assign n65028 = pi19 ? n65023 : n65027;
  assign n65029 = pi18 ? n41157 : n65028;
  assign n65030 = pi17 ? n32 : n65029;
  assign n65031 = pi16 ? n32 : n65030;
  assign n65032 = pi15 ? n65021 : n65031;
  assign n65033 = pi20 ? n38754 : n51280;
  assign n65034 = pi19 ? n38377 : n65033;
  assign n65035 = pi21 ? n47220 : n33792;
  assign n65036 = pi20 ? n53326 : n65035;
  assign n65037 = pi22 ? n139 : n61844;
  assign n65038 = pi22 ? n51564 : n54563;
  assign n65039 = pi21 ? n65037 : n65038;
  assign n65040 = pi20 ? n65039 : n32;
  assign n65041 = pi19 ? n65036 : n65040;
  assign n65042 = pi18 ? n65034 : n65041;
  assign n65043 = pi17 ? n32 : n65042;
  assign n65044 = pi16 ? n32 : n65043;
  assign n65045 = pi20 ? n56630 : n51280;
  assign n65046 = pi19 ? n38377 : n65045;
  assign n65047 = pi21 ? n47360 : n33792;
  assign n65048 = pi20 ? n41578 : n65047;
  assign n65049 = pi23 ? n64587 : n204;
  assign n65050 = pi22 ? n36659 : n65049;
  assign n65051 = pi21 ? n65050 : n58470;
  assign n65052 = pi20 ? n65051 : n32;
  assign n65053 = pi19 ? n65048 : n65052;
  assign n65054 = pi18 ? n65046 : n65053;
  assign n65055 = pi17 ? n32 : n65054;
  assign n65056 = pi16 ? n32 : n65055;
  assign n65057 = pi15 ? n65044 : n65056;
  assign n65058 = pi14 ? n65032 : n65057;
  assign n65059 = pi13 ? n65013 : n65058;
  assign n65060 = pi20 ? n55020 : n54450;
  assign n65061 = pi19 ? n56687 : n65060;
  assign n65062 = pi20 ? n20563 : n47361;
  assign n65063 = pi24 ? n36659 : n204;
  assign n65064 = pi23 ? n65063 : n43198;
  assign n65065 = pi22 ? n36659 : n65064;
  assign n65066 = pi22 ? n56622 : n32;
  assign n65067 = pi21 ? n65065 : n65066;
  assign n65068 = pi20 ? n65067 : n32;
  assign n65069 = pi19 ? n65062 : n65068;
  assign n65070 = pi18 ? n65061 : n65069;
  assign n65071 = pi17 ? n32 : n65070;
  assign n65072 = pi16 ? n32 : n65071;
  assign n65073 = pi24 ? n36781 : n233;
  assign n65074 = pi23 ? n65073 : n233;
  assign n65075 = pi22 ? n36781 : n65074;
  assign n65076 = pi21 ? n65075 : n59342;
  assign n65077 = pi20 ? n65076 : n32;
  assign n65078 = pi19 ? n56631 : n65077;
  assign n65079 = pi18 ? n47056 : n65078;
  assign n65080 = pi17 ? n32 : n65079;
  assign n65081 = pi16 ? n32 : n65080;
  assign n65082 = pi15 ? n65072 : n65081;
  assign n65083 = pi23 ? n52672 : n32;
  assign n65084 = pi22 ? n65083 : n32;
  assign n65085 = pi21 ? n58999 : n65084;
  assign n65086 = pi20 ? n65085 : n32;
  assign n65087 = pi19 ? n63239 : n65086;
  assign n65088 = pi18 ? n47056 : n65087;
  assign n65089 = pi17 ? n32 : n65088;
  assign n65090 = pi16 ? n32 : n65089;
  assign n65091 = pi22 ? n36798 : n316;
  assign n65092 = pi21 ? n65091 : n59357;
  assign n65093 = pi20 ? n65092 : n32;
  assign n65094 = pi19 ? n63239 : n65093;
  assign n65095 = pi18 ? n41168 : n65094;
  assign n65096 = pi17 ? n32 : n65095;
  assign n65097 = pi16 ? n32 : n65096;
  assign n65098 = pi15 ? n65090 : n65097;
  assign n65099 = pi14 ? n65082 : n65098;
  assign n65100 = pi21 ? n20563 : n36798;
  assign n65101 = pi20 ? n20563 : n65100;
  assign n65102 = pi21 ? n57733 : n37639;
  assign n65103 = pi20 ? n65102 : n32;
  assign n65104 = pi19 ? n65101 : n65103;
  assign n65105 = pi18 ? n41168 : n65104;
  assign n65106 = pi17 ? n32 : n65105;
  assign n65107 = pi16 ? n32 : n65106;
  assign n65108 = pi21 ? n61251 : n32;
  assign n65109 = pi20 ? n65108 : n32;
  assign n65110 = pi19 ? n65101 : n65109;
  assign n65111 = pi18 ? n41168 : n65110;
  assign n65112 = pi17 ? n32 : n65111;
  assign n65113 = pi16 ? n32 : n65112;
  assign n65114 = pi15 ? n65107 : n65113;
  assign n65115 = pi22 ? n14626 : n625;
  assign n65116 = pi21 ? n65115 : n32;
  assign n65117 = pi20 ? n65116 : n32;
  assign n65118 = pi19 ? n65101 : n65117;
  assign n65119 = pi18 ? n41168 : n65118;
  assign n65120 = pi17 ? n32 : n65119;
  assign n65121 = pi16 ? n32 : n65120;
  assign n65122 = pi23 ? n20563 : n20627;
  assign n65123 = pi22 ? n37 : n65122;
  assign n65124 = pi21 ? n65123 : n59774;
  assign n65125 = pi20 ? n20563 : n65124;
  assign n65126 = pi21 ? n63010 : n32;
  assign n65127 = pi20 ? n65126 : n32;
  assign n65128 = pi19 ? n65125 : n65127;
  assign n65129 = pi18 ? n40023 : n65128;
  assign n65130 = pi17 ? n32 : n65129;
  assign n65131 = pi16 ? n32 : n65130;
  assign n65132 = pi15 ? n65121 : n65131;
  assign n65133 = pi14 ? n65114 : n65132;
  assign n65134 = pi13 ? n65099 : n65133;
  assign n65135 = pi12 ? n65059 : n65134;
  assign n65136 = pi19 ? n62374 : n60490;
  assign n65137 = pi23 ? n30868 : n3491;
  assign n65138 = pi22 ? n30868 : n65137;
  assign n65139 = pi21 ? n65138 : n55708;
  assign n65140 = pi20 ? n30868 : n65139;
  assign n65141 = pi19 ? n65140 : n64209;
  assign n65142 = pi18 ? n65136 : n65141;
  assign n65143 = pi17 ? n32 : n65142;
  assign n65144 = pi16 ? n32 : n65143;
  assign n65145 = pi21 ? n64224 : n39801;
  assign n65146 = pi20 ? n32 : n65145;
  assign n65147 = pi19 ? n65146 : n30868;
  assign n65148 = pi24 ? n33792 : n36798;
  assign n65149 = pi23 ? n65148 : n36798;
  assign n65150 = pi22 ? n65149 : n51564;
  assign n65151 = pi21 ? n33792 : n65150;
  assign n65152 = pi20 ? n30868 : n65151;
  assign n65153 = pi19 ? n65152 : n64209;
  assign n65154 = pi18 ? n65147 : n65153;
  assign n65155 = pi17 ? n32 : n65154;
  assign n65156 = pi16 ? n32 : n65155;
  assign n65157 = pi15 ? n65144 : n65156;
  assign n65158 = pi19 ? n62355 : n60490;
  assign n65159 = pi24 ? n36659 : n51564;
  assign n65160 = pi23 ? n65159 : n14626;
  assign n65161 = pi22 ? n65160 : n13481;
  assign n65162 = pi21 ? n64518 : n65161;
  assign n65163 = pi20 ? n30868 : n65162;
  assign n65164 = pi21 ? n59785 : n32;
  assign n65165 = pi20 ? n65164 : n32;
  assign n65166 = pi19 ? n65163 : n65165;
  assign n65167 = pi18 ? n65158 : n65166;
  assign n65168 = pi17 ? n32 : n65167;
  assign n65169 = pi16 ? n32 : n65168;
  assign n65170 = pi24 ? n36659 : n13481;
  assign n65171 = pi23 ? n65170 : n14626;
  assign n65172 = pi22 ? n65171 : n56186;
  assign n65173 = pi21 ? n42146 : n65172;
  assign n65174 = pi20 ? n30868 : n65173;
  assign n65175 = pi19 ? n65174 : n37641;
  assign n65176 = pi18 ? n59644 : n65175;
  assign n65177 = pi17 ? n32 : n65176;
  assign n65178 = pi16 ? n32 : n65177;
  assign n65179 = pi15 ? n65169 : n65178;
  assign n65180 = pi14 ? n65157 : n65179;
  assign n65181 = pi19 ? n37321 : n60490;
  assign n65182 = pi23 ? n65073 : n51564;
  assign n65183 = pi23 ? n13481 : n63008;
  assign n65184 = pi22 ? n65182 : n65183;
  assign n65185 = pi21 ? n40002 : n65184;
  assign n65186 = pi20 ? n56662 : n65185;
  assign n65187 = pi19 ? n65186 : n32;
  assign n65188 = pi18 ? n65181 : n65187;
  assign n65189 = pi17 ? n32 : n65188;
  assign n65190 = pi16 ? n32 : n65189;
  assign n65191 = pi23 ? n65073 : n14626;
  assign n65192 = pi22 ? n65191 : n59672;
  assign n65193 = pi21 ? n38901 : n65192;
  assign n65194 = pi20 ? n56662 : n65193;
  assign n65195 = pi19 ? n65194 : n32;
  assign n65196 = pi18 ? n65181 : n65195;
  assign n65197 = pi17 ? n32 : n65196;
  assign n65198 = pi16 ? n32 : n65197;
  assign n65199 = pi15 ? n65190 : n65198;
  assign n65200 = pi21 ? n32 : n36489;
  assign n65201 = pi20 ? n32 : n65200;
  assign n65202 = pi20 ? n42005 : n30868;
  assign n65203 = pi19 ? n65201 : n65202;
  assign n65204 = pi21 ? n30868 : n43198;
  assign n65205 = pi22 ? n43198 : n49412;
  assign n65206 = pi24 ? n36798 : n685;
  assign n65207 = pi23 ? n65206 : n51564;
  assign n65208 = pi22 ? n65207 : n59672;
  assign n65209 = pi21 ? n65205 : n65208;
  assign n65210 = pi20 ? n65204 : n65209;
  assign n65211 = pi19 ? n65210 : n32;
  assign n65212 = pi18 ? n65203 : n65211;
  assign n65213 = pi17 ? n32 : n65212;
  assign n65214 = pi16 ? n32 : n65213;
  assign n65215 = pi21 ? n32 : n47220;
  assign n65216 = pi20 ? n32 : n65215;
  assign n65217 = pi19 ? n65216 : n33792;
  assign n65218 = pi23 ? n61508 : n51564;
  assign n65219 = pi22 ? n65218 : n56665;
  assign n65220 = pi21 ? n56207 : n65219;
  assign n65221 = pi20 ? n55729 : n65220;
  assign n65222 = pi19 ? n65221 : n32;
  assign n65223 = pi18 ? n65217 : n65222;
  assign n65224 = pi17 ? n32 : n65223;
  assign n65225 = pi16 ? n32 : n65224;
  assign n65226 = pi15 ? n65214 : n65225;
  assign n65227 = pi14 ? n65199 : n65226;
  assign n65228 = pi13 ? n65180 : n65227;
  assign n65229 = pi19 ? n62446 : n33792;
  assign n65230 = pi24 ? n43198 : n316;
  assign n65231 = pi23 ? n65230 : n13481;
  assign n65232 = pi22 ? n65231 : n706;
  assign n65233 = pi21 ? n43198 : n65232;
  assign n65234 = pi20 ? n55729 : n65233;
  assign n65235 = pi19 ? n65234 : n32;
  assign n65236 = pi18 ? n65229 : n65235;
  assign n65237 = pi17 ? n32 : n65236;
  assign n65238 = pi16 ? n32 : n65237;
  assign n65239 = pi21 ? n61930 : n2678;
  assign n65240 = pi20 ? n55729 : n65239;
  assign n65241 = pi19 ? n65240 : n32;
  assign n65242 = pi18 ? n65229 : n65241;
  assign n65243 = pi17 ? n32 : n65242;
  assign n65244 = pi16 ? n32 : n65243;
  assign n65245 = pi15 ? n65238 : n65244;
  assign n65246 = pi19 ? n50811 : n59742;
  assign n65247 = pi22 ? n63009 : n32;
  assign n65248 = pi21 ? n51564 : n65247;
  assign n65249 = pi20 ? n43198 : n65248;
  assign n65250 = pi19 ? n65249 : n32;
  assign n65251 = pi18 ? n65246 : n65250;
  assign n65252 = pi17 ? n32 : n65251;
  assign n65253 = pi16 ? n32 : n65252;
  assign n65254 = pi22 ? n43198 : n38284;
  assign n65255 = pi21 ? n32 : n65254;
  assign n65256 = pi20 ? n32 : n65255;
  assign n65257 = pi19 ? n65256 : n43198;
  assign n65258 = pi18 ? n65257 : n64310;
  assign n65259 = pi17 ? n32 : n65258;
  assign n65260 = pi16 ? n32 : n65259;
  assign n65261 = pi15 ? n65253 : n65260;
  assign n65262 = pi14 ? n65245 : n65261;
  assign n65263 = pi22 ? n32 : n36781;
  assign n65264 = pi21 ? n32 : n65263;
  assign n65265 = pi20 ? n32 : n65264;
  assign n65266 = pi20 ? n52447 : n54009;
  assign n65267 = pi19 ? n65265 : n65266;
  assign n65268 = pi21 ? n63423 : n53983;
  assign n65269 = pi20 ? n46284 : n65268;
  assign n65270 = pi19 ? n65269 : n32;
  assign n65271 = pi18 ? n65267 : n65270;
  assign n65272 = pi17 ? n32 : n65271;
  assign n65273 = pi16 ? n32 : n65272;
  assign n65274 = pi22 ? n14626 : n49412;
  assign n65275 = pi21 ? n32 : n65274;
  assign n65276 = pi20 ? n32 : n65275;
  assign n65277 = pi19 ? n65276 : n14626;
  assign n65278 = pi20 ? n14626 : n64336;
  assign n65279 = pi19 ? n65278 : n32;
  assign n65280 = pi18 ? n65277 : n65279;
  assign n65281 = pi17 ? n32 : n65280;
  assign n65282 = pi16 ? n32 : n65281;
  assign n65283 = pi15 ? n65273 : n65282;
  assign n65284 = pi22 ? n32 : n53550;
  assign n65285 = pi21 ? n32 : n65284;
  assign n65286 = pi20 ? n32 : n65285;
  assign n65287 = pi21 ? n14626 : n58777;
  assign n65288 = pi20 ? n65287 : n14626;
  assign n65289 = pi19 ? n65286 : n65288;
  assign n65290 = pi18 ? n65289 : n63439;
  assign n65291 = pi17 ? n32 : n65290;
  assign n65292 = pi16 ? n32 : n65291;
  assign n65293 = pi20 ? n43198 : n14626;
  assign n65294 = pi19 ? n48858 : n65293;
  assign n65295 = pi20 ? n14626 : n64354;
  assign n65296 = pi19 ? n65295 : n32;
  assign n65297 = pi18 ? n65294 : n65296;
  assign n65298 = pi17 ? n32 : n65297;
  assign n65299 = pi16 ? n32 : n65298;
  assign n65300 = pi15 ? n65292 : n65299;
  assign n65301 = pi14 ? n65283 : n65300;
  assign n65302 = pi13 ? n65262 : n65301;
  assign n65303 = pi12 ? n65228 : n65302;
  assign n65304 = pi11 ? n65135 : n65303;
  assign n65305 = pi10 ? n64982 : n65304;
  assign n65306 = pi09 ? n64805 : n65305;
  assign n65307 = pi18 ? n40056 : n64789;
  assign n65308 = pi17 ? n32 : n65307;
  assign n65309 = pi16 ? n32 : n65308;
  assign n65310 = pi15 ? n32 : n65309;
  assign n65311 = pi18 ? n38999 : n62955;
  assign n65312 = pi17 ? n32 : n65311;
  assign n65313 = pi16 ? n32 : n65312;
  assign n65314 = pi18 ? n37322 : n62955;
  assign n65315 = pi17 ? n32 : n65314;
  assign n65316 = pi16 ? n32 : n65315;
  assign n65317 = pi15 ? n65313 : n65316;
  assign n65318 = pi14 ? n65310 : n65317;
  assign n65319 = pi13 ? n32 : n65318;
  assign n65320 = pi12 ? n32 : n65319;
  assign n65321 = pi11 ? n32 : n65320;
  assign n65322 = pi10 ? n32 : n65321;
  assign n65323 = pi18 ? n37335 : n62955;
  assign n65324 = pi17 ? n32 : n65323;
  assign n65325 = pi16 ? n32 : n65324;
  assign n65326 = pi18 ? n38378 : n62955;
  assign n65327 = pi17 ? n32 : n65326;
  assign n65328 = pi16 ? n32 : n65327;
  assign n65329 = pi15 ? n65325 : n65328;
  assign n65330 = pi18 ? n38378 : n62976;
  assign n65331 = pi17 ? n32 : n65330;
  assign n65332 = pi16 ? n32 : n65331;
  assign n65333 = pi18 ? n39455 : n62976;
  assign n65334 = pi17 ? n32 : n65333;
  assign n65335 = pi16 ? n32 : n65334;
  assign n65336 = pi15 ? n65332 : n65335;
  assign n65337 = pi14 ? n65329 : n65336;
  assign n65338 = pi15 ? n65335 : n64823;
  assign n65339 = pi18 ? n43222 : n62976;
  assign n65340 = pi17 ? n32 : n65339;
  assign n65341 = pi16 ? n32 : n65340;
  assign n65342 = pi15 ? n65341 : n64389;
  assign n65343 = pi14 ? n65338 : n65342;
  assign n65344 = pi13 ? n65337 : n65343;
  assign n65345 = pi14 ? n64389 : n63465;
  assign n65346 = pi18 ? n44273 : n59296;
  assign n65347 = pi17 ? n32 : n65346;
  assign n65348 = pi16 ? n32 : n65347;
  assign n65349 = pi18 ? n48623 : n59307;
  assign n65350 = pi17 ? n32 : n65349;
  assign n65351 = pi16 ? n32 : n65350;
  assign n65352 = pi15 ? n65348 : n65351;
  assign n65353 = pi24 ? n99 : n14626;
  assign n65354 = pi23 ? n65353 : n14626;
  assign n65355 = pi22 ? n65354 : n14626;
  assign n65356 = pi22 ? n14626 : n688;
  assign n65357 = pi21 ? n65355 : n65356;
  assign n65358 = pi20 ? n38754 : n65357;
  assign n65359 = pi19 ? n20563 : n65358;
  assign n65360 = pi18 ? n42644 : n65359;
  assign n65361 = pi17 ? n32 : n65360;
  assign n65362 = pi16 ? n32 : n65361;
  assign n65363 = pi18 ? n42644 : n64850;
  assign n65364 = pi17 ? n32 : n65363;
  assign n65365 = pi16 ? n32 : n65364;
  assign n65366 = pi15 ? n65362 : n65365;
  assign n65367 = pi14 ? n65352 : n65366;
  assign n65368 = pi13 ? n65345 : n65367;
  assign n65369 = pi12 ? n65344 : n65368;
  assign n65370 = pi18 ? n42644 : n64861;
  assign n65371 = pi17 ? n32 : n65370;
  assign n65372 = pi16 ? n32 : n65371;
  assign n65373 = pi18 ? n42654 : n64443;
  assign n65374 = pi17 ? n32 : n65373;
  assign n65375 = pi16 ? n32 : n65374;
  assign n65376 = pi15 ? n65372 : n65375;
  assign n65377 = pi18 ? n42654 : n64870;
  assign n65378 = pi17 ? n32 : n65377;
  assign n65379 = pi16 ? n32 : n65378;
  assign n65380 = pi18 ? n42680 : n64875;
  assign n65381 = pi17 ? n32 : n65380;
  assign n65382 = pi16 ? n32 : n65381;
  assign n65383 = pi15 ? n65379 : n65382;
  assign n65384 = pi14 ? n65376 : n65383;
  assign n65385 = pi18 ? n42680 : n64883;
  assign n65386 = pi17 ? n32 : n65385;
  assign n65387 = pi16 ? n32 : n65386;
  assign n65388 = pi18 ? n42193 : n64890;
  assign n65389 = pi17 ? n32 : n65388;
  assign n65390 = pi16 ? n32 : n65389;
  assign n65391 = pi15 ? n65387 : n65390;
  assign n65392 = pi18 ? n42193 : n64898;
  assign n65393 = pi17 ? n32 : n65392;
  assign n65394 = pi16 ? n32 : n65393;
  assign n65395 = pi18 ? n42193 : n64905;
  assign n65396 = pi17 ? n32 : n65395;
  assign n65397 = pi16 ? n32 : n65396;
  assign n65398 = pi15 ? n65394 : n65397;
  assign n65399 = pi14 ? n65391 : n65398;
  assign n65400 = pi13 ? n65384 : n65399;
  assign n65401 = pi23 ? n204 : n63008;
  assign n65402 = pi22 ? n204 : n65401;
  assign n65403 = pi21 ? n65402 : n32;
  assign n65404 = pi20 ? n64913 : n65403;
  assign n65405 = pi19 ? n20563 : n65404;
  assign n65406 = pi18 ? n43254 : n65405;
  assign n65407 = pi17 ? n32 : n65406;
  assign n65408 = pi16 ? n32 : n65407;
  assign n65409 = pi18 ? n43254 : n64922;
  assign n65410 = pi17 ? n32 : n65409;
  assign n65411 = pi16 ? n32 : n65410;
  assign n65412 = pi15 ? n65408 : n65411;
  assign n65413 = pi18 ? n42200 : n64933;
  assign n65414 = pi17 ? n32 : n65413;
  assign n65415 = pi16 ? n32 : n65414;
  assign n65416 = pi18 ? n42200 : n64940;
  assign n65417 = pi17 ? n32 : n65416;
  assign n65418 = pi16 ? n32 : n65417;
  assign n65419 = pi15 ? n65415 : n65418;
  assign n65420 = pi14 ? n65412 : n65419;
  assign n65421 = pi22 ? n33792 : n63328;
  assign n65422 = pi21 ? n30868 : n65421;
  assign n65423 = pi20 ? n65422 : n54547;
  assign n65424 = pi19 ? n20563 : n65423;
  assign n65425 = pi18 ? n43261 : n65424;
  assign n65426 = pi17 ? n32 : n65425;
  assign n65427 = pi16 ? n32 : n65426;
  assign n65428 = pi18 ? n43261 : n64956;
  assign n65429 = pi17 ? n32 : n65428;
  assign n65430 = pi16 ? n32 : n65429;
  assign n65431 = pi15 ? n65427 : n65430;
  assign n65432 = pi23 ? n14626 : n63008;
  assign n65433 = pi22 ? n65432 : n32;
  assign n65434 = pi21 ? n65433 : n32;
  assign n65435 = pi20 ? n64962 : n65434;
  assign n65436 = pi19 ? n20563 : n65435;
  assign n65437 = pi18 ? n43261 : n65436;
  assign n65438 = pi17 ? n32 : n65437;
  assign n65439 = pi16 ? n32 : n65438;
  assign n65440 = pi18 ? n43261 : n64974;
  assign n65441 = pi17 ? n32 : n65440;
  assign n65442 = pi16 ? n32 : n65441;
  assign n65443 = pi15 ? n65439 : n65442;
  assign n65444 = pi14 ? n65431 : n65443;
  assign n65445 = pi13 ? n65420 : n65444;
  assign n65446 = pi12 ? n65400 : n65445;
  assign n65447 = pi11 ? n65369 : n65446;
  assign n65448 = pi18 ? n48120 : n64984;
  assign n65449 = pi17 ? n32 : n65448;
  assign n65450 = pi16 ? n32 : n65449;
  assign n65451 = pi18 ? n48120 : n64991;
  assign n65452 = pi17 ? n32 : n65451;
  assign n65453 = pi16 ? n32 : n65452;
  assign n65454 = pi15 ? n65450 : n65453;
  assign n65455 = pi18 ? n42687 : n64999;
  assign n65456 = pi17 ? n32 : n65455;
  assign n65457 = pi16 ? n32 : n65456;
  assign n65458 = pi22 ? n43579 : n335;
  assign n65459 = pi21 ? n65458 : n55597;
  assign n65460 = pi20 ? n65459 : n20953;
  assign n65461 = pi19 ? n20563 : n65460;
  assign n65462 = pi18 ? n41641 : n65461;
  assign n65463 = pi17 ? n32 : n65462;
  assign n65464 = pi16 ? n32 : n65463;
  assign n65465 = pi15 ? n65457 : n65464;
  assign n65466 = pi14 ? n65454 : n65465;
  assign n65467 = pi24 ? n30868 : n363;
  assign n65468 = pi23 ? n65467 : n363;
  assign n65469 = pi22 ? n30868 : n65468;
  assign n65470 = pi23 ? n233 : n63008;
  assign n65471 = pi22 ? n63317 : n65470;
  assign n65472 = pi21 ? n65469 : n65471;
  assign n65473 = pi20 ? n65472 : n32;
  assign n65474 = pi19 ? n65014 : n65473;
  assign n65475 = pi18 ? n41641 : n65474;
  assign n65476 = pi17 ? n32 : n65475;
  assign n65477 = pi16 ? n32 : n65476;
  assign n65478 = pi22 ? n51564 : n54520;
  assign n65479 = pi21 ? n65024 : n65478;
  assign n65480 = pi20 ? n65479 : n32;
  assign n65481 = pi19 ? n65023 : n65480;
  assign n65482 = pi18 ? n41641 : n65481;
  assign n65483 = pi17 ? n32 : n65482;
  assign n65484 = pi16 ? n32 : n65483;
  assign n65485 = pi15 ? n65477 : n65484;
  assign n65486 = pi19 ? n37956 : n65033;
  assign n65487 = pi22 ? n139 : n65149;
  assign n65488 = pi21 ? n65487 : n65038;
  assign n65489 = pi20 ? n65488 : n32;
  assign n65490 = pi19 ? n65036 : n65489;
  assign n65491 = pi18 ? n65486 : n65490;
  assign n65492 = pi17 ? n32 : n65491;
  assign n65493 = pi16 ? n32 : n65492;
  assign n65494 = pi19 ? n37956 : n65045;
  assign n65495 = pi18 ? n65494 : n65053;
  assign n65496 = pi17 ? n32 : n65495;
  assign n65497 = pi16 ? n32 : n65496;
  assign n65498 = pi15 ? n65493 : n65497;
  assign n65499 = pi14 ? n65485 : n65498;
  assign n65500 = pi13 ? n65466 : n65499;
  assign n65501 = pi22 ? n45597 : n56111;
  assign n65502 = pi21 ? n32 : n65501;
  assign n65503 = pi20 ? n32 : n65502;
  assign n65504 = pi20 ? n55020 : n54155;
  assign n65505 = pi19 ? n65503 : n65504;
  assign n65506 = pi23 ? n64129 : n43198;
  assign n65507 = pi22 ? n36659 : n65506;
  assign n65508 = pi21 ? n65507 : n65066;
  assign n65509 = pi20 ? n65508 : n32;
  assign n65510 = pi19 ? n65062 : n65509;
  assign n65511 = pi18 ? n65505 : n65510;
  assign n65512 = pi17 ? n32 : n65511;
  assign n65513 = pi16 ? n32 : n65512;
  assign n65514 = pi18 ? n42699 : n65078;
  assign n65515 = pi17 ? n32 : n65514;
  assign n65516 = pi16 ? n32 : n65515;
  assign n65517 = pi15 ? n65513 : n65516;
  assign n65518 = pi18 ? n42699 : n65087;
  assign n65519 = pi17 ? n32 : n65518;
  assign n65520 = pi16 ? n32 : n65519;
  assign n65521 = pi18 ? n42699 : n65094;
  assign n65522 = pi17 ? n32 : n65521;
  assign n65523 = pi16 ? n32 : n65522;
  assign n65524 = pi15 ? n65520 : n65523;
  assign n65525 = pi14 ? n65517 : n65524;
  assign n65526 = pi18 ? n42699 : n65104;
  assign n65527 = pi17 ? n32 : n65526;
  assign n65528 = pi16 ? n32 : n65527;
  assign n65529 = pi18 ? n42699 : n65110;
  assign n65530 = pi17 ? n32 : n65529;
  assign n65531 = pi16 ? n32 : n65530;
  assign n65532 = pi15 ? n65528 : n65531;
  assign n65533 = pi22 ? n20563 : n63260;
  assign n65534 = pi21 ? n65533 : n36798;
  assign n65535 = pi20 ? n20563 : n65534;
  assign n65536 = pi19 ? n65535 : n65117;
  assign n65537 = pi18 ? n42699 : n65536;
  assign n65538 = pi17 ? n32 : n65537;
  assign n65539 = pi16 ? n32 : n65538;
  assign n65540 = pi23 ? n37 : n56987;
  assign n65541 = pi22 ? n65540 : n37809;
  assign n65542 = pi21 ? n65541 : n59774;
  assign n65543 = pi20 ? n20563 : n65542;
  assign n65544 = pi22 ? n64606 : n688;
  assign n65545 = pi21 ? n65544 : n32;
  assign n65546 = pi20 ? n65545 : n32;
  assign n65547 = pi19 ? n65543 : n65546;
  assign n65548 = pi18 ? n46997 : n65547;
  assign n65549 = pi17 ? n32 : n65548;
  assign n65550 = pi16 ? n32 : n65549;
  assign n65551 = pi15 ? n65539 : n65550;
  assign n65552 = pi14 ? n65532 : n65551;
  assign n65553 = pi13 ? n65525 : n65552;
  assign n65554 = pi12 ? n65500 : n65553;
  assign n65555 = pi19 ? n48790 : n60490;
  assign n65556 = pi21 ? n64663 : n55708;
  assign n65557 = pi20 ? n30868 : n65556;
  assign n65558 = pi19 ? n65557 : n64209;
  assign n65559 = pi18 ? n65555 : n65558;
  assign n65560 = pi17 ? n32 : n65559;
  assign n65561 = pi16 ? n32 : n65560;
  assign n65562 = pi19 ? n60024 : n30868;
  assign n65563 = pi22 ? n52451 : n51564;
  assign n65564 = pi21 ? n33792 : n65563;
  assign n65565 = pi20 ? n30868 : n65564;
  assign n65566 = pi21 ? n58778 : n32;
  assign n65567 = pi20 ? n65566 : n32;
  assign n65568 = pi19 ? n65565 : n65567;
  assign n65569 = pi18 ? n65562 : n65568;
  assign n65570 = pi17 ? n32 : n65569;
  assign n65571 = pi16 ? n32 : n65570;
  assign n65572 = pi15 ? n65561 : n65571;
  assign n65573 = pi19 ? n60024 : n60490;
  assign n65574 = pi22 ? n53930 : n13481;
  assign n65575 = pi21 ? n64518 : n65574;
  assign n65576 = pi20 ? n30868 : n65575;
  assign n65577 = pi19 ? n65576 : n10012;
  assign n65578 = pi18 ? n65573 : n65577;
  assign n65579 = pi17 ? n32 : n65578;
  assign n65580 = pi16 ? n32 : n65579;
  assign n65581 = pi19 ? n37934 : n30868;
  assign n65582 = pi23 ? n65063 : n14626;
  assign n65583 = pi23 ? n51564 : n63008;
  assign n65584 = pi22 ? n65582 : n65583;
  assign n65585 = pi21 ? n42146 : n65584;
  assign n65586 = pi20 ? n30868 : n65585;
  assign n65587 = pi19 ? n65586 : n32;
  assign n65588 = pi18 ? n65581 : n65587;
  assign n65589 = pi17 ? n32 : n65588;
  assign n65590 = pi16 ? n32 : n65589;
  assign n65591 = pi15 ? n65580 : n65590;
  assign n65592 = pi14 ? n65572 : n65591;
  assign n65593 = pi19 ? n37934 : n60490;
  assign n65594 = pi22 ? n57197 : n65183;
  assign n65595 = pi21 ? n40002 : n65594;
  assign n65596 = pi20 ? n56662 : n65595;
  assign n65597 = pi19 ? n65596 : n32;
  assign n65598 = pi18 ? n65593 : n65597;
  assign n65599 = pi17 ? n32 : n65598;
  assign n65600 = pi16 ? n32 : n65599;
  assign n65601 = pi24 ? n14626 : n685;
  assign n65602 = pi23 ? n65601 : n51565;
  assign n65603 = pi22 ? n64140 : n65602;
  assign n65604 = pi21 ? n38901 : n65603;
  assign n65605 = pi20 ? n56662 : n65604;
  assign n65606 = pi19 ? n65605 : n32;
  assign n65607 = pi18 ? n65593 : n65606;
  assign n65608 = pi17 ? n32 : n65607;
  assign n65609 = pi16 ? n32 : n65608;
  assign n65610 = pi15 ? n65600 : n65609;
  assign n65611 = pi19 ? n46062 : n65202;
  assign n65612 = pi21 ? n65205 : n64706;
  assign n65613 = pi20 ? n65204 : n65612;
  assign n65614 = pi19 ? n65613 : n32;
  assign n65615 = pi18 ? n65611 : n65614;
  assign n65616 = pi17 ? n32 : n65615;
  assign n65617 = pi16 ? n32 : n65616;
  assign n65618 = pi19 ? n54445 : n33792;
  assign n65619 = pi21 ? n56207 : n62849;
  assign n65620 = pi20 ? n55729 : n65619;
  assign n65621 = pi19 ? n65620 : n32;
  assign n65622 = pi18 ? n65618 : n65621;
  assign n65623 = pi17 ? n32 : n65622;
  assign n65624 = pi16 ? n32 : n65623;
  assign n65625 = pi15 ? n65617 : n65624;
  assign n65626 = pi14 ? n65610 : n65625;
  assign n65627 = pi13 ? n65592 : n65626;
  assign n65628 = pi21 ? n43198 : n56129;
  assign n65629 = pi20 ? n55729 : n65628;
  assign n65630 = pi19 ? n65629 : n32;
  assign n65631 = pi18 ? n65618 : n65630;
  assign n65632 = pi17 ? n32 : n65631;
  assign n65633 = pi16 ? n32 : n65632;
  assign n65634 = pi18 ? n65618 : n65241;
  assign n65635 = pi17 ? n32 : n65634;
  assign n65636 = pi16 ? n32 : n65635;
  assign n65637 = pi15 ? n65633 : n65636;
  assign n65638 = pi19 ? n48858 : n59742;
  assign n65639 = pi18 ? n65638 : n63417;
  assign n65640 = pi17 ? n32 : n65639;
  assign n65641 = pi16 ? n32 : n65640;
  assign n65642 = pi19 ? n32 : n43198;
  assign n65643 = pi18 ? n65642 : n64749;
  assign n65644 = pi17 ? n32 : n65643;
  assign n65645 = pi16 ? n32 : n65644;
  assign n65646 = pi15 ? n65641 : n65645;
  assign n65647 = pi14 ? n65637 : n65646;
  assign n65648 = pi19 ? n32 : n65266;
  assign n65649 = pi20 ? n46284 : n63424;
  assign n65650 = pi19 ? n65649 : n32;
  assign n65651 = pi18 ? n65648 : n65650;
  assign n65652 = pi17 ? n32 : n65651;
  assign n65653 = pi16 ? n32 : n65652;
  assign n65654 = pi19 ? n32 : n14626;
  assign n65655 = pi18 ? n65654 : n63439;
  assign n65656 = pi17 ? n32 : n65655;
  assign n65657 = pi16 ? n32 : n65656;
  assign n65658 = pi15 ? n65653 : n65657;
  assign n65659 = pi19 ? n32 : n65288;
  assign n65660 = pi20 ? n14626 : n60045;
  assign n65661 = pi19 ? n65660 : n32;
  assign n65662 = pi18 ? n65659 : n65661;
  assign n65663 = pi17 ? n32 : n65662;
  assign n65664 = pi16 ? n32 : n65663;
  assign n65665 = pi19 ? n32 : n65293;
  assign n65666 = pi21 ? n59342 : n32;
  assign n65667 = pi20 ? n14626 : n65666;
  assign n65668 = pi19 ? n65667 : n32;
  assign n65669 = pi18 ? n65665 : n65668;
  assign n65670 = pi17 ? n32 : n65669;
  assign n65671 = pi16 ? n32 : n65670;
  assign n65672 = pi15 ? n65664 : n65671;
  assign n65673 = pi14 ? n65658 : n65672;
  assign n65674 = pi13 ? n65647 : n65673;
  assign n65675 = pi12 ? n65627 : n65674;
  assign n65676 = pi11 ? n65554 : n65675;
  assign n65677 = pi10 ? n65447 : n65676;
  assign n65678 = pi09 ? n65322 : n65677;
  assign n65679 = pi08 ? n65306 : n65678;
  assign n65680 = pi19 ? n38315 : n64788;
  assign n65681 = pi18 ? n32 : n65680;
  assign n65682 = pi17 ? n32 : n65681;
  assign n65683 = pi16 ? n32 : n65682;
  assign n65684 = pi15 ? n32 : n65683;
  assign n65685 = pi18 ? n40056 : n62955;
  assign n65686 = pi17 ? n32 : n65685;
  assign n65687 = pi16 ? n32 : n65686;
  assign n65688 = pi18 ? n37935 : n62955;
  assign n65689 = pi17 ? n32 : n65688;
  assign n65690 = pi16 ? n32 : n65689;
  assign n65691 = pi15 ? n65687 : n65690;
  assign n65692 = pi14 ? n65684 : n65691;
  assign n65693 = pi13 ? n32 : n65692;
  assign n65694 = pi12 ? n32 : n65693;
  assign n65695 = pi11 ? n32 : n65694;
  assign n65696 = pi10 ? n32 : n65695;
  assign n65697 = pi18 ? n37957 : n62955;
  assign n65698 = pi17 ? n32 : n65697;
  assign n65699 = pi16 ? n32 : n65698;
  assign n65700 = pi15 ? n65690 : n65699;
  assign n65701 = pi18 ? n37957 : n62976;
  assign n65702 = pi17 ? n32 : n65701;
  assign n65703 = pi16 ? n32 : n65702;
  assign n65704 = pi18 ? n38999 : n62976;
  assign n65705 = pi17 ? n32 : n65704;
  assign n65706 = pi16 ? n32 : n65705;
  assign n65707 = pi15 ? n65703 : n65706;
  assign n65708 = pi14 ? n65700 : n65707;
  assign n65709 = pi18 ? n28159 : n62976;
  assign n65710 = pi17 ? n32 : n65709;
  assign n65711 = pi16 ? n32 : n65710;
  assign n65712 = pi15 ? n65706 : n65711;
  assign n65713 = pi18 ? n30119 : n62976;
  assign n65714 = pi17 ? n32 : n65713;
  assign n65715 = pi16 ? n32 : n65714;
  assign n65716 = pi15 ? n65715 : n64815;
  assign n65717 = pi14 ? n65712 : n65716;
  assign n65718 = pi13 ? n65708 : n65717;
  assign n65719 = pi18 ? n31315 : n62955;
  assign n65720 = pi17 ? n32 : n65719;
  assign n65721 = pi16 ? n32 : n65720;
  assign n65722 = pi14 ? n64815 : n65721;
  assign n65723 = pi18 ? n44246 : n59296;
  assign n65724 = pi17 ? n32 : n65723;
  assign n65725 = pi16 ? n32 : n65724;
  assign n65726 = pi18 ? n43222 : n59307;
  assign n65727 = pi17 ? n32 : n65726;
  assign n65728 = pi16 ? n32 : n65727;
  assign n65729 = pi15 ? n65725 : n65728;
  assign n65730 = pi18 ? n43226 : n65359;
  assign n65731 = pi17 ? n32 : n65730;
  assign n65732 = pi16 ? n32 : n65731;
  assign n65733 = pi18 ? n43226 : n64850;
  assign n65734 = pi17 ? n32 : n65733;
  assign n65735 = pi16 ? n32 : n65734;
  assign n65736 = pi15 ? n65732 : n65735;
  assign n65737 = pi14 ? n65729 : n65736;
  assign n65738 = pi13 ? n65722 : n65737;
  assign n65739 = pi12 ? n65718 : n65738;
  assign n65740 = pi22 ? n20563 : n37218;
  assign n65741 = pi21 ? n20563 : n65740;
  assign n65742 = pi20 ? n65741 : n64441;
  assign n65743 = pi19 ? n20563 : n65742;
  assign n65744 = pi18 ? n43226 : n65743;
  assign n65745 = pi17 ? n32 : n65744;
  assign n65746 = pi16 ? n32 : n65745;
  assign n65747 = pi18 ? n43247 : n65743;
  assign n65748 = pi17 ? n32 : n65747;
  assign n65749 = pi16 ? n32 : n65748;
  assign n65750 = pi15 ? n65746 : n65749;
  assign n65751 = pi23 ? n20563 : n335;
  assign n65752 = pi22 ? n20563 : n65751;
  assign n65753 = pi21 ? n20563 : n65752;
  assign n65754 = pi20 ? n65753 : n59343;
  assign n65755 = pi19 ? n20563 : n65754;
  assign n65756 = pi18 ? n43247 : n65755;
  assign n65757 = pi17 ? n32 : n65756;
  assign n65758 = pi16 ? n32 : n65757;
  assign n65759 = pi22 ? n20563 : n37783;
  assign n65760 = pi21 ? n20563 : n65759;
  assign n65761 = pi20 ? n65760 : n23203;
  assign n65762 = pi19 ? n20563 : n65761;
  assign n65763 = pi18 ? n44273 : n65762;
  assign n65764 = pi17 ? n32 : n65763;
  assign n65765 = pi16 ? n32 : n65764;
  assign n65766 = pi15 ? n65758 : n65765;
  assign n65767 = pi14 ? n65750 : n65766;
  assign n65768 = pi22 ? n30868 : n57380;
  assign n65769 = pi21 ? n20563 : n65768;
  assign n65770 = pi20 ? n65769 : n14723;
  assign n65771 = pi19 ? n20563 : n65770;
  assign n65772 = pi18 ? n44273 : n65771;
  assign n65773 = pi17 ? n32 : n65772;
  assign n65774 = pi16 ? n32 : n65773;
  assign n65775 = pi23 ? n20563 : n157;
  assign n65776 = pi22 ? n30868 : n65775;
  assign n65777 = pi21 ? n20563 : n65776;
  assign n65778 = pi20 ? n65777 : n14723;
  assign n65779 = pi19 ? n20563 : n65778;
  assign n65780 = pi18 ? n48623 : n65779;
  assign n65781 = pi17 ? n32 : n65780;
  assign n65782 = pi16 ? n32 : n65781;
  assign n65783 = pi15 ? n65774 : n65782;
  assign n65784 = pi22 ? n33792 : n65775;
  assign n65785 = pi21 ? n30868 : n65784;
  assign n65786 = pi20 ? n65785 : n1010;
  assign n65787 = pi19 ? n20563 : n65786;
  assign n65788 = pi18 ? n48623 : n65787;
  assign n65789 = pi17 ? n32 : n65788;
  assign n65790 = pi16 ? n32 : n65789;
  assign n65791 = pi23 ? n20563 : n204;
  assign n65792 = pi22 ? n33792 : n65791;
  assign n65793 = pi21 ? n45016 : n65792;
  assign n65794 = pi20 ? n65793 : n1010;
  assign n65795 = pi19 ? n20563 : n65794;
  assign n65796 = pi18 ? n48623 : n65795;
  assign n65797 = pi17 ? n32 : n65796;
  assign n65798 = pi16 ? n32 : n65797;
  assign n65799 = pi15 ? n65790 : n65798;
  assign n65800 = pi14 ? n65783 : n65799;
  assign n65801 = pi13 ? n65767 : n65800;
  assign n65802 = pi23 ? n30868 : n204;
  assign n65803 = pi22 ? n20563 : n65802;
  assign n65804 = pi21 ? n20563 : n65803;
  assign n65805 = pi20 ? n65804 : n65403;
  assign n65806 = pi19 ? n20563 : n65805;
  assign n65807 = pi18 ? n42644 : n65806;
  assign n65808 = pi17 ? n32 : n65807;
  assign n65809 = pi16 ? n32 : n65808;
  assign n65810 = pi22 ? n30868 : n63091;
  assign n65811 = pi21 ? n20563 : n65810;
  assign n65812 = pi20 ? n65811 : n17510;
  assign n65813 = pi19 ? n20563 : n65812;
  assign n65814 = pi18 ? n42644 : n65813;
  assign n65815 = pi17 ? n32 : n65814;
  assign n65816 = pi16 ? n32 : n65815;
  assign n65817 = pi15 ? n65809 : n65816;
  assign n65818 = pi23 ? n33792 : n14626;
  assign n65819 = pi22 ? n30868 : n65818;
  assign n65820 = pi21 ? n20563 : n65819;
  assign n65821 = pi21 ? n63197 : n32;
  assign n65822 = pi20 ? n65820 : n65821;
  assign n65823 = pi19 ? n20563 : n65822;
  assign n65824 = pi18 ? n42654 : n65823;
  assign n65825 = pi17 ? n32 : n65824;
  assign n65826 = pi16 ? n32 : n65825;
  assign n65827 = pi23 ? n139 : n51564;
  assign n65828 = pi22 ? n33792 : n65827;
  assign n65829 = pi21 ? n20563 : n65828;
  assign n65830 = pi22 ? n51564 : n19696;
  assign n65831 = pi21 ? n65830 : n32;
  assign n65832 = pi20 ? n65829 : n65831;
  assign n65833 = pi19 ? n20563 : n65832;
  assign n65834 = pi18 ? n42654 : n65833;
  assign n65835 = pi17 ? n32 : n65834;
  assign n65836 = pi16 ? n32 : n65835;
  assign n65837 = pi15 ? n65826 : n65836;
  assign n65838 = pi14 ? n65817 : n65837;
  assign n65839 = pi21 ? n30868 : n61192;
  assign n65840 = pi20 ? n65839 : n4008;
  assign n65841 = pi19 ? n20563 : n65840;
  assign n65842 = pi18 ? n42680 : n65841;
  assign n65843 = pi17 ? n32 : n65842;
  assign n65844 = pi16 ? n32 : n65843;
  assign n65845 = pi21 ? n45016 : n63130;
  assign n65846 = pi20 ? n65845 : n55668;
  assign n65847 = pi19 ? n20563 : n65846;
  assign n65848 = pi18 ? n42680 : n65847;
  assign n65849 = pi17 ? n32 : n65848;
  assign n65850 = pi16 ? n32 : n65849;
  assign n65851 = pi15 ? n65844 : n65850;
  assign n65852 = pi18 ? n42680 : n65436;
  assign n65853 = pi17 ? n32 : n65852;
  assign n65854 = pi16 ? n32 : n65853;
  assign n65855 = pi23 ? n139 : n61843;
  assign n65856 = pi22 ? n65855 : n14626;
  assign n65857 = pi21 ? n40986 : n65856;
  assign n65858 = pi20 ? n65857 : n4116;
  assign n65859 = pi19 ? n20563 : n65858;
  assign n65860 = pi18 ? n42680 : n65859;
  assign n65861 = pi17 ? n32 : n65860;
  assign n65862 = pi16 ? n32 : n65861;
  assign n65863 = pi15 ? n65854 : n65862;
  assign n65864 = pi14 ? n65851 : n65863;
  assign n65865 = pi13 ? n65838 : n65864;
  assign n65866 = pi12 ? n65801 : n65865;
  assign n65867 = pi11 ? n65739 : n65866;
  assign n65868 = pi23 ? n139 : n64110;
  assign n65869 = pi22 ? n65868 : n62803;
  assign n65870 = pi21 ? n40986 : n65869;
  assign n65871 = pi20 ? n65870 : n51568;
  assign n65872 = pi19 ? n40792 : n65871;
  assign n65873 = pi18 ? n42680 : n65872;
  assign n65874 = pi17 ? n32 : n65873;
  assign n65875 = pi16 ? n32 : n65874;
  assign n65876 = pi23 ? n335 : n64110;
  assign n65877 = pi22 ? n65876 : n62473;
  assign n65878 = pi21 ? n45016 : n65877;
  assign n65879 = pi20 ? n65878 : n10011;
  assign n65880 = pi19 ? n40792 : n65879;
  assign n65881 = pi18 ? n42193 : n65880;
  assign n65882 = pi17 ? n32 : n65881;
  assign n65883 = pi16 ? n32 : n65882;
  assign n65884 = pi15 ? n65875 : n65883;
  assign n65885 = pi24 ? n51564 : n43198;
  assign n65886 = pi23 ? n36659 : n65885;
  assign n65887 = pi22 ? n65886 : n56186;
  assign n65888 = pi21 ? n40986 : n65887;
  assign n65889 = pi20 ? n65888 : n53984;
  assign n65890 = pi19 ? n59458 : n65889;
  assign n65891 = pi18 ? n42193 : n65890;
  assign n65892 = pi17 ? n32 : n65891;
  assign n65893 = pi16 ? n32 : n65892;
  assign n65894 = pi22 ? n14626 : n65432;
  assign n65895 = pi21 ? n55685 : n65894;
  assign n65896 = pi20 ? n65895 : n32;
  assign n65897 = pi19 ? n54543 : n65896;
  assign n65898 = pi18 ? n43254 : n65897;
  assign n65899 = pi17 ? n32 : n65898;
  assign n65900 = pi16 ? n32 : n65899;
  assign n65901 = pi15 ? n65893 : n65900;
  assign n65902 = pi14 ? n65884 : n65901;
  assign n65903 = pi22 ? n37173 : n30868;
  assign n65904 = pi21 ? n65903 : n20563;
  assign n65905 = pi20 ? n65904 : n48184;
  assign n65906 = pi21 ? n51313 : n65894;
  assign n65907 = pi20 ? n65906 : n32;
  assign n65908 = pi19 ? n65905 : n65907;
  assign n65909 = pi18 ? n43254 : n65908;
  assign n65910 = pi17 ? n32 : n65909;
  assign n65911 = pi16 ? n32 : n65910;
  assign n65912 = pi21 ? n30155 : n40960;
  assign n65913 = pi20 ? n65912 : n20563;
  assign n65914 = pi19 ? n32 : n65913;
  assign n65915 = pi21 ? n54446 : n20563;
  assign n65916 = pi21 ? n45016 : n30868;
  assign n65917 = pi20 ? n65915 : n65916;
  assign n65918 = pi23 ? n3145 : n157;
  assign n65919 = pi22 ? n33792 : n65918;
  assign n65920 = pi21 ? n65919 : n64706;
  assign n65921 = pi20 ? n65920 : n32;
  assign n65922 = pi19 ? n65917 : n65921;
  assign n65923 = pi18 ? n65914 : n65922;
  assign n65924 = pi17 ? n32 : n65923;
  assign n65925 = pi16 ? n32 : n65924;
  assign n65926 = pi15 ? n65911 : n65925;
  assign n65927 = pi22 ? n20563 : n43571;
  assign n65928 = pi21 ? n30155 : n65927;
  assign n65929 = pi20 ? n65928 : n51280;
  assign n65930 = pi19 ? n32 : n65929;
  assign n65931 = pi21 ? n51762 : n33792;
  assign n65932 = pi20 ? n65931 : n65035;
  assign n65933 = pi23 ? n64570 : n204;
  assign n65934 = pi22 ? n33792 : n65933;
  assign n65935 = pi23 ? n204 : n51564;
  assign n65936 = pi22 ? n65935 : n55688;
  assign n65937 = pi21 ? n65934 : n65936;
  assign n65938 = pi20 ? n65937 : n32;
  assign n65939 = pi19 ? n65932 : n65938;
  assign n65940 = pi18 ? n65930 : n65939;
  assign n65941 = pi17 ? n32 : n65940;
  assign n65942 = pi16 ? n32 : n65941;
  assign n65943 = pi21 ? n45092 : n36659;
  assign n65944 = pi20 ? n65943 : n51280;
  assign n65945 = pi19 ? n51757 : n65944;
  assign n65946 = pi23 ? n233 : n51564;
  assign n65947 = pi22 ? n65946 : n14363;
  assign n65948 = pi21 ? n65050 : n65947;
  assign n65949 = pi20 ? n65948 : n32;
  assign n65950 = pi19 ? n65048 : n65949;
  assign n65951 = pi18 ? n65945 : n65950;
  assign n65952 = pi17 ? n32 : n65951;
  assign n65953 = pi16 ? n32 : n65952;
  assign n65954 = pi15 ? n65942 : n65953;
  assign n65955 = pi14 ? n65926 : n65954;
  assign n65956 = pi13 ? n65902 : n65955;
  assign n65957 = pi23 ? n36781 : n20563;
  assign n65958 = pi22 ? n55502 : n65957;
  assign n65959 = pi21 ? n30866 : n65958;
  assign n65960 = pi20 ? n65959 : n38754;
  assign n65961 = pi19 ? n32 : n65960;
  assign n65962 = pi22 ? n30869 : n20563;
  assign n65963 = pi21 ? n20563 : n65962;
  assign n65964 = pi20 ? n65963 : n47361;
  assign n65965 = pi24 ? n363 : n43198;
  assign n65966 = pi23 ? n65965 : n233;
  assign n65967 = pi22 ? n36659 : n65966;
  assign n65968 = pi21 ? n65967 : n59342;
  assign n65969 = pi20 ? n65968 : n32;
  assign n65970 = pi19 ? n65964 : n65969;
  assign n65971 = pi18 ? n65961 : n65970;
  assign n65972 = pi17 ? n32 : n65971;
  assign n65973 = pi16 ? n32 : n65972;
  assign n65974 = pi24 ? n157 : n14626;
  assign n65975 = pi23 ? n65974 : n14626;
  assign n65976 = pi22 ? n36781 : n65975;
  assign n65977 = pi21 ? n65976 : n2637;
  assign n65978 = pi20 ? n65977 : n32;
  assign n65979 = pi19 ? n56631 : n65978;
  assign n65980 = pi18 ? n42206 : n65979;
  assign n65981 = pi17 ? n32 : n65980;
  assign n65982 = pi16 ? n32 : n65981;
  assign n65983 = pi15 ? n65973 : n65982;
  assign n65984 = pi21 ? n57698 : n65084;
  assign n65985 = pi20 ? n65984 : n32;
  assign n65986 = pi19 ? n63239 : n65985;
  assign n65987 = pi18 ? n42206 : n65986;
  assign n65988 = pi17 ? n32 : n65987;
  assign n65989 = pi16 ? n32 : n65988;
  assign n65990 = pi21 ? n65091 : n928;
  assign n65991 = pi20 ? n65990 : n32;
  assign n65992 = pi19 ? n63239 : n65991;
  assign n65993 = pi18 ? n42206 : n65992;
  assign n65994 = pi17 ? n32 : n65993;
  assign n65995 = pi16 ? n32 : n65994;
  assign n65996 = pi15 ? n65989 : n65995;
  assign n65997 = pi14 ? n65983 : n65996;
  assign n65998 = pi18 ? n42206 : n65104;
  assign n65999 = pi17 ? n32 : n65998;
  assign n66000 = pi16 ? n32 : n65999;
  assign n66001 = pi20 ? n61941 : n32;
  assign n66002 = pi19 ? n65101 : n66001;
  assign n66003 = pi18 ? n42206 : n66002;
  assign n66004 = pi17 ? n32 : n66003;
  assign n66005 = pi16 ? n32 : n66004;
  assign n66006 = pi15 ? n66000 : n66005;
  assign n66007 = pi23 ? n30868 : n56987;
  assign n66008 = pi22 ? n20563 : n66007;
  assign n66009 = pi21 ? n66008 : n36798;
  assign n66010 = pi20 ? n20563 : n66009;
  assign n66011 = pi21 ? n64842 : n32;
  assign n66012 = pi20 ? n66011 : n32;
  assign n66013 = pi19 ? n66010 : n66012;
  assign n66014 = pi18 ? n42206 : n66013;
  assign n66015 = pi17 ? n32 : n66014;
  assign n66016 = pi16 ? n32 : n66015;
  assign n66017 = pi22 ? n39190 : n42106;
  assign n66018 = pi21 ? n66017 : n59774;
  assign n66019 = pi20 ? n20563 : n66018;
  assign n66020 = pi21 ? n65356 : n32;
  assign n66021 = pi20 ? n66020 : n32;
  assign n66022 = pi19 ? n66019 : n66021;
  assign n66023 = pi18 ? n41630 : n66022;
  assign n66024 = pi17 ? n32 : n66023;
  assign n66025 = pi16 ? n32 : n66024;
  assign n66026 = pi15 ? n66016 : n66025;
  assign n66027 = pi14 ? n66006 : n66026;
  assign n66028 = pi13 ? n65997 : n66027;
  assign n66029 = pi12 ? n65956 : n66028;
  assign n66030 = pi19 ? n46062 : n60490;
  assign n66031 = pi24 ? n36798 : n14626;
  assign n66032 = pi23 ? n157 : n66031;
  assign n66033 = pi22 ? n36798 : n66032;
  assign n66034 = pi21 ? n64663 : n66033;
  assign n66035 = pi20 ? n30868 : n66034;
  assign n66036 = pi19 ? n66035 : n64209;
  assign n66037 = pi18 ? n66030 : n66036;
  assign n66038 = pi17 ? n32 : n66037;
  assign n66039 = pi16 ? n32 : n66038;
  assign n66040 = pi21 ? n33792 : n59681;
  assign n66041 = pi20 ? n30868 : n66040;
  assign n66042 = pi23 ? n13481 : n51564;
  assign n66043 = pi22 ? n66042 : n706;
  assign n66044 = pi21 ? n66043 : n32;
  assign n66045 = pi20 ? n66044 : n32;
  assign n66046 = pi19 ? n66041 : n66045;
  assign n66047 = pi18 ? n66030 : n66046;
  assign n66048 = pi17 ? n32 : n66047;
  assign n66049 = pi16 ? n32 : n66048;
  assign n66050 = pi15 ? n66039 : n66049;
  assign n66051 = pi19 ? n32 : n60503;
  assign n66052 = pi21 ? n37878 : n57760;
  assign n66053 = pi20 ? n30868 : n66052;
  assign n66054 = pi19 ? n66053 : n57717;
  assign n66055 = pi18 ? n66051 : n66054;
  assign n66056 = pi17 ? n32 : n66055;
  assign n66057 = pi16 ? n32 : n66056;
  assign n66058 = pi22 ? n36781 : n37276;
  assign n66059 = pi22 ? n43198 : n65432;
  assign n66060 = pi21 ? n66058 : n66059;
  assign n66061 = pi20 ? n30868 : n66060;
  assign n66062 = pi19 ? n66061 : n32;
  assign n66063 = pi18 ? n66051 : n66062;
  assign n66064 = pi17 ? n32 : n66063;
  assign n66065 = pi16 ? n32 : n66064;
  assign n66066 = pi15 ? n66057 : n66065;
  assign n66067 = pi14 ? n66050 : n66066;
  assign n66068 = pi19 ? n32 : n60490;
  assign n66069 = pi22 ? n13481 : n65432;
  assign n66070 = pi21 ? n39972 : n66069;
  assign n66071 = pi20 ? n56662 : n66070;
  assign n66072 = pi19 ? n66071 : n32;
  assign n66073 = pi18 ? n66068 : n66072;
  assign n66074 = pi17 ? n32 : n66073;
  assign n66075 = pi16 ? n32 : n66074;
  assign n66076 = pi22 ? n57197 : n65602;
  assign n66077 = pi21 ? n53551 : n66076;
  assign n66078 = pi20 ? n56662 : n66077;
  assign n66079 = pi19 ? n66078 : n32;
  assign n66080 = pi18 ? n66068 : n66079;
  assign n66081 = pi17 ? n32 : n66080;
  assign n66082 = pi16 ? n32 : n66081;
  assign n66083 = pi15 ? n66075 : n66082;
  assign n66084 = pi22 ? n56186 : n59672;
  assign n66085 = pi21 ? n43198 : n66084;
  assign n66086 = pi20 ? n65204 : n66085;
  assign n66087 = pi19 ? n66086 : n32;
  assign n66088 = pi18 ? n49322 : n66087;
  assign n66089 = pi17 ? n32 : n66088;
  assign n66090 = pi16 ? n32 : n66089;
  assign n66091 = pi20 ? n65035 : n33792;
  assign n66092 = pi19 ? n32 : n66091;
  assign n66093 = pi21 ? n43198 : n64278;
  assign n66094 = pi20 ? n55729 : n66093;
  assign n66095 = pi19 ? n66094 : n32;
  assign n66096 = pi18 ? n66092 : n66095;
  assign n66097 = pi17 ? n32 : n66096;
  assign n66098 = pi16 ? n32 : n66097;
  assign n66099 = pi15 ? n66090 : n66098;
  assign n66100 = pi14 ? n66083 : n66099;
  assign n66101 = pi13 ? n66067 : n66100;
  assign n66102 = pi19 ? n32 : n33792;
  assign n66103 = pi18 ? n66102 : n65630;
  assign n66104 = pi17 ? n32 : n66103;
  assign n66105 = pi16 ? n32 : n66104;
  assign n66106 = pi21 ? n56760 : n65247;
  assign n66107 = pi20 ? n55729 : n66106;
  assign n66108 = pi19 ? n66107 : n32;
  assign n66109 = pi18 ? n66102 : n66108;
  assign n66110 = pi17 ? n32 : n66109;
  assign n66111 = pi16 ? n32 : n66110;
  assign n66112 = pi15 ? n66105 : n66111;
  assign n66113 = pi22 ? n32 : n43199;
  assign n66114 = pi21 ? n66113 : n43198;
  assign n66115 = pi20 ? n66114 : n43198;
  assign n66116 = pi19 ? n32 : n66115;
  assign n66117 = pi18 ? n66116 : n64749;
  assign n66118 = pi17 ? n32 : n66117;
  assign n66119 = pi16 ? n32 : n66118;
  assign n66120 = pi21 ? n57760 : n53983;
  assign n66121 = pi20 ? n43198 : n66120;
  assign n66122 = pi19 ? n66121 : n32;
  assign n66123 = pi18 ? n66116 : n66122;
  assign n66124 = pi17 ? n32 : n66123;
  assign n66125 = pi16 ? n32 : n66124;
  assign n66126 = pi15 ? n66119 : n66125;
  assign n66127 = pi14 ? n66112 : n66126;
  assign n66128 = pi21 ? n46727 : n64332;
  assign n66129 = pi21 ? n58725 : n64333;
  assign n66130 = pi20 ? n66128 : n66129;
  assign n66131 = pi19 ? n32 : n66130;
  assign n66132 = pi22 ? n64325 : n49412;
  assign n66133 = pi21 ? n66132 : n43198;
  assign n66134 = pi20 ? n66133 : n58439;
  assign n66135 = pi19 ? n66134 : n32;
  assign n66136 = pi18 ? n66131 : n66135;
  assign n66137 = pi17 ? n32 : n66136;
  assign n66138 = pi16 ? n32 : n66137;
  assign n66139 = pi22 ? n32 : n55641;
  assign n66140 = pi21 ? n66139 : n14626;
  assign n66141 = pi20 ? n66140 : n14626;
  assign n66142 = pi19 ? n32 : n66141;
  assign n66143 = pi18 ? n66142 : n63439;
  assign n66144 = pi17 ? n32 : n66143;
  assign n66145 = pi16 ? n32 : n66144;
  assign n66146 = pi15 ? n66138 : n66145;
  assign n66147 = pi21 ? n48856 : n55708;
  assign n66148 = pi20 ? n66147 : n14626;
  assign n66149 = pi19 ? n32 : n66148;
  assign n66150 = pi21 ? n65066 : n32;
  assign n66151 = pi20 ? n14626 : n66150;
  assign n66152 = pi19 ? n66151 : n32;
  assign n66153 = pi18 ? n66149 : n66152;
  assign n66154 = pi17 ? n32 : n66153;
  assign n66155 = pi16 ? n32 : n66154;
  assign n66156 = pi20 ? n64753 : n14626;
  assign n66157 = pi19 ? n32 : n66156;
  assign n66158 = pi21 ? n14626 : n57746;
  assign n66159 = pi20 ? n66158 : n65666;
  assign n66160 = pi19 ? n66159 : n32;
  assign n66161 = pi18 ? n66157 : n66160;
  assign n66162 = pi17 ? n32 : n66161;
  assign n66163 = pi16 ? n32 : n66162;
  assign n66164 = pi15 ? n66155 : n66163;
  assign n66165 = pi14 ? n66146 : n66164;
  assign n66166 = pi13 ? n66127 : n66165;
  assign n66167 = pi12 ? n66101 : n66166;
  assign n66168 = pi11 ? n66029 : n66167;
  assign n66169 = pi10 ? n65867 : n66168;
  assign n66170 = pi09 ? n65696 : n66169;
  assign n66171 = pi19 ? n39396 : n64788;
  assign n66172 = pi18 ? n32 : n66171;
  assign n66173 = pi17 ? n32 : n66172;
  assign n66174 = pi16 ? n32 : n66173;
  assign n66175 = pi15 ? n32 : n66174;
  assign n66176 = pi19 ? n38315 : n62954;
  assign n66177 = pi18 ? n32 : n66176;
  assign n66178 = pi17 ? n32 : n66177;
  assign n66179 = pi16 ? n32 : n66178;
  assign n66180 = pi18 ? n32 : n62955;
  assign n66181 = pi17 ? n32 : n66180;
  assign n66182 = pi16 ? n32 : n66181;
  assign n66183 = pi15 ? n66179 : n66182;
  assign n66184 = pi14 ? n66175 : n66183;
  assign n66185 = pi13 ? n32 : n66184;
  assign n66186 = pi12 ? n32 : n66185;
  assign n66187 = pi11 ? n32 : n66186;
  assign n66188 = pi10 ? n32 : n66187;
  assign n66189 = pi18 ? n37928 : n62955;
  assign n66190 = pi17 ? n32 : n66189;
  assign n66191 = pi16 ? n32 : n66190;
  assign n66192 = pi15 ? n66182 : n66191;
  assign n66193 = pi18 ? n37928 : n62976;
  assign n66194 = pi17 ? n32 : n66193;
  assign n66195 = pi16 ? n32 : n66194;
  assign n66196 = pi18 ? n40056 : n62976;
  assign n66197 = pi17 ? n32 : n66196;
  assign n66198 = pi16 ? n32 : n66197;
  assign n66199 = pi15 ? n66195 : n66198;
  assign n66200 = pi14 ? n66192 : n66199;
  assign n66201 = pi18 ? n37935 : n62976;
  assign n66202 = pi17 ? n32 : n66201;
  assign n66203 = pi16 ? n32 : n66202;
  assign n66204 = pi18 ? n37322 : n62976;
  assign n66205 = pi17 ? n32 : n66204;
  assign n66206 = pi16 ? n32 : n66205;
  assign n66207 = pi15 ? n66203 : n66206;
  assign n66208 = pi18 ? n37335 : n62976;
  assign n66209 = pi17 ? n32 : n66208;
  assign n66210 = pi16 ? n32 : n66209;
  assign n66211 = pi15 ? n66210 : n65332;
  assign n66212 = pi14 ? n66207 : n66211;
  assign n66213 = pi13 ? n66200 : n66212;
  assign n66214 = pi14 ? n65332 : n64796;
  assign n66215 = pi18 ? n28159 : n59296;
  assign n66216 = pi17 ? n32 : n66215;
  assign n66217 = pi16 ? n32 : n66216;
  assign n66218 = pi18 ? n30119 : n59307;
  assign n66219 = pi17 ? n32 : n66218;
  assign n66220 = pi16 ? n32 : n66219;
  assign n66221 = pi15 ? n66217 : n66220;
  assign n66222 = pi18 ? n31265 : n65359;
  assign n66223 = pi17 ? n32 : n66222;
  assign n66224 = pi16 ? n32 : n66223;
  assign n66225 = pi18 ? n31265 : n64850;
  assign n66226 = pi17 ? n32 : n66225;
  assign n66227 = pi16 ? n32 : n66226;
  assign n66228 = pi15 ? n66224 : n66227;
  assign n66229 = pi14 ? n66221 : n66228;
  assign n66230 = pi13 ? n66214 : n66229;
  assign n66231 = pi12 ? n66213 : n66230;
  assign n66232 = pi18 ? n31265 : n65743;
  assign n66233 = pi17 ? n32 : n66232;
  assign n66234 = pi16 ? n32 : n66233;
  assign n66235 = pi18 ? n31315 : n65743;
  assign n66236 = pi17 ? n32 : n66235;
  assign n66237 = pi16 ? n32 : n66236;
  assign n66238 = pi15 ? n66234 : n66237;
  assign n66239 = pi18 ? n31315 : n65755;
  assign n66240 = pi17 ? n32 : n66239;
  assign n66241 = pi16 ? n32 : n66240;
  assign n66242 = pi18 ? n44246 : n65762;
  assign n66243 = pi17 ? n32 : n66242;
  assign n66244 = pi16 ? n32 : n66243;
  assign n66245 = pi15 ? n66241 : n66244;
  assign n66246 = pi14 ? n66238 : n66245;
  assign n66247 = pi18 ? n44246 : n65771;
  assign n66248 = pi17 ? n32 : n66247;
  assign n66249 = pi16 ? n32 : n66248;
  assign n66250 = pi18 ? n43222 : n65779;
  assign n66251 = pi17 ? n32 : n66250;
  assign n66252 = pi16 ? n32 : n66251;
  assign n66253 = pi15 ? n66249 : n66252;
  assign n66254 = pi18 ? n43222 : n65787;
  assign n66255 = pi17 ? n32 : n66254;
  assign n66256 = pi16 ? n32 : n66255;
  assign n66257 = pi18 ? n43222 : n65795;
  assign n66258 = pi17 ? n32 : n66257;
  assign n66259 = pi16 ? n32 : n66258;
  assign n66260 = pi15 ? n66256 : n66259;
  assign n66261 = pi14 ? n66253 : n66260;
  assign n66262 = pi13 ? n66246 : n66261;
  assign n66263 = pi18 ? n43226 : n65806;
  assign n66264 = pi17 ? n32 : n66263;
  assign n66265 = pi16 ? n32 : n66264;
  assign n66266 = pi18 ? n43226 : n65813;
  assign n66267 = pi17 ? n32 : n66266;
  assign n66268 = pi16 ? n32 : n66267;
  assign n66269 = pi15 ? n66265 : n66268;
  assign n66270 = pi18 ? n43247 : n65823;
  assign n66271 = pi17 ? n32 : n66270;
  assign n66272 = pi16 ? n32 : n66271;
  assign n66273 = pi18 ? n43247 : n65833;
  assign n66274 = pi17 ? n32 : n66273;
  assign n66275 = pi16 ? n32 : n66274;
  assign n66276 = pi15 ? n66272 : n66275;
  assign n66277 = pi14 ? n66269 : n66276;
  assign n66278 = pi18 ? n44273 : n65841;
  assign n66279 = pi17 ? n32 : n66278;
  assign n66280 = pi16 ? n32 : n66279;
  assign n66281 = pi20 ? n65845 : n56130;
  assign n66282 = pi19 ? n20563 : n66281;
  assign n66283 = pi18 ? n44273 : n66282;
  assign n66284 = pi17 ? n32 : n66283;
  assign n66285 = pi16 ? n32 : n66284;
  assign n66286 = pi15 ? n66280 : n66285;
  assign n66287 = pi18 ? n44273 : n65436;
  assign n66288 = pi17 ? n32 : n66287;
  assign n66289 = pi16 ? n32 : n66288;
  assign n66290 = pi22 ? n861 : n14626;
  assign n66291 = pi21 ? n40986 : n66290;
  assign n66292 = pi20 ? n66291 : n4116;
  assign n66293 = pi19 ? n20563 : n66292;
  assign n66294 = pi18 ? n44273 : n66293;
  assign n66295 = pi17 ? n32 : n66294;
  assign n66296 = pi16 ? n32 : n66295;
  assign n66297 = pi15 ? n66289 : n66296;
  assign n66298 = pi14 ? n66286 : n66297;
  assign n66299 = pi13 ? n66277 : n66298;
  assign n66300 = pi12 ? n66262 : n66299;
  assign n66301 = pi11 ? n66231 : n66300;
  assign n66302 = pi23 ? n65206 : n685;
  assign n66303 = pi22 ? n861 : n66302;
  assign n66304 = pi21 ? n40986 : n66303;
  assign n66305 = pi20 ? n66304 : n10011;
  assign n66306 = pi19 ? n40792 : n66305;
  assign n66307 = pi18 ? n44273 : n66306;
  assign n66308 = pi17 ? n32 : n66307;
  assign n66309 = pi16 ? n32 : n66308;
  assign n66310 = pi23 ? n61520 : n316;
  assign n66311 = pi22 ? n448 : n66310;
  assign n66312 = pi21 ? n45016 : n66311;
  assign n66313 = pi20 ? n66312 : n32257;
  assign n66314 = pi19 ? n40792 : n66313;
  assign n66315 = pi18 ? n48623 : n66314;
  assign n66316 = pi17 ? n32 : n66315;
  assign n66317 = pi16 ? n32 : n66316;
  assign n66318 = pi15 ? n66309 : n66317;
  assign n66319 = pi22 ? n59412 : n63543;
  assign n66320 = pi21 ? n40986 : n66319;
  assign n66321 = pi20 ? n66320 : n20953;
  assign n66322 = pi19 ? n59458 : n66321;
  assign n66323 = pi18 ? n48623 : n66322;
  assign n66324 = pi17 ? n32 : n66323;
  assign n66325 = pi16 ? n32 : n66324;
  assign n66326 = pi23 ? n56987 : n30868;
  assign n66327 = pi22 ? n20563 : n66326;
  assign n66328 = pi21 ? n38375 : n66327;
  assign n66329 = pi20 ? n66328 : n20563;
  assign n66330 = pi19 ? n32 : n66329;
  assign n66331 = pi18 ? n66330 : n65897;
  assign n66332 = pi17 ? n32 : n66331;
  assign n66333 = pi16 ? n32 : n66332;
  assign n66334 = pi15 ? n66325 : n66333;
  assign n66335 = pi14 ? n66318 : n66334;
  assign n66336 = pi23 ? n62332 : n33792;
  assign n66337 = pi22 ? n20563 : n66336;
  assign n66338 = pi21 ? n38375 : n66337;
  assign n66339 = pi20 ? n66338 : n20563;
  assign n66340 = pi19 ? n32 : n66339;
  assign n66341 = pi21 ? n51313 : n64248;
  assign n66342 = pi20 ? n66341 : n32;
  assign n66343 = pi19 ? n65905 : n66342;
  assign n66344 = pi18 ? n66340 : n66343;
  assign n66345 = pi17 ? n32 : n66344;
  assign n66346 = pi16 ? n32 : n66345;
  assign n66347 = pi21 ? n38375 : n45016;
  assign n66348 = pi20 ? n66347 : n20563;
  assign n66349 = pi19 ? n32 : n66348;
  assign n66350 = pi20 ? n51280 : n65916;
  assign n66351 = pi21 ? n65919 : n65038;
  assign n66352 = pi20 ? n66351 : n32;
  assign n66353 = pi19 ? n66350 : n66352;
  assign n66354 = pi18 ? n66349 : n66353;
  assign n66355 = pi17 ? n32 : n66354;
  assign n66356 = pi16 ? n32 : n66355;
  assign n66357 = pi15 ? n66346 : n66356;
  assign n66358 = pi21 ? n38375 : n40986;
  assign n66359 = pi20 ? n66358 : n51280;
  assign n66360 = pi19 ? n32 : n66359;
  assign n66361 = pi20 ? n41578 : n65035;
  assign n66362 = pi22 ? n33792 : n65049;
  assign n66363 = pi22 ? n2299 : n56665;
  assign n66364 = pi21 ? n66362 : n66363;
  assign n66365 = pi20 ? n66364 : n32;
  assign n66366 = pi19 ? n66361 : n66365;
  assign n66367 = pi18 ? n66360 : n66366;
  assign n66368 = pi17 ? n32 : n66367;
  assign n66369 = pi16 ? n32 : n66368;
  assign n66370 = pi21 ? n38375 : n36659;
  assign n66371 = pi20 ? n66370 : n51280;
  assign n66372 = pi19 ? n32 : n66371;
  assign n66373 = pi23 ? n65063 : n204;
  assign n66374 = pi22 ? n36659 : n66373;
  assign n66375 = pi22 ? n57659 : n14363;
  assign n66376 = pi21 ? n66374 : n66375;
  assign n66377 = pi20 ? n66376 : n32;
  assign n66378 = pi19 ? n65048 : n66377;
  assign n66379 = pi18 ? n66372 : n66378;
  assign n66380 = pi17 ? n32 : n66379;
  assign n66381 = pi16 ? n32 : n66380;
  assign n66382 = pi15 ? n66369 : n66381;
  assign n66383 = pi14 ? n66357 : n66382;
  assign n66384 = pi13 ? n66335 : n66383;
  assign n66385 = pi24 ? n36781 : n20563;
  assign n66386 = pi23 ? n36781 : n66385;
  assign n66387 = pi22 ? n40386 : n66386;
  assign n66388 = pi21 ? n39394 : n66387;
  assign n66389 = pi21 ? n20563 : n52632;
  assign n66390 = pi20 ? n66388 : n66389;
  assign n66391 = pi19 ? n32 : n66390;
  assign n66392 = pi22 ? n36781 : n20563;
  assign n66393 = pi21 ? n66392 : n36249;
  assign n66394 = pi20 ? n66393 : n47361;
  assign n66395 = pi23 ? n24414 : n233;
  assign n66396 = pi22 ? n36659 : n66395;
  assign n66397 = pi21 ? n66396 : n59342;
  assign n66398 = pi20 ? n66397 : n32;
  assign n66399 = pi19 ? n66394 : n66398;
  assign n66400 = pi18 ? n66391 : n66399;
  assign n66401 = pi17 ? n32 : n66400;
  assign n66402 = pi16 ? n32 : n66401;
  assign n66403 = pi18 ? n42200 : n65979;
  assign n66404 = pi17 ? n32 : n66403;
  assign n66405 = pi16 ? n32 : n66404;
  assign n66406 = pi15 ? n66402 : n66405;
  assign n66407 = pi21 ? n57698 : n5370;
  assign n66408 = pi20 ? n66407 : n32;
  assign n66409 = pi19 ? n63239 : n66408;
  assign n66410 = pi18 ? n42200 : n66409;
  assign n66411 = pi17 ? n32 : n66410;
  assign n66412 = pi16 ? n32 : n66411;
  assign n66413 = pi18 ? n42200 : n65992;
  assign n66414 = pi17 ? n32 : n66413;
  assign n66415 = pi16 ? n32 : n66414;
  assign n66416 = pi15 ? n66412 : n66415;
  assign n66417 = pi14 ? n66406 : n66416;
  assign n66418 = pi21 ? n57733 : n1009;
  assign n66419 = pi20 ? n66418 : n32;
  assign n66420 = pi19 ? n65101 : n66419;
  assign n66421 = pi18 ? n42654 : n66420;
  assign n66422 = pi17 ? n32 : n66421;
  assign n66423 = pi16 ? n32 : n66422;
  assign n66424 = pi22 ? n43198 : n63009;
  assign n66425 = pi21 ? n66424 : n32;
  assign n66426 = pi20 ? n66425 : n32;
  assign n66427 = pi19 ? n65101 : n66426;
  assign n66428 = pi18 ? n42654 : n66427;
  assign n66429 = pi17 ? n32 : n66428;
  assign n66430 = pi16 ? n32 : n66429;
  assign n66431 = pi15 ? n66423 : n66430;
  assign n66432 = pi23 ? n30868 : n36798;
  assign n66433 = pi22 ? n20563 : n66432;
  assign n66434 = pi21 ? n66433 : n36798;
  assign n66435 = pi20 ? n20563 : n66434;
  assign n66436 = pi19 ? n66435 : n66012;
  assign n66437 = pi18 ? n42654 : n66436;
  assign n66438 = pi17 ? n32 : n66437;
  assign n66439 = pi16 ? n32 : n66438;
  assign n66440 = pi21 ? n59539 : n32;
  assign n66441 = pi20 ? n66440 : n32;
  assign n66442 = pi19 ? n66019 : n66441;
  assign n66443 = pi18 ? n42680 : n66442;
  assign n66444 = pi17 ? n32 : n66443;
  assign n66445 = pi16 ? n32 : n66444;
  assign n66446 = pi15 ? n66439 : n66445;
  assign n66447 = pi14 ? n66431 : n66446;
  assign n66448 = pi13 ? n66417 : n66447;
  assign n66449 = pi12 ? n66384 : n66448;
  assign n66450 = pi23 ? n55567 : n33792;
  assign n66451 = pi22 ? n30868 : n66450;
  assign n66452 = pi22 ? n36798 : n1457;
  assign n66453 = pi21 ? n66451 : n66452;
  assign n66454 = pi20 ? n30868 : n66453;
  assign n66455 = pi21 ? n57563 : n32;
  assign n66456 = pi20 ? n66455 : n32;
  assign n66457 = pi19 ? n66454 : n66456;
  assign n66458 = pi18 ? n60868 : n66457;
  assign n66459 = pi17 ? n32 : n66458;
  assign n66460 = pi16 ? n32 : n66459;
  assign n66461 = pi19 ? n66041 : n56131;
  assign n66462 = pi18 ? n60868 : n66461;
  assign n66463 = pi17 ? n32 : n66462;
  assign n66464 = pi16 ? n32 : n66463;
  assign n66465 = pi15 ? n66460 : n66464;
  assign n66466 = pi19 ? n66053 : n60046;
  assign n66467 = pi18 ? n60868 : n66466;
  assign n66468 = pi17 ? n32 : n66467;
  assign n66469 = pi16 ? n32 : n66468;
  assign n66470 = pi18 ? n60868 : n66062;
  assign n66471 = pi17 ? n32 : n66470;
  assign n66472 = pi16 ? n32 : n66471;
  assign n66473 = pi15 ? n66469 : n66472;
  assign n66474 = pi14 ? n66465 : n66473;
  assign n66475 = pi22 ? n13481 : n59395;
  assign n66476 = pi21 ? n39972 : n66475;
  assign n66477 = pi20 ? n56662 : n66476;
  assign n66478 = pi19 ? n66477 : n32;
  assign n66479 = pi18 ? n60868 : n66478;
  assign n66480 = pi17 ? n32 : n66479;
  assign n66481 = pi16 ? n32 : n66480;
  assign n66482 = pi22 ? n57197 : n54563;
  assign n66483 = pi21 ? n53551 : n66482;
  assign n66484 = pi20 ? n56662 : n66483;
  assign n66485 = pi19 ? n66484 : n32;
  assign n66486 = pi18 ? n60868 : n66485;
  assign n66487 = pi17 ? n32 : n66486;
  assign n66488 = pi16 ? n32 : n66487;
  assign n66489 = pi15 ? n66481 : n66488;
  assign n66490 = pi22 ? n56186 : n55688;
  assign n66491 = pi21 ? n43198 : n66490;
  assign n66492 = pi20 ? n65204 : n66491;
  assign n66493 = pi19 ? n66492 : n32;
  assign n66494 = pi18 ? n49789 : n66493;
  assign n66495 = pi17 ? n32 : n66494;
  assign n66496 = pi16 ? n32 : n66495;
  assign n66497 = pi19 ? n32 : n52261;
  assign n66498 = pi21 ? n43198 : n59648;
  assign n66499 = pi20 ? n55729 : n66498;
  assign n66500 = pi19 ? n66499 : n32;
  assign n66501 = pi18 ? n66497 : n66500;
  assign n66502 = pi17 ? n32 : n66501;
  assign n66503 = pi16 ? n32 : n66502;
  assign n66504 = pi15 ? n66496 : n66503;
  assign n66505 = pi14 ? n66489 : n66504;
  assign n66506 = pi13 ? n66474 : n66505;
  assign n66507 = pi19 ? n32 : n63796;
  assign n66508 = pi21 ? n43198 : n57097;
  assign n66509 = pi20 ? n55729 : n66508;
  assign n66510 = pi19 ? n66509 : n32;
  assign n66511 = pi18 ? n66507 : n66510;
  assign n66512 = pi17 ? n32 : n66511;
  assign n66513 = pi16 ? n32 : n66512;
  assign n66514 = pi18 ? n66507 : n66108;
  assign n66515 = pi17 ? n32 : n66514;
  assign n66516 = pi16 ? n32 : n66515;
  assign n66517 = pi15 ? n66513 : n66516;
  assign n66518 = pi18 ? n60908 : n64749;
  assign n66519 = pi17 ? n32 : n66518;
  assign n66520 = pi16 ? n32 : n66519;
  assign n66521 = pi21 ? n57760 : n20952;
  assign n66522 = pi20 ? n43198 : n66521;
  assign n66523 = pi19 ? n66522 : n32;
  assign n66524 = pi18 ? n60908 : n66523;
  assign n66525 = pi17 ? n32 : n66524;
  assign n66526 = pi16 ? n32 : n66525;
  assign n66527 = pi15 ? n66520 : n66526;
  assign n66528 = pi14 ? n66517 : n66527;
  assign n66529 = pi22 ? n14626 : n63317;
  assign n66530 = pi21 ? n32 : n66529;
  assign n66531 = pi21 ? n64326 : n64333;
  assign n66532 = pi20 ? n66530 : n66531;
  assign n66533 = pi19 ? n32 : n66532;
  assign n66534 = pi22 ? n14626 : n62510;
  assign n66535 = pi21 ? n66534 : n43198;
  assign n66536 = pi20 ? n66535 : n58439;
  assign n66537 = pi19 ? n66536 : n32;
  assign n66538 = pi18 ? n66533 : n66537;
  assign n66539 = pi17 ? n32 : n66538;
  assign n66540 = pi16 ? n32 : n66539;
  assign n66541 = pi21 ? n32 : n14626;
  assign n66542 = pi20 ? n66541 : n14626;
  assign n66543 = pi19 ? n32 : n66542;
  assign n66544 = pi20 ? n14626 : n59649;
  assign n66545 = pi19 ? n66544 : n32;
  assign n66546 = pi18 ? n66543 : n66545;
  assign n66547 = pi17 ? n32 : n66546;
  assign n66548 = pi16 ? n32 : n66547;
  assign n66549 = pi15 ? n66540 : n66548;
  assign n66550 = pi19 ? n32 : n63831;
  assign n66551 = pi18 ? n66550 : n66152;
  assign n66552 = pi17 ? n32 : n66551;
  assign n66553 = pi16 ? n32 : n66552;
  assign n66554 = pi20 ? n48857 : n14626;
  assign n66555 = pi19 ? n32 : n66554;
  assign n66556 = pi20 ? n66158 : n59466;
  assign n66557 = pi19 ? n66556 : n32;
  assign n66558 = pi18 ? n66555 : n66557;
  assign n66559 = pi17 ? n32 : n66558;
  assign n66560 = pi16 ? n32 : n66559;
  assign n66561 = pi15 ? n66553 : n66560;
  assign n66562 = pi14 ? n66549 : n66561;
  assign n66563 = pi13 ? n66528 : n66562;
  assign n66564 = pi12 ? n66506 : n66563;
  assign n66565 = pi11 ? n66449 : n66564;
  assign n66566 = pi10 ? n66301 : n66565;
  assign n66567 = pi09 ? n66188 : n66566;
  assign n66568 = pi08 ? n66170 : n66567;
  assign n66569 = pi07 ? n65679 : n66568;
  assign n66570 = pi06 ? n64786 : n66569;
  assign n66571 = pi20 ? n31266 : n12225;
  assign n66572 = pi19 ? n39396 : n66571;
  assign n66573 = pi18 ? n32 : n66572;
  assign n66574 = pi17 ? n32 : n66573;
  assign n66575 = pi16 ? n32 : n66574;
  assign n66576 = pi15 ? n32 : n66575;
  assign n66577 = pi21 ? n29133 : n1618;
  assign n66578 = pi20 ? n36250 : n66577;
  assign n66579 = pi19 ? n39396 : n66578;
  assign n66580 = pi18 ? n32 : n66579;
  assign n66581 = pi17 ? n32 : n66580;
  assign n66582 = pi16 ? n32 : n66581;
  assign n66583 = pi19 ? n40549 : n62975;
  assign n66584 = pi18 ? n32 : n66583;
  assign n66585 = pi17 ? n32 : n66584;
  assign n66586 = pi16 ? n32 : n66585;
  assign n66587 = pi15 ? n66582 : n66586;
  assign n66588 = pi14 ? n66576 : n66587;
  assign n66589 = pi13 ? n32 : n66588;
  assign n66590 = pi12 ? n32 : n66589;
  assign n66591 = pi11 ? n32 : n66590;
  assign n66592 = pi10 ? n32 : n66591;
  assign n66593 = pi20 ? n48905 : n1619;
  assign n66594 = pi19 ? n42192 : n66593;
  assign n66595 = pi18 ? n32 : n66594;
  assign n66596 = pi17 ? n32 : n66595;
  assign n66597 = pi16 ? n32 : n66596;
  assign n66598 = pi15 ? n66586 : n66597;
  assign n66599 = pi20 ? n31263 : n31266;
  assign n66600 = pi19 ? n66599 : n66593;
  assign n66601 = pi18 ? n32 : n66600;
  assign n66602 = pi17 ? n32 : n66601;
  assign n66603 = pi16 ? n32 : n66602;
  assign n66604 = pi18 ? n32 : n62976;
  assign n66605 = pi17 ? n32 : n66604;
  assign n66606 = pi16 ? n32 : n66605;
  assign n66607 = pi15 ? n66603 : n66606;
  assign n66608 = pi14 ? n66598 : n66607;
  assign n66609 = pi15 ? n66182 : n65690;
  assign n66610 = pi18 ? n36869 : n62976;
  assign n66611 = pi17 ? n32 : n66610;
  assign n66612 = pi16 ? n32 : n66611;
  assign n66613 = pi14 ? n66609 : n66612;
  assign n66614 = pi13 ? n66608 : n66613;
  assign n66615 = pi20 ? n31913 : n1619;
  assign n66616 = pi19 ? n20563 : n66615;
  assign n66617 = pi18 ? n37957 : n66616;
  assign n66618 = pi17 ? n32 : n66617;
  assign n66619 = pi16 ? n32 : n66618;
  assign n66620 = pi20 ? n36977 : n1619;
  assign n66621 = pi19 ? n20563 : n66620;
  assign n66622 = pi18 ? n37957 : n66621;
  assign n66623 = pi17 ? n32 : n66622;
  assign n66624 = pi16 ? n32 : n66623;
  assign n66625 = pi15 ? n66619 : n66624;
  assign n66626 = pi20 ? n31913 : n61008;
  assign n66627 = pi19 ? n20563 : n66626;
  assign n66628 = pi18 ? n38999 : n66627;
  assign n66629 = pi17 ? n32 : n66628;
  assign n66630 = pi16 ? n32 : n66629;
  assign n66631 = pi15 ? n66630 : n65313;
  assign n66632 = pi14 ? n66625 : n66631;
  assign n66633 = pi23 ? n11117 : n43198;
  assign n66634 = pi22 ? n66633 : n43198;
  assign n66635 = pi22 ? n43198 : n532;
  assign n66636 = pi21 ? n66634 : n66635;
  assign n66637 = pi20 ? n43010 : n66636;
  assign n66638 = pi19 ? n20563 : n66637;
  assign n66639 = pi18 ? n37322 : n66638;
  assign n66640 = pi17 ? n32 : n66639;
  assign n66641 = pi16 ? n32 : n66640;
  assign n66642 = pi21 ? n30868 : n36249;
  assign n66643 = pi20 ? n66642 : n59305;
  assign n66644 = pi19 ? n20563 : n66643;
  assign n66645 = pi18 ? n37335 : n66644;
  assign n66646 = pi17 ? n32 : n66645;
  assign n66647 = pi16 ? n32 : n66646;
  assign n66648 = pi15 ? n66641 : n66647;
  assign n66649 = pi23 ? n65353 : n685;
  assign n66650 = pi22 ? n66649 : n685;
  assign n66651 = pi21 ? n66650 : n696;
  assign n66652 = pi20 ? n40791 : n66651;
  assign n66653 = pi19 ? n20563 : n66652;
  assign n66654 = pi18 ? n38378 : n66653;
  assign n66655 = pi17 ? n32 : n66654;
  assign n66656 = pi16 ? n32 : n66655;
  assign n66657 = pi20 ? n56488 : n64422;
  assign n66658 = pi19 ? n20563 : n66657;
  assign n66659 = pi18 ? n38378 : n66658;
  assign n66660 = pi17 ? n32 : n66659;
  assign n66661 = pi16 ? n32 : n66660;
  assign n66662 = pi15 ? n66656 : n66661;
  assign n66663 = pi14 ? n66648 : n66662;
  assign n66664 = pi13 ? n66632 : n66663;
  assign n66665 = pi12 ? n66614 : n66664;
  assign n66666 = pi22 ? n37 : n49800;
  assign n66667 = pi21 ? n20563 : n66666;
  assign n66668 = pi20 ? n66667 : n64441;
  assign n66669 = pi19 ? n20563 : n66668;
  assign n66670 = pi18 ? n38378 : n66669;
  assign n66671 = pi17 ? n32 : n66670;
  assign n66672 = pi16 ? n32 : n66671;
  assign n66673 = pi22 ? n57349 : n13481;
  assign n66674 = pi21 ? n66673 : n55560;
  assign n66675 = pi20 ? n55475 : n66674;
  assign n66676 = pi19 ? n20563 : n66675;
  assign n66677 = pi18 ? n39455 : n66676;
  assign n66678 = pi17 ? n32 : n66677;
  assign n66679 = pi16 ? n32 : n66678;
  assign n66680 = pi15 ? n66672 : n66679;
  assign n66681 = pi20 ? n65760 : n61108;
  assign n66682 = pi19 ? n20563 : n66681;
  assign n66683 = pi18 ? n39455 : n66682;
  assign n66684 = pi17 ? n32 : n66683;
  assign n66685 = pi16 ? n32 : n66684;
  assign n66686 = pi22 ? n20563 : n58428;
  assign n66687 = pi21 ? n20563 : n66686;
  assign n66688 = pi20 ? n66687 : n59351;
  assign n66689 = pi19 ? n20563 : n66688;
  assign n66690 = pi18 ? n28159 : n66689;
  assign n66691 = pi17 ? n32 : n66690;
  assign n66692 = pi16 ? n32 : n66691;
  assign n66693 = pi15 ? n66685 : n66692;
  assign n66694 = pi14 ? n66680 : n66693;
  assign n66695 = pi21 ? n33792 : n66686;
  assign n66696 = pi20 ? n66695 : n980;
  assign n66697 = pi19 ? n20563 : n66696;
  assign n66698 = pi18 ? n28159 : n66697;
  assign n66699 = pi17 ? n32 : n66698;
  assign n66700 = pi16 ? n32 : n66699;
  assign n66701 = pi22 ? n20563 : n62321;
  assign n66702 = pi21 ? n33792 : n66701;
  assign n66703 = pi20 ? n66702 : n980;
  assign n66704 = pi19 ? n20563 : n66703;
  assign n66705 = pi18 ? n30119 : n66704;
  assign n66706 = pi17 ? n32 : n66705;
  assign n66707 = pi16 ? n32 : n66706;
  assign n66708 = pi15 ? n66700 : n66707;
  assign n66709 = pi21 ? n30868 : n66701;
  assign n66710 = pi20 ? n66709 : n59388;
  assign n66711 = pi19 ? n20563 : n66710;
  assign n66712 = pi18 ? n30119 : n66711;
  assign n66713 = pi17 ? n32 : n66712;
  assign n66714 = pi16 ? n32 : n66713;
  assign n66715 = pi22 ? n30868 : n62127;
  assign n66716 = pi21 ? n36489 : n66715;
  assign n66717 = pi20 ? n66716 : n59388;
  assign n66718 = pi19 ? n20563 : n66717;
  assign n66719 = pi18 ? n30119 : n66718;
  assign n66720 = pi17 ? n32 : n66719;
  assign n66721 = pi16 ? n32 : n66720;
  assign n66722 = pi15 ? n66714 : n66721;
  assign n66723 = pi14 ? n66708 : n66722;
  assign n66724 = pi13 ? n66694 : n66723;
  assign n66725 = pi23 ? n30868 : n43198;
  assign n66726 = pi22 ? n112 : n66725;
  assign n66727 = pi21 ? n20563 : n66726;
  assign n66728 = pi23 ? n43198 : n63008;
  assign n66729 = pi22 ? n14626 : n66728;
  assign n66730 = pi21 ? n66729 : n32;
  assign n66731 = pi20 ? n66727 : n66730;
  assign n66732 = pi19 ? n20563 : n66731;
  assign n66733 = pi18 ? n31265 : n66732;
  assign n66734 = pi17 ? n32 : n66733;
  assign n66735 = pi16 ? n32 : n66734;
  assign n66736 = pi22 ? n685 : n59395;
  assign n66737 = pi21 ? n66736 : n32;
  assign n66738 = pi20 ? n63101 : n66737;
  assign n66739 = pi19 ? n20563 : n66738;
  assign n66740 = pi18 ? n31265 : n66739;
  assign n66741 = pi17 ? n32 : n66740;
  assign n66742 = pi16 ? n32 : n66741;
  assign n66743 = pi15 ? n66735 : n66742;
  assign n66744 = pi23 ? n33792 : n51564;
  assign n66745 = pi22 ? n33792 : n66744;
  assign n66746 = pi21 ? n30868 : n66745;
  assign n66747 = pi22 ? n51564 : n2192;
  assign n66748 = pi21 ? n66747 : n32;
  assign n66749 = pi20 ? n66746 : n66748;
  assign n66750 = pi19 ? n20563 : n66749;
  assign n66751 = pi18 ? n43217 : n66750;
  assign n66752 = pi17 ? n32 : n66751;
  assign n66753 = pi16 ? n32 : n66752;
  assign n66754 = pi22 ? n36659 : n66744;
  assign n66755 = pi21 ? n30868 : n66754;
  assign n66756 = pi22 ? n13481 : n19696;
  assign n66757 = pi21 ? n66756 : n32;
  assign n66758 = pi20 ? n66755 : n66757;
  assign n66759 = pi19 ? n20563 : n66758;
  assign n66760 = pi18 ? n43217 : n66759;
  assign n66761 = pi17 ? n32 : n66760;
  assign n66762 = pi16 ? n32 : n66761;
  assign n66763 = pi15 ? n66753 : n66762;
  assign n66764 = pi14 ? n66743 : n66763;
  assign n66765 = pi23 ? n36659 : n13481;
  assign n66766 = pi22 ? n363 : n66765;
  assign n66767 = pi21 ? n36659 : n66766;
  assign n66768 = pi20 ? n66767 : n55668;
  assign n66769 = pi19 ? n20563 : n66768;
  assign n66770 = pi18 ? n44246 : n66769;
  assign n66771 = pi17 ? n32 : n66770;
  assign n66772 = pi16 ? n32 : n66771;
  assign n66773 = pi23 ? n64129 : n13481;
  assign n66774 = pi22 ? n36781 : n66773;
  assign n66775 = pi21 ? n36659 : n66774;
  assign n66776 = pi20 ? n66775 : n56130;
  assign n66777 = pi19 ? n20563 : n66776;
  assign n66778 = pi18 ? n44246 : n66777;
  assign n66779 = pi17 ? n32 : n66778;
  assign n66780 = pi16 ? n32 : n66779;
  assign n66781 = pi15 ? n66772 : n66780;
  assign n66782 = pi22 ? n157 : n14626;
  assign n66783 = pi21 ? n45016 : n66782;
  assign n66784 = pi23 ? n685 : n63008;
  assign n66785 = pi22 ? n66784 : n32;
  assign n66786 = pi21 ? n66785 : n32;
  assign n66787 = pi20 ? n66783 : n66786;
  assign n66788 = pi19 ? n20563 : n66787;
  assign n66789 = pi18 ? n44246 : n66788;
  assign n66790 = pi17 ? n32 : n66789;
  assign n66791 = pi16 ? n32 : n66790;
  assign n66792 = pi21 ? n40986 : n55708;
  assign n66793 = pi20 ? n66792 : n58168;
  assign n66794 = pi19 ? n20563 : n66793;
  assign n66795 = pi18 ? n44246 : n66794;
  assign n66796 = pi17 ? n32 : n66795;
  assign n66797 = pi16 ? n32 : n66796;
  assign n66798 = pi15 ? n66791 : n66797;
  assign n66799 = pi14 ? n66781 : n66798;
  assign n66800 = pi13 ? n66764 : n66799;
  assign n66801 = pi12 ? n66724 : n66800;
  assign n66802 = pi11 ? n66665 : n66801;
  assign n66803 = pi21 ? n47220 : n59691;
  assign n66804 = pi20 ? n66803 : n10011;
  assign n66805 = pi19 ? n51301 : n66804;
  assign n66806 = pi18 ? n44246 : n66805;
  assign n66807 = pi17 ? n32 : n66806;
  assign n66808 = pi16 ? n32 : n66807;
  assign n66809 = pi20 ? n20563 : n48278;
  assign n66810 = pi21 ? n47360 : n59691;
  assign n66811 = pi20 ? n66810 : n32257;
  assign n66812 = pi19 ? n66809 : n66811;
  assign n66813 = pi18 ? n43222 : n66812;
  assign n66814 = pi17 ? n32 : n66813;
  assign n66815 = pi16 ? n32 : n66814;
  assign n66816 = pi15 ? n66808 : n66815;
  assign n66817 = pi22 ? n14626 : n62427;
  assign n66818 = pi21 ? n39952 : n66817;
  assign n66819 = pi20 ? n66818 : n20953;
  assign n66820 = pi19 ? n59458 : n66819;
  assign n66821 = pi18 ? n43222 : n66820;
  assign n66822 = pi17 ? n32 : n66821;
  assign n66823 = pi16 ? n32 : n66822;
  assign n66824 = pi22 ? n685 : n65432;
  assign n66825 = pi21 ? n37878 : n66824;
  assign n66826 = pi20 ? n66825 : n32;
  assign n66827 = pi19 ? n20563 : n66826;
  assign n66828 = pi18 ? n43226 : n66827;
  assign n66829 = pi17 ? n32 : n66828;
  assign n66830 = pi16 ? n32 : n66829;
  assign n66831 = pi15 ? n66823 : n66830;
  assign n66832 = pi14 ? n66816 : n66831;
  assign n66833 = pi22 ? n30154 : n39190;
  assign n66834 = pi21 ? n32 : n66833;
  assign n66835 = pi20 ? n66834 : n41912;
  assign n66836 = pi19 ? n32 : n66835;
  assign n66837 = pi20 ? n52244 : n49246;
  assign n66838 = pi22 ? n51564 : n59449;
  assign n66839 = pi21 ? n61446 : n66838;
  assign n66840 = pi20 ? n66839 : n32;
  assign n66841 = pi19 ? n66837 : n66840;
  assign n66842 = pi18 ? n66836 : n66841;
  assign n66843 = pi17 ? n32 : n66842;
  assign n66844 = pi16 ? n32 : n66843;
  assign n66845 = pi21 ? n65903 : n33792;
  assign n66846 = pi20 ? n53326 : n66845;
  assign n66847 = pi22 ? n33792 : n65149;
  assign n66848 = pi21 ? n66847 : n54648;
  assign n66849 = pi20 ? n66848 : n32;
  assign n66850 = pi19 ? n66846 : n66849;
  assign n66851 = pi18 ? n66836 : n66850;
  assign n66852 = pi17 ? n32 : n66851;
  assign n66853 = pi16 ? n32 : n66852;
  assign n66854 = pi15 ? n66844 : n66853;
  assign n66855 = pi22 ? n30154 : n37173;
  assign n66856 = pi21 ? n32 : n66855;
  assign n66857 = pi20 ? n66856 : n45017;
  assign n66858 = pi19 ? n32 : n66857;
  assign n66859 = pi21 ? n36659 : n47360;
  assign n66860 = pi21 ? n54446 : n36659;
  assign n66861 = pi20 ? n66859 : n66860;
  assign n66862 = pi22 ? n33792 : n65506;
  assign n66863 = pi21 ? n66862 : n66756;
  assign n66864 = pi20 ? n66863 : n32;
  assign n66865 = pi19 ? n66861 : n66864;
  assign n66866 = pi18 ? n66858 : n66865;
  assign n66867 = pi17 ? n32 : n66866;
  assign n66868 = pi16 ? n32 : n66867;
  assign n66869 = pi22 ? n36659 : n20563;
  assign n66870 = pi21 ? n36659 : n66869;
  assign n66871 = pi22 ? n37783 : n33792;
  assign n66872 = pi21 ? n66871 : n36781;
  assign n66873 = pi20 ? n66870 : n66872;
  assign n66874 = pi22 ? n36781 : n65506;
  assign n66875 = pi22 ? n56622 : n14363;
  assign n66876 = pi21 ? n66874 : n66875;
  assign n66877 = pi20 ? n66876 : n32;
  assign n66878 = pi19 ? n66873 : n66877;
  assign n66879 = pi18 ? n66858 : n66878;
  assign n66880 = pi17 ? n32 : n66879;
  assign n66881 = pi16 ? n32 : n66880;
  assign n66882 = pi15 ? n66868 : n66881;
  assign n66883 = pi14 ? n66854 : n66882;
  assign n66884 = pi13 ? n66832 : n66883;
  assign n66885 = pi21 ? n64141 : n59342;
  assign n66886 = pi20 ? n66885 : n32;
  assign n66887 = pi19 ? n63239 : n66886;
  assign n66888 = pi18 ? n42654 : n66887;
  assign n66889 = pi17 ? n32 : n66888;
  assign n66890 = pi16 ? n32 : n66889;
  assign n66891 = pi23 ? n66031 : n14626;
  assign n66892 = pi22 ? n36781 : n66891;
  assign n66893 = pi21 ? n66892 : n59357;
  assign n66894 = pi20 ? n66893 : n32;
  assign n66895 = pi19 ? n63239 : n66894;
  assign n66896 = pi18 ? n43247 : n66895;
  assign n66897 = pi17 ? n32 : n66896;
  assign n66898 = pi16 ? n32 : n66897;
  assign n66899 = pi15 ? n66890 : n66898;
  assign n66900 = pi21 ? n20563 : n39972;
  assign n66901 = pi20 ? n20563 : n66900;
  assign n66902 = pi22 ? n14626 : n66302;
  assign n66903 = pi21 ? n66902 : n5370;
  assign n66904 = pi20 ? n66903 : n32;
  assign n66905 = pi19 ? n66901 : n66904;
  assign n66906 = pi18 ? n43247 : n66905;
  assign n66907 = pi17 ? n32 : n66906;
  assign n66908 = pi16 ? n32 : n66907;
  assign n66909 = pi21 ? n59774 : n37639;
  assign n66910 = pi20 ? n66909 : n32;
  assign n66911 = pi19 ? n63239 : n66910;
  assign n66912 = pi18 ? n43247 : n66911;
  assign n66913 = pi17 ? n32 : n66912;
  assign n66914 = pi16 ? n32 : n66913;
  assign n66915 = pi15 ? n66908 : n66914;
  assign n66916 = pi14 ? n66899 : n66915;
  assign n66917 = pi21 ? n57760 : n1009;
  assign n66918 = pi20 ? n66917 : n32;
  assign n66919 = pi19 ? n65101 : n66918;
  assign n66920 = pi18 ? n43247 : n66919;
  assign n66921 = pi17 ? n32 : n66920;
  assign n66922 = pi16 ? n32 : n66921;
  assign n66923 = pi22 ? n56622 : n63009;
  assign n66924 = pi21 ? n66923 : n32;
  assign n66925 = pi20 ? n66924 : n32;
  assign n66926 = pi19 ? n55656 : n66925;
  assign n66927 = pi18 ? n43247 : n66926;
  assign n66928 = pi17 ? n32 : n66927;
  assign n66929 = pi16 ? n32 : n66928;
  assign n66930 = pi15 ? n66922 : n66929;
  assign n66931 = pi21 ? n45016 : n36798;
  assign n66932 = pi20 ? n20563 : n66931;
  assign n66933 = pi22 ? n13481 : n63009;
  assign n66934 = pi21 ? n66933 : n32;
  assign n66935 = pi20 ? n66934 : n32;
  assign n66936 = pi19 ? n66932 : n66935;
  assign n66937 = pi18 ? n43247 : n66936;
  assign n66938 = pi17 ? n32 : n66937;
  assign n66939 = pi16 ? n32 : n66938;
  assign n66940 = pi21 ? n47220 : n59681;
  assign n66941 = pi20 ? n20563 : n66940;
  assign n66942 = pi22 ? n64689 : n53982;
  assign n66943 = pi21 ? n66942 : n32;
  assign n66944 = pi20 ? n66943 : n32;
  assign n66945 = pi19 ? n66941 : n66944;
  assign n66946 = pi18 ? n44273 : n66945;
  assign n66947 = pi17 ? n32 : n66946;
  assign n66948 = pi16 ? n32 : n66947;
  assign n66949 = pi15 ? n66939 : n66948;
  assign n66950 = pi14 ? n66930 : n66949;
  assign n66951 = pi13 ? n66916 : n66950;
  assign n66952 = pi12 ? n66884 : n66951;
  assign n66953 = pi21 ? n32 : n48173;
  assign n66954 = pi20 ? n66953 : n30868;
  assign n66955 = pi19 ? n32 : n66954;
  assign n66956 = pi23 ? n55567 : n36659;
  assign n66957 = pi22 ? n30868 : n66956;
  assign n66958 = pi21 ? n66957 : n59774;
  assign n66959 = pi20 ? n30868 : n66958;
  assign n66960 = pi19 ? n66959 : n56131;
  assign n66961 = pi18 ? n66955 : n66960;
  assign n66962 = pi17 ? n32 : n66961;
  assign n66963 = pi16 ? n32 : n66962;
  assign n66964 = pi20 ? n47192 : n48184;
  assign n66965 = pi19 ? n32 : n66964;
  assign n66966 = pi20 ? n30868 : n53489;
  assign n66967 = pi19 ? n66966 : n56131;
  assign n66968 = pi18 ? n66965 : n66967;
  assign n66969 = pi17 ? n32 : n66968;
  assign n66970 = pi16 ? n32 : n66969;
  assign n66971 = pi15 ? n66963 : n66970;
  assign n66972 = pi20 ? n60023 : n48184;
  assign n66973 = pi19 ? n32 : n66972;
  assign n66974 = pi23 ? n64129 : n14626;
  assign n66975 = pi22 ? n66974 : n13481;
  assign n66976 = pi21 ? n39952 : n66975;
  assign n66977 = pi20 ? n30868 : n66976;
  assign n66978 = pi19 ? n66977 : n60046;
  assign n66979 = pi18 ? n66973 : n66978;
  assign n66980 = pi17 ? n32 : n66979;
  assign n66981 = pi16 ? n32 : n66980;
  assign n66982 = pi20 ? n37933 : n40791;
  assign n66983 = pi19 ? n32 : n66982;
  assign n66984 = pi24 ? n36781 : n43198;
  assign n66985 = pi23 ? n66984 : n51564;
  assign n66986 = pi22 ? n66985 : n65432;
  assign n66987 = pi21 ? n61412 : n66986;
  assign n66988 = pi20 ? n63363 : n66987;
  assign n66989 = pi19 ? n66988 : n32;
  assign n66990 = pi18 ? n66983 : n66989;
  assign n66991 = pi17 ? n32 : n66990;
  assign n66992 = pi16 ? n32 : n66991;
  assign n66993 = pi15 ? n66981 : n66992;
  assign n66994 = pi14 ? n66971 : n66993;
  assign n66995 = pi19 ? n32 : n64239;
  assign n66996 = pi23 ? n66031 : n13481;
  assign n66997 = pi22 ? n66996 : n59672;
  assign n66998 = pi21 ? n46260 : n66997;
  assign n66999 = pi20 ? n63363 : n66998;
  assign n67000 = pi19 ? n66999 : n32;
  assign n67001 = pi18 ? n66995 : n67000;
  assign n67002 = pi17 ? n32 : n67001;
  assign n67003 = pi16 ? n32 : n67002;
  assign n67004 = pi20 ? n37933 : n39805;
  assign n67005 = pi19 ? n32 : n67004;
  assign n67006 = pi21 ? n30868 : n61446;
  assign n67007 = pi22 ? n56622 : n56665;
  assign n67008 = pi21 ? n46283 : n67007;
  assign n67009 = pi20 ? n67006 : n67008;
  assign n67010 = pi19 ? n67009 : n32;
  assign n67011 = pi18 ? n67005 : n67010;
  assign n67012 = pi17 ? n32 : n67011;
  assign n67013 = pi16 ? n32 : n67012;
  assign n67014 = pi15 ? n67003 : n67013;
  assign n67015 = pi22 ? n66725 : n43198;
  assign n67016 = pi21 ? n30868 : n67015;
  assign n67017 = pi22 ? n62473 : n56665;
  assign n67018 = pi21 ? n43198 : n67017;
  assign n67019 = pi20 ? n67016 : n67018;
  assign n67020 = pi19 ? n67019 : n32;
  assign n67021 = pi18 ? n61454 : n67020;
  assign n67022 = pi17 ? n32 : n67021;
  assign n67023 = pi16 ? n32 : n67022;
  assign n67024 = pi21 ? n33792 : n47220;
  assign n67025 = pi20 ? n46061 : n67024;
  assign n67026 = pi19 ? n32 : n67025;
  assign n67027 = pi21 ? n61930 : n59648;
  assign n67028 = pi20 ? n61480 : n67027;
  assign n67029 = pi19 ? n67028 : n32;
  assign n67030 = pi18 ? n67026 : n67029;
  assign n67031 = pi17 ? n32 : n67030;
  assign n67032 = pi16 ? n32 : n67031;
  assign n67033 = pi15 ? n67023 : n67032;
  assign n67034 = pi14 ? n67014 : n67033;
  assign n67035 = pi13 ? n66994 : n67034;
  assign n67036 = pi21 ? n61930 : n55689;
  assign n67037 = pi20 ? n55729 : n67036;
  assign n67038 = pi19 ? n67037 : n32;
  assign n67039 = pi18 ? n61468 : n67038;
  assign n67040 = pi17 ? n32 : n67039;
  assign n67041 = pi16 ? n32 : n67040;
  assign n67042 = pi21 ? n59691 : n53983;
  assign n67043 = pi20 ? n55729 : n67042;
  assign n67044 = pi19 ? n67043 : n32;
  assign n67045 = pi18 ? n61468 : n67044;
  assign n67046 = pi17 ? n32 : n67045;
  assign n67047 = pi16 ? n32 : n67046;
  assign n67048 = pi15 ? n67041 : n67047;
  assign n67049 = pi20 ? n48857 : n56165;
  assign n67050 = pi19 ? n32 : n67049;
  assign n67051 = pi22 ? n55641 : n13481;
  assign n67052 = pi21 ? n67051 : n20952;
  assign n67053 = pi20 ? n43198 : n67052;
  assign n67054 = pi19 ? n67053 : n32;
  assign n67055 = pi18 ? n67050 : n67054;
  assign n67056 = pi17 ? n32 : n67055;
  assign n67057 = pi16 ? n32 : n67056;
  assign n67058 = pi21 ? n58721 : n46280;
  assign n67059 = pi20 ? n32 : n67058;
  assign n67060 = pi19 ? n32 : n67059;
  assign n67061 = pi20 ? n54655 : n58439;
  assign n67062 = pi19 ? n67061 : n32;
  assign n67063 = pi18 ? n67060 : n67062;
  assign n67064 = pi17 ? n32 : n67063;
  assign n67065 = pi16 ? n32 : n67064;
  assign n67066 = pi15 ? n67057 : n67065;
  assign n67067 = pi14 ? n67048 : n67066;
  assign n67068 = pi22 ? n49412 : n14626;
  assign n67069 = pi21 ? n67068 : n14626;
  assign n67070 = pi20 ? n63830 : n67069;
  assign n67071 = pi19 ? n32 : n67070;
  assign n67072 = pi22 ? n57197 : n21502;
  assign n67073 = pi21 ? n67072 : n32;
  assign n67074 = pi20 ? n14626 : n67073;
  assign n67075 = pi19 ? n67074 : n32;
  assign n67076 = pi18 ? n67071 : n67075;
  assign n67077 = pi17 ? n32 : n67076;
  assign n67078 = pi16 ? n32 : n67077;
  assign n67079 = pi21 ? n55708 : n63443;
  assign n67080 = pi20 ? n32 : n67079;
  assign n67081 = pi19 ? n32 : n67080;
  assign n67082 = pi20 ? n14626 : n56130;
  assign n67083 = pi19 ? n67082 : n32;
  assign n67084 = pi18 ? n67081 : n67083;
  assign n67085 = pi17 ? n32 : n67084;
  assign n67086 = pi16 ? n32 : n67085;
  assign n67087 = pi15 ? n67078 : n67086;
  assign n67088 = pi21 ? n63434 : n64333;
  assign n67089 = pi20 ? n32 : n67088;
  assign n67090 = pi19 ? n32 : n67089;
  assign n67091 = pi21 ? n14626 : n63779;
  assign n67092 = pi20 ? n67091 : n60045;
  assign n67093 = pi19 ? n67092 : n32;
  assign n67094 = pi18 ? n67090 : n67093;
  assign n67095 = pi17 ? n32 : n67094;
  assign n67096 = pi16 ? n32 : n67095;
  assign n67097 = pi20 ? n32 : n64329;
  assign n67098 = pi19 ? n32 : n67097;
  assign n67099 = pi20 ? n67091 : n37640;
  assign n67100 = pi19 ? n67099 : n32;
  assign n67101 = pi18 ? n67098 : n67100;
  assign n67102 = pi17 ? n32 : n67101;
  assign n67103 = pi16 ? n32 : n67102;
  assign n67104 = pi15 ? n67096 : n67103;
  assign n67105 = pi14 ? n67087 : n67104;
  assign n67106 = pi13 ? n67067 : n67105;
  assign n67107 = pi12 ? n67035 : n67106;
  assign n67108 = pi11 ? n66952 : n67107;
  assign n67109 = pi10 ? n66802 : n67108;
  assign n67110 = pi09 ? n66592 : n67109;
  assign n67111 = pi19 ? n43246 : n66571;
  assign n67112 = pi18 ? n32 : n67111;
  assign n67113 = pi17 ? n32 : n67112;
  assign n67114 = pi16 ? n32 : n67113;
  assign n67115 = pi15 ? n32 : n67114;
  assign n67116 = pi19 ? n43246 : n66578;
  assign n67117 = pi18 ? n32 : n67116;
  assign n67118 = pi17 ? n32 : n67117;
  assign n67119 = pi16 ? n32 : n67118;
  assign n67120 = pi19 ? n38947 : n62975;
  assign n67121 = pi18 ? n32 : n67120;
  assign n67122 = pi17 ? n32 : n67121;
  assign n67123 = pi16 ? n32 : n67122;
  assign n67124 = pi15 ? n67119 : n67123;
  assign n67125 = pi14 ? n67115 : n67124;
  assign n67126 = pi13 ? n32 : n67125;
  assign n67127 = pi12 ? n32 : n67126;
  assign n67128 = pi11 ? n32 : n67127;
  assign n67129 = pi10 ? n32 : n67128;
  assign n67130 = pi19 ? n40044 : n66593;
  assign n67131 = pi18 ? n32 : n67130;
  assign n67132 = pi17 ? n32 : n67131;
  assign n67133 = pi16 ? n32 : n67132;
  assign n67134 = pi15 ? n67123 : n67133;
  assign n67135 = pi20 ? n39395 : n31266;
  assign n67136 = pi19 ? n67135 : n66593;
  assign n67137 = pi18 ? n32 : n67136;
  assign n67138 = pi17 ? n32 : n67137;
  assign n67139 = pi16 ? n32 : n67138;
  assign n67140 = pi15 ? n67139 : n66586;
  assign n67141 = pi14 ? n67134 : n67140;
  assign n67142 = pi19 ? n40549 : n62954;
  assign n67143 = pi18 ? n32 : n67142;
  assign n67144 = pi17 ? n32 : n67143;
  assign n67145 = pi16 ? n32 : n67144;
  assign n67146 = pi15 ? n67145 : n66182;
  assign n67147 = pi14 ? n67146 : n66195;
  assign n67148 = pi13 ? n67141 : n67147;
  assign n67149 = pi22 ? n20563 : n65540;
  assign n67150 = pi21 ? n20563 : n67149;
  assign n67151 = pi20 ? n67150 : n1619;
  assign n67152 = pi19 ? n20563 : n67151;
  assign n67153 = pi18 ? n37928 : n67152;
  assign n67154 = pi17 ? n32 : n67153;
  assign n67155 = pi16 ? n32 : n67154;
  assign n67156 = pi22 ? n37 : n65540;
  assign n67157 = pi21 ? n20563 : n67156;
  assign n67158 = pi20 ? n67157 : n1619;
  assign n67159 = pi19 ? n20563 : n67158;
  assign n67160 = pi18 ? n37928 : n67159;
  assign n67161 = pi17 ? n32 : n67160;
  assign n67162 = pi16 ? n32 : n67161;
  assign n67163 = pi15 ? n67155 : n67162;
  assign n67164 = pi23 ? n37 : n62332;
  assign n67165 = pi22 ? n20563 : n67164;
  assign n67166 = pi21 ? n20563 : n67165;
  assign n67167 = pi20 ? n67166 : n61008;
  assign n67168 = pi19 ? n20563 : n67167;
  assign n67169 = pi18 ? n40056 : n67168;
  assign n67170 = pi17 ? n32 : n67169;
  assign n67171 = pi16 ? n32 : n67170;
  assign n67172 = pi22 ? n20563 : n62333;
  assign n67173 = pi21 ? n20563 : n67172;
  assign n67174 = pi20 ? n67173 : n61008;
  assign n67175 = pi19 ? n20563 : n67174;
  assign n67176 = pi18 ? n37935 : n67175;
  assign n67177 = pi17 ? n32 : n67176;
  assign n67178 = pi16 ? n32 : n67177;
  assign n67179 = pi15 ? n67171 : n67178;
  assign n67180 = pi14 ? n67163 : n67179;
  assign n67181 = pi20 ? n43010 : n61066;
  assign n67182 = pi19 ? n20563 : n67181;
  assign n67183 = pi18 ? n37935 : n67182;
  assign n67184 = pi17 ? n32 : n67183;
  assign n67185 = pi16 ? n32 : n67184;
  assign n67186 = pi23 ? n64839 : n233;
  assign n67187 = pi22 ? n67186 : n233;
  assign n67188 = pi21 ? n67187 : n650;
  assign n67189 = pi20 ? n66642 : n67188;
  assign n67190 = pi19 ? n20563 : n67189;
  assign n67191 = pi18 ? n36869 : n67190;
  assign n67192 = pi17 ? n32 : n67191;
  assign n67193 = pi16 ? n32 : n67192;
  assign n67194 = pi15 ? n67185 : n67193;
  assign n67195 = pi21 ? n64421 : n696;
  assign n67196 = pi20 ? n40791 : n67195;
  assign n67197 = pi19 ? n20563 : n67196;
  assign n67198 = pi18 ? n36869 : n67197;
  assign n67199 = pi17 ? n32 : n67198;
  assign n67200 = pi16 ? n32 : n67199;
  assign n67201 = pi22 ? n63531 : n685;
  assign n67202 = pi21 ? n67201 : n8486;
  assign n67203 = pi20 ? n56488 : n67202;
  assign n67204 = pi19 ? n20563 : n67203;
  assign n67205 = pi18 ? n37957 : n67204;
  assign n67206 = pi17 ? n32 : n67205;
  assign n67207 = pi16 ? n32 : n67206;
  assign n67208 = pi15 ? n67200 : n67207;
  assign n67209 = pi14 ? n67194 : n67208;
  assign n67210 = pi13 ? n67180 : n67209;
  assign n67211 = pi12 ? n67148 : n67210;
  assign n67212 = pi18 ? n37957 : n66669;
  assign n67213 = pi17 ? n32 : n67212;
  assign n67214 = pi16 ? n32 : n67213;
  assign n67215 = pi24 ? n33792 : n316;
  assign n67216 = pi23 ? n67215 : n316;
  assign n67217 = pi22 ? n67216 : n13481;
  assign n67218 = pi21 ? n67217 : n55560;
  assign n67219 = pi20 ? n55475 : n67218;
  assign n67220 = pi19 ? n20563 : n67219;
  assign n67221 = pi18 ? n38999 : n67220;
  assign n67222 = pi17 ? n32 : n67221;
  assign n67223 = pi16 ? n32 : n67222;
  assign n67224 = pi15 ? n67214 : n67223;
  assign n67225 = pi18 ? n38999 : n66682;
  assign n67226 = pi17 ? n32 : n67225;
  assign n67227 = pi16 ? n32 : n67226;
  assign n67228 = pi18 ? n37322 : n66689;
  assign n67229 = pi17 ? n32 : n67228;
  assign n67230 = pi16 ? n32 : n67229;
  assign n67231 = pi15 ? n67227 : n67230;
  assign n67232 = pi14 ? n67224 : n67231;
  assign n67233 = pi18 ? n37322 : n66697;
  assign n67234 = pi17 ? n32 : n67233;
  assign n67235 = pi16 ? n32 : n67234;
  assign n67236 = pi18 ? n37335 : n66704;
  assign n67237 = pi17 ? n32 : n67236;
  assign n67238 = pi16 ? n32 : n67237;
  assign n67239 = pi15 ? n67235 : n67238;
  assign n67240 = pi18 ? n37335 : n66711;
  assign n67241 = pi17 ? n32 : n67240;
  assign n67242 = pi16 ? n32 : n67241;
  assign n67243 = pi18 ? n37335 : n66718;
  assign n67244 = pi17 ? n32 : n67243;
  assign n67245 = pi16 ? n32 : n67244;
  assign n67246 = pi15 ? n67242 : n67245;
  assign n67247 = pi14 ? n67239 : n67246;
  assign n67248 = pi13 ? n67232 : n67247;
  assign n67249 = pi23 ? n43198 : n687;
  assign n67250 = pi22 ? n14626 : n67249;
  assign n67251 = pi21 ? n67250 : n32;
  assign n67252 = pi20 ? n66727 : n67251;
  assign n67253 = pi19 ? n20563 : n67252;
  assign n67254 = pi18 ? n38378 : n67253;
  assign n67255 = pi17 ? n32 : n67254;
  assign n67256 = pi16 ? n32 : n67255;
  assign n67257 = pi18 ? n38378 : n66739;
  assign n67258 = pi17 ? n32 : n67257;
  assign n67259 = pi16 ? n32 : n67258;
  assign n67260 = pi15 ? n67256 : n67259;
  assign n67261 = pi18 ? n39455 : n66750;
  assign n67262 = pi17 ? n32 : n67261;
  assign n67263 = pi16 ? n32 : n67262;
  assign n67264 = pi23 ? n33792 : n62637;
  assign n67265 = pi22 ? n36659 : n67264;
  assign n67266 = pi21 ? n30868 : n67265;
  assign n67267 = pi20 ? n67266 : n66757;
  assign n67268 = pi19 ? n20563 : n67267;
  assign n67269 = pi18 ? n39455 : n67268;
  assign n67270 = pi17 ? n32 : n67269;
  assign n67271 = pi16 ? n32 : n67270;
  assign n67272 = pi15 ? n67263 : n67271;
  assign n67273 = pi14 ? n67260 : n67272;
  assign n67274 = pi18 ? n28159 : n66769;
  assign n67275 = pi17 ? n32 : n67274;
  assign n67276 = pi16 ? n32 : n67275;
  assign n67277 = pi21 ? n36659 : n46283;
  assign n67278 = pi22 ? n65183 : n32;
  assign n67279 = pi21 ? n67278 : n32;
  assign n67280 = pi20 ? n67277 : n67279;
  assign n67281 = pi19 ? n20563 : n67280;
  assign n67282 = pi18 ? n28159 : n67281;
  assign n67283 = pi17 ? n32 : n67282;
  assign n67284 = pi16 ? n32 : n67283;
  assign n67285 = pi15 ? n67276 : n67284;
  assign n67286 = pi20 ? n66783 : n4116;
  assign n67287 = pi19 ? n20563 : n67286;
  assign n67288 = pi18 ? n28159 : n67287;
  assign n67289 = pi17 ? n32 : n67288;
  assign n67290 = pi16 ? n32 : n67289;
  assign n67291 = pi22 ? n39190 : n36659;
  assign n67292 = pi21 ? n67291 : n55708;
  assign n67293 = pi20 ? n67292 : n5830;
  assign n67294 = pi19 ? n20563 : n67293;
  assign n67295 = pi18 ? n28159 : n67294;
  assign n67296 = pi17 ? n32 : n67295;
  assign n67297 = pi16 ? n32 : n67296;
  assign n67298 = pi15 ? n67290 : n67297;
  assign n67299 = pi14 ? n67285 : n67298;
  assign n67300 = pi13 ? n67273 : n67299;
  assign n67301 = pi12 ? n67248 : n67300;
  assign n67302 = pi11 ? n67211 : n67301;
  assign n67303 = pi18 ? n28159 : n66805;
  assign n67304 = pi17 ? n32 : n67303;
  assign n67305 = pi16 ? n32 : n67304;
  assign n67306 = pi20 ? n66810 : n2653;
  assign n67307 = pi19 ? n66809 : n67306;
  assign n67308 = pi18 ? n43683 : n67307;
  assign n67309 = pi17 ? n32 : n67308;
  assign n67310 = pi16 ? n32 : n67309;
  assign n67311 = pi15 ? n67305 : n67310;
  assign n67312 = pi23 ? n56987 : n20563;
  assign n67313 = pi22 ? n20563 : n67312;
  assign n67314 = pi21 ? n20563 : n67313;
  assign n67315 = pi20 ? n67314 : n53326;
  assign n67316 = pi21 ? n39952 : n66729;
  assign n67317 = pi20 ? n67316 : n32;
  assign n67318 = pi19 ? n67315 : n67317;
  assign n67319 = pi18 ? n43683 : n67318;
  assign n67320 = pi17 ? n32 : n67319;
  assign n67321 = pi16 ? n32 : n67320;
  assign n67322 = pi18 ? n44686 : n66827;
  assign n67323 = pi17 ? n32 : n67322;
  assign n67324 = pi16 ? n32 : n67323;
  assign n67325 = pi15 ? n67321 : n67324;
  assign n67326 = pi14 ? n67311 : n67325;
  assign n67327 = pi20 ? n47848 : n41912;
  assign n67328 = pi19 ? n32 : n67327;
  assign n67329 = pi18 ? n67328 : n66841;
  assign n67330 = pi17 ? n32 : n67329;
  assign n67331 = pi16 ? n32 : n67330;
  assign n67332 = pi18 ? n67328 : n66850;
  assign n67333 = pi17 ? n32 : n67332;
  assign n67334 = pi16 ? n32 : n67333;
  assign n67335 = pi15 ? n67331 : n67334;
  assign n67336 = pi20 ? n51731 : n45017;
  assign n67337 = pi19 ? n32 : n67336;
  assign n67338 = pi21 ? n66862 : n59634;
  assign n67339 = pi20 ? n67338 : n32;
  assign n67340 = pi19 ? n66861 : n67339;
  assign n67341 = pi18 ? n67337 : n67340;
  assign n67342 = pi17 ? n32 : n67341;
  assign n67343 = pi16 ? n32 : n67342;
  assign n67344 = pi23 ? n66385 : n20563;
  assign n67345 = pi22 ? n36659 : n67344;
  assign n67346 = pi21 ? n36659 : n67345;
  assign n67347 = pi20 ? n67346 : n66872;
  assign n67348 = pi23 ? n66984 : n43198;
  assign n67349 = pi22 ? n36781 : n67348;
  assign n67350 = pi21 ? n67349 : n59342;
  assign n67351 = pi20 ? n67350 : n32;
  assign n67352 = pi19 ? n67347 : n67351;
  assign n67353 = pi18 ? n67337 : n67352;
  assign n67354 = pi17 ? n32 : n67353;
  assign n67355 = pi16 ? n32 : n67354;
  assign n67356 = pi15 ? n67343 : n67355;
  assign n67357 = pi14 ? n67335 : n67356;
  assign n67358 = pi13 ? n67326 : n67357;
  assign n67359 = pi18 ? n43217 : n66887;
  assign n67360 = pi17 ? n32 : n67359;
  assign n67361 = pi16 ? n32 : n67360;
  assign n67362 = pi23 ? n60075 : n14626;
  assign n67363 = pi22 ? n36781 : n67362;
  assign n67364 = pi21 ? n67363 : n59357;
  assign n67365 = pi20 ? n67364 : n32;
  assign n67366 = pi19 ? n63239 : n67365;
  assign n67367 = pi18 ? n43217 : n67366;
  assign n67368 = pi17 ? n32 : n67367;
  assign n67369 = pi16 ? n32 : n67368;
  assign n67370 = pi15 ? n67361 : n67369;
  assign n67371 = pi22 ? n14626 : n65207;
  assign n67372 = pi21 ? n67371 : n928;
  assign n67373 = pi20 ? n67372 : n32;
  assign n67374 = pi19 ? n66901 : n67373;
  assign n67375 = pi18 ? n43217 : n67374;
  assign n67376 = pi17 ? n32 : n67375;
  assign n67377 = pi16 ? n32 : n67376;
  assign n67378 = pi18 ? n43217 : n66911;
  assign n67379 = pi17 ? n32 : n67378;
  assign n67380 = pi16 ? n32 : n67379;
  assign n67381 = pi15 ? n67377 : n67380;
  assign n67382 = pi14 ? n67370 : n67381;
  assign n67383 = pi20 ? n66521 : n32;
  assign n67384 = pi19 ? n65101 : n67383;
  assign n67385 = pi18 ? n43217 : n67384;
  assign n67386 = pi17 ? n32 : n67385;
  assign n67387 = pi16 ? n32 : n67386;
  assign n67388 = pi21 ? n66875 : n32;
  assign n67389 = pi20 ? n67388 : n32;
  assign n67390 = pi19 ? n55656 : n67389;
  assign n67391 = pi18 ? n43217 : n67390;
  assign n67392 = pi17 ? n32 : n67391;
  assign n67393 = pi16 ? n32 : n67392;
  assign n67394 = pi15 ? n67387 : n67393;
  assign n67395 = pi19 ? n66932 : n56131;
  assign n67396 = pi18 ? n43217 : n67395;
  assign n67397 = pi17 ? n32 : n67396;
  assign n67398 = pi16 ? n32 : n67397;
  assign n67399 = pi22 ? n66007 : n33792;
  assign n67400 = pi21 ? n67399 : n59681;
  assign n67401 = pi20 ? n20563 : n67400;
  assign n67402 = pi19 ? n67401 : n65567;
  assign n67403 = pi18 ? n44246 : n67402;
  assign n67404 = pi17 ? n32 : n67403;
  assign n67405 = pi16 ? n32 : n67404;
  assign n67406 = pi15 ? n67398 : n67405;
  assign n67407 = pi14 ? n67394 : n67406;
  assign n67408 = pi13 ? n67382 : n67407;
  assign n67409 = pi12 ? n67358 : n67408;
  assign n67410 = pi21 ? n61264 : n59774;
  assign n67411 = pi20 ? n30868 : n67410;
  assign n67412 = pi19 ? n67411 : n55669;
  assign n67413 = pi18 ? n61454 : n67412;
  assign n67414 = pi17 ? n32 : n67413;
  assign n67415 = pi16 ? n32 : n67414;
  assign n67416 = pi20 ? n46061 : n48184;
  assign n67417 = pi19 ? n32 : n67416;
  assign n67418 = pi19 ? n66966 : n60046;
  assign n67419 = pi18 ? n67417 : n67418;
  assign n67420 = pi17 ? n32 : n67419;
  assign n67421 = pi16 ? n32 : n67420;
  assign n67422 = pi15 ? n67415 : n67421;
  assign n67423 = pi20 ? n32 : n48184;
  assign n67424 = pi19 ? n32 : n67423;
  assign n67425 = pi23 ? n64148 : n14626;
  assign n67426 = pi22 ? n67425 : n13481;
  assign n67427 = pi21 ? n39952 : n67426;
  assign n67428 = pi20 ? n30868 : n67427;
  assign n67429 = pi19 ? n67428 : n35482;
  assign n67430 = pi18 ? n67424 : n67429;
  assign n67431 = pi17 ? n32 : n67430;
  assign n67432 = pi16 ? n32 : n67431;
  assign n67433 = pi20 ? n32 : n40791;
  assign n67434 = pi19 ? n32 : n67433;
  assign n67435 = pi22 ? n56664 : n65432;
  assign n67436 = pi21 ? n61412 : n67435;
  assign n67437 = pi20 ? n63363 : n67436;
  assign n67438 = pi19 ? n67437 : n32;
  assign n67439 = pi18 ? n67434 : n67438;
  assign n67440 = pi17 ? n32 : n67439;
  assign n67441 = pi16 ? n32 : n67440;
  assign n67442 = pi15 ? n67432 : n67441;
  assign n67443 = pi14 ? n67422 : n67442;
  assign n67444 = pi19 ? n32 : n59109;
  assign n67445 = pi22 ? n62411 : n59672;
  assign n67446 = pi21 ? n46260 : n67445;
  assign n67447 = pi20 ? n63363 : n67446;
  assign n67448 = pi19 ? n67447 : n32;
  assign n67449 = pi18 ? n67444 : n67448;
  assign n67450 = pi17 ? n32 : n67449;
  assign n67451 = pi16 ? n32 : n67450;
  assign n67452 = pi20 ? n32 : n39805;
  assign n67453 = pi19 ? n32 : n67452;
  assign n67454 = pi22 ? n66432 : n43198;
  assign n67455 = pi21 ? n30868 : n67454;
  assign n67456 = pi22 ? n62888 : n56665;
  assign n67457 = pi21 ? n46283 : n67456;
  assign n67458 = pi20 ? n67455 : n67457;
  assign n67459 = pi19 ? n67458 : n32;
  assign n67460 = pi18 ? n67453 : n67459;
  assign n67461 = pi17 ? n32 : n67460;
  assign n67462 = pi16 ? n32 : n67461;
  assign n67463 = pi15 ? n67451 : n67462;
  assign n67464 = pi21 ? n30868 : n53471;
  assign n67465 = pi24 ? n43198 : n685;
  assign n67466 = pi23 ? n67465 : n316;
  assign n67467 = pi22 ? n67466 : n56665;
  assign n67468 = pi21 ? n43198 : n67467;
  assign n67469 = pi20 ? n67464 : n67468;
  assign n67470 = pi19 ? n67469 : n32;
  assign n67471 = pi18 ? n61860 : n67470;
  assign n67472 = pi17 ? n32 : n67471;
  assign n67473 = pi16 ? n32 : n67472;
  assign n67474 = pi20 ? n32 : n67024;
  assign n67475 = pi19 ? n32 : n67474;
  assign n67476 = pi21 ? n33792 : n55727;
  assign n67477 = pi21 ? n61930 : n55560;
  assign n67478 = pi20 ? n67476 : n67477;
  assign n67479 = pi19 ? n67478 : n32;
  assign n67480 = pi18 ? n67475 : n67479;
  assign n67481 = pi17 ? n32 : n67480;
  assign n67482 = pi16 ? n32 : n67481;
  assign n67483 = pi15 ? n67473 : n67482;
  assign n67484 = pi14 ? n67463 : n67483;
  assign n67485 = pi13 ? n67443 : n67484;
  assign n67486 = pi19 ? n32 : n53306;
  assign n67487 = pi21 ? n58777 : n55689;
  assign n67488 = pi20 ? n55729 : n67487;
  assign n67489 = pi19 ? n67488 : n32;
  assign n67490 = pi18 ? n67486 : n67489;
  assign n67491 = pi17 ? n32 : n67490;
  assign n67492 = pi16 ? n32 : n67491;
  assign n67493 = pi18 ? n67486 : n67044;
  assign n67494 = pi17 ? n32 : n67493;
  assign n67495 = pi16 ? n32 : n67494;
  assign n67496 = pi15 ? n67492 : n67495;
  assign n67497 = pi22 ? n64297 : n13481;
  assign n67498 = pi21 ? n67497 : n20952;
  assign n67499 = pi20 ? n43198 : n67498;
  assign n67500 = pi19 ? n67499 : n32;
  assign n67501 = pi18 ? n61903 : n67500;
  assign n67502 = pi17 ? n32 : n67501;
  assign n67503 = pi16 ? n32 : n67502;
  assign n67504 = pi20 ? n32 : n51903;
  assign n67505 = pi19 ? n32 : n67504;
  assign n67506 = pi21 ? n47396 : n61522;
  assign n67507 = pi20 ? n67506 : n58439;
  assign n67508 = pi19 ? n67507 : n32;
  assign n67509 = pi18 ? n67505 : n67508;
  assign n67510 = pi17 ? n32 : n67509;
  assign n67511 = pi16 ? n32 : n67510;
  assign n67512 = pi15 ? n67503 : n67511;
  assign n67513 = pi14 ? n67496 : n67512;
  assign n67514 = pi19 ? n32 : n64761;
  assign n67515 = pi18 ? n67514 : n67075;
  assign n67516 = pi17 ? n32 : n67515;
  assign n67517 = pi16 ? n32 : n67516;
  assign n67518 = pi21 ? n63829 : n63443;
  assign n67519 = pi20 ? n32 : n67518;
  assign n67520 = pi19 ? n32 : n67519;
  assign n67521 = pi22 ? n14626 : n63307;
  assign n67522 = pi21 ? n14626 : n67521;
  assign n67523 = pi20 ? n67522 : n56130;
  assign n67524 = pi19 ? n67523 : n32;
  assign n67525 = pi18 ? n67520 : n67524;
  assign n67526 = pi17 ? n32 : n67525;
  assign n67527 = pi16 ? n32 : n67526;
  assign n67528 = pi15 ? n67517 : n67527;
  assign n67529 = pi21 ? n63829 : n64333;
  assign n67530 = pi20 ? n32 : n67529;
  assign n67531 = pi19 ? n32 : n67530;
  assign n67532 = pi18 ? n67531 : n67093;
  assign n67533 = pi17 ? n32 : n67532;
  assign n67534 = pi16 ? n32 : n67533;
  assign n67535 = pi19 ? n32 : n64754;
  assign n67536 = pi20 ? n67091 : n20953;
  assign n67537 = pi19 ? n67536 : n32;
  assign n67538 = pi18 ? n67535 : n67537;
  assign n67539 = pi17 ? n32 : n67538;
  assign n67540 = pi16 ? n32 : n67539;
  assign n67541 = pi15 ? n67534 : n67540;
  assign n67542 = pi14 ? n67528 : n67541;
  assign n67543 = pi13 ? n67513 : n67542;
  assign n67544 = pi12 ? n67485 : n67543;
  assign n67545 = pi11 ? n67409 : n67544;
  assign n67546 = pi10 ? n67302 : n67545;
  assign n67547 = pi09 ? n67129 : n67546;
  assign n67548 = pi08 ? n67110 : n67547;
  assign n67549 = pi20 ? n31220 : n12225;
  assign n67550 = pi19 ? n40509 : n67549;
  assign n67551 = pi18 ? n32 : n67550;
  assign n67552 = pi17 ? n32 : n67551;
  assign n67553 = pi16 ? n32 : n67552;
  assign n67554 = pi15 ? n32 : n67553;
  assign n67555 = pi19 ? n40509 : n61569;
  assign n67556 = pi18 ? n32 : n67555;
  assign n67557 = pi17 ? n32 : n67556;
  assign n67558 = pi16 ? n32 : n67557;
  assign n67559 = pi19 ? n40531 : n62975;
  assign n67560 = pi18 ? n32 : n67559;
  assign n67561 = pi17 ? n32 : n67560;
  assign n67562 = pi16 ? n32 : n67561;
  assign n67563 = pi15 ? n67558 : n67562;
  assign n67564 = pi14 ? n67554 : n67563;
  assign n67565 = pi13 ? n32 : n67564;
  assign n67566 = pi12 ? n32 : n67565;
  assign n67567 = pi11 ? n32 : n67566;
  assign n67568 = pi10 ? n32 : n67567;
  assign n67569 = pi21 ? n29133 : n31924;
  assign n67570 = pi20 ? n38997 : n67569;
  assign n67571 = pi19 ? n67570 : n66593;
  assign n67572 = pi18 ? n32 : n67571;
  assign n67573 = pi17 ? n32 : n67572;
  assign n67574 = pi16 ? n32 : n67573;
  assign n67575 = pi15 ? n67562 : n67574;
  assign n67576 = pi20 ? n37320 : n31925;
  assign n67577 = pi19 ? n67576 : n66593;
  assign n67578 = pi18 ? n32 : n67577;
  assign n67579 = pi17 ? n32 : n67578;
  assign n67580 = pi16 ? n32 : n67579;
  assign n67581 = pi15 ? n67580 : n67123;
  assign n67582 = pi14 ? n67575 : n67581;
  assign n67583 = pi19 ? n40549 : n66626;
  assign n67584 = pi18 ? n32 : n67583;
  assign n67585 = pi17 ? n32 : n67584;
  assign n67586 = pi16 ? n32 : n67585;
  assign n67587 = pi15 ? n67145 : n67586;
  assign n67588 = pi19 ? n42192 : n62975;
  assign n67589 = pi18 ? n32 : n67588;
  assign n67590 = pi17 ? n32 : n67589;
  assign n67591 = pi16 ? n32 : n67590;
  assign n67592 = pi14 ? n67587 : n67591;
  assign n67593 = pi13 ? n67582 : n67592;
  assign n67594 = pi19 ? n42192 : n61976;
  assign n67595 = pi18 ? n32 : n67594;
  assign n67596 = pi17 ? n32 : n67595;
  assign n67597 = pi16 ? n32 : n67596;
  assign n67598 = pi20 ? n31263 : n38028;
  assign n67599 = pi21 ? n37 : n57500;
  assign n67600 = pi20 ? n67599 : n1619;
  assign n67601 = pi19 ? n67598 : n67600;
  assign n67602 = pi18 ? n32 : n67601;
  assign n67603 = pi17 ? n32 : n67602;
  assign n67604 = pi16 ? n32 : n67603;
  assign n67605 = pi15 ? n67597 : n67604;
  assign n67606 = pi20 ? n31266 : n61008;
  assign n67607 = pi19 ? n20563 : n67606;
  assign n67608 = pi18 ? n32 : n67607;
  assign n67609 = pi17 ? n32 : n67608;
  assign n67610 = pi16 ? n32 : n67609;
  assign n67611 = pi20 ? n52131 : n61008;
  assign n67612 = pi19 ? n20563 : n67611;
  assign n67613 = pi18 ? n32 : n67612;
  assign n67614 = pi17 ? n32 : n67613;
  assign n67615 = pi16 ? n32 : n67614;
  assign n67616 = pi15 ? n67610 : n67615;
  assign n67617 = pi14 ? n67605 : n67616;
  assign n67618 = pi20 ? n47751 : n61066;
  assign n67619 = pi19 ? n20563 : n67618;
  assign n67620 = pi18 ? n32 : n67619;
  assign n67621 = pi17 ? n32 : n67620;
  assign n67622 = pi16 ? n32 : n67621;
  assign n67623 = pi21 ? n30868 : n56487;
  assign n67624 = pi20 ? n67623 : n67188;
  assign n67625 = pi19 ? n20563 : n67624;
  assign n67626 = pi18 ? n37928 : n67625;
  assign n67627 = pi17 ? n32 : n67626;
  assign n67628 = pi16 ? n32 : n67627;
  assign n67629 = pi15 ? n67622 : n67628;
  assign n67630 = pi18 ? n37928 : n67197;
  assign n67631 = pi17 ? n32 : n67630;
  assign n67632 = pi16 ? n32 : n67631;
  assign n67633 = pi20 ? n58628 : n67202;
  assign n67634 = pi19 ? n20563 : n67633;
  assign n67635 = pi18 ? n37928 : n67634;
  assign n67636 = pi17 ? n32 : n67635;
  assign n67637 = pi16 ? n32 : n67636;
  assign n67638 = pi15 ? n67632 : n67637;
  assign n67639 = pi14 ? n67629 : n67638;
  assign n67640 = pi13 ? n67617 : n67639;
  assign n67641 = pi12 ? n67593 : n67640;
  assign n67642 = pi22 ? n67216 : n316;
  assign n67643 = pi21 ? n67642 : n2320;
  assign n67644 = pi20 ? n58628 : n67643;
  assign n67645 = pi19 ? n20563 : n67644;
  assign n67646 = pi18 ? n37928 : n67645;
  assign n67647 = pi17 ? n32 : n67646;
  assign n67648 = pi16 ? n32 : n67647;
  assign n67649 = pi23 ? n1991 : n13481;
  assign n67650 = pi22 ? n67649 : n13481;
  assign n67651 = pi21 ? n67650 : n55560;
  assign n67652 = pi20 ? n55475 : n67651;
  assign n67653 = pi19 ? n20563 : n67652;
  assign n67654 = pi18 ? n40056 : n67653;
  assign n67655 = pi17 ? n32 : n67654;
  assign n67656 = pi16 ? n32 : n67655;
  assign n67657 = pi15 ? n67648 : n67656;
  assign n67658 = pi20 ? n31913 : n61108;
  assign n67659 = pi19 ? n20563 : n67658;
  assign n67660 = pi18 ? n37935 : n67659;
  assign n67661 = pi17 ? n32 : n67660;
  assign n67662 = pi16 ? n32 : n67661;
  assign n67663 = pi18 ? n37935 : n66689;
  assign n67664 = pi17 ? n32 : n67663;
  assign n67665 = pi16 ? n32 : n67664;
  assign n67666 = pi15 ? n67662 : n67665;
  assign n67667 = pi14 ? n67657 : n67666;
  assign n67668 = pi21 ? n33792 : n63072;
  assign n67669 = pi20 ? n67668 : n980;
  assign n67670 = pi19 ? n20563 : n67669;
  assign n67671 = pi18 ? n37935 : n67670;
  assign n67672 = pi17 ? n32 : n67671;
  assign n67673 = pi16 ? n32 : n67672;
  assign n67674 = pi20 ? n67668 : n63066;
  assign n67675 = pi19 ? n20563 : n67674;
  assign n67676 = pi18 ? n37935 : n67675;
  assign n67677 = pi17 ? n32 : n67676;
  assign n67678 = pi16 ? n32 : n67677;
  assign n67679 = pi15 ? n67673 : n67678;
  assign n67680 = pi23 ? n37 : n43198;
  assign n67681 = pi22 ? n20563 : n67680;
  assign n67682 = pi21 ? n30868 : n67681;
  assign n67683 = pi20 ? n67682 : n59388;
  assign n67684 = pi19 ? n20563 : n67683;
  assign n67685 = pi18 ? n36869 : n67684;
  assign n67686 = pi17 ? n32 : n67685;
  assign n67687 = pi16 ? n32 : n67686;
  assign n67688 = pi23 ? n99 : n43198;
  assign n67689 = pi22 ? n30868 : n67688;
  assign n67690 = pi21 ? n36489 : n67689;
  assign n67691 = pi20 ? n67690 : n58439;
  assign n67692 = pi19 ? n20563 : n67691;
  assign n67693 = pi18 ? n36869 : n67692;
  assign n67694 = pi17 ? n32 : n67693;
  assign n67695 = pi16 ? n32 : n67694;
  assign n67696 = pi15 ? n67687 : n67695;
  assign n67697 = pi14 ? n67679 : n67696;
  assign n67698 = pi13 ? n67667 : n67697;
  assign n67699 = pi23 ? n99 : n14626;
  assign n67700 = pi22 ? n112 : n67699;
  assign n67701 = pi21 ? n20563 : n67700;
  assign n67702 = pi21 ? n64248 : n32;
  assign n67703 = pi20 ? n67701 : n67702;
  assign n67704 = pi19 ? n20563 : n67703;
  assign n67705 = pi18 ? n37957 : n67704;
  assign n67706 = pi17 ? n32 : n67705;
  assign n67707 = pi16 ? n32 : n67706;
  assign n67708 = pi23 ? n30868 : n685;
  assign n67709 = pi22 ? n30869 : n67708;
  assign n67710 = pi21 ? n20563 : n67709;
  assign n67711 = pi22 ? n685 : n54520;
  assign n67712 = pi21 ? n67711 : n32;
  assign n67713 = pi20 ? n67710 : n67712;
  assign n67714 = pi19 ? n20563 : n67713;
  assign n67715 = pi18 ? n37957 : n67714;
  assign n67716 = pi17 ? n32 : n67715;
  assign n67717 = pi16 ? n32 : n67716;
  assign n67718 = pi15 ? n67707 : n67717;
  assign n67719 = pi21 ? n65038 : n32;
  assign n67720 = pi20 ? n66746 : n67719;
  assign n67721 = pi19 ? n20563 : n67720;
  assign n67722 = pi18 ? n38999 : n67721;
  assign n67723 = pi17 ? n32 : n67722;
  assign n67724 = pi16 ? n32 : n67723;
  assign n67725 = pi23 ? n33792 : n316;
  assign n67726 = pi22 ? n36659 : n67725;
  assign n67727 = pi21 ? n30868 : n67726;
  assign n67728 = pi21 ? n64278 : n32;
  assign n67729 = pi20 ? n67727 : n67728;
  assign n67730 = pi19 ? n20563 : n67729;
  assign n67731 = pi18 ? n38999 : n67730;
  assign n67732 = pi17 ? n32 : n67731;
  assign n67733 = pi16 ? n32 : n67732;
  assign n67734 = pi15 ? n67724 : n67733;
  assign n67735 = pi14 ? n67718 : n67734;
  assign n67736 = pi23 ? n363 : n13481;
  assign n67737 = pi22 ? n363 : n67736;
  assign n67738 = pi21 ? n36659 : n67737;
  assign n67739 = pi20 ? n67738 : n56130;
  assign n67740 = pi19 ? n20563 : n67739;
  assign n67741 = pi18 ? n37322 : n67740;
  assign n67742 = pi17 ? n32 : n67741;
  assign n67743 = pi16 ? n32 : n67742;
  assign n67744 = pi22 ? n36781 : n60291;
  assign n67745 = pi21 ? n36659 : n67744;
  assign n67746 = pi20 ? n67745 : n59658;
  assign n67747 = pi19 ? n20563 : n67746;
  assign n67748 = pi18 ? n37322 : n67747;
  assign n67749 = pi17 ? n32 : n67748;
  assign n67750 = pi16 ? n32 : n67749;
  assign n67751 = pi15 ? n67743 : n67750;
  assign n67752 = pi21 ? n45016 : n20460;
  assign n67753 = pi20 ? n67752 : n4116;
  assign n67754 = pi19 ? n20563 : n67753;
  assign n67755 = pi18 ? n37322 : n67754;
  assign n67756 = pi17 ? n32 : n67755;
  assign n67757 = pi16 ? n32 : n67756;
  assign n67758 = pi21 ? n40986 : n59681;
  assign n67759 = pi20 ? n67758 : n54565;
  assign n67760 = pi19 ? n20563 : n67759;
  assign n67761 = pi18 ? n37322 : n67760;
  assign n67762 = pi17 ? n32 : n67761;
  assign n67763 = pi16 ? n32 : n67762;
  assign n67764 = pi15 ? n67757 : n67763;
  assign n67765 = pi14 ? n67751 : n67764;
  assign n67766 = pi13 ? n67735 : n67765;
  assign n67767 = pi12 ? n67698 : n67766;
  assign n67768 = pi11 ? n67641 : n67767;
  assign n67769 = pi21 ? n45016 : n59691;
  assign n67770 = pi20 ? n67769 : n57716;
  assign n67771 = pi19 ? n51301 : n67770;
  assign n67772 = pi18 ? n37322 : n67771;
  assign n67773 = pi17 ? n32 : n67772;
  assign n67774 = pi16 ? n32 : n67773;
  assign n67775 = pi21 ? n40986 : n59691;
  assign n67776 = pi20 ? n67775 : n37640;
  assign n67777 = pi19 ? n66809 : n67776;
  assign n67778 = pi18 ? n37335 : n67777;
  assign n67779 = pi17 ? n32 : n67778;
  assign n67780 = pi16 ? n32 : n67779;
  assign n67781 = pi15 ? n67774 : n67780;
  assign n67782 = pi20 ? n51202 : n53326;
  assign n67783 = pi22 ? n14626 : n6415;
  assign n67784 = pi21 ? n51313 : n67783;
  assign n67785 = pi20 ? n67784 : n32;
  assign n67786 = pi19 ? n67782 : n67785;
  assign n67787 = pi18 ? n37335 : n67786;
  assign n67788 = pi17 ? n32 : n67787;
  assign n67789 = pi16 ? n32 : n67788;
  assign n67790 = pi22 ? n56111 : n20563;
  assign n67791 = pi21 ? n67790 : n20563;
  assign n67792 = pi20 ? n20563 : n67791;
  assign n67793 = pi21 ? n51313 : n2147;
  assign n67794 = pi20 ? n67793 : n32;
  assign n67795 = pi19 ? n67792 : n67794;
  assign n67796 = pi18 ? n38378 : n67795;
  assign n67797 = pi17 ? n32 : n67796;
  assign n67798 = pi16 ? n32 : n67797;
  assign n67799 = pi15 ? n67789 : n67798;
  assign n67800 = pi14 ? n67781 : n67799;
  assign n67801 = pi21 ? n38375 : n36489;
  assign n67802 = pi20 ? n32 : n67801;
  assign n67803 = pi19 ? n32 : n67802;
  assign n67804 = pi22 ? n66450 : n43198;
  assign n67805 = pi21 ? n67804 : n66747;
  assign n67806 = pi20 ? n67805 : n32;
  assign n67807 = pi19 ? n50136 : n67806;
  assign n67808 = pi18 ? n67803 : n67807;
  assign n67809 = pi17 ? n32 : n67808;
  assign n67810 = pi16 ? n32 : n67809;
  assign n67811 = pi22 ? n33792 : n30868;
  assign n67812 = pi21 ? n67811 : n33792;
  assign n67813 = pi20 ? n53326 : n67812;
  assign n67814 = pi22 ? n13481 : n55688;
  assign n67815 = pi21 ? n53471 : n67814;
  assign n67816 = pi20 ? n67815 : n32;
  assign n67817 = pi19 ? n67813 : n67816;
  assign n67818 = pi18 ? n67803 : n67817;
  assign n67819 = pi17 ? n32 : n67818;
  assign n67820 = pi16 ? n32 : n67819;
  assign n67821 = pi15 ? n67810 : n67820;
  assign n67822 = pi20 ? n32 : n66347;
  assign n67823 = pi19 ? n32 : n67822;
  assign n67824 = pi21 ? n33792 : n36659;
  assign n67825 = pi20 ? n41578 : n67824;
  assign n67826 = pi21 ? n64961 : n59648;
  assign n67827 = pi20 ? n67826 : n32;
  assign n67828 = pi19 ? n67825 : n67827;
  assign n67829 = pi18 ? n67823 : n67828;
  assign n67830 = pi17 ? n32 : n67829;
  assign n67831 = pi16 ? n32 : n67830;
  assign n67832 = pi22 ? n36659 : n33792;
  assign n67833 = pi21 ? n67832 : n36781;
  assign n67834 = pi20 ? n36659 : n67833;
  assign n67835 = pi21 ? n63253 : n2637;
  assign n67836 = pi20 ? n67835 : n32;
  assign n67837 = pi19 ? n67834 : n67836;
  assign n67838 = pi18 ? n67823 : n67837;
  assign n67839 = pi17 ? n32 : n67838;
  assign n67840 = pi16 ? n32 : n67839;
  assign n67841 = pi15 ? n67831 : n67840;
  assign n67842 = pi14 ? n67821 : n67841;
  assign n67843 = pi13 ? n67800 : n67842;
  assign n67844 = pi19 ? n63239 : n67836;
  assign n67845 = pi18 ? n31315 : n67844;
  assign n67846 = pi17 ? n32 : n67845;
  assign n67847 = pi16 ? n32 : n67846;
  assign n67848 = pi21 ? n59681 : n928;
  assign n67849 = pi20 ? n67848 : n32;
  assign n67850 = pi19 ? n63239 : n67849;
  assign n67851 = pi18 ? n31315 : n67850;
  assign n67852 = pi17 ? n32 : n67851;
  assign n67853 = pi16 ? n32 : n67852;
  assign n67854 = pi15 ? n67847 : n67853;
  assign n67855 = pi22 ? n36798 : n57674;
  assign n67856 = pi21 ? n67855 : n37639;
  assign n67857 = pi20 ? n67856 : n32;
  assign n67858 = pi19 ? n66901 : n67857;
  assign n67859 = pi18 ? n31315 : n67858;
  assign n67860 = pi17 ? n32 : n67859;
  assign n67861 = pi16 ? n32 : n67860;
  assign n67862 = pi20 ? n60614 : n32;
  assign n67863 = pi19 ? n63239 : n67862;
  assign n67864 = pi18 ? n31315 : n67863;
  assign n67865 = pi17 ? n32 : n67864;
  assign n67866 = pi16 ? n32 : n67865;
  assign n67867 = pi15 ? n67861 : n67866;
  assign n67868 = pi14 ? n67854 : n67867;
  assign n67869 = pi21 ? n51270 : n36798;
  assign n67870 = pi20 ? n20563 : n67869;
  assign n67871 = pi21 ? n57746 : n20952;
  assign n67872 = pi20 ? n67871 : n32;
  assign n67873 = pi19 ? n67870 : n67872;
  assign n67874 = pi18 ? n31315 : n67873;
  assign n67875 = pi17 ? n32 : n67874;
  assign n67876 = pi16 ? n32 : n67875;
  assign n67877 = pi21 ? n61352 : n36798;
  assign n67878 = pi20 ? n20563 : n67877;
  assign n67879 = pi22 ? n57197 : n688;
  assign n67880 = pi21 ? n67879 : n32;
  assign n67881 = pi20 ? n67880 : n32;
  assign n67882 = pi19 ? n67878 : n67881;
  assign n67883 = pi18 ? n31315 : n67882;
  assign n67884 = pi17 ? n32 : n67883;
  assign n67885 = pi16 ? n32 : n67884;
  assign n67886 = pi15 ? n67876 : n67885;
  assign n67887 = pi19 ? n67878 : n64209;
  assign n67888 = pi18 ? n39455 : n67887;
  assign n67889 = pi17 ? n32 : n67888;
  assign n67890 = pi16 ? n32 : n67889;
  assign n67891 = pi20 ? n32 : n46600;
  assign n67892 = pi19 ? n32 : n67891;
  assign n67893 = pi22 ? n57085 : n52395;
  assign n67894 = pi23 ? n43198 : n57517;
  assign n67895 = pi22 ? n36798 : n67894;
  assign n67896 = pi21 ? n67893 : n67895;
  assign n67897 = pi20 ? n54417 : n67896;
  assign n67898 = pi22 ? n56186 : n706;
  assign n67899 = pi21 ? n67898 : n32;
  assign n67900 = pi20 ? n67899 : n32;
  assign n67901 = pi19 ? n67897 : n67900;
  assign n67902 = pi18 ? n67892 : n67901;
  assign n67903 = pi17 ? n32 : n67902;
  assign n67904 = pi16 ? n32 : n67903;
  assign n67905 = pi15 ? n67890 : n67904;
  assign n67906 = pi14 ? n67886 : n67905;
  assign n67907 = pi13 ? n67868 : n67906;
  assign n67908 = pi12 ? n67843 : n67907;
  assign n67909 = pi22 ? n30868 : n52395;
  assign n67910 = pi21 ? n67909 : n58777;
  assign n67911 = pi20 ? n30868 : n67910;
  assign n67912 = pi19 ? n67911 : n56131;
  assign n67913 = pi18 ? n62375 : n67912;
  assign n67914 = pi17 ? n32 : n67913;
  assign n67915 = pi16 ? n32 : n67914;
  assign n67916 = pi22 ? n64662 : n36798;
  assign n67917 = pi21 ? n67916 : n13481;
  assign n67918 = pi20 ? n30868 : n67917;
  assign n67919 = pi19 ? n67918 : n60046;
  assign n67920 = pi18 ? n62375 : n67919;
  assign n67921 = pi17 ? n32 : n67920;
  assign n67922 = pi16 ? n32 : n67921;
  assign n67923 = pi15 ? n67915 : n67922;
  assign n67924 = pi21 ? n64224 : n30868;
  assign n67925 = pi20 ? n32 : n67924;
  assign n67926 = pi19 ? n32 : n67925;
  assign n67927 = pi24 ? n36798 : n33792;
  assign n67928 = pi23 ? n36781 : n67927;
  assign n67929 = pi22 ? n67928 : n36781;
  assign n67930 = pi21 ? n67929 : n57746;
  assign n67931 = pi20 ? n30868 : n67930;
  assign n67932 = pi19 ? n67931 : n35482;
  assign n67933 = pi18 ? n67926 : n67932;
  assign n67934 = pi17 ? n32 : n67933;
  assign n67935 = pi16 ? n32 : n67934;
  assign n67936 = pi22 ? n57782 : n36798;
  assign n67937 = pi21 ? n67936 : n64706;
  assign n67938 = pi20 ? n63363 : n67937;
  assign n67939 = pi19 ? n67938 : n32;
  assign n67940 = pi18 ? n67926 : n67939;
  assign n67941 = pi17 ? n32 : n67940;
  assign n67942 = pi16 ? n32 : n67941;
  assign n67943 = pi15 ? n67935 : n67942;
  assign n67944 = pi14 ? n67923 : n67943;
  assign n67945 = pi19 ? n32 : n59643;
  assign n67946 = pi22 ? n63717 : n43198;
  assign n67947 = pi21 ? n67946 : n62849;
  assign n67948 = pi20 ? n63363 : n67947;
  assign n67949 = pi19 ? n67948 : n32;
  assign n67950 = pi18 ? n67945 : n67949;
  assign n67951 = pi17 ? n32 : n67950;
  assign n67952 = pi16 ? n32 : n67951;
  assign n67953 = pi21 ? n61930 : n64278;
  assign n67954 = pi20 ? n67006 : n67953;
  assign n67955 = pi19 ? n67954 : n32;
  assign n67956 = pi18 ? n62387 : n67955;
  assign n67957 = pi17 ? n32 : n67956;
  assign n67958 = pi16 ? n32 : n67957;
  assign n67959 = pi15 ? n67952 : n67958;
  assign n67960 = pi21 ? n52259 : n30868;
  assign n67961 = pi20 ? n32 : n67960;
  assign n67962 = pi19 ? n32 : n67961;
  assign n67963 = pi21 ? n47220 : n53471;
  assign n67964 = pi22 ? n56186 : n32;
  assign n67965 = pi21 ? n62420 : n67964;
  assign n67966 = pi20 ? n67963 : n67965;
  assign n67967 = pi19 ? n67966 : n32;
  assign n67968 = pi18 ? n67962 : n67967;
  assign n67969 = pi17 ? n32 : n67968;
  assign n67970 = pi16 ? n32 : n67969;
  assign n67971 = pi21 ? n52259 : n47220;
  assign n67972 = pi20 ? n32 : n67971;
  assign n67973 = pi19 ? n32 : n67972;
  assign n67974 = pi20 ? n61480 : n62494;
  assign n67975 = pi19 ? n67974 : n32;
  assign n67976 = pi18 ? n67973 : n67975;
  assign n67977 = pi17 ? n32 : n67976;
  assign n67978 = pi16 ? n32 : n67977;
  assign n67979 = pi15 ? n67970 : n67978;
  assign n67980 = pi14 ? n67959 : n67979;
  assign n67981 = pi13 ? n67944 : n67980;
  assign n67982 = pi21 ? n59691 : n57097;
  assign n67983 = pi20 ? n55729 : n67982;
  assign n67984 = pi19 ? n67983 : n32;
  assign n67985 = pi18 ? n62447 : n67984;
  assign n67986 = pi17 ? n32 : n67985;
  assign n67987 = pi16 ? n32 : n67986;
  assign n67988 = pi20 ? n55729 : n62822;
  assign n67989 = pi19 ? n67988 : n32;
  assign n67990 = pi18 ? n62447 : n67989;
  assign n67991 = pi17 ? n32 : n67990;
  assign n67992 = pi16 ? n32 : n67991;
  assign n67993 = pi15 ? n67987 : n67992;
  assign n67994 = pi21 ? n32 : n55792;
  assign n67995 = pi20 ? n32 : n67994;
  assign n67996 = pi19 ? n32 : n67995;
  assign n67997 = pi21 ? n61485 : n32;
  assign n67998 = pi20 ? n43198 : n67997;
  assign n67999 = pi19 ? n67998 : n32;
  assign n68000 = pi18 ? n67996 : n67999;
  assign n68001 = pi17 ? n32 : n68000;
  assign n68002 = pi16 ? n32 : n68001;
  assign n68003 = pi22 ? n55641 : n14626;
  assign n68004 = pi21 ? n32 : n68003;
  assign n68005 = pi20 ? n32 : n68004;
  assign n68006 = pi19 ? n32 : n68005;
  assign n68007 = pi20 ? n58777 : n64354;
  assign n68008 = pi19 ? n68007 : n32;
  assign n68009 = pi18 ? n68006 : n68008;
  assign n68010 = pi17 ? n32 : n68009;
  assign n68011 = pi16 ? n32 : n68010;
  assign n68012 = pi15 ? n68002 : n68011;
  assign n68013 = pi14 ? n67993 : n68012;
  assign n68014 = pi21 ? n32 : n46280;
  assign n68015 = pi20 ? n32 : n68014;
  assign n68016 = pi19 ? n32 : n68015;
  assign n68017 = pi20 ? n66158 : n56130;
  assign n68018 = pi19 ? n68017 : n32;
  assign n68019 = pi18 ? n68016 : n68018;
  assign n68020 = pi17 ? n32 : n68019;
  assign n68021 = pi16 ? n32 : n68020;
  assign n68022 = pi21 ? n32 : n63443;
  assign n68023 = pi20 ? n32 : n68022;
  assign n68024 = pi19 ? n32 : n68023;
  assign n68025 = pi20 ? n66158 : n60045;
  assign n68026 = pi19 ? n68025 : n32;
  assign n68027 = pi18 ? n68024 : n68026;
  assign n68028 = pi17 ? n32 : n68027;
  assign n68029 = pi16 ? n32 : n68028;
  assign n68030 = pi15 ? n68021 : n68029;
  assign n68031 = pi20 ? n66158 : n32;
  assign n68032 = pi19 ? n68031 : n32;
  assign n68033 = pi18 ? n51332 : n68032;
  assign n68034 = pi17 ? n32 : n68033;
  assign n68035 = pi16 ? n32 : n68034;
  assign n68036 = pi22 ? n56622 : n55688;
  assign n68037 = pi21 ? n14626 : n68036;
  assign n68038 = pi20 ? n68037 : n32;
  assign n68039 = pi19 ? n68038 : n32;
  assign n68040 = pi18 ? n51351 : n68039;
  assign n68041 = pi17 ? n32 : n68040;
  assign n68042 = pi16 ? n32 : n68041;
  assign n68043 = pi15 ? n68035 : n68042;
  assign n68044 = pi14 ? n68030 : n68043;
  assign n68045 = pi13 ? n68013 : n68044;
  assign n68046 = pi12 ? n67981 : n68045;
  assign n68047 = pi11 ? n67908 : n68046;
  assign n68048 = pi10 ? n67768 : n68047;
  assign n68049 = pi09 ? n67568 : n68048;
  assign n68050 = pi19 ? n41681 : n67549;
  assign n68051 = pi18 ? n32 : n68050;
  assign n68052 = pi17 ? n32 : n68051;
  assign n68053 = pi16 ? n32 : n68052;
  assign n68054 = pi15 ? n32 : n68053;
  assign n68055 = pi19 ? n41681 : n61569;
  assign n68056 = pi18 ? n32 : n68055;
  assign n68057 = pi17 ? n32 : n68056;
  assign n68058 = pi16 ? n32 : n68057;
  assign n68059 = pi19 ? n41681 : n62975;
  assign n68060 = pi18 ? n32 : n68059;
  assign n68061 = pi17 ? n32 : n68060;
  assign n68062 = pi16 ? n32 : n68061;
  assign n68063 = pi15 ? n68058 : n68062;
  assign n68064 = pi14 ? n68054 : n68063;
  assign n68065 = pi13 ? n32 : n68064;
  assign n68066 = pi12 ? n32 : n68065;
  assign n68067 = pi11 ? n32 : n68066;
  assign n68068 = pi10 ? n32 : n68067;
  assign n68069 = pi20 ? n37933 : n67569;
  assign n68070 = pi19 ? n68069 : n66593;
  assign n68071 = pi18 ? n32 : n68070;
  assign n68072 = pi17 ? n32 : n68071;
  assign n68073 = pi16 ? n32 : n68072;
  assign n68074 = pi15 ? n68062 : n68073;
  assign n68075 = pi20 ? n37933 : n31925;
  assign n68076 = pi19 ? n68075 : n66593;
  assign n68077 = pi18 ? n32 : n68076;
  assign n68078 = pi17 ? n32 : n68077;
  assign n68079 = pi16 ? n32 : n68078;
  assign n68080 = pi19 ? n39372 : n62975;
  assign n68081 = pi18 ? n32 : n68080;
  assign n68082 = pi17 ? n32 : n68081;
  assign n68083 = pi16 ? n32 : n68082;
  assign n68084 = pi15 ? n68079 : n68083;
  assign n68085 = pi14 ? n68074 : n68084;
  assign n68086 = pi19 ? n38947 : n62954;
  assign n68087 = pi18 ? n32 : n68086;
  assign n68088 = pi17 ? n32 : n68087;
  assign n68089 = pi16 ? n32 : n68088;
  assign n68090 = pi19 ? n38947 : n66626;
  assign n68091 = pi18 ? n32 : n68090;
  assign n68092 = pi17 ? n32 : n68091;
  assign n68093 = pi16 ? n32 : n68092;
  assign n68094 = pi15 ? n68089 : n68093;
  assign n68095 = pi19 ? n38956 : n62975;
  assign n68096 = pi18 ? n32 : n68095;
  assign n68097 = pi17 ? n32 : n68096;
  assign n68098 = pi16 ? n32 : n68097;
  assign n68099 = pi14 ? n68094 : n68098;
  assign n68100 = pi13 ? n68085 : n68099;
  assign n68101 = pi19 ? n40044 : n61976;
  assign n68102 = pi18 ? n32 : n68101;
  assign n68103 = pi17 ? n32 : n68102;
  assign n68104 = pi16 ? n32 : n68103;
  assign n68105 = pi20 ? n39395 : n38028;
  assign n68106 = pi19 ? n68105 : n67600;
  assign n68107 = pi18 ? n32 : n68106;
  assign n68108 = pi17 ? n32 : n68107;
  assign n68109 = pi16 ? n32 : n68108;
  assign n68110 = pi15 ? n68104 : n68109;
  assign n68111 = pi19 ? n40549 : n67606;
  assign n68112 = pi18 ? n32 : n68111;
  assign n68113 = pi17 ? n32 : n68112;
  assign n68114 = pi16 ? n32 : n68113;
  assign n68115 = pi19 ? n40549 : n67611;
  assign n68116 = pi18 ? n32 : n68115;
  assign n68117 = pi17 ? n32 : n68116;
  assign n68118 = pi16 ? n32 : n68117;
  assign n68119 = pi15 ? n68114 : n68118;
  assign n68120 = pi14 ? n68110 : n68119;
  assign n68121 = pi19 ? n40549 : n67618;
  assign n68122 = pi18 ? n32 : n68121;
  assign n68123 = pi17 ? n32 : n68122;
  assign n68124 = pi16 ? n32 : n68123;
  assign n68125 = pi23 ? n234 : n233;
  assign n68126 = pi22 ? n68125 : n233;
  assign n68127 = pi21 ? n68126 : n650;
  assign n68128 = pi20 ? n67623 : n68127;
  assign n68129 = pi19 ? n42192 : n68128;
  assign n68130 = pi18 ? n32 : n68129;
  assign n68131 = pi17 ? n32 : n68130;
  assign n68132 = pi16 ? n32 : n68131;
  assign n68133 = pi15 ? n68124 : n68132;
  assign n68134 = pi19 ? n42192 : n67196;
  assign n68135 = pi18 ? n32 : n68134;
  assign n68136 = pi17 ? n32 : n68135;
  assign n68137 = pi16 ? n32 : n68136;
  assign n68138 = pi23 ? n1748 : n685;
  assign n68139 = pi22 ? n68138 : n685;
  assign n68140 = pi21 ? n68139 : n8486;
  assign n68141 = pi20 ? n58628 : n68140;
  assign n68142 = pi19 ? n42192 : n68141;
  assign n68143 = pi18 ? n32 : n68142;
  assign n68144 = pi17 ? n32 : n68143;
  assign n68145 = pi16 ? n32 : n68144;
  assign n68146 = pi15 ? n68137 : n68145;
  assign n68147 = pi14 ? n68133 : n68146;
  assign n68148 = pi13 ? n68120 : n68147;
  assign n68149 = pi12 ? n68100 : n68148;
  assign n68150 = pi19 ? n43253 : n67644;
  assign n68151 = pi18 ? n32 : n68150;
  assign n68152 = pi17 ? n32 : n68151;
  assign n68153 = pi16 ? n32 : n68152;
  assign n68154 = pi23 ? n65170 : n13481;
  assign n68155 = pi22 ? n68154 : n13481;
  assign n68156 = pi21 ? n68155 : n55560;
  assign n68157 = pi20 ? n55475 : n68156;
  assign n68158 = pi19 ? n20563 : n68157;
  assign n68159 = pi18 ? n32 : n68158;
  assign n68160 = pi17 ? n32 : n68159;
  assign n68161 = pi16 ? n32 : n68160;
  assign n68162 = pi15 ? n68153 : n68161;
  assign n68163 = pi20 ? n63057 : n61108;
  assign n68164 = pi19 ? n20563 : n68163;
  assign n68165 = pi18 ? n32 : n68164;
  assign n68166 = pi17 ? n32 : n68165;
  assign n68167 = pi16 ? n32 : n68166;
  assign n68168 = pi18 ? n32 : n66689;
  assign n68169 = pi17 ? n32 : n68168;
  assign n68170 = pi16 ? n32 : n68169;
  assign n68171 = pi15 ? n68167 : n68170;
  assign n68172 = pi14 ? n68162 : n68171;
  assign n68173 = pi18 ? n32 : n67670;
  assign n68174 = pi17 ? n32 : n68173;
  assign n68175 = pi16 ? n32 : n68174;
  assign n68176 = pi18 ? n32 : n67675;
  assign n68177 = pi17 ? n32 : n68176;
  assign n68178 = pi16 ? n32 : n68177;
  assign n68179 = pi15 ? n68175 : n68178;
  assign n68180 = pi20 ? n67682 : n58439;
  assign n68181 = pi19 ? n20563 : n68180;
  assign n68182 = pi18 ? n32 : n68181;
  assign n68183 = pi17 ? n32 : n68182;
  assign n68184 = pi16 ? n32 : n68183;
  assign n68185 = pi18 ? n32 : n67692;
  assign n68186 = pi17 ? n32 : n68185;
  assign n68187 = pi16 ? n32 : n68186;
  assign n68188 = pi15 ? n68184 : n68187;
  assign n68189 = pi14 ? n68179 : n68188;
  assign n68190 = pi13 ? n68172 : n68189;
  assign n68191 = pi18 ? n38983 : n67704;
  assign n68192 = pi17 ? n32 : n68191;
  assign n68193 = pi16 ? n32 : n68192;
  assign n68194 = pi22 ? n295 : n3472;
  assign n68195 = pi21 ? n20563 : n68194;
  assign n68196 = pi20 ? n68195 : n67712;
  assign n68197 = pi19 ? n20563 : n68196;
  assign n68198 = pi18 ? n40056 : n68197;
  assign n68199 = pi17 ? n32 : n68198;
  assign n68200 = pi16 ? n32 : n68199;
  assign n68201 = pi15 ? n68193 : n68200;
  assign n68202 = pi20 ? n66746 : n58666;
  assign n68203 = pi19 ? n20563 : n68202;
  assign n68204 = pi18 ? n40056 : n68203;
  assign n68205 = pi17 ? n32 : n68204;
  assign n68206 = pi16 ? n32 : n68205;
  assign n68207 = pi23 ? n335 : n13481;
  assign n68208 = pi22 ? n36659 : n68207;
  assign n68209 = pi21 ? n30868 : n68208;
  assign n68210 = pi20 ? n68209 : n67728;
  assign n68211 = pi19 ? n20563 : n68210;
  assign n68212 = pi18 ? n40056 : n68211;
  assign n68213 = pi17 ? n32 : n68212;
  assign n68214 = pi16 ? n32 : n68213;
  assign n68215 = pi15 ? n68206 : n68214;
  assign n68216 = pi14 ? n68201 : n68215;
  assign n68217 = pi18 ? n40056 : n67740;
  assign n68218 = pi17 ? n32 : n68217;
  assign n68219 = pi16 ? n32 : n68218;
  assign n68220 = pi18 ? n37935 : n67747;
  assign n68221 = pi17 ? n32 : n68220;
  assign n68222 = pi16 ? n32 : n68221;
  assign n68223 = pi15 ? n68219 : n68222;
  assign n68224 = pi20 ? n67752 : n58168;
  assign n68225 = pi19 ? n20563 : n68224;
  assign n68226 = pi18 ? n37935 : n68225;
  assign n68227 = pi17 ? n32 : n68226;
  assign n68228 = pi16 ? n32 : n68227;
  assign n68229 = pi20 ? n67758 : n58504;
  assign n68230 = pi19 ? n20563 : n68229;
  assign n68231 = pi18 ? n37935 : n68230;
  assign n68232 = pi17 ? n32 : n68231;
  assign n68233 = pi16 ? n32 : n68232;
  assign n68234 = pi15 ? n68228 : n68233;
  assign n68235 = pi14 ? n68223 : n68234;
  assign n68236 = pi13 ? n68216 : n68235;
  assign n68237 = pi12 ? n68190 : n68236;
  assign n68238 = pi11 ? n68149 : n68237;
  assign n68239 = pi18 ? n37935 : n67771;
  assign n68240 = pi17 ? n32 : n68239;
  assign n68241 = pi16 ? n32 : n68240;
  assign n68242 = pi18 ? n36869 : n67777;
  assign n68243 = pi17 ? n32 : n68242;
  assign n68244 = pi16 ? n32 : n68243;
  assign n68245 = pi15 ? n68241 : n68244;
  assign n68246 = pi18 ? n36869 : n67786;
  assign n68247 = pi17 ? n32 : n68246;
  assign n68248 = pi16 ? n32 : n68247;
  assign n68249 = pi19 ? n20563 : n67794;
  assign n68250 = pi18 ? n37957 : n68249;
  assign n68251 = pi17 ? n32 : n68250;
  assign n68252 = pi16 ? n32 : n68251;
  assign n68253 = pi15 ? n68248 : n68252;
  assign n68254 = pi14 ? n68245 : n68253;
  assign n68255 = pi22 ? n30154 : n30868;
  assign n68256 = pi21 ? n32 : n68255;
  assign n68257 = pi20 ? n32 : n68256;
  assign n68258 = pi19 ? n32 : n68257;
  assign n68259 = pi22 ? n66336 : n20563;
  assign n68260 = pi21 ? n68259 : n30868;
  assign n68261 = pi20 ? n68260 : n43010;
  assign n68262 = pi22 ? n51564 : n52251;
  assign n68263 = pi21 ? n67804 : n68262;
  assign n68264 = pi20 ? n68263 : n32;
  assign n68265 = pi19 ? n68261 : n68264;
  assign n68266 = pi18 ? n68258 : n68265;
  assign n68267 = pi17 ? n32 : n68266;
  assign n68268 = pi16 ? n32 : n68267;
  assign n68269 = pi22 ? n33792 : n39291;
  assign n68270 = pi21 ? n20563 : n68269;
  assign n68271 = pi20 ? n68270 : n67812;
  assign n68272 = pi21 ? n53471 : n64278;
  assign n68273 = pi20 ? n68272 : n32;
  assign n68274 = pi19 ? n68271 : n68273;
  assign n68275 = pi18 ? n68258 : n68274;
  assign n68276 = pi17 ? n32 : n68275;
  assign n68277 = pi16 ? n32 : n68276;
  assign n68278 = pi15 ? n68268 : n68277;
  assign n68279 = pi22 ? n30154 : n33792;
  assign n68280 = pi21 ? n32 : n68279;
  assign n68281 = pi20 ? n32 : n68280;
  assign n68282 = pi19 ? n32 : n68281;
  assign n68283 = pi21 ? n36659 : n40955;
  assign n68284 = pi20 ? n68283 : n67824;
  assign n68285 = pi19 ? n68284 : n67827;
  assign n68286 = pi18 ? n68282 : n68285;
  assign n68287 = pi17 ? n32 : n68286;
  assign n68288 = pi16 ? n32 : n68287;
  assign n68289 = pi22 ? n36659 : n43571;
  assign n68290 = pi21 ? n36659 : n68289;
  assign n68291 = pi20 ? n68290 : n67833;
  assign n68292 = pi19 ? n68291 : n67836;
  assign n68293 = pi18 ? n68282 : n68292;
  assign n68294 = pi17 ? n32 : n68293;
  assign n68295 = pi16 ? n32 : n68294;
  assign n68296 = pi15 ? n68288 : n68295;
  assign n68297 = pi14 ? n68278 : n68296;
  assign n68298 = pi13 ? n68254 : n68297;
  assign n68299 = pi18 ? n39455 : n67844;
  assign n68300 = pi17 ? n32 : n68299;
  assign n68301 = pi16 ? n32 : n68300;
  assign n68302 = pi22 ? n57782 : n51564;
  assign n68303 = pi21 ? n68302 : n928;
  assign n68304 = pi20 ? n68303 : n32;
  assign n68305 = pi19 ? n63239 : n68304;
  assign n68306 = pi18 ? n39455 : n68305;
  assign n68307 = pi17 ? n32 : n68306;
  assign n68308 = pi16 ? n32 : n68307;
  assign n68309 = pi15 ? n68301 : n68308;
  assign n68310 = pi18 ? n38999 : n67858;
  assign n68311 = pi17 ? n32 : n68310;
  assign n68312 = pi16 ? n32 : n68311;
  assign n68313 = pi22 ? n62321 : n20563;
  assign n68314 = pi21 ? n68313 : n36781;
  assign n68315 = pi20 ? n20563 : n68314;
  assign n68316 = pi19 ? n68315 : n63720;
  assign n68317 = pi18 ? n38999 : n68316;
  assign n68318 = pi17 ? n32 : n68317;
  assign n68319 = pi16 ? n32 : n68318;
  assign n68320 = pi15 ? n68312 : n68319;
  assign n68321 = pi14 ? n68309 : n68320;
  assign n68322 = pi22 ? n62321 : n36781;
  assign n68323 = pi21 ? n68322 : n36798;
  assign n68324 = pi20 ? n20563 : n68323;
  assign n68325 = pi22 ? n14626 : n21502;
  assign n68326 = pi21 ? n68325 : n32;
  assign n68327 = pi20 ? n68326 : n32;
  assign n68328 = pi19 ? n68324 : n68327;
  assign n68329 = pi18 ? n38999 : n68328;
  assign n68330 = pi17 ? n32 : n68329;
  assign n68331 = pi16 ? n32 : n68330;
  assign n68332 = pi18 ? n38999 : n67882;
  assign n68333 = pi17 ? n32 : n68332;
  assign n68334 = pi16 ? n32 : n68333;
  assign n68335 = pi15 ? n68331 : n68334;
  assign n68336 = pi18 ? n38999 : n67887;
  assign n68337 = pi17 ? n32 : n68336;
  assign n68338 = pi16 ? n32 : n68337;
  assign n68339 = pi21 ? n32 : n57086;
  assign n68340 = pi20 ? n32 : n68339;
  assign n68341 = pi19 ? n32 : n68340;
  assign n68342 = pi23 ? n55567 : n36781;
  assign n68343 = pi22 ? n39190 : n68342;
  assign n68344 = pi21 ? n68343 : n47397;
  assign n68345 = pi20 ? n54417 : n68344;
  assign n68346 = pi19 ? n68345 : n56700;
  assign n68347 = pi18 ? n68341 : n68346;
  assign n68348 = pi17 ? n32 : n68347;
  assign n68349 = pi16 ? n32 : n68348;
  assign n68350 = pi15 ? n68338 : n68349;
  assign n68351 = pi14 ? n68335 : n68350;
  assign n68352 = pi13 ? n68321 : n68351;
  assign n68353 = pi12 ? n68298 : n68352;
  assign n68354 = pi22 ? n30868 : n64074;
  assign n68355 = pi21 ? n68354 : n58777;
  assign n68356 = pi20 ? n30868 : n68355;
  assign n68357 = pi19 ? n68356 : n56131;
  assign n68358 = pi18 ? n51289 : n68357;
  assign n68359 = pi17 ? n32 : n68358;
  assign n68360 = pi16 ? n32 : n68359;
  assign n68361 = pi23 ? n30868 : n36781;
  assign n68362 = pi22 ? n68361 : n36798;
  assign n68363 = pi21 ? n68362 : n13481;
  assign n68364 = pi20 ? n30868 : n68363;
  assign n68365 = pi19 ? n68364 : n37641;
  assign n68366 = pi18 ? n51289 : n68365;
  assign n68367 = pi17 ? n32 : n68366;
  assign n68368 = pi16 ? n32 : n68367;
  assign n68369 = pi15 ? n68360 : n68368;
  assign n68370 = pi22 ? n38284 : n49412;
  assign n68371 = pi21 ? n68370 : n57746;
  assign n68372 = pi20 ? n30868 : n68371;
  assign n68373 = pi19 ? n68372 : n35482;
  assign n68374 = pi18 ? n51289 : n68373;
  assign n68375 = pi17 ? n32 : n68374;
  assign n68376 = pi16 ? n32 : n68375;
  assign n68377 = pi22 ? n49412 : n53550;
  assign n68378 = pi21 ? n68377 : n64706;
  assign n68379 = pi20 ? n63363 : n68378;
  assign n68380 = pi19 ? n68379 : n32;
  assign n68381 = pi18 ? n51289 : n68380;
  assign n68382 = pi17 ? n32 : n68381;
  assign n68383 = pi16 ? n32 : n68382;
  assign n68384 = pi15 ? n68376 : n68383;
  assign n68385 = pi14 ? n68369 : n68384;
  assign n68386 = pi21 ? n55715 : n62849;
  assign n68387 = pi20 ? n63363 : n68386;
  assign n68388 = pi19 ? n68387 : n32;
  assign n68389 = pi18 ? n37935 : n68388;
  assign n68390 = pi17 ? n32 : n68389;
  assign n68391 = pi16 ? n32 : n68390;
  assign n68392 = pi22 ? n53550 : n55641;
  assign n68393 = pi21 ? n68392 : n64278;
  assign n68394 = pi20 ? n67006 : n68393;
  assign n68395 = pi19 ? n68394 : n32;
  assign n68396 = pi18 ? n46063 : n68395;
  assign n68397 = pi17 ? n32 : n68396;
  assign n68398 = pi16 ? n32 : n68397;
  assign n68399 = pi15 ? n68391 : n68398;
  assign n68400 = pi18 ? n46063 : n67967;
  assign n68401 = pi17 ? n32 : n68400;
  assign n68402 = pi16 ? n32 : n68401;
  assign n68403 = pi18 ? n62906 : n67975;
  assign n68404 = pi17 ? n32 : n68403;
  assign n68405 = pi16 ? n32 : n68404;
  assign n68406 = pi15 ? n68402 : n68405;
  assign n68407 = pi14 ? n68399 : n68406;
  assign n68408 = pi13 ? n68385 : n68407;
  assign n68409 = pi18 ? n62906 : n67984;
  assign n68410 = pi17 ? n32 : n68409;
  assign n68411 = pi16 ? n32 : n68410;
  assign n68412 = pi21 ? n57746 : n32;
  assign n68413 = pi20 ? n55729 : n68412;
  assign n68414 = pi19 ? n68413 : n32;
  assign n68415 = pi18 ? n62906 : n68414;
  assign n68416 = pi17 ? n32 : n68415;
  assign n68417 = pi16 ? n32 : n68416;
  assign n68418 = pi15 ? n68411 : n68417;
  assign n68419 = pi22 ? n56186 : n21502;
  assign n68420 = pi21 ? n68419 : n32;
  assign n68421 = pi20 ? n43198 : n68420;
  assign n68422 = pi19 ? n68421 : n32;
  assign n68423 = pi18 ? n51351 : n68422;
  assign n68424 = pi17 ? n32 : n68423;
  assign n68425 = pi16 ? n32 : n68424;
  assign n68426 = pi20 ? n32 : n63830;
  assign n68427 = pi19 ? n32 : n68426;
  assign n68428 = pi20 ? n58777 : n68420;
  assign n68429 = pi19 ? n68428 : n32;
  assign n68430 = pi18 ? n68427 : n68429;
  assign n68431 = pi17 ? n32 : n68430;
  assign n68432 = pi16 ? n32 : n68431;
  assign n68433 = pi15 ? n68425 : n68432;
  assign n68434 = pi14 ? n68418 : n68433;
  assign n68435 = pi18 ? n32 : n68018;
  assign n68436 = pi17 ? n32 : n68435;
  assign n68437 = pi16 ? n32 : n68436;
  assign n68438 = pi18 ? n32 : n68026;
  assign n68439 = pi17 ? n32 : n68438;
  assign n68440 = pi16 ? n32 : n68439;
  assign n68441 = pi15 ? n68437 : n68440;
  assign n68442 = pi18 ? n32 : n68032;
  assign n68443 = pi17 ? n32 : n68442;
  assign n68444 = pi16 ? n32 : n68443;
  assign n68445 = pi21 ? n14626 : n67007;
  assign n68446 = pi20 ? n68445 : n32;
  assign n68447 = pi19 ? n68446 : n32;
  assign n68448 = pi18 ? n32 : n68447;
  assign n68449 = pi17 ? n32 : n68448;
  assign n68450 = pi16 ? n32 : n68449;
  assign n68451 = pi15 ? n68444 : n68450;
  assign n68452 = pi14 ? n68441 : n68451;
  assign n68453 = pi13 ? n68434 : n68452;
  assign n68454 = pi12 ? n68408 : n68453;
  assign n68455 = pi11 ? n68353 : n68454;
  assign n68456 = pi10 ? n68238 : n68455;
  assign n68457 = pi09 ? n68068 : n68456;
  assign n68458 = pi08 ? n68049 : n68457;
  assign n68459 = pi07 ? n67548 : n68458;
  assign n68460 = pi21 ? n30843 : n29133;
  assign n68461 = pi20 ? n68460 : n13040;
  assign n68462 = pi19 ? n43672 : n68461;
  assign n68463 = pi18 ? n32 : n68462;
  assign n68464 = pi17 ? n32 : n68463;
  assign n68465 = pi16 ? n32 : n68464;
  assign n68466 = pi15 ? n32 : n68465;
  assign n68467 = pi20 ? n38028 : n1619;
  assign n68468 = pi19 ? n43672 : n68467;
  assign n68469 = pi18 ? n32 : n68468;
  assign n68470 = pi17 ? n32 : n68469;
  assign n68471 = pi16 ? n32 : n68470;
  assign n68472 = pi19 ? n43672 : n62975;
  assign n68473 = pi18 ? n32 : n68472;
  assign n68474 = pi17 ? n32 : n68473;
  assign n68475 = pi16 ? n32 : n68474;
  assign n68476 = pi15 ? n68471 : n68475;
  assign n68477 = pi14 ? n68466 : n68476;
  assign n68478 = pi13 ? n32 : n68477;
  assign n68479 = pi12 ? n32 : n68478;
  assign n68480 = pi11 ? n32 : n68479;
  assign n68481 = pi10 ? n32 : n68480;
  assign n68482 = pi20 ? n32 : n31913;
  assign n68483 = pi22 ? n54738 : n37;
  assign n68484 = pi21 ? n68483 : n20563;
  assign n68485 = pi20 ? n68484 : n1619;
  assign n68486 = pi19 ? n68482 : n68485;
  assign n68487 = pi18 ? n32 : n68486;
  assign n68488 = pi17 ? n32 : n68487;
  assign n68489 = pi16 ? n32 : n68488;
  assign n68490 = pi20 ? n52962 : n1619;
  assign n68491 = pi19 ? n40496 : n68490;
  assign n68492 = pi18 ? n32 : n68491;
  assign n68493 = pi17 ? n32 : n68492;
  assign n68494 = pi16 ? n32 : n68493;
  assign n68495 = pi15 ? n68489 : n68494;
  assign n68496 = pi19 ? n40496 : n62975;
  assign n68497 = pi18 ? n32 : n68496;
  assign n68498 = pi17 ? n32 : n68497;
  assign n68499 = pi16 ? n32 : n68498;
  assign n68500 = pi14 ? n68495 : n68499;
  assign n68501 = pi20 ? n37 : n61008;
  assign n68502 = pi19 ? n68075 : n68501;
  assign n68503 = pi18 ? n32 : n68502;
  assign n68504 = pi17 ? n32 : n68503;
  assign n68505 = pi16 ? n32 : n68504;
  assign n68506 = pi20 ? n37933 : n31924;
  assign n68507 = pi19 ? n68506 : n68501;
  assign n68508 = pi18 ? n32 : n68507;
  assign n68509 = pi17 ? n32 : n68508;
  assign n68510 = pi16 ? n32 : n68509;
  assign n68511 = pi15 ? n68505 : n68510;
  assign n68512 = pi19 ? n41707 : n62975;
  assign n68513 = pi18 ? n32 : n68512;
  assign n68514 = pi17 ? n32 : n68513;
  assign n68515 = pi16 ? n32 : n68514;
  assign n68516 = pi14 ? n68511 : n68515;
  assign n68517 = pi13 ? n68500 : n68516;
  assign n68518 = pi20 ? n38997 : n31924;
  assign n68519 = pi20 ? n54040 : n1619;
  assign n68520 = pi19 ? n68518 : n68519;
  assign n68521 = pi18 ? n32 : n68520;
  assign n68522 = pi17 ? n32 : n68521;
  assign n68523 = pi16 ? n32 : n68522;
  assign n68524 = pi19 ? n67576 : n68490;
  assign n68525 = pi18 ? n32 : n68524;
  assign n68526 = pi17 ? n32 : n68525;
  assign n68527 = pi16 ? n32 : n68526;
  assign n68528 = pi15 ? n68523 : n68527;
  assign n68529 = pi14 ? n68528 : n67123;
  assign n68530 = pi20 ? n31266 : n67188;
  assign n68531 = pi19 ? n38947 : n68530;
  assign n68532 = pi18 ? n32 : n68531;
  assign n68533 = pi17 ? n32 : n68532;
  assign n68534 = pi16 ? n32 : n68533;
  assign n68535 = pi20 ? n37333 : n38754;
  assign n68536 = pi20 ? n38754 : n68127;
  assign n68537 = pi19 ? n68535 : n68536;
  assign n68538 = pi18 ? n32 : n68537;
  assign n68539 = pi17 ? n32 : n68538;
  assign n68540 = pi16 ? n32 : n68539;
  assign n68541 = pi15 ? n68534 : n68540;
  assign n68542 = pi21 ? n67201 : n696;
  assign n68543 = pi20 ? n40791 : n68542;
  assign n68544 = pi19 ? n68535 : n68543;
  assign n68545 = pi18 ? n32 : n68544;
  assign n68546 = pi17 ? n32 : n68545;
  assign n68547 = pi16 ? n32 : n68546;
  assign n68548 = pi24 ? n33792 : n685;
  assign n68549 = pi23 ? n68548 : n685;
  assign n68550 = pi22 ? n68549 : n51564;
  assign n68551 = pi21 ? n68550 : n58778;
  assign n68552 = pi20 ? n47158 : n68551;
  assign n68553 = pi19 ? n40044 : n68552;
  assign n68554 = pi18 ? n32 : n68553;
  assign n68555 = pi17 ? n32 : n68554;
  assign n68556 = pi16 ? n32 : n68555;
  assign n68557 = pi15 ? n68547 : n68556;
  assign n68558 = pi14 ? n68541 : n68557;
  assign n68559 = pi13 ? n68529 : n68558;
  assign n68560 = pi12 ? n68517 : n68559;
  assign n68561 = pi21 ? n30843 : n31924;
  assign n68562 = pi20 ? n39395 : n68561;
  assign n68563 = pi21 ? n31200 : n53366;
  assign n68564 = pi23 ? n1991 : n316;
  assign n68565 = pi22 ? n68564 : n316;
  assign n68566 = pi21 ? n68565 : n2320;
  assign n68567 = pi20 ? n68563 : n68566;
  assign n68568 = pi19 ? n68562 : n68567;
  assign n68569 = pi18 ? n32 : n68568;
  assign n68570 = pi17 ? n32 : n68569;
  assign n68571 = pi16 ? n32 : n68570;
  assign n68572 = pi19 ? n40549 : n68157;
  assign n68573 = pi18 ? n32 : n68572;
  assign n68574 = pi17 ? n32 : n68573;
  assign n68575 = pi16 ? n32 : n68574;
  assign n68576 = pi15 ? n68571 : n68575;
  assign n68577 = pi21 ? n30868 : n53385;
  assign n68578 = pi22 ? n66395 : n233;
  assign n68579 = pi21 ? n68578 : n2637;
  assign n68580 = pi20 ? n68577 : n68579;
  assign n68581 = pi19 ? n40549 : n68580;
  assign n68582 = pi18 ? n32 : n68581;
  assign n68583 = pi17 ? n32 : n68582;
  assign n68584 = pi16 ? n32 : n68583;
  assign n68585 = pi20 ? n28157 : n47432;
  assign n68586 = pi21 ? n30868 : n63064;
  assign n68587 = pi20 ? n68586 : n27076;
  assign n68588 = pi19 ? n68585 : n68587;
  assign n68589 = pi18 ? n32 : n68588;
  assign n68590 = pi17 ? n32 : n68589;
  assign n68591 = pi16 ? n32 : n68590;
  assign n68592 = pi15 ? n68584 : n68591;
  assign n68593 = pi14 ? n68576 : n68592;
  assign n68594 = pi20 ? n28157 : n38754;
  assign n68595 = pi22 ? n40386 : n61145;
  assign n68596 = pi21 ? n33792 : n68595;
  assign n68597 = pi20 ? n68596 : n980;
  assign n68598 = pi19 ? n68594 : n68597;
  assign n68599 = pi18 ? n32 : n68598;
  assign n68600 = pi17 ? n32 : n68599;
  assign n68601 = pi16 ? n32 : n68600;
  assign n68602 = pi22 ? n40386 : n33792;
  assign n68603 = pi21 ? n20563 : n68602;
  assign n68604 = pi20 ? n28157 : n68603;
  assign n68605 = pi22 ? n30868 : n61145;
  assign n68606 = pi21 ? n33792 : n68605;
  assign n68607 = pi20 ? n68606 : n63066;
  assign n68608 = pi19 ? n68604 : n68607;
  assign n68609 = pi18 ? n32 : n68608;
  assign n68610 = pi17 ? n32 : n68609;
  assign n68611 = pi16 ? n32 : n68610;
  assign n68612 = pi15 ? n68601 : n68611;
  assign n68613 = pi20 ? n28157 : n54998;
  assign n68614 = pi22 ? n36615 : n62127;
  assign n68615 = pi21 ? n30868 : n68614;
  assign n68616 = pi20 ? n68615 : n58439;
  assign n68617 = pi19 ? n68613 : n68616;
  assign n68618 = pi18 ? n32 : n68617;
  assign n68619 = pi17 ? n32 : n68618;
  assign n68620 = pi16 ? n32 : n68619;
  assign n68621 = pi20 ? n30117 : n55014;
  assign n68622 = pi22 ? n39190 : n11047;
  assign n68623 = pi21 ? n30868 : n68622;
  assign n68624 = pi22 ? n233 : n65470;
  assign n68625 = pi21 ? n68624 : n32;
  assign n68626 = pi20 ? n68623 : n68625;
  assign n68627 = pi19 ? n68621 : n68626;
  assign n68628 = pi18 ? n32 : n68627;
  assign n68629 = pi17 ? n32 : n68628;
  assign n68630 = pi16 ? n32 : n68629;
  assign n68631 = pi15 ? n68620 : n68630;
  assign n68632 = pi14 ? n68612 : n68631;
  assign n68633 = pi13 ? n68593 : n68632;
  assign n68634 = pi22 ? n39190 : n63099;
  assign n68635 = pi21 ? n20563 : n68634;
  assign n68636 = pi20 ? n68635 : n11695;
  assign n68637 = pi19 ? n38315 : n68636;
  assign n68638 = pi18 ? n32 : n68637;
  assign n68639 = pi17 ? n32 : n68638;
  assign n68640 = pi16 ? n32 : n68639;
  assign n68641 = pi20 ? n31313 : n40791;
  assign n68642 = pi23 ? n33792 : n685;
  assign n68643 = pi22 ? n36617 : n68642;
  assign n68644 = pi21 ? n30868 : n68643;
  assign n68645 = pi20 ? n68644 : n66748;
  assign n68646 = pi19 ? n68641 : n68645;
  assign n68647 = pi18 ? n32 : n68646;
  assign n68648 = pi17 ? n32 : n68647;
  assign n68649 = pi16 ? n32 : n68648;
  assign n68650 = pi15 ? n68640 : n68649;
  assign n68651 = pi22 ? n37783 : n448;
  assign n68652 = pi21 ? n30868 : n68651;
  assign n68653 = pi21 ? n50346 : n32;
  assign n68654 = pi20 ? n68652 : n68653;
  assign n68655 = pi19 ? n68641 : n68654;
  assign n68656 = pi18 ? n32 : n68655;
  assign n68657 = pi17 ? n32 : n68656;
  assign n68658 = pi16 ? n32 : n68657;
  assign n68659 = pi20 ? n31313 : n54068;
  assign n68660 = pi22 ? n36659 : n66765;
  assign n68661 = pi21 ? n33792 : n68660;
  assign n68662 = pi20 ? n68661 : n59649;
  assign n68663 = pi19 ? n68659 : n68662;
  assign n68664 = pi18 ? n32 : n68663;
  assign n68665 = pi17 ? n32 : n68664;
  assign n68666 = pi16 ? n32 : n68665;
  assign n68667 = pi15 ? n68658 : n68666;
  assign n68668 = pi14 ? n68650 : n68667;
  assign n68669 = pi22 ? n36781 : n673;
  assign n68670 = pi21 ? n36659 : n68669;
  assign n68671 = pi22 ? n65470 : n32;
  assign n68672 = pi21 ? n68671 : n32;
  assign n68673 = pi20 ? n68670 : n68672;
  assign n68674 = pi19 ? n38315 : n68673;
  assign n68675 = pi18 ? n32 : n68674;
  assign n68676 = pi17 ? n32 : n68675;
  assign n68677 = pi16 ? n32 : n68676;
  assign n68678 = pi22 ? n36798 : n59423;
  assign n68679 = pi21 ? n36659 : n68678;
  assign n68680 = pi20 ? n68679 : n4116;
  assign n68681 = pi19 ? n38315 : n68680;
  assign n68682 = pi18 ? n32 : n68681;
  assign n68683 = pi17 ? n32 : n68682;
  assign n68684 = pi16 ? n32 : n68683;
  assign n68685 = pi15 ? n68677 : n68684;
  assign n68686 = pi22 ? n36798 : n57632;
  assign n68687 = pi21 ? n36659 : n68686;
  assign n68688 = pi20 ? n68687 : n5830;
  assign n68689 = pi19 ? n57682 : n68688;
  assign n68690 = pi18 ? n32 : n68689;
  assign n68691 = pi17 ? n32 : n68690;
  assign n68692 = pi16 ? n32 : n68691;
  assign n68693 = pi22 ? n43198 : n61191;
  assign n68694 = pi21 ? n36659 : n68693;
  assign n68695 = pi20 ? n68694 : n32257;
  assign n68696 = pi19 ? n20563 : n68695;
  assign n68697 = pi18 ? n32 : n68696;
  assign n68698 = pi17 ? n32 : n68697;
  assign n68699 = pi16 ? n32 : n68698;
  assign n68700 = pi15 ? n68692 : n68699;
  assign n68701 = pi14 ? n68685 : n68700;
  assign n68702 = pi13 ? n68668 : n68701;
  assign n68703 = pi12 ? n68633 : n68702;
  assign n68704 = pi11 ? n68560 : n68703;
  assign n68705 = pi20 ? n38754 : n40915;
  assign n68706 = pi22 ? n50339 : n13481;
  assign n68707 = pi21 ? n51564 : n68706;
  assign n68708 = pi20 ? n68707 : n37640;
  assign n68709 = pi19 ? n68705 : n68708;
  assign n68710 = pi18 ? n37928 : n68709;
  assign n68711 = pi17 ? n32 : n68710;
  assign n68712 = pi16 ? n32 : n68711;
  assign n68713 = pi22 ? n39190 : n36781;
  assign n68714 = pi22 ? n14626 : n65470;
  assign n68715 = pi21 ? n68713 : n68714;
  assign n68716 = pi20 ? n68715 : n32;
  assign n68717 = pi19 ? n60490 : n68716;
  assign n68718 = pi18 ? n37928 : n68717;
  assign n68719 = pi17 ? n32 : n68718;
  assign n68720 = pi16 ? n32 : n68719;
  assign n68721 = pi15 ? n68712 : n68720;
  assign n68722 = pi21 ? n48173 : n45016;
  assign n68723 = pi20 ? n68722 : n47223;
  assign n68724 = pi22 ? n42109 : n43198;
  assign n68725 = pi22 ? n63317 : n59395;
  assign n68726 = pi21 ? n68724 : n68725;
  assign n68727 = pi20 ? n68726 : n32;
  assign n68728 = pi19 ? n68723 : n68727;
  assign n68729 = pi18 ? n37928 : n68728;
  assign n68730 = pi17 ? n32 : n68729;
  assign n68731 = pi16 ? n32 : n68730;
  assign n68732 = pi22 ? n46172 : n43198;
  assign n68733 = pi21 ? n68732 : n65478;
  assign n68734 = pi20 ? n68733 : n32;
  assign n68735 = pi19 ? n20563 : n68734;
  assign n68736 = pi18 ? n51823 : n68735;
  assign n68737 = pi17 ? n32 : n68736;
  assign n68738 = pi16 ? n32 : n68737;
  assign n68739 = pi15 ? n68731 : n68738;
  assign n68740 = pi14 ? n68721 : n68739;
  assign n68741 = pi20 ? n52339 : n41912;
  assign n68742 = pi22 ? n58710 : n14626;
  assign n68743 = pi21 ? n68742 : n63376;
  assign n68744 = pi20 ? n68743 : n32;
  assign n68745 = pi19 ? n68741 : n68744;
  assign n68746 = pi18 ? n51703 : n68745;
  assign n68747 = pi17 ? n32 : n68746;
  assign n68748 = pi16 ? n32 : n68747;
  assign n68749 = pi20 ? n61280 : n39805;
  assign n68750 = pi23 ? n8184 : n36781;
  assign n68751 = pi22 ? n68750 : n14626;
  assign n68752 = pi21 ? n68751 : n64278;
  assign n68753 = pi20 ? n68752 : n32;
  assign n68754 = pi19 ? n68749 : n68753;
  assign n68755 = pi18 ? n51733 : n68754;
  assign n68756 = pi17 ? n32 : n68755;
  assign n68757 = pi16 ? n32 : n68756;
  assign n68758 = pi15 ? n68748 : n68757;
  assign n68759 = pi21 ? n67832 : n36489;
  assign n68760 = pi21 ? n67811 : n47220;
  assign n68761 = pi20 ? n68759 : n68760;
  assign n68762 = pi22 ? n38284 : n51564;
  assign n68763 = pi21 ? n68762 : n64353;
  assign n68764 = pi20 ? n68763 : n32;
  assign n68765 = pi19 ? n68761 : n68764;
  assign n68766 = pi18 ? n51733 : n68765;
  assign n68767 = pi17 ? n32 : n68766;
  assign n68768 = pi16 ? n32 : n68767;
  assign n68769 = pi21 ? n33792 : n40986;
  assign n68770 = pi20 ? n51712 : n68769;
  assign n68771 = pi19 ? n68770 : n67836;
  assign n68772 = pi18 ? n51758 : n68771;
  assign n68773 = pi17 ? n32 : n68772;
  assign n68774 = pi16 ? n32 : n68773;
  assign n68775 = pi15 ? n68768 : n68774;
  assign n68776 = pi14 ? n68758 : n68775;
  assign n68777 = pi13 ? n68740 : n68776;
  assign n68778 = pi21 ? n20563 : n47360;
  assign n68779 = pi20 ? n20563 : n68778;
  assign n68780 = pi22 ? n49412 : n51564;
  assign n68781 = pi21 ? n68780 : n59357;
  assign n68782 = pi20 ? n68781 : n32;
  assign n68783 = pi19 ? n68779 : n68782;
  assign n68784 = pi18 ? n40056 : n68783;
  assign n68785 = pi17 ? n32 : n68784;
  assign n68786 = pi16 ? n32 : n68785;
  assign n68787 = pi21 ? n40986 : n38901;
  assign n68788 = pi20 ? n20563 : n68787;
  assign n68789 = pi19 ? n68788 : n67862;
  assign n68790 = pi18 ? n40056 : n68789;
  assign n68791 = pi17 ? n32 : n68790;
  assign n68792 = pi16 ? n32 : n68791;
  assign n68793 = pi15 ? n68786 : n68792;
  assign n68794 = pi21 ? n36798 : n37878;
  assign n68795 = pi20 ? n20563 : n68794;
  assign n68796 = pi22 ? n55622 : n57674;
  assign n68797 = pi21 ? n68796 : n37639;
  assign n68798 = pi20 ? n68797 : n32;
  assign n68799 = pi19 ? n68795 : n68798;
  assign n68800 = pi18 ? n40056 : n68799;
  assign n68801 = pi17 ? n32 : n68800;
  assign n68802 = pi16 ? n32 : n68801;
  assign n68803 = pi20 ? n20563 : n39973;
  assign n68804 = pi19 ? n68803 : n67383;
  assign n68805 = pi18 ? n40056 : n68804;
  assign n68806 = pi17 ? n32 : n68805;
  assign n68807 = pi16 ? n32 : n68806;
  assign n68808 = pi15 ? n68802 : n68807;
  assign n68809 = pi14 ? n68793 : n68808;
  assign n68810 = pi21 ? n62322 : n39972;
  assign n68811 = pi20 ? n20563 : n68810;
  assign n68812 = pi19 ? n68811 : n59650;
  assign n68813 = pi18 ? n40056 : n68812;
  assign n68814 = pi17 ? n32 : n68813;
  assign n68815 = pi16 ? n32 : n68814;
  assign n68816 = pi21 ? n61352 : n60591;
  assign n68817 = pi20 ? n20563 : n68816;
  assign n68818 = pi20 ? n61185 : n32;
  assign n68819 = pi19 ? n68817 : n68818;
  assign n68820 = pi18 ? n40056 : n68819;
  assign n68821 = pi17 ? n32 : n68820;
  assign n68822 = pi16 ? n32 : n68821;
  assign n68823 = pi15 ? n68815 : n68822;
  assign n68824 = pi22 ? n36798 : n62510;
  assign n68825 = pi21 ? n59524 : n68824;
  assign n68826 = pi20 ? n60502 : n68825;
  assign n68827 = pi19 ? n68826 : n56131;
  assign n68828 = pi18 ? n40056 : n68827;
  assign n68829 = pi17 ? n32 : n68828;
  assign n68830 = pi16 ? n32 : n68829;
  assign n68831 = pi22 ? n13481 : n14626;
  assign n68832 = pi21 ? n59524 : n68831;
  assign n68833 = pi20 ? n20563 : n68832;
  assign n68834 = pi19 ? n68833 : n56131;
  assign n68835 = pi18 ? n37935 : n68834;
  assign n68836 = pi17 ? n32 : n68835;
  assign n68837 = pi16 ? n32 : n68836;
  assign n68838 = pi15 ? n68830 : n68837;
  assign n68839 = pi14 ? n68823 : n68838;
  assign n68840 = pi13 ? n68809 : n68839;
  assign n68841 = pi12 ? n68777 : n68840;
  assign n68842 = pi22 ? n66956 : n13481;
  assign n68843 = pi21 ? n68842 : n13481;
  assign n68844 = pi20 ? n40791 : n68843;
  assign n68845 = pi19 ? n68844 : n37641;
  assign n68846 = pi18 ? n46063 : n68845;
  assign n68847 = pi17 ? n32 : n68846;
  assign n68848 = pi16 ? n32 : n68847;
  assign n68849 = pi22 ? n58710 : n51564;
  assign n68850 = pi21 ? n68849 : n51564;
  assign n68851 = pi20 ? n40791 : n68850;
  assign n68852 = pi19 ? n68851 : n35482;
  assign n68853 = pi18 ? n46063 : n68852;
  assign n68854 = pi17 ? n32 : n68853;
  assign n68855 = pi16 ? n32 : n68854;
  assign n68856 = pi15 ? n68848 : n68855;
  assign n68857 = pi22 ? n38284 : n13481;
  assign n68858 = pi21 ? n68857 : n57760;
  assign n68859 = pi20 ? n40791 : n68858;
  assign n68860 = pi19 ? n68859 : n35482;
  assign n68861 = pi18 ? n32 : n68860;
  assign n68862 = pi17 ? n32 : n68861;
  assign n68863 = pi16 ? n32 : n68862;
  assign n68864 = pi21 ? n36489 : n51313;
  assign n68865 = pi22 ? n36781 : n62389;
  assign n68866 = pi21 ? n68865 : n64278;
  assign n68867 = pi20 ? n68864 : n68866;
  assign n68868 = pi19 ? n68867 : n32;
  assign n68869 = pi18 ? n32 : n68868;
  assign n68870 = pi17 ? n32 : n68869;
  assign n68871 = pi16 ? n32 : n68870;
  assign n68872 = pi15 ? n68863 : n68871;
  assign n68873 = pi14 ? n68856 : n68872;
  assign n68874 = pi21 ? n36489 : n59524;
  assign n68875 = pi21 ? n47397 : n55560;
  assign n68876 = pi20 ? n68874 : n68875;
  assign n68877 = pi19 ? n68876 : n32;
  assign n68878 = pi18 ? n32 : n68877;
  assign n68879 = pi17 ? n32 : n68878;
  assign n68880 = pi16 ? n32 : n68879;
  assign n68881 = pi21 ? n48173 : n36798;
  assign n68882 = pi22 ? n36798 : n61484;
  assign n68883 = pi21 ? n68882 : n55560;
  assign n68884 = pi20 ? n68881 : n68883;
  assign n68885 = pi19 ? n68884 : n32;
  assign n68886 = pi18 ? n32 : n68885;
  assign n68887 = pi17 ? n32 : n68886;
  assign n68888 = pi16 ? n32 : n68887;
  assign n68889 = pi15 ? n68880 : n68888;
  assign n68890 = pi22 ? n52395 : n43198;
  assign n68891 = pi21 ? n47220 : n68890;
  assign n68892 = pi21 ? n61495 : n57097;
  assign n68893 = pi20 ? n68891 : n68892;
  assign n68894 = pi19 ? n68893 : n32;
  assign n68895 = pi18 ? n32 : n68894;
  assign n68896 = pi17 ? n32 : n68895;
  assign n68897 = pi16 ? n32 : n68896;
  assign n68898 = pi21 ? n42109 : n43198;
  assign n68899 = pi21 ? n67051 : n37639;
  assign n68900 = pi20 ? n68898 : n68899;
  assign n68901 = pi19 ? n68900 : n32;
  assign n68902 = pi18 ? n32 : n68901;
  assign n68903 = pi17 ? n32 : n68902;
  assign n68904 = pi16 ? n32 : n68903;
  assign n68905 = pi15 ? n68897 : n68904;
  assign n68906 = pi14 ? n68889 : n68905;
  assign n68907 = pi13 ? n68873 : n68906;
  assign n68908 = pi21 ? n33792 : n47397;
  assign n68909 = pi21 ? n63376 : n32;
  assign n68910 = pi20 ? n68908 : n68909;
  assign n68911 = pi19 ? n68910 : n32;
  assign n68912 = pi18 ? n32 : n68911;
  assign n68913 = pi17 ? n32 : n68912;
  assign n68914 = pi16 ? n32 : n68913;
  assign n68915 = pi22 ? n65218 : n21502;
  assign n68916 = pi21 ? n68915 : n32;
  assign n68917 = pi20 ? n68908 : n68916;
  assign n68918 = pi19 ? n68917 : n32;
  assign n68919 = pi18 ? n32 : n68918;
  assign n68920 = pi17 ? n32 : n68919;
  assign n68921 = pi16 ? n32 : n68920;
  assign n68922 = pi15 ? n68914 : n68921;
  assign n68923 = pi22 ? n32 : n49412;
  assign n68924 = pi21 ? n68923 : n61930;
  assign n68925 = pi20 ? n68924 : n68420;
  assign n68926 = pi19 ? n68925 : n32;
  assign n68927 = pi18 ? n32 : n68926;
  assign n68928 = pi17 ? n32 : n68927;
  assign n68929 = pi16 ? n32 : n68928;
  assign n68930 = pi21 ? n46727 : n14626;
  assign n68931 = pi20 ? n68930 : n56130;
  assign n68932 = pi19 ? n68931 : n32;
  assign n68933 = pi18 ? n32 : n68932;
  assign n68934 = pi17 ? n32 : n68933;
  assign n68935 = pi16 ? n32 : n68934;
  assign n68936 = pi15 ? n68929 : n68935;
  assign n68937 = pi14 ? n68922 : n68936;
  assign n68938 = pi22 ? n14626 : n57197;
  assign n68939 = pi21 ? n65284 : n68938;
  assign n68940 = pi20 ? n68939 : n60045;
  assign n68941 = pi19 ? n68940 : n32;
  assign n68942 = pi18 ? n32 : n68941;
  assign n68943 = pi17 ? n32 : n68942;
  assign n68944 = pi16 ? n32 : n68943;
  assign n68945 = pi21 ? n48856 : n57746;
  assign n68946 = pi20 ? n68945 : n20953;
  assign n68947 = pi19 ? n68946 : n32;
  assign n68948 = pi18 ? n32 : n68947;
  assign n68949 = pi17 ? n32 : n68948;
  assign n68950 = pi16 ? n32 : n68949;
  assign n68951 = pi15 ? n68944 : n68950;
  assign n68952 = pi21 ? n66139 : n62515;
  assign n68953 = pi20 ? n68952 : n32;
  assign n68954 = pi19 ? n68953 : n32;
  assign n68955 = pi18 ? n32 : n68954;
  assign n68956 = pi17 ? n32 : n68955;
  assign n68957 = pi16 ? n32 : n68956;
  assign n68958 = pi21 ? n63829 : n67007;
  assign n68959 = pi20 ? n68958 : n32;
  assign n68960 = pi19 ? n68959 : n32;
  assign n68961 = pi18 ? n32 : n68960;
  assign n68962 = pi17 ? n32 : n68961;
  assign n68963 = pi16 ? n32 : n68962;
  assign n68964 = pi15 ? n68957 : n68963;
  assign n68965 = pi14 ? n68951 : n68964;
  assign n68966 = pi13 ? n68937 : n68965;
  assign n68967 = pi12 ? n68907 : n68966;
  assign n68968 = pi11 ? n68841 : n68967;
  assign n68969 = pi10 ? n68704 : n68968;
  assign n68970 = pi09 ? n68481 : n68969;
  assign n68971 = pi20 ? n29133 : n13040;
  assign n68972 = pi19 ? n31264 : n68971;
  assign n68973 = pi18 ? n32 : n68972;
  assign n68974 = pi17 ? n32 : n68973;
  assign n68975 = pi16 ? n32 : n68974;
  assign n68976 = pi15 ? n32 : n68975;
  assign n68977 = pi19 ? n31264 : n61976;
  assign n68978 = pi18 ? n32 : n68977;
  assign n68979 = pi17 ? n32 : n68978;
  assign n68980 = pi16 ? n32 : n68979;
  assign n68981 = pi19 ? n31264 : n62975;
  assign n68982 = pi18 ? n32 : n68981;
  assign n68983 = pi17 ? n32 : n68982;
  assign n68984 = pi16 ? n32 : n68983;
  assign n68985 = pi15 ? n68980 : n68984;
  assign n68986 = pi14 ? n68976 : n68985;
  assign n68987 = pi13 ? n32 : n68986;
  assign n68988 = pi12 ? n32 : n68987;
  assign n68989 = pi11 ? n32 : n68988;
  assign n68990 = pi10 ? n32 : n68989;
  assign n68991 = pi20 ? n38477 : n1619;
  assign n68992 = pi19 ? n32401 : n68991;
  assign n68993 = pi18 ? n32 : n68992;
  assign n68994 = pi17 ? n32 : n68993;
  assign n68995 = pi16 ? n32 : n68994;
  assign n68996 = pi19 ? n43672 : n68490;
  assign n68997 = pi18 ? n32 : n68996;
  assign n68998 = pi17 ? n32 : n68997;
  assign n68999 = pi16 ? n32 : n68998;
  assign n69000 = pi15 ? n68995 : n68999;
  assign n69001 = pi14 ? n69000 : n68475;
  assign n69002 = pi22 ? n20563 : n60973;
  assign n69003 = pi21 ? n20563 : n69002;
  assign n69004 = pi20 ? n40054 : n69003;
  assign n69005 = pi19 ? n69004 : n68501;
  assign n69006 = pi18 ? n32 : n69005;
  assign n69007 = pi17 ? n32 : n69006;
  assign n69008 = pi16 ? n32 : n69007;
  assign n69009 = pi20 ? n36879 : n61008;
  assign n69010 = pi19 ? n40509 : n69009;
  assign n69011 = pi18 ? n32 : n69010;
  assign n69012 = pi17 ? n32 : n69011;
  assign n69013 = pi16 ? n32 : n69012;
  assign n69014 = pi15 ? n69008 : n69013;
  assign n69015 = pi19 ? n40509 : n62975;
  assign n69016 = pi18 ? n32 : n69015;
  assign n69017 = pi17 ? n32 : n69016;
  assign n69018 = pi16 ? n32 : n69017;
  assign n69019 = pi14 ? n69014 : n69018;
  assign n69020 = pi13 ? n69001 : n69019;
  assign n69021 = pi19 ? n39372 : n68519;
  assign n69022 = pi18 ? n32 : n69021;
  assign n69023 = pi17 ? n32 : n69022;
  assign n69024 = pi16 ? n32 : n69023;
  assign n69025 = pi19 ? n39372 : n68490;
  assign n69026 = pi18 ? n32 : n69025;
  assign n69027 = pi17 ? n32 : n69026;
  assign n69028 = pi16 ? n32 : n69027;
  assign n69029 = pi15 ? n69024 : n69028;
  assign n69030 = pi14 ? n69029 : n68083;
  assign n69031 = pi19 ? n39372 : n68530;
  assign n69032 = pi18 ? n32 : n69031;
  assign n69033 = pi17 ? n32 : n69032;
  assign n69034 = pi16 ? n32 : n69033;
  assign n69035 = pi20 ? n37955 : n38754;
  assign n69036 = pi19 ? n69035 : n68536;
  assign n69037 = pi18 ? n32 : n69036;
  assign n69038 = pi17 ? n32 : n69037;
  assign n69039 = pi16 ? n32 : n69038;
  assign n69040 = pi15 ? n69034 : n69039;
  assign n69041 = pi19 ? n69035 : n68543;
  assign n69042 = pi18 ? n32 : n69041;
  assign n69043 = pi17 ? n32 : n69042;
  assign n69044 = pi16 ? n32 : n69043;
  assign n69045 = pi22 ? n17226 : n51564;
  assign n69046 = pi21 ? n69045 : n58778;
  assign n69047 = pi20 ? n47158 : n69046;
  assign n69048 = pi19 ? n43246 : n69047;
  assign n69049 = pi18 ? n32 : n69048;
  assign n69050 = pi17 ? n32 : n69049;
  assign n69051 = pi16 ? n32 : n69050;
  assign n69052 = pi15 ? n69044 : n69051;
  assign n69053 = pi14 ? n69040 : n69052;
  assign n69054 = pi13 ? n69030 : n69053;
  assign n69055 = pi12 ? n69020 : n69054;
  assign n69056 = pi20 ? n37320 : n67569;
  assign n69057 = pi21 ? n31889 : n53366;
  assign n69058 = pi20 ? n69057 : n68566;
  assign n69059 = pi19 ? n69056 : n69058;
  assign n69060 = pi18 ? n32 : n69059;
  assign n69061 = pi17 ? n32 : n69060;
  assign n69062 = pi16 ? n32 : n69061;
  assign n69063 = pi24 ? n363 : n13481;
  assign n69064 = pi23 ? n69063 : n13481;
  assign n69065 = pi22 ? n69064 : n13481;
  assign n69066 = pi21 ? n69065 : n55560;
  assign n69067 = pi20 ? n55475 : n69066;
  assign n69068 = pi19 ? n38947 : n69067;
  assign n69069 = pi18 ? n32 : n69068;
  assign n69070 = pi17 ? n32 : n69069;
  assign n69071 = pi16 ? n32 : n69070;
  assign n69072 = pi15 ? n69062 : n69071;
  assign n69073 = pi19 ? n38947 : n68580;
  assign n69074 = pi18 ? n32 : n69073;
  assign n69075 = pi17 ? n32 : n69074;
  assign n69076 = pi16 ? n32 : n69075;
  assign n69077 = pi21 ? n30868 : n66686;
  assign n69078 = pi20 ? n69077 : n27076;
  assign n69079 = pi19 ? n38947 : n69078;
  assign n69080 = pi18 ? n32 : n69079;
  assign n69081 = pi17 ? n32 : n69080;
  assign n69082 = pi16 ? n32 : n69081;
  assign n69083 = pi15 ? n69076 : n69082;
  assign n69084 = pi14 ? n69072 : n69083;
  assign n69085 = pi20 ? n37320 : n38754;
  assign n69086 = pi19 ? n69085 : n68597;
  assign n69087 = pi18 ? n32 : n69086;
  assign n69088 = pi17 ? n32 : n69087;
  assign n69089 = pi16 ? n32 : n69088;
  assign n69090 = pi20 ? n37320 : n68603;
  assign n69091 = pi19 ? n69090 : n68607;
  assign n69092 = pi18 ? n32 : n69091;
  assign n69093 = pi17 ? n32 : n69092;
  assign n69094 = pi16 ? n32 : n69093;
  assign n69095 = pi15 ? n69089 : n69094;
  assign n69096 = pi20 ? n37333 : n54998;
  assign n69097 = pi19 ? n69096 : n68616;
  assign n69098 = pi18 ? n32 : n69097;
  assign n69099 = pi17 ? n32 : n69098;
  assign n69100 = pi16 ? n32 : n69099;
  assign n69101 = pi20 ? n38376 : n55014;
  assign n69102 = pi20 ? n68623 : n17510;
  assign n69103 = pi19 ? n69101 : n69102;
  assign n69104 = pi18 ? n32 : n69103;
  assign n69105 = pi17 ? n32 : n69104;
  assign n69106 = pi16 ? n32 : n69105;
  assign n69107 = pi15 ? n69100 : n69106;
  assign n69108 = pi14 ? n69095 : n69107;
  assign n69109 = pi13 ? n69084 : n69108;
  assign n69110 = pi19 ? n39396 : n68636;
  assign n69111 = pi18 ? n32 : n69110;
  assign n69112 = pi17 ? n32 : n69111;
  assign n69113 = pi16 ? n32 : n69112;
  assign n69114 = pi20 ? n39395 : n40791;
  assign n69115 = pi19 ? n69114 : n68645;
  assign n69116 = pi18 ? n32 : n69115;
  assign n69117 = pi17 ? n32 : n69116;
  assign n69118 = pi16 ? n32 : n69117;
  assign n69119 = pi15 ? n69113 : n69118;
  assign n69120 = pi19 ? n69114 : n68654;
  assign n69121 = pi18 ? n32 : n69120;
  assign n69122 = pi17 ? n32 : n69121;
  assign n69123 = pi16 ? n32 : n69122;
  assign n69124 = pi19 ? n39396 : n68662;
  assign n69125 = pi18 ? n32 : n69124;
  assign n69126 = pi17 ? n32 : n69125;
  assign n69127 = pi16 ? n32 : n69126;
  assign n69128 = pi15 ? n69123 : n69127;
  assign n69129 = pi14 ? n69119 : n69128;
  assign n69130 = pi20 ? n68670 : n6417;
  assign n69131 = pi19 ? n39396 : n69130;
  assign n69132 = pi18 ? n32 : n69131;
  assign n69133 = pi17 ? n32 : n69132;
  assign n69134 = pi16 ? n32 : n69133;
  assign n69135 = pi19 ? n39396 : n68680;
  assign n69136 = pi18 ? n32 : n69135;
  assign n69137 = pi17 ? n32 : n69136;
  assign n69138 = pi16 ? n32 : n69137;
  assign n69139 = pi15 ? n69134 : n69138;
  assign n69140 = pi19 ? n68594 : n68688;
  assign n69141 = pi18 ? n32 : n69140;
  assign n69142 = pi17 ? n32 : n69141;
  assign n69143 = pi16 ? n32 : n69142;
  assign n69144 = pi19 ? n42192 : n68695;
  assign n69145 = pi18 ? n32 : n69144;
  assign n69146 = pi17 ? n32 : n69145;
  assign n69147 = pi16 ? n32 : n69146;
  assign n69148 = pi15 ? n69143 : n69147;
  assign n69149 = pi14 ? n69139 : n69148;
  assign n69150 = pi13 ? n69129 : n69149;
  assign n69151 = pi12 ? n69109 : n69150;
  assign n69152 = pi11 ? n69055 : n69151;
  assign n69153 = pi21 ? n30116 : n36489;
  assign n69154 = pi20 ? n69153 : n40915;
  assign n69155 = pi19 ? n69154 : n68708;
  assign n69156 = pi18 ? n32 : n69155;
  assign n69157 = pi17 ? n32 : n69156;
  assign n69158 = pi16 ? n32 : n69157;
  assign n69159 = pi22 ? n37240 : n36781;
  assign n69160 = pi21 ? n69159 : n68714;
  assign n69161 = pi20 ? n69160 : n32;
  assign n69162 = pi19 ? n46700 : n69161;
  assign n69163 = pi18 ? n32 : n69162;
  assign n69164 = pi17 ? n32 : n69163;
  assign n69165 = pi16 ? n32 : n69164;
  assign n69166 = pi15 ? n69158 : n69165;
  assign n69167 = pi21 ? n46166 : n45016;
  assign n69168 = pi20 ? n69167 : n47223;
  assign n69169 = pi19 ? n69168 : n68727;
  assign n69170 = pi18 ? n32 : n69169;
  assign n69171 = pi17 ? n32 : n69170;
  assign n69172 = pi16 ? n32 : n69171;
  assign n69173 = pi21 ? n54400 : n20563;
  assign n69174 = pi20 ? n69173 : n20563;
  assign n69175 = pi21 ? n60543 : n65478;
  assign n69176 = pi20 ? n69175 : n32;
  assign n69177 = pi19 ? n69174 : n69176;
  assign n69178 = pi18 ? n32 : n69177;
  assign n69179 = pi17 ? n32 : n69178;
  assign n69180 = pi16 ? n32 : n69179;
  assign n69181 = pi15 ? n69172 : n69180;
  assign n69182 = pi14 ? n69166 : n69181;
  assign n69183 = pi21 ? n54427 : n39801;
  assign n69184 = pi20 ? n69183 : n41912;
  assign n69185 = pi23 ? n56478 : n36659;
  assign n69186 = pi22 ? n69185 : n14626;
  assign n69187 = pi21 ? n69186 : n63376;
  assign n69188 = pi20 ? n69187 : n32;
  assign n69189 = pi19 ? n69184 : n69188;
  assign n69190 = pi18 ? n32 : n69189;
  assign n69191 = pi17 ? n32 : n69190;
  assign n69192 = pi16 ? n32 : n69191;
  assign n69193 = pi22 ? n46757 : n33792;
  assign n69194 = pi21 ? n69193 : n37768;
  assign n69195 = pi20 ? n69194 : n39805;
  assign n69196 = pi22 ? n58519 : n14626;
  assign n69197 = pi21 ? n69196 : n59648;
  assign n69198 = pi20 ? n69197 : n32;
  assign n69199 = pi19 ? n69195 : n69198;
  assign n69200 = pi18 ? n32 : n69199;
  assign n69201 = pi17 ? n32 : n69200;
  assign n69202 = pi16 ? n32 : n69201;
  assign n69203 = pi15 ? n69192 : n69202;
  assign n69204 = pi22 ? n51754 : n33792;
  assign n69205 = pi21 ? n69204 : n64086;
  assign n69206 = pi20 ? n69205 : n68760;
  assign n69207 = pi23 ? n63194 : n36781;
  assign n69208 = pi22 ? n69207 : n51564;
  assign n69209 = pi21 ? n69208 : n57458;
  assign n69210 = pi20 ? n69209 : n32;
  assign n69211 = pi19 ? n69206 : n69210;
  assign n69212 = pi18 ? n32 : n69211;
  assign n69213 = pi17 ? n32 : n69212;
  assign n69214 = pi16 ? n32 : n69213;
  assign n69215 = pi20 ? n36490 : n68769;
  assign n69216 = pi21 ? n68780 : n2637;
  assign n69217 = pi20 ? n69216 : n32;
  assign n69218 = pi19 ? n69215 : n69217;
  assign n69219 = pi18 ? n32 : n69218;
  assign n69220 = pi17 ? n32 : n69219;
  assign n69221 = pi16 ? n32 : n69220;
  assign n69222 = pi15 ? n69214 : n69221;
  assign n69223 = pi14 ? n69203 : n69222;
  assign n69224 = pi13 ? n69182 : n69223;
  assign n69225 = pi20 ? n31313 : n68778;
  assign n69226 = pi21 ? n59681 : n59357;
  assign n69227 = pi20 ? n69226 : n32;
  assign n69228 = pi19 ? n69225 : n69227;
  assign n69229 = pi18 ? n32 : n69228;
  assign n69230 = pi17 ? n32 : n69229;
  assign n69231 = pi16 ? n32 : n69230;
  assign n69232 = pi20 ? n31313 : n68787;
  assign n69233 = pi19 ? n69232 : n67862;
  assign n69234 = pi18 ? n32 : n69233;
  assign n69235 = pi17 ? n32 : n69234;
  assign n69236 = pi16 ? n32 : n69235;
  assign n69237 = pi15 ? n69231 : n69236;
  assign n69238 = pi20 ? n31313 : n68794;
  assign n69239 = pi22 ? n55641 : n57674;
  assign n69240 = pi21 ? n69239 : n37639;
  assign n69241 = pi20 ? n69240 : n32;
  assign n69242 = pi19 ? n69238 : n69241;
  assign n69243 = pi18 ? n32 : n69242;
  assign n69244 = pi17 ? n32 : n69243;
  assign n69245 = pi16 ? n32 : n69244;
  assign n69246 = pi20 ? n31313 : n39973;
  assign n69247 = pi19 ? n69246 : n62851;
  assign n69248 = pi18 ? n32 : n69247;
  assign n69249 = pi17 ? n32 : n69248;
  assign n69250 = pi16 ? n32 : n69249;
  assign n69251 = pi15 ? n69245 : n69250;
  assign n69252 = pi14 ? n69237 : n69251;
  assign n69253 = pi20 ? n31313 : n68810;
  assign n69254 = pi19 ? n69253 : n59650;
  assign n69255 = pi18 ? n32 : n69254;
  assign n69256 = pi17 ? n32 : n69255;
  assign n69257 = pi16 ? n32 : n69256;
  assign n69258 = pi22 ? n36798 : n55766;
  assign n69259 = pi21 ? n61352 : n69258;
  assign n69260 = pi20 ? n30117 : n69259;
  assign n69261 = pi19 ? n69260 : n68818;
  assign n69262 = pi18 ? n32 : n69261;
  assign n69263 = pi17 ? n32 : n69262;
  assign n69264 = pi16 ? n32 : n69263;
  assign n69265 = pi15 ? n69257 : n69264;
  assign n69266 = pi21 ? n59524 : n55708;
  assign n69267 = pi20 ? n37806 : n69266;
  assign n69268 = pi19 ? n69267 : n56131;
  assign n69269 = pi18 ? n32 : n69268;
  assign n69270 = pi17 ? n32 : n69269;
  assign n69271 = pi16 ? n32 : n69270;
  assign n69272 = pi22 ? n13481 : n62803;
  assign n69273 = pi21 ? n59524 : n69272;
  assign n69274 = pi20 ? n69173 : n69273;
  assign n69275 = pi19 ? n69274 : n56131;
  assign n69276 = pi18 ? n32 : n69275;
  assign n69277 = pi17 ? n32 : n69276;
  assign n69278 = pi16 ? n32 : n69277;
  assign n69279 = pi15 ? n69271 : n69278;
  assign n69280 = pi14 ? n69265 : n69279;
  assign n69281 = pi13 ? n69252 : n69280;
  assign n69282 = pi12 ? n69224 : n69281;
  assign n69283 = pi21 ? n54400 : n30868;
  assign n69284 = pi23 ? n56064 : n36659;
  assign n69285 = pi22 ? n69284 : n13481;
  assign n69286 = pi21 ? n69285 : n13481;
  assign n69287 = pi20 ? n69283 : n69286;
  assign n69288 = pi19 ? n69287 : n37641;
  assign n69289 = pi18 ? n32 : n69288;
  assign n69290 = pi17 ? n32 : n69289;
  assign n69291 = pi16 ? n32 : n69290;
  assign n69292 = pi22 ? n36659 : n51564;
  assign n69293 = pi22 ? n51564 : n56186;
  assign n69294 = pi21 ? n69292 : n69293;
  assign n69295 = pi20 ? n62373 : n69294;
  assign n69296 = pi19 ? n69295 : n35482;
  assign n69297 = pi18 ? n32 : n69296;
  assign n69298 = pi17 ? n32 : n69297;
  assign n69299 = pi16 ? n32 : n69298;
  assign n69300 = pi15 ? n69291 : n69299;
  assign n69301 = pi22 ? n36781 : n13481;
  assign n69302 = pi21 ? n69301 : n57760;
  assign n69303 = pi20 ? n62373 : n69302;
  assign n69304 = pi19 ? n69303 : n35482;
  assign n69305 = pi18 ? n32 : n69304;
  assign n69306 = pi17 ? n32 : n69305;
  assign n69307 = pi16 ? n32 : n69306;
  assign n69308 = pi21 ? n46060 : n51313;
  assign n69309 = pi21 ? n68865 : n59648;
  assign n69310 = pi20 ? n69308 : n69309;
  assign n69311 = pi19 ? n69310 : n32;
  assign n69312 = pi18 ? n32 : n69311;
  assign n69313 = pi17 ? n32 : n69312;
  assign n69314 = pi16 ? n32 : n69313;
  assign n69315 = pi15 ? n69307 : n69314;
  assign n69316 = pi14 ? n69300 : n69315;
  assign n69317 = pi21 ? n46060 : n59524;
  assign n69318 = pi22 ? n36798 : n54664;
  assign n69319 = pi21 ? n69318 : n55560;
  assign n69320 = pi20 ? n69317 : n69319;
  assign n69321 = pi19 ? n69320 : n32;
  assign n69322 = pi18 ? n32 : n69321;
  assign n69323 = pi17 ? n32 : n69322;
  assign n69324 = pi16 ? n32 : n69323;
  assign n69325 = pi22 ? n32 : n42109;
  assign n69326 = pi21 ? n69325 : n36798;
  assign n69327 = pi22 ? n36798 : n56622;
  assign n69328 = pi21 ? n69327 : n55560;
  assign n69329 = pi20 ? n69326 : n69328;
  assign n69330 = pi19 ? n69329 : n32;
  assign n69331 = pi18 ? n32 : n69330;
  assign n69332 = pi17 ? n32 : n69331;
  assign n69333 = pi16 ? n32 : n69332;
  assign n69334 = pi15 ? n69324 : n69333;
  assign n69335 = pi21 ? n52259 : n68890;
  assign n69336 = pi21 ? n63771 : n57097;
  assign n69337 = pi20 ? n69335 : n69336;
  assign n69338 = pi19 ? n69337 : n32;
  assign n69339 = pi18 ? n32 : n69338;
  assign n69340 = pi17 ? n32 : n69339;
  assign n69341 = pi16 ? n32 : n69340;
  assign n69342 = pi23 ? n13481 : n14626;
  assign n69343 = pi22 ? n69342 : n13481;
  assign n69344 = pi21 ? n69343 : n37639;
  assign n69345 = pi20 ? n46791 : n69344;
  assign n69346 = pi19 ? n69345 : n32;
  assign n69347 = pi18 ? n32 : n69346;
  assign n69348 = pi17 ? n32 : n69347;
  assign n69349 = pi16 ? n32 : n69348;
  assign n69350 = pi15 ? n69341 : n69349;
  assign n69351 = pi14 ? n69334 : n69350;
  assign n69352 = pi13 ? n69316 : n69351;
  assign n69353 = pi21 ? n46276 : n47397;
  assign n69354 = pi22 ? n66042 : n57647;
  assign n69355 = pi21 ? n69354 : n32;
  assign n69356 = pi20 ? n69353 : n69355;
  assign n69357 = pi19 ? n69356 : n32;
  assign n69358 = pi18 ? n32 : n69357;
  assign n69359 = pi17 ? n32 : n69358;
  assign n69360 = pi16 ? n32 : n69359;
  assign n69361 = pi21 ? n32 : n47397;
  assign n69362 = pi22 ? n66042 : n21502;
  assign n69363 = pi21 ? n69362 : n32;
  assign n69364 = pi20 ? n69361 : n69363;
  assign n69365 = pi19 ? n69364 : n32;
  assign n69366 = pi18 ? n32 : n69365;
  assign n69367 = pi17 ? n32 : n69366;
  assign n69368 = pi16 ? n32 : n69367;
  assign n69369 = pi15 ? n69360 : n69368;
  assign n69370 = pi21 ? n63433 : n61930;
  assign n69371 = pi23 ? n63306 : n13481;
  assign n69372 = pi22 ? n69371 : n21502;
  assign n69373 = pi21 ? n69372 : n32;
  assign n69374 = pi20 ? n69370 : n69373;
  assign n69375 = pi19 ? n69374 : n32;
  assign n69376 = pi18 ? n32 : n69375;
  assign n69377 = pi17 ? n32 : n69376;
  assign n69378 = pi16 ? n32 : n69377;
  assign n69379 = pi20 ? n66541 : n60045;
  assign n69380 = pi19 ? n69379 : n32;
  assign n69381 = pi18 ? n32 : n69380;
  assign n69382 = pi17 ? n32 : n69381;
  assign n69383 = pi16 ? n32 : n69382;
  assign n69384 = pi15 ? n69378 : n69383;
  assign n69385 = pi14 ? n69369 : n69384;
  assign n69386 = pi21 ? n32 : n59595;
  assign n69387 = pi20 ? n69386 : n37640;
  assign n69388 = pi19 ? n69387 : n32;
  assign n69389 = pi18 ? n32 : n69388;
  assign n69390 = pi17 ? n32 : n69389;
  assign n69391 = pi16 ? n32 : n69390;
  assign n69392 = pi22 ? n56622 : n13481;
  assign n69393 = pi21 ? n32 : n69392;
  assign n69394 = pi20 ? n69393 : n20953;
  assign n69395 = pi19 ? n69394 : n32;
  assign n69396 = pi18 ? n32 : n69395;
  assign n69397 = pi17 ? n32 : n69396;
  assign n69398 = pi16 ? n32 : n69397;
  assign n69399 = pi15 ? n69391 : n69398;
  assign n69400 = pi24 ? n32 : n13481;
  assign n69401 = pi23 ? n32 : n69400;
  assign n69402 = pi22 ? n69401 : n13481;
  assign n69403 = pi21 ? n32 : n69402;
  assign n69404 = pi20 ? n69403 : n32;
  assign n69405 = pi19 ? n69404 : n32;
  assign n69406 = pi18 ? n32 : n69405;
  assign n69407 = pi17 ? n32 : n69406;
  assign n69408 = pi16 ? n32 : n69407;
  assign n69409 = pi22 ? n32 : n56665;
  assign n69410 = pi21 ? n32 : n69409;
  assign n69411 = pi20 ? n69410 : n32;
  assign n69412 = pi19 ? n69411 : n32;
  assign n69413 = pi18 ? n32 : n69412;
  assign n69414 = pi17 ? n32 : n69413;
  assign n69415 = pi16 ? n32 : n69414;
  assign n69416 = pi15 ? n69408 : n69415;
  assign n69417 = pi14 ? n69399 : n69416;
  assign n69418 = pi13 ? n69385 : n69417;
  assign n69419 = pi12 ? n69352 : n69418;
  assign n69420 = pi11 ? n69282 : n69419;
  assign n69421 = pi10 ? n69152 : n69420;
  assign n69422 = pi09 ? n68990 : n69421;
  assign n69423 = pi08 ? n68970 : n69422;
  assign n69424 = pi20 ? n31266 : n13040;
  assign n69425 = pi19 ? n39454 : n69424;
  assign n69426 = pi18 ? n32 : n69425;
  assign n69427 = pi17 ? n32 : n69426;
  assign n69428 = pi16 ? n32 : n69427;
  assign n69429 = pi15 ? n32 : n69428;
  assign n69430 = pi19 ? n39454 : n61976;
  assign n69431 = pi18 ? n32 : n69430;
  assign n69432 = pi17 ? n32 : n69431;
  assign n69433 = pi16 ? n32 : n69432;
  assign n69434 = pi19 ? n39454 : n62975;
  assign n69435 = pi18 ? n32 : n69434;
  assign n69436 = pi17 ? n32 : n69435;
  assign n69437 = pi16 ? n32 : n69436;
  assign n69438 = pi15 ? n69433 : n69437;
  assign n69439 = pi14 ? n69429 : n69438;
  assign n69440 = pi13 ? n32 : n69439;
  assign n69441 = pi12 ? n32 : n69440;
  assign n69442 = pi11 ? n32 : n69441;
  assign n69443 = pi10 ? n32 : n69442;
  assign n69444 = pi19 ? n28158 : n62975;
  assign n69445 = pi18 ? n32 : n69444;
  assign n69446 = pi17 ? n32 : n69445;
  assign n69447 = pi16 ? n32 : n69446;
  assign n69448 = pi19 ? n30118 : n62975;
  assign n69449 = pi18 ? n32 : n69448;
  assign n69450 = pi17 ? n32 : n69449;
  assign n69451 = pi16 ? n32 : n69450;
  assign n69452 = pi15 ? n69447 : n69451;
  assign n69453 = pi14 ? n69452 : n68984;
  assign n69454 = pi21 ? n68483 : n29133;
  assign n69455 = pi20 ? n69454 : n61008;
  assign n69456 = pi19 ? n40496 : n69455;
  assign n69457 = pi18 ? n32 : n69456;
  assign n69458 = pi17 ? n32 : n69457;
  assign n69459 = pi16 ? n32 : n69458;
  assign n69460 = pi19 ? n40496 : n67606;
  assign n69461 = pi18 ? n32 : n69460;
  assign n69462 = pi17 ? n32 : n69461;
  assign n69463 = pi16 ? n32 : n69462;
  assign n69464 = pi15 ? n69459 : n69463;
  assign n69465 = pi14 ? n69464 : n68499;
  assign n69466 = pi13 ? n69453 : n69465;
  assign n69467 = pi15 ? n68499 : n68062;
  assign n69468 = pi14 ? n68499 : n69467;
  assign n69469 = pi20 ? n31266 : n59305;
  assign n69470 = pi19 ? n40509 : n69469;
  assign n69471 = pi18 ? n32 : n69470;
  assign n69472 = pi17 ? n32 : n69471;
  assign n69473 = pi16 ? n32 : n69472;
  assign n69474 = pi24 ? n30868 : n233;
  assign n69475 = pi23 ? n69474 : n233;
  assign n69476 = pi22 ? n69475 : n233;
  assign n69477 = pi21 ? n69476 : n650;
  assign n69478 = pi20 ? n38754 : n69477;
  assign n69479 = pi19 ? n56095 : n69478;
  assign n69480 = pi18 ? n32 : n69479;
  assign n69481 = pi17 ? n32 : n69480;
  assign n69482 = pi16 ? n32 : n69481;
  assign n69483 = pi15 ? n69473 : n69482;
  assign n69484 = pi21 ? n68139 : n696;
  assign n69485 = pi20 ? n40791 : n69484;
  assign n69486 = pi19 ? n56095 : n69485;
  assign n69487 = pi18 ? n32 : n69486;
  assign n69488 = pi17 ? n32 : n69487;
  assign n69489 = pi16 ? n32 : n69488;
  assign n69490 = pi24 ? n335 : n51564;
  assign n69491 = pi23 ? n69490 : n51564;
  assign n69492 = pi22 ? n69491 : n51564;
  assign n69493 = pi21 ? n69492 : n58778;
  assign n69494 = pi20 ? n47158 : n69493;
  assign n69495 = pi19 ? n40509 : n69494;
  assign n69496 = pi18 ? n32 : n69495;
  assign n69497 = pi17 ? n32 : n69496;
  assign n69498 = pi16 ? n32 : n69497;
  assign n69499 = pi15 ? n69489 : n69498;
  assign n69500 = pi14 ? n69483 : n69499;
  assign n69501 = pi13 ? n69468 : n69500;
  assign n69502 = pi12 ? n69466 : n69501;
  assign n69503 = pi21 ? n36249 : n53366;
  assign n69504 = pi20 ? n69503 : n68566;
  assign n69505 = pi19 ? n39372 : n69504;
  assign n69506 = pi18 ? n32 : n69505;
  assign n69507 = pi17 ? n32 : n69506;
  assign n69508 = pi16 ? n32 : n69507;
  assign n69509 = pi19 ? n39372 : n69067;
  assign n69510 = pi18 ? n32 : n69509;
  assign n69511 = pi17 ? n32 : n69510;
  assign n69512 = pi16 ? n32 : n69511;
  assign n69513 = pi15 ? n69508 : n69512;
  assign n69514 = pi19 ? n39372 : n68580;
  assign n69515 = pi18 ? n32 : n69514;
  assign n69516 = pi17 ? n32 : n69515;
  assign n69517 = pi16 ? n32 : n69516;
  assign n69518 = pi21 ? n30868 : n65740;
  assign n69519 = pi20 ? n69518 : n63941;
  assign n69520 = pi19 ? n39372 : n69519;
  assign n69521 = pi18 ? n32 : n69520;
  assign n69522 = pi17 ? n32 : n69521;
  assign n69523 = pi16 ? n32 : n69522;
  assign n69524 = pi15 ? n69517 : n69523;
  assign n69525 = pi14 ? n69513 : n69524;
  assign n69526 = pi20 ? n37933 : n38754;
  assign n69527 = pi19 ? n69526 : n67669;
  assign n69528 = pi18 ? n32 : n69527;
  assign n69529 = pi17 ? n32 : n69528;
  assign n69530 = pi16 ? n32 : n69529;
  assign n69531 = pi20 ? n36867 : n47158;
  assign n69532 = pi21 ? n33792 : n65752;
  assign n69533 = pi20 ? n69532 : n63066;
  assign n69534 = pi19 ? n69531 : n69533;
  assign n69535 = pi18 ? n32 : n69534;
  assign n69536 = pi17 ? n32 : n69535;
  assign n69537 = pi16 ? n32 : n69536;
  assign n69538 = pi15 ? n69530 : n69537;
  assign n69539 = pi23 ? n30868 : n363;
  assign n69540 = pi22 ? n30868 : n69539;
  assign n69541 = pi21 ? n30868 : n69540;
  assign n69542 = pi20 ? n69541 : n58439;
  assign n69543 = pi19 ? n40531 : n69542;
  assign n69544 = pi18 ? n32 : n69543;
  assign n69545 = pi17 ? n32 : n69544;
  assign n69546 = pi16 ? n32 : n69545;
  assign n69547 = pi23 ? n33792 : n233;
  assign n69548 = pi22 ? n30869 : n69547;
  assign n69549 = pi21 ? n30868 : n69548;
  assign n69550 = pi20 ? n69549 : n17510;
  assign n69551 = pi19 ? n41707 : n69550;
  assign n69552 = pi18 ? n32 : n69551;
  assign n69553 = pi17 ? n32 : n69552;
  assign n69554 = pi16 ? n32 : n69553;
  assign n69555 = pi15 ? n69546 : n69554;
  assign n69556 = pi14 ? n69538 : n69555;
  assign n69557 = pi13 ? n69525 : n69556;
  assign n69558 = pi23 ? n33792 : n157;
  assign n69559 = pi22 ? n36617 : n69558;
  assign n69560 = pi21 ? n20563 : n69559;
  assign n69561 = pi20 ? n69560 : n67712;
  assign n69562 = pi19 ? n43246 : n69561;
  assign n69563 = pi18 ? n32 : n69562;
  assign n69564 = pi17 ? n32 : n69563;
  assign n69565 = pi16 ? n32 : n69564;
  assign n69566 = pi20 ? n38997 : n40791;
  assign n69567 = pi24 ? n37 : n33792;
  assign n69568 = pi23 ? n20563 : n69567;
  assign n69569 = pi22 ? n69568 : n66744;
  assign n69570 = pi21 ? n30868 : n69569;
  assign n69571 = pi20 ? n69570 : n67719;
  assign n69572 = pi19 ? n69566 : n69571;
  assign n69573 = pi18 ? n32 : n69572;
  assign n69574 = pi17 ? n32 : n69573;
  assign n69575 = pi16 ? n32 : n69574;
  assign n69576 = pi15 ? n69565 : n69575;
  assign n69577 = pi23 ? n36659 : n204;
  assign n69578 = pi22 ? n37783 : n69577;
  assign n69579 = pi21 ? n30868 : n69578;
  assign n69580 = pi20 ? n69579 : n68653;
  assign n69581 = pi19 ? n69566 : n69580;
  assign n69582 = pi18 ? n32 : n69581;
  assign n69583 = pi17 ? n32 : n69582;
  assign n69584 = pi16 ? n32 : n69583;
  assign n69585 = pi20 ? n38997 : n51223;
  assign n69586 = pi22 ? n46172 : n67736;
  assign n69587 = pi21 ? n33792 : n69586;
  assign n69588 = pi20 ? n69587 : n59649;
  assign n69589 = pi19 ? n69585 : n69588;
  assign n69590 = pi18 ? n32 : n69589;
  assign n69591 = pi17 ? n32 : n69590;
  assign n69592 = pi16 ? n32 : n69591;
  assign n69593 = pi15 ? n69584 : n69592;
  assign n69594 = pi14 ? n69576 : n69593;
  assign n69595 = pi23 ? n36781 : n233;
  assign n69596 = pi22 ? n69539 : n69595;
  assign n69597 = pi21 ? n36659 : n69596;
  assign n69598 = pi20 ? n69597 : n6417;
  assign n69599 = pi19 ? n43246 : n69598;
  assign n69600 = pi18 ? n32 : n69599;
  assign n69601 = pi17 ? n32 : n69600;
  assign n69602 = pi16 ? n32 : n69601;
  assign n69603 = pi22 ? n59056 : n20563;
  assign n69604 = pi21 ? n20563 : n69603;
  assign n69605 = pi20 ? n38997 : n69604;
  assign n69606 = pi22 ? n54574 : n57632;
  assign n69607 = pi21 ? n36659 : n69606;
  assign n69608 = pi20 ? n69607 : n58168;
  assign n69609 = pi19 ? n69605 : n69608;
  assign n69610 = pi18 ? n32 : n69609;
  assign n69611 = pi17 ? n32 : n69610;
  assign n69612 = pi16 ? n32 : n69611;
  assign n69613 = pi15 ? n69602 : n69612;
  assign n69614 = pi23 ? n37 : n55501;
  assign n69615 = pi22 ? n69614 : n20563;
  assign n69616 = pi21 ? n20563 : n69615;
  assign n69617 = pi20 ? n37320 : n69616;
  assign n69618 = pi21 ? n36659 : n63329;
  assign n69619 = pi20 ? n69618 : n54565;
  assign n69620 = pi19 ? n69617 : n69619;
  assign n69621 = pi18 ? n32 : n69620;
  assign n69622 = pi17 ? n32 : n69621;
  assign n69623 = pi16 ? n32 : n69622;
  assign n69624 = pi22 ? n50339 : n62880;
  assign n69625 = pi21 ? n36659 : n69624;
  assign n69626 = pi20 ? n69625 : n32257;
  assign n69627 = pi19 ? n38956 : n69626;
  assign n69628 = pi18 ? n32 : n69627;
  assign n69629 = pi17 ? n32 : n69628;
  assign n69630 = pi16 ? n32 : n69629;
  assign n69631 = pi15 ? n69623 : n69630;
  assign n69632 = pi14 ? n69613 : n69631;
  assign n69633 = pi13 ? n69594 : n69632;
  assign n69634 = pi12 ? n69557 : n69633;
  assign n69635 = pi11 ? n69502 : n69634;
  assign n69636 = pi20 ? n59665 : n41463;
  assign n69637 = pi22 ? n69595 : n13481;
  assign n69638 = pi21 ? n51564 : n69637;
  assign n69639 = pi20 ? n69638 : n37640;
  assign n69640 = pi19 ? n69636 : n69639;
  assign n69641 = pi18 ? n32 : n69640;
  assign n69642 = pi17 ? n32 : n69641;
  assign n69643 = pi16 ? n32 : n69642;
  assign n69644 = pi20 ? n59665 : n30868;
  assign n69645 = pi22 ? n69595 : n59395;
  assign n69646 = pi21 ? n37878 : n69645;
  assign n69647 = pi20 ? n69646 : n32;
  assign n69648 = pi19 ? n69644 : n69647;
  assign n69649 = pi18 ? n32 : n69648;
  assign n69650 = pi17 ? n32 : n69649;
  assign n69651 = pi16 ? n32 : n69650;
  assign n69652 = pi15 ? n69643 : n69651;
  assign n69653 = pi21 ? n47321 : n68602;
  assign n69654 = pi22 ? n33792 : n42106;
  assign n69655 = pi21 ? n30868 : n69654;
  assign n69656 = pi20 ? n69653 : n69655;
  assign n69657 = pi22 ? n63328 : n59672;
  assign n69658 = pi21 ? n64961 : n69657;
  assign n69659 = pi20 ? n69658 : n32;
  assign n69660 = pi19 ? n69656 : n69659;
  assign n69661 = pi18 ? n32 : n69660;
  assign n69662 = pi17 ? n32 : n69661;
  assign n69663 = pi16 ? n32 : n69662;
  assign n69664 = pi23 ? n20563 : n66385;
  assign n69665 = pi22 ? n69664 : n39190;
  assign n69666 = pi21 ? n20563 : n69665;
  assign n69667 = pi20 ? n55483 : n69666;
  assign n69668 = pi21 ? n63253 : n65038;
  assign n69669 = pi20 ? n69668 : n32;
  assign n69670 = pi19 ? n69667 : n69669;
  assign n69671 = pi18 ? n32 : n69670;
  assign n69672 = pi17 ? n32 : n69671;
  assign n69673 = pi16 ? n32 : n69672;
  assign n69674 = pi15 ? n69663 : n69673;
  assign n69675 = pi14 ? n69652 : n69674;
  assign n69676 = pi21 ? n55516 : n36489;
  assign n69677 = pi20 ? n69676 : n56604;
  assign n69678 = pi22 ? n60841 : n51564;
  assign n69679 = pi21 ? n69678 : n64278;
  assign n69680 = pi20 ? n69679 : n32;
  assign n69681 = pi19 ? n69677 : n69680;
  assign n69682 = pi18 ? n32 : n69681;
  assign n69683 = pi17 ? n32 : n69682;
  assign n69684 = pi16 ? n32 : n69683;
  assign n69685 = pi21 ? n46758 : n36489;
  assign n69686 = pi22 ? n20563 : n46172;
  assign n69687 = pi21 ? n48173 : n69686;
  assign n69688 = pi20 ? n69685 : n69687;
  assign n69689 = pi23 ? n55580 : n36798;
  assign n69690 = pi22 ? n69689 : n14626;
  assign n69691 = pi21 ? n69690 : n59648;
  assign n69692 = pi20 ? n69691 : n32;
  assign n69693 = pi19 ? n69688 : n69692;
  assign n69694 = pi18 ? n32 : n69693;
  assign n69695 = pi17 ? n32 : n69694;
  assign n69696 = pi16 ? n32 : n69695;
  assign n69697 = pi15 ? n69684 : n69696;
  assign n69698 = pi22 ? n20563 : n68361;
  assign n69699 = pi21 ? n51755 : n69698;
  assign n69700 = pi21 ? n48173 : n61264;
  assign n69701 = pi20 ? n69699 : n69700;
  assign n69702 = pi23 ? n63194 : n36798;
  assign n69703 = pi22 ? n69702 : n51564;
  assign n69704 = pi21 ? n69703 : n54564;
  assign n69705 = pi20 ? n69704 : n32;
  assign n69706 = pi19 ? n69701 : n69705;
  assign n69707 = pi18 ? n32 : n69706;
  assign n69708 = pi17 ? n32 : n69707;
  assign n69709 = pi16 ? n32 : n69708;
  assign n69710 = pi22 ? n58428 : n36781;
  assign n69711 = pi21 ? n45016 : n69710;
  assign n69712 = pi20 ? n39395 : n69711;
  assign n69713 = pi22 ? n43199 : n51564;
  assign n69714 = pi21 ? n69713 : n59357;
  assign n69715 = pi20 ? n69714 : n32;
  assign n69716 = pi19 ? n69712 : n69715;
  assign n69717 = pi18 ? n32 : n69716;
  assign n69718 = pi17 ? n32 : n69717;
  assign n69719 = pi16 ? n32 : n69718;
  assign n69720 = pi15 ? n69709 : n69719;
  assign n69721 = pi14 ? n69697 : n69720;
  assign n69722 = pi13 ? n69675 : n69721;
  assign n69723 = pi20 ? n39395 : n59602;
  assign n69724 = pi24 ? n51564 : n13481;
  assign n69725 = pi23 ? n14626 : n69724;
  assign n69726 = pi22 ? n62300 : n69725;
  assign n69727 = pi21 ? n69726 : n37639;
  assign n69728 = pi20 ? n69727 : n32;
  assign n69729 = pi19 ? n69723 : n69728;
  assign n69730 = pi18 ? n32 : n69729;
  assign n69731 = pi17 ? n32 : n69730;
  assign n69732 = pi16 ? n32 : n69731;
  assign n69733 = pi21 ? n40986 : n36798;
  assign n69734 = pi20 ? n39395 : n69733;
  assign n69735 = pi20 ? n68899 : n32;
  assign n69736 = pi19 ? n69734 : n69735;
  assign n69737 = pi18 ? n32 : n69736;
  assign n69738 = pi17 ? n32 : n69737;
  assign n69739 = pi16 ? n32 : n69738;
  assign n69740 = pi15 ? n69732 : n69739;
  assign n69741 = pi21 ? n36798 : n46260;
  assign n69742 = pi20 ? n39395 : n69741;
  assign n69743 = pi23 ? n52672 : n14362;
  assign n69744 = pi22 ? n62803 : n69743;
  assign n69745 = pi21 ? n69744 : n32;
  assign n69746 = pi20 ? n69745 : n32;
  assign n69747 = pi19 ? n69742 : n69746;
  assign n69748 = pi18 ? n32 : n69747;
  assign n69749 = pi17 ? n32 : n69748;
  assign n69750 = pi16 ? n32 : n69749;
  assign n69751 = pi21 ? n36798 : n56695;
  assign n69752 = pi20 ? n39395 : n69751;
  assign n69753 = pi19 ? n69752 : n61415;
  assign n69754 = pi18 ? n32 : n69753;
  assign n69755 = pi17 ? n32 : n69754;
  assign n69756 = pi16 ? n32 : n69755;
  assign n69757 = pi15 ? n69750 : n69756;
  assign n69758 = pi14 ? n69740 : n69757;
  assign n69759 = pi21 ? n62322 : n58794;
  assign n69760 = pi20 ? n37333 : n69759;
  assign n69761 = pi19 ? n69760 : n59650;
  assign n69762 = pi18 ? n32 : n69761;
  assign n69763 = pi17 ? n32 : n69762;
  assign n69764 = pi16 ? n32 : n69763;
  assign n69765 = pi21 ? n63401 : n59681;
  assign n69766 = pi20 ? n37333 : n69765;
  assign n69767 = pi19 ? n69766 : n56131;
  assign n69768 = pi18 ? n32 : n69767;
  assign n69769 = pi17 ? n32 : n69768;
  assign n69770 = pi16 ? n32 : n69769;
  assign n69771 = pi15 ? n69764 : n69770;
  assign n69772 = pi21 ? n47321 : n36489;
  assign n69773 = pi22 ? n36798 : n64161;
  assign n69774 = pi21 ? n68362 : n69773;
  assign n69775 = pi20 ? n69772 : n69774;
  assign n69776 = pi19 ? n69775 : n37641;
  assign n69777 = pi18 ? n32 : n69776;
  assign n69778 = pi17 ? n32 : n69777;
  assign n69779 = pi16 ? n32 : n69778;
  assign n69780 = pi22 ? n49412 : n36798;
  assign n69781 = pi21 ? n69780 : n13481;
  assign n69782 = pi20 ? n55483 : n69781;
  assign n69783 = pi19 ? n69782 : n37641;
  assign n69784 = pi18 ? n32 : n69783;
  assign n69785 = pi17 ? n32 : n69784;
  assign n69786 = pi16 ? n32 : n69785;
  assign n69787 = pi15 ? n69779 : n69786;
  assign n69788 = pi14 ? n69771 : n69787;
  assign n69789 = pi13 ? n69758 : n69788;
  assign n69790 = pi12 ? n69722 : n69789;
  assign n69791 = pi22 ? n49412 : n13481;
  assign n69792 = pi21 ? n69791 : n13481;
  assign n69793 = pi20 ? n69772 : n69792;
  assign n69794 = pi19 ? n69793 : n35482;
  assign n69795 = pi18 ? n32 : n69794;
  assign n69796 = pi17 ? n32 : n69795;
  assign n69797 = pi16 ? n32 : n69796;
  assign n69798 = pi21 ? n61930 : n57760;
  assign n69799 = pi20 ? n65200 : n69798;
  assign n69800 = pi19 ? n69799 : n32;
  assign n69801 = pi18 ? n32 : n69800;
  assign n69802 = pi17 ? n32 : n69801;
  assign n69803 = pi16 ? n32 : n69802;
  assign n69804 = pi15 ? n69797 : n69803;
  assign n69805 = pi22 ? n30868 : n46172;
  assign n69806 = pi21 ? n32 : n69805;
  assign n69807 = pi21 ? n59774 : n57563;
  assign n69808 = pi20 ? n69806 : n69807;
  assign n69809 = pi19 ? n69808 : n32;
  assign n69810 = pi18 ? n32 : n69809;
  assign n69811 = pi17 ? n32 : n69810;
  assign n69812 = pi16 ? n32 : n69811;
  assign n69813 = pi21 ? n32 : n59524;
  assign n69814 = pi22 ? n55799 : n63328;
  assign n69815 = pi21 ? n69814 : n55560;
  assign n69816 = pi20 ? n69813 : n69815;
  assign n69817 = pi19 ? n69816 : n32;
  assign n69818 = pi18 ? n32 : n69817;
  assign n69819 = pi17 ? n32 : n69818;
  assign n69820 = pi16 ? n32 : n69819;
  assign n69821 = pi15 ? n69812 : n69820;
  assign n69822 = pi14 ? n69804 : n69821;
  assign n69823 = pi22 ? n56712 : n36798;
  assign n69824 = pi21 ? n32 : n69823;
  assign n69825 = pi21 ? n62420 : n55560;
  assign n69826 = pi20 ? n69824 : n69825;
  assign n69827 = pi19 ? n69826 : n32;
  assign n69828 = pi18 ? n32 : n69827;
  assign n69829 = pi17 ? n32 : n69828;
  assign n69830 = pi16 ? n32 : n69829;
  assign n69831 = pi21 ? n32 : n56211;
  assign n69832 = pi21 ? n67051 : n57097;
  assign n69833 = pi20 ? n69831 : n69832;
  assign n69834 = pi19 ? n69833 : n32;
  assign n69835 = pi18 ? n32 : n69834;
  assign n69836 = pi17 ? n32 : n69835;
  assign n69837 = pi16 ? n32 : n69836;
  assign n69838 = pi15 ? n69830 : n69837;
  assign n69839 = pi22 ? n45160 : n49412;
  assign n69840 = pi21 ? n32 : n69839;
  assign n69841 = pi21 ? n62515 : n37639;
  assign n69842 = pi20 ? n69840 : n69841;
  assign n69843 = pi19 ? n69842 : n32;
  assign n69844 = pi18 ? n32 : n69843;
  assign n69845 = pi17 ? n32 : n69844;
  assign n69846 = pi16 ? n32 : n69845;
  assign n69847 = pi22 ? n46789 : n43199;
  assign n69848 = pi21 ? n32 : n69847;
  assign n69849 = pi20 ? n69848 : n62850;
  assign n69850 = pi19 ? n69849 : n32;
  assign n69851 = pi18 ? n32 : n69850;
  assign n69852 = pi17 ? n32 : n69851;
  assign n69853 = pi16 ? n32 : n69852;
  assign n69854 = pi15 ? n69846 : n69853;
  assign n69855 = pi14 ? n69838 : n69854;
  assign n69856 = pi13 ? n69822 : n69855;
  assign n69857 = pi20 ? n63812 : n67728;
  assign n69858 = pi19 ? n69857 : n32;
  assign n69859 = pi18 ? n32 : n69858;
  assign n69860 = pi17 ? n32 : n69859;
  assign n69861 = pi16 ? n32 : n69860;
  assign n69862 = pi20 ? n65285 : n59649;
  assign n69863 = pi19 ? n69862 : n32;
  assign n69864 = pi18 ? n32 : n69863;
  assign n69865 = pi17 ? n32 : n69864;
  assign n69866 = pi16 ? n32 : n69865;
  assign n69867 = pi15 ? n69861 : n69866;
  assign n69868 = pi22 ? n63432 : n55641;
  assign n69869 = pi21 ? n32 : n69868;
  assign n69870 = pi20 ? n69869 : n60045;
  assign n69871 = pi19 ? n69870 : n32;
  assign n69872 = pi18 ? n32 : n69871;
  assign n69873 = pi17 ? n32 : n69872;
  assign n69874 = pi16 ? n32 : n69873;
  assign n69875 = pi20 ? n63830 : n37640;
  assign n69876 = pi19 ? n69875 : n32;
  assign n69877 = pi18 ? n32 : n69876;
  assign n69878 = pi17 ? n32 : n69877;
  assign n69879 = pi16 ? n32 : n69878;
  assign n69880 = pi15 ? n69874 : n69879;
  assign n69881 = pi14 ? n69867 : n69880;
  assign n69882 = pi23 ? n63008 : n13481;
  assign n69883 = pi22 ? n32 : n69882;
  assign n69884 = pi21 ? n32 : n69883;
  assign n69885 = pi20 ? n69884 : n20953;
  assign n69886 = pi19 ? n69885 : n32;
  assign n69887 = pi18 ? n32 : n69886;
  assign n69888 = pi17 ? n32 : n69887;
  assign n69889 = pi16 ? n32 : n69888;
  assign n69890 = pi23 ? n32 : n13481;
  assign n69891 = pi22 ? n32 : n69890;
  assign n69892 = pi21 ? n32 : n69891;
  assign n69893 = pi20 ? n69892 : n20953;
  assign n69894 = pi19 ? n69893 : n32;
  assign n69895 = pi18 ? n32 : n69894;
  assign n69896 = pi17 ? n32 : n69895;
  assign n69897 = pi16 ? n32 : n69896;
  assign n69898 = pi15 ? n69889 : n69897;
  assign n69899 = pi14 ? n69898 : n32;
  assign n69900 = pi13 ? n69881 : n69899;
  assign n69901 = pi12 ? n69856 : n69900;
  assign n69902 = pi11 ? n69790 : n69901;
  assign n69903 = pi10 ? n69635 : n69902;
  assign n69904 = pi09 ? n69443 : n69903;
  assign n69905 = pi19 ? n37334 : n69424;
  assign n69906 = pi18 ? n32 : n69905;
  assign n69907 = pi17 ? n32 : n69906;
  assign n69908 = pi16 ? n32 : n69907;
  assign n69909 = pi15 ? n32 : n69908;
  assign n69910 = pi19 ? n37334 : n61976;
  assign n69911 = pi18 ? n32 : n69910;
  assign n69912 = pi17 ? n32 : n69911;
  assign n69913 = pi16 ? n32 : n69912;
  assign n69914 = pi19 ? n37334 : n62975;
  assign n69915 = pi18 ? n32 : n69914;
  assign n69916 = pi17 ? n32 : n69915;
  assign n69917 = pi16 ? n32 : n69916;
  assign n69918 = pi15 ? n69913 : n69917;
  assign n69919 = pi14 ? n69909 : n69918;
  assign n69920 = pi13 ? n32 : n69919;
  assign n69921 = pi12 ? n32 : n69920;
  assign n69922 = pi11 ? n32 : n69921;
  assign n69923 = pi10 ? n32 : n69922;
  assign n69924 = pi19 ? n38377 : n62975;
  assign n69925 = pi18 ? n32 : n69924;
  assign n69926 = pi17 ? n32 : n69925;
  assign n69927 = pi16 ? n32 : n69926;
  assign n69928 = pi15 ? n69927 : n69437;
  assign n69929 = pi15 ? n69437 : n68984;
  assign n69930 = pi14 ? n69928 : n69929;
  assign n69931 = pi20 ? n68460 : n61008;
  assign n69932 = pi19 ? n31314 : n69931;
  assign n69933 = pi18 ? n32 : n69932;
  assign n69934 = pi17 ? n32 : n69933;
  assign n69935 = pi16 ? n32 : n69934;
  assign n69936 = pi19 ? n31314 : n67606;
  assign n69937 = pi18 ? n32 : n69936;
  assign n69938 = pi17 ? n32 : n69937;
  assign n69939 = pi16 ? n32 : n69938;
  assign n69940 = pi15 ? n69935 : n69939;
  assign n69941 = pi19 ? n31314 : n62975;
  assign n69942 = pi18 ? n32 : n69941;
  assign n69943 = pi17 ? n32 : n69942;
  assign n69944 = pi16 ? n32 : n69943;
  assign n69945 = pi14 ? n69940 : n69944;
  assign n69946 = pi13 ? n69930 : n69945;
  assign n69947 = pi19 ? n40496 : n69469;
  assign n69948 = pi18 ? n32 : n69947;
  assign n69949 = pi17 ? n32 : n69948;
  assign n69950 = pi16 ? n32 : n69949;
  assign n69951 = pi20 ? n37926 : n38754;
  assign n69952 = pi20 ? n38754 : n59305;
  assign n69953 = pi19 ? n69951 : n69952;
  assign n69954 = pi18 ? n32 : n69953;
  assign n69955 = pi17 ? n32 : n69954;
  assign n69956 = pi16 ? n32 : n69955;
  assign n69957 = pi15 ? n69950 : n69956;
  assign n69958 = pi19 ? n69951 : n69485;
  assign n69959 = pi18 ? n32 : n69958;
  assign n69960 = pi17 ? n32 : n69959;
  assign n69961 = pi16 ? n32 : n69960;
  assign n69962 = pi19 ? n40496 : n69494;
  assign n69963 = pi18 ? n32 : n69962;
  assign n69964 = pi17 ? n32 : n69963;
  assign n69965 = pi16 ? n32 : n69964;
  assign n69966 = pi15 ? n69961 : n69965;
  assign n69967 = pi14 ? n69957 : n69966;
  assign n69968 = pi13 ? n68475 : n69967;
  assign n69969 = pi12 ? n69946 : n69968;
  assign n69970 = pi19 ? n40496 : n69504;
  assign n69971 = pi18 ? n32 : n69970;
  assign n69972 = pi17 ? n32 : n69971;
  assign n69973 = pi16 ? n32 : n69972;
  assign n69974 = pi23 ? n24414 : n13481;
  assign n69975 = pi22 ? n69974 : n13481;
  assign n69976 = pi21 ? n69975 : n37639;
  assign n69977 = pi20 ? n55475 : n69976;
  assign n69978 = pi19 ? n40496 : n69977;
  assign n69979 = pi18 ? n32 : n69978;
  assign n69980 = pi17 ? n32 : n69979;
  assign n69981 = pi16 ? n32 : n69980;
  assign n69982 = pi15 ? n69973 : n69981;
  assign n69983 = pi19 ? n40496 : n68580;
  assign n69984 = pi18 ? n32 : n69983;
  assign n69985 = pi17 ? n32 : n69984;
  assign n69986 = pi16 ? n32 : n69985;
  assign n69987 = pi19 ? n41681 : n69519;
  assign n69988 = pi18 ? n32 : n69987;
  assign n69989 = pi17 ? n32 : n69988;
  assign n69990 = pi16 ? n32 : n69989;
  assign n69991 = pi15 ? n69986 : n69990;
  assign n69992 = pi14 ? n69982 : n69991;
  assign n69993 = pi20 ? n38981 : n38754;
  assign n69994 = pi19 ? n69993 : n67669;
  assign n69995 = pi18 ? n32 : n69994;
  assign n69996 = pi17 ? n32 : n69995;
  assign n69997 = pi16 ? n32 : n69996;
  assign n69998 = pi20 ? n38981 : n47158;
  assign n69999 = pi20 ? n69532 : n1010;
  assign n70000 = pi19 ? n69998 : n69999;
  assign n70001 = pi18 ? n32 : n70000;
  assign n70002 = pi17 ? n32 : n70001;
  assign n70003 = pi16 ? n32 : n70002;
  assign n70004 = pi15 ? n69997 : n70003;
  assign n70005 = pi23 ? n62332 : n20563;
  assign n70006 = pi22 ? n20563 : n70005;
  assign n70007 = pi21 ? n20563 : n70006;
  assign n70008 = pi20 ? n38981 : n70007;
  assign n70009 = pi23 ? n13481 : n624;
  assign n70010 = pi22 ? n13481 : n70009;
  assign n70011 = pi21 ? n70010 : n32;
  assign n70012 = pi20 ? n69541 : n70011;
  assign n70013 = pi19 ? n70008 : n70012;
  assign n70014 = pi18 ? n32 : n70013;
  assign n70015 = pi17 ? n32 : n70014;
  assign n70016 = pi16 ? n32 : n70015;
  assign n70017 = pi22 ? n295 : n69547;
  assign n70018 = pi21 ? n30868 : n70017;
  assign n70019 = pi20 ? n70018 : n17510;
  assign n70020 = pi19 ? n41681 : n70019;
  assign n70021 = pi18 ? n32 : n70020;
  assign n70022 = pi17 ? n32 : n70021;
  assign n70023 = pi16 ? n32 : n70022;
  assign n70024 = pi15 ? n70016 : n70023;
  assign n70025 = pi14 ? n70004 : n70024;
  assign n70026 = pi13 ? n69992 : n70025;
  assign n70027 = pi22 ? n13624 : n69558;
  assign n70028 = pi21 ? n20563 : n70027;
  assign n70029 = pi20 ? n70028 : n67712;
  assign n70030 = pi19 ? n40509 : n70029;
  assign n70031 = pi18 ? n32 : n70030;
  assign n70032 = pi17 ? n32 : n70031;
  assign n70033 = pi16 ? n32 : n70032;
  assign n70034 = pi20 ? n40054 : n40791;
  assign n70035 = pi23 ? n20563 : n65003;
  assign n70036 = pi23 ? n335 : n51564;
  assign n70037 = pi22 ? n70035 : n70036;
  assign n70038 = pi21 ? n30868 : n70037;
  assign n70039 = pi20 ? n70038 : n67719;
  assign n70040 = pi19 ? n70034 : n70039;
  assign n70041 = pi18 ? n32 : n70040;
  assign n70042 = pi17 ? n32 : n70041;
  assign n70043 = pi16 ? n32 : n70042;
  assign n70044 = pi15 ? n70033 : n70043;
  assign n70045 = pi22 ? n62742 : n69577;
  assign n70046 = pi21 ? n30868 : n70045;
  assign n70047 = pi20 ? n70046 : n5667;
  assign n70048 = pi19 ? n70034 : n70047;
  assign n70049 = pi18 ? n32 : n70048;
  assign n70050 = pi17 ? n32 : n70049;
  assign n70051 = pi16 ? n32 : n70050;
  assign n70052 = pi20 ? n40054 : n51223;
  assign n70053 = pi23 ? n30868 : n65467;
  assign n70054 = pi22 ? n70053 : n67736;
  assign n70055 = pi21 ? n33792 : n70054;
  assign n70056 = pi22 ? n70009 : n32;
  assign n70057 = pi21 ? n70056 : n32;
  assign n70058 = pi20 ? n70055 : n70057;
  assign n70059 = pi19 ? n70052 : n70058;
  assign n70060 = pi18 ? n32 : n70059;
  assign n70061 = pi17 ? n32 : n70060;
  assign n70062 = pi16 ? n32 : n70061;
  assign n70063 = pi15 ? n70051 : n70062;
  assign n70064 = pi14 ? n70044 : n70063;
  assign n70065 = pi23 ? n33792 : n363;
  assign n70066 = pi22 ? n70065 : n69595;
  assign n70067 = pi21 ? n36659 : n70066;
  assign n70068 = pi20 ? n70067 : n6417;
  assign n70069 = pi19 ? n40509 : n70068;
  assign n70070 = pi18 ? n32 : n70069;
  assign n70071 = pi17 ? n32 : n70070;
  assign n70072 = pi16 ? n32 : n70071;
  assign n70073 = pi20 ? n37933 : n38961;
  assign n70074 = pi22 ? n45675 : n57632;
  assign n70075 = pi21 ? n36659 : n70074;
  assign n70076 = pi20 ? n70075 : n58168;
  assign n70077 = pi19 ? n70073 : n70076;
  assign n70078 = pi18 ? n32 : n70077;
  assign n70079 = pi17 ? n32 : n70078;
  assign n70080 = pi16 ? n32 : n70079;
  assign n70081 = pi15 ? n70072 : n70080;
  assign n70082 = pi19 ? n70073 : n69619;
  assign n70083 = pi18 ? n32 : n70082;
  assign n70084 = pi17 ? n32 : n70083;
  assign n70085 = pi16 ? n32 : n70084;
  assign n70086 = pi23 ? n363 : n43198;
  assign n70087 = pi22 ? n70086 : n62880;
  assign n70088 = pi21 ? n36659 : n70087;
  assign n70089 = pi20 ? n70088 : n32257;
  assign n70090 = pi19 ? n40531 : n70089;
  assign n70091 = pi18 ? n32 : n70090;
  assign n70092 = pi17 ? n32 : n70091;
  assign n70093 = pi16 ? n32 : n70092;
  assign n70094 = pi15 ? n70085 : n70093;
  assign n70095 = pi14 ? n70081 : n70094;
  assign n70096 = pi13 ? n70064 : n70095;
  assign n70097 = pi12 ? n70026 : n70096;
  assign n70098 = pi11 ? n69969 : n70097;
  assign n70099 = pi20 ? n60055 : n41463;
  assign n70100 = pi22 ? n63317 : n13481;
  assign n70101 = pi21 ? n51564 : n70100;
  assign n70102 = pi20 ? n70101 : n37640;
  assign n70103 = pi19 ? n70099 : n70102;
  assign n70104 = pi18 ? n32 : n70103;
  assign n70105 = pi17 ? n32 : n70104;
  assign n70106 = pi16 ? n32 : n70105;
  assign n70107 = pi20 ? n60055 : n30868;
  assign n70108 = pi22 ? n62300 : n59395;
  assign n70109 = pi21 ? n37878 : n70108;
  assign n70110 = pi20 ? n70109 : n32;
  assign n70111 = pi19 ? n70107 : n70110;
  assign n70112 = pi18 ? n32 : n70111;
  assign n70113 = pi17 ? n32 : n70112;
  assign n70114 = pi16 ? n32 : n70113;
  assign n70115 = pi15 ? n70106 : n70114;
  assign n70116 = pi22 ? n46165 : n33792;
  assign n70117 = pi21 ? n32 : n70116;
  assign n70118 = pi20 ? n70117 : n69655;
  assign n70119 = pi19 ? n70118 : n69659;
  assign n70120 = pi18 ? n32 : n70119;
  assign n70121 = pi17 ? n32 : n70120;
  assign n70122 = pi16 ? n32 : n70121;
  assign n70123 = pi23 ? n64063 : n30868;
  assign n70124 = pi22 ? n20563 : n70123;
  assign n70125 = pi21 ? n40954 : n70124;
  assign n70126 = pi20 ? n54401 : n70125;
  assign n70127 = pi19 ? n70126 : n69669;
  assign n70128 = pi18 ? n32 : n70127;
  assign n70129 = pi17 ? n32 : n70128;
  assign n70130 = pi16 ? n32 : n70129;
  assign n70131 = pi15 ? n70122 : n70130;
  assign n70132 = pi14 ? n70115 : n70131;
  assign n70133 = pi23 ? n56064 : n20563;
  assign n70134 = pi22 ? n70133 : n20563;
  assign n70135 = pi22 ? n20563 : n58736;
  assign n70136 = pi21 ? n70134 : n70135;
  assign n70137 = pi20 ? n54428 : n70136;
  assign n70138 = pi21 ? n68762 : n64278;
  assign n70139 = pi20 ? n70138 : n32;
  assign n70140 = pi19 ? n70137 : n70139;
  assign n70141 = pi18 ? n32 : n70140;
  assign n70142 = pi17 ? n32 : n70141;
  assign n70143 = pi16 ? n32 : n70142;
  assign n70144 = pi22 ? n46757 : n30868;
  assign n70145 = pi21 ? n32 : n70144;
  assign n70146 = pi23 ? n55580 : n30868;
  assign n70147 = pi22 ? n70146 : n30868;
  assign n70148 = pi22 ? n20563 : n37288;
  assign n70149 = pi21 ? n70147 : n70148;
  assign n70150 = pi20 ? n70145 : n70149;
  assign n70151 = pi21 ? n67068 : n55560;
  assign n70152 = pi20 ? n70151 : n32;
  assign n70153 = pi19 ? n70150 : n70152;
  assign n70154 = pi18 ? n32 : n70153;
  assign n70155 = pi17 ? n32 : n70154;
  assign n70156 = pi16 ? n32 : n70155;
  assign n70157 = pi15 ? n70143 : n70156;
  assign n70158 = pi22 ? n51754 : n40386;
  assign n70159 = pi21 ? n32 : n70158;
  assign n70160 = pi23 ? n56079 : n30868;
  assign n70161 = pi22 ? n70160 : n30868;
  assign n70162 = pi24 ? n36781 : n36659;
  assign n70163 = pi23 ? n70162 : n36659;
  assign n70164 = pi22 ? n30868 : n70163;
  assign n70165 = pi21 ? n70161 : n70164;
  assign n70166 = pi20 ? n70159 : n70165;
  assign n70167 = pi21 ? n68780 : n54564;
  assign n70168 = pi20 ? n70167 : n32;
  assign n70169 = pi19 ? n70166 : n70168;
  assign n70170 = pi18 ? n32 : n70169;
  assign n70171 = pi17 ? n32 : n70170;
  assign n70172 = pi16 ? n32 : n70171;
  assign n70173 = pi22 ? n57085 : n36781;
  assign n70174 = pi21 ? n45016 : n70173;
  assign n70175 = pi20 ? n38997 : n70174;
  assign n70176 = pi23 ? n8310 : n43198;
  assign n70177 = pi22 ? n70176 : n51564;
  assign n70178 = pi21 ? n70177 : n59357;
  assign n70179 = pi20 ? n70178 : n32;
  assign n70180 = pi19 ? n70175 : n70179;
  assign n70181 = pi18 ? n32 : n70180;
  assign n70182 = pi17 ? n32 : n70181;
  assign n70183 = pi16 ? n32 : n70182;
  assign n70184 = pi15 ? n70172 : n70183;
  assign n70185 = pi14 ? n70157 : n70184;
  assign n70186 = pi13 ? n70132 : n70185;
  assign n70187 = pi20 ? n38997 : n59602;
  assign n70188 = pi22 ? n62300 : n56622;
  assign n70189 = pi21 ? n70188 : n37639;
  assign n70190 = pi20 ? n70189 : n32;
  assign n70191 = pi19 ? n70187 : n70190;
  assign n70192 = pi18 ? n32 : n70191;
  assign n70193 = pi17 ? n32 : n70192;
  assign n70194 = pi16 ? n32 : n70193;
  assign n70195 = pi20 ? n38997 : n69733;
  assign n70196 = pi19 ? n70195 : n69735;
  assign n70197 = pi18 ? n32 : n70196;
  assign n70198 = pi17 ? n32 : n70197;
  assign n70199 = pi16 ? n32 : n70198;
  assign n70200 = pi15 ? n70194 : n70199;
  assign n70201 = pi20 ? n38997 : n69741;
  assign n70202 = pi22 ? n57197 : n57647;
  assign n70203 = pi21 ? n70202 : n32;
  assign n70204 = pi20 ? n70203 : n32;
  assign n70205 = pi19 ? n70201 : n70204;
  assign n70206 = pi18 ? n32 : n70205;
  assign n70207 = pi17 ? n32 : n70206;
  assign n70208 = pi16 ? n32 : n70207;
  assign n70209 = pi22 ? n36781 : n61543;
  assign n70210 = pi21 ? n36798 : n70209;
  assign n70211 = pi20 ? n38997 : n70210;
  assign n70212 = pi19 ? n70211 : n61415;
  assign n70213 = pi18 ? n32 : n70212;
  assign n70214 = pi17 ? n32 : n70213;
  assign n70215 = pi16 ? n32 : n70214;
  assign n70216 = pi15 ? n70208 : n70215;
  assign n70217 = pi14 ? n70200 : n70216;
  assign n70218 = pi22 ? n36781 : n64689;
  assign n70219 = pi21 ? n62322 : n70218;
  assign n70220 = pi20 ? n36867 : n70219;
  assign n70221 = pi19 ? n70220 : n59650;
  assign n70222 = pi18 ? n32 : n70221;
  assign n70223 = pi17 ? n32 : n70222;
  assign n70224 = pi16 ? n32 : n70223;
  assign n70225 = pi23 ? n56987 : n36798;
  assign n70226 = pi22 ? n70225 : n36798;
  assign n70227 = pi21 ? n70226 : n59681;
  assign n70228 = pi20 ? n36867 : n70227;
  assign n70229 = pi19 ? n70228 : n60046;
  assign n70230 = pi18 ? n32 : n70229;
  assign n70231 = pi17 ? n32 : n70230;
  assign n70232 = pi16 ? n32 : n70231;
  assign n70233 = pi15 ? n70224 : n70232;
  assign n70234 = pi22 ? n36798 : n66042;
  assign n70235 = pi21 ? n68362 : n70234;
  assign n70236 = pi20 ? n46167 : n70235;
  assign n70237 = pi19 ? n70236 : n37641;
  assign n70238 = pi18 ? n32 : n70237;
  assign n70239 = pi17 ? n32 : n70238;
  assign n70240 = pi16 ? n32 : n70239;
  assign n70241 = pi23 ? n56064 : n36798;
  assign n70242 = pi22 ? n70241 : n36798;
  assign n70243 = pi21 ? n70242 : n13481;
  assign n70244 = pi20 ? n54401 : n70243;
  assign n70245 = pi19 ? n70244 : n37641;
  assign n70246 = pi18 ? n32 : n70245;
  assign n70247 = pi17 ? n32 : n70246;
  assign n70248 = pi16 ? n32 : n70247;
  assign n70249 = pi15 ? n70240 : n70248;
  assign n70250 = pi14 ? n70233 : n70249;
  assign n70251 = pi13 ? n70217 : n70250;
  assign n70252 = pi12 ? n70186 : n70251;
  assign n70253 = pi22 ? n70241 : n13481;
  assign n70254 = pi21 ? n70253 : n13481;
  assign n70255 = pi20 ? n46167 : n70254;
  assign n70256 = pi19 ? n70255 : n35482;
  assign n70257 = pi18 ? n32 : n70256;
  assign n70258 = pi17 ? n32 : n70257;
  assign n70259 = pi16 ? n32 : n70258;
  assign n70260 = pi20 ? n46061 : n69798;
  assign n70261 = pi19 ? n70260 : n32;
  assign n70262 = pi18 ? n32 : n70261;
  assign n70263 = pi17 ? n32 : n70262;
  assign n70264 = pi16 ? n32 : n70263;
  assign n70265 = pi15 ? n70259 : n70264;
  assign n70266 = pi22 ? n32 : n46172;
  assign n70267 = pi21 ? n32 : n70266;
  assign n70268 = pi22 ? n56606 : n13481;
  assign n70269 = pi21 ? n70268 : n57563;
  assign n70270 = pi20 ? n70267 : n70269;
  assign n70271 = pi19 ? n70270 : n32;
  assign n70272 = pi18 ? n32 : n70271;
  assign n70273 = pi17 ? n32 : n70272;
  assign n70274 = pi16 ? n32 : n70273;
  assign n70275 = pi23 ? n36798 : n55783;
  assign n70276 = pi22 ? n70275 : n56607;
  assign n70277 = pi21 ? n70276 : n55560;
  assign n70278 = pi20 ? n48822 : n70277;
  assign n70279 = pi19 ? n70278 : n32;
  assign n70280 = pi18 ? n32 : n70279;
  assign n70281 = pi17 ? n32 : n70280;
  assign n70282 = pi16 ? n32 : n70281;
  assign n70283 = pi15 ? n70274 : n70282;
  assign n70284 = pi14 ? n70265 : n70283;
  assign n70285 = pi21 ? n56760 : n55560;
  assign n70286 = pi20 ? n48822 : n70285;
  assign n70287 = pi19 ? n70286 : n32;
  assign n70288 = pi18 ? n32 : n70287;
  assign n70289 = pi17 ? n32 : n70288;
  assign n70290 = pi16 ? n32 : n70289;
  assign n70291 = pi20 ? n48857 : n68899;
  assign n70292 = pi19 ? n70291 : n32;
  assign n70293 = pi18 ? n32 : n70292;
  assign n70294 = pi17 ? n32 : n70293;
  assign n70295 = pi16 ? n32 : n70294;
  assign n70296 = pi15 ? n70290 : n70295;
  assign n70297 = pi21 ? n32 : n46772;
  assign n70298 = pi22 ? n57197 : n13481;
  assign n70299 = pi21 ? n70298 : n32;
  assign n70300 = pi20 ? n70297 : n70299;
  assign n70301 = pi19 ? n70300 : n32;
  assign n70302 = pi18 ? n32 : n70301;
  assign n70303 = pi17 ? n32 : n70302;
  assign n70304 = pi16 ? n32 : n70303;
  assign n70305 = pi20 ? n52918 : n62850;
  assign n70306 = pi19 ? n70305 : n32;
  assign n70307 = pi18 ? n32 : n70306;
  assign n70308 = pi17 ? n32 : n70307;
  assign n70309 = pi16 ? n32 : n70308;
  assign n70310 = pi15 ? n70304 : n70309;
  assign n70311 = pi14 ? n70296 : n70310;
  assign n70312 = pi13 ? n70284 : n70311;
  assign n70313 = pi22 ? n32 : n69401;
  assign n70314 = pi21 ? n32 : n70313;
  assign n70315 = pi20 ? n70314 : n67728;
  assign n70316 = pi19 ? n70315 : n32;
  assign n70317 = pi18 ? n32 : n70316;
  assign n70318 = pi17 ? n32 : n70317;
  assign n70319 = pi16 ? n32 : n70318;
  assign n70320 = pi20 ? n32 : n59649;
  assign n70321 = pi19 ? n70320 : n32;
  assign n70322 = pi18 ? n32 : n70321;
  assign n70323 = pi17 ? n32 : n70322;
  assign n70324 = pi16 ? n32 : n70323;
  assign n70325 = pi15 ? n70319 : n70324;
  assign n70326 = pi20 ? n32 : n60045;
  assign n70327 = pi19 ? n70326 : n32;
  assign n70328 = pi18 ? n32 : n70327;
  assign n70329 = pi17 ? n32 : n70328;
  assign n70330 = pi16 ? n32 : n70329;
  assign n70331 = pi20 ? n32 : n37640;
  assign n70332 = pi19 ? n70331 : n32;
  assign n70333 = pi18 ? n32 : n70332;
  assign n70334 = pi17 ? n32 : n70333;
  assign n70335 = pi16 ? n32 : n70334;
  assign n70336 = pi15 ? n70330 : n70335;
  assign n70337 = pi14 ? n70325 : n70336;
  assign n70338 = pi13 ? n70337 : n32;
  assign n70339 = pi12 ? n70312 : n70338;
  assign n70340 = pi11 ? n70252 : n70339;
  assign n70341 = pi10 ? n70098 : n70340;
  assign n70342 = pi09 ? n69923 : n70341;
  assign n70343 = pi08 ? n69904 : n70342;
  assign n70344 = pi07 ? n69423 : n70343;
  assign n70345 = pi06 ? n68459 : n70344;
  assign n70346 = pi05 ? n66570 : n70345;
  assign n70347 = pi04 ? n62947 : n70346;
  assign n70348 = pi20 ? n20563 : n13040;
  assign n70349 = pi19 ? n38998 : n70348;
  assign n70350 = pi18 ? n32 : n70349;
  assign n70351 = pi17 ? n32 : n70350;
  assign n70352 = pi16 ? n32 : n70351;
  assign n70353 = pi15 ? n32 : n70352;
  assign n70354 = pi20 ? n40791 : n1619;
  assign n70355 = pi19 ? n38998 : n70354;
  assign n70356 = pi18 ? n32 : n70355;
  assign n70357 = pi17 ? n32 : n70356;
  assign n70358 = pi16 ? n32 : n70357;
  assign n70359 = pi14 ? n70353 : n70358;
  assign n70360 = pi13 ? n32 : n70359;
  assign n70361 = pi12 ? n32 : n70360;
  assign n70362 = pi11 ? n32 : n70361;
  assign n70363 = pi10 ? n32 : n70362;
  assign n70364 = pi19 ? n37321 : n62975;
  assign n70365 = pi18 ? n32 : n70364;
  assign n70366 = pi17 ? n32 : n70365;
  assign n70367 = pi16 ? n32 : n70366;
  assign n70368 = pi15 ? n70367 : n69917;
  assign n70369 = pi15 ? n69917 : n69437;
  assign n70370 = pi14 ? n70368 : n70369;
  assign n70371 = pi19 ? n28158 : n62954;
  assign n70372 = pi18 ? n32 : n70371;
  assign n70373 = pi17 ? n32 : n70372;
  assign n70374 = pi16 ? n32 : n70373;
  assign n70375 = pi14 ? n69447 : n70374;
  assign n70376 = pi13 ? n70370 : n70375;
  assign n70377 = pi19 ? n30118 : n62954;
  assign n70378 = pi18 ? n32 : n70377;
  assign n70379 = pi17 ? n32 : n70378;
  assign n70380 = pi16 ? n32 : n70379;
  assign n70381 = pi19 ? n31264 : n62954;
  assign n70382 = pi18 ? n32 : n70381;
  assign n70383 = pi17 ? n32 : n70382;
  assign n70384 = pi16 ? n32 : n70383;
  assign n70385 = pi14 ? n70380 : n70384;
  assign n70386 = pi19 ? n31314 : n59306;
  assign n70387 = pi18 ? n32 : n70386;
  assign n70388 = pi17 ? n32 : n70387;
  assign n70389 = pi16 ? n32 : n70388;
  assign n70390 = pi23 ? n11127 : n14626;
  assign n70391 = pi22 ? n70390 : n14626;
  assign n70392 = pi21 ? n70391 : n65115;
  assign n70393 = pi20 ? n20563 : n70392;
  assign n70394 = pi19 ? n31314 : n70393;
  assign n70395 = pi18 ? n32 : n70394;
  assign n70396 = pi17 ? n32 : n70395;
  assign n70397 = pi16 ? n32 : n70396;
  assign n70398 = pi15 ? n70389 : n70397;
  assign n70399 = pi20 ? n53356 : n69484;
  assign n70400 = pi19 ? n31314 : n70399;
  assign n70401 = pi18 ? n32 : n70400;
  assign n70402 = pi17 ? n32 : n70401;
  assign n70403 = pi16 ? n32 : n70402;
  assign n70404 = pi22 ? n69491 : n316;
  assign n70405 = pi21 ? n70404 : n3523;
  assign n70406 = pi20 ? n20563 : n70405;
  assign n70407 = pi19 ? n31314 : n70406;
  assign n70408 = pi18 ? n32 : n70407;
  assign n70409 = pi17 ? n32 : n70408;
  assign n70410 = pi16 ? n32 : n70409;
  assign n70411 = pi15 ? n70403 : n70410;
  assign n70412 = pi14 ? n70398 : n70411;
  assign n70413 = pi13 ? n70385 : n70412;
  assign n70414 = pi12 ? n70376 : n70413;
  assign n70415 = pi20 ? n53367 : n68566;
  assign n70416 = pi19 ? n43672 : n70415;
  assign n70417 = pi18 ? n32 : n70416;
  assign n70418 = pi17 ? n32 : n70417;
  assign n70419 = pi16 ? n32 : n70418;
  assign n70420 = pi21 ? n68578 : n59342;
  assign n70421 = pi20 ? n38754 : n70420;
  assign n70422 = pi19 ? n43672 : n70421;
  assign n70423 = pi18 ? n32 : n70422;
  assign n70424 = pi17 ? n32 : n70423;
  assign n70425 = pi16 ? n32 : n70424;
  assign n70426 = pi15 ? n70419 : n70425;
  assign n70427 = pi22 ? n64606 : n14626;
  assign n70428 = pi21 ? n70427 : n2637;
  assign n70429 = pi20 ? n56539 : n70428;
  assign n70430 = pi19 ? n43672 : n70429;
  assign n70431 = pi18 ? n32 : n70430;
  assign n70432 = pi17 ? n32 : n70431;
  assign n70433 = pi16 ? n32 : n70432;
  assign n70434 = pi20 ? n47158 : n63941;
  assign n70435 = pi19 ? n43672 : n70434;
  assign n70436 = pi18 ? n32 : n70435;
  assign n70437 = pi17 ? n32 : n70436;
  assign n70438 = pi16 ? n32 : n70437;
  assign n70439 = pi15 ? n70433 : n70438;
  assign n70440 = pi14 ? n70426 : n70439;
  assign n70441 = pi21 ? n13481 : n928;
  assign n70442 = pi20 ? n65753 : n70441;
  assign n70443 = pi19 ? n43672 : n70442;
  assign n70444 = pi18 ? n32 : n70443;
  assign n70445 = pi17 ? n32 : n70444;
  assign n70446 = pi16 ? n32 : n70445;
  assign n70447 = pi20 ? n32 : n67791;
  assign n70448 = pi22 ? n20563 : n65791;
  assign n70449 = pi21 ? n20563 : n70448;
  assign n70450 = pi20 ? n70449 : n59388;
  assign n70451 = pi19 ? n70447 : n70450;
  assign n70452 = pi18 ? n32 : n70451;
  assign n70453 = pi17 ? n32 : n70452;
  assign n70454 = pi16 ? n32 : n70453;
  assign n70455 = pi15 ? n70446 : n70454;
  assign n70456 = pi23 ? n55534 : n20563;
  assign n70457 = pi22 ? n70456 : n20563;
  assign n70458 = pi21 ? n70457 : n20563;
  assign n70459 = pi20 ? n32 : n70458;
  assign n70460 = pi22 ? n30868 : n68361;
  assign n70461 = pi21 ? n30868 : n70460;
  assign n70462 = pi20 ? n70461 : n10297;
  assign n70463 = pi19 ? n70459 : n70462;
  assign n70464 = pi18 ? n32 : n70463;
  assign n70465 = pi17 ? n32 : n70464;
  assign n70466 = pi16 ? n32 : n70465;
  assign n70467 = pi22 ? n70456 : n40386;
  assign n70468 = pi21 ? n70467 : n20563;
  assign n70469 = pi20 ? n32 : n70468;
  assign n70470 = pi22 ? n33792 : n233;
  assign n70471 = pi21 ? n30868 : n70470;
  assign n70472 = pi21 ? n67783 : n32;
  assign n70473 = pi20 ? n70471 : n70472;
  assign n70474 = pi19 ? n70469 : n70473;
  assign n70475 = pi18 ? n32 : n70474;
  assign n70476 = pi17 ? n32 : n70475;
  assign n70477 = pi16 ? n32 : n70476;
  assign n70478 = pi15 ? n70466 : n70477;
  assign n70479 = pi14 ? n70455 : n70478;
  assign n70480 = pi13 ? n70440 : n70479;
  assign n70481 = pi22 ? n69568 : n54574;
  assign n70482 = pi21 ? n20563 : n70481;
  assign n70483 = pi21 ? n65478 : n32;
  assign n70484 = pi20 ? n70482 : n70483;
  assign n70485 = pi19 ? n43672 : n70484;
  assign n70486 = pi18 ? n32 : n70485;
  assign n70487 = pi17 ? n32 : n70486;
  assign n70488 = pi16 ? n32 : n70487;
  assign n70489 = pi20 ? n32 : n36489;
  assign n70490 = pi23 ? n30868 : n64063;
  assign n70491 = pi23 ? n36659 : n51564;
  assign n70492 = pi22 ? n70490 : n70491;
  assign n70493 = pi21 ? n20563 : n70492;
  assign n70494 = pi22 ? n316 : n54563;
  assign n70495 = pi21 ? n70494 : n32;
  assign n70496 = pi20 ? n70493 : n70495;
  assign n70497 = pi19 ? n70489 : n70496;
  assign n70498 = pi18 ? n32 : n70497;
  assign n70499 = pi17 ? n32 : n70498;
  assign n70500 = pi16 ? n32 : n70499;
  assign n70501 = pi15 ? n70488 : n70500;
  assign n70502 = pi21 ? n41489 : n45016;
  assign n70503 = pi20 ? n32 : n70502;
  assign n70504 = pi23 ? n33792 : n56478;
  assign n70505 = pi22 ? n70504 : n50339;
  assign n70506 = pi21 ? n33792 : n70505;
  assign n70507 = pi20 ? n70506 : n59635;
  assign n70508 = pi19 ? n70503 : n70507;
  assign n70509 = pi18 ? n32 : n70508;
  assign n70510 = pi17 ? n32 : n70509;
  assign n70511 = pi16 ? n32 : n70510;
  assign n70512 = pi20 ? n37926 : n40986;
  assign n70513 = pi23 ? n33792 : n3134;
  assign n70514 = pi22 ? n70513 : n69595;
  assign n70515 = pi21 ? n36659 : n70514;
  assign n70516 = pi20 ? n70515 : n4110;
  assign n70517 = pi19 ? n70512 : n70516;
  assign n70518 = pi18 ? n32 : n70517;
  assign n70519 = pi17 ? n32 : n70518;
  assign n70520 = pi16 ? n32 : n70519;
  assign n70521 = pi15 ? n70511 : n70520;
  assign n70522 = pi14 ? n70501 : n70521;
  assign n70523 = pi21 ? n65759 : n40986;
  assign n70524 = pi20 ? n37926 : n70523;
  assign n70525 = pi22 ? n38284 : n55622;
  assign n70526 = pi21 ? n36659 : n70525;
  assign n70527 = pi20 ? n70526 : n59658;
  assign n70528 = pi19 ? n70524 : n70527;
  assign n70529 = pi18 ? n32 : n70528;
  assign n70530 = pi17 ? n32 : n70529;
  assign n70531 = pi16 ? n32 : n70530;
  assign n70532 = pi20 ? n37926 : n55475;
  assign n70533 = pi22 ? n37276 : n65935;
  assign n70534 = pi21 ? n36659 : n70533;
  assign n70535 = pi20 ? n70534 : n59674;
  assign n70536 = pi19 ? n70532 : n70535;
  assign n70537 = pi18 ? n32 : n70536;
  assign n70538 = pi17 ? n32 : n70537;
  assign n70539 = pi16 ? n32 : n70538;
  assign n70540 = pi15 ? n70531 : n70539;
  assign n70541 = pi22 ? n50339 : n56607;
  assign n70542 = pi21 ? n36659 : n70541;
  assign n70543 = pi20 ? n70542 : n54565;
  assign n70544 = pi19 ? n40496 : n70543;
  assign n70545 = pi18 ? n32 : n70544;
  assign n70546 = pi17 ? n32 : n70545;
  assign n70547 = pi16 ? n32 : n70546;
  assign n70548 = pi22 ? n43199 : n57659;
  assign n70549 = pi21 ? n36659 : n70548;
  assign n70550 = pi20 ? n70549 : n37640;
  assign n70551 = pi19 ? n40496 : n70550;
  assign n70552 = pi18 ? n32 : n70551;
  assign n70553 = pi17 ? n32 : n70552;
  assign n70554 = pi16 ? n32 : n70553;
  assign n70555 = pi15 ? n70547 : n70554;
  assign n70556 = pi14 ? n70540 : n70555;
  assign n70557 = pi13 ? n70522 : n70556;
  assign n70558 = pi12 ? n70480 : n70557;
  assign n70559 = pi11 ? n70414 : n70558;
  assign n70560 = pi21 ? n36489 : n40917;
  assign n70561 = pi20 ? n37926 : n70560;
  assign n70562 = pi22 ? n64689 : n64963;
  assign n70563 = pi21 ? n36781 : n70562;
  assign n70564 = pi20 ? n70563 : n32;
  assign n70565 = pi19 ? n70561 : n70564;
  assign n70566 = pi18 ? n32 : n70565;
  assign n70567 = pi17 ? n32 : n70566;
  assign n70568 = pi16 ? n32 : n70567;
  assign n70569 = pi20 ? n37926 : n42006;
  assign n70570 = pi21 ? n39972 : n64697;
  assign n70571 = pi20 ? n70570 : n32;
  assign n70572 = pi19 ? n70569 : n70571;
  assign n70573 = pi18 ? n32 : n70572;
  assign n70574 = pi17 ? n32 : n70573;
  assign n70575 = pi16 ? n32 : n70574;
  assign n70576 = pi15 ? n70568 : n70575;
  assign n70577 = pi22 ? n20563 : n42106;
  assign n70578 = pi21 ? n45016 : n70577;
  assign n70579 = pi20 ? n37926 : n70578;
  assign n70580 = pi22 ? n56607 : n59672;
  assign n70581 = pi21 ? n39972 : n70580;
  assign n70582 = pi20 ? n70581 : n32;
  assign n70583 = pi19 ? n70579 : n70582;
  assign n70584 = pi18 ? n32 : n70583;
  assign n70585 = pi17 ? n32 : n70584;
  assign n70586 = pi16 ? n32 : n70585;
  assign n70587 = pi21 ? n40986 : n45016;
  assign n70588 = pi20 ? n37926 : n70587;
  assign n70589 = pi21 ? n14626 : n62849;
  assign n70590 = pi20 ? n70589 : n32;
  assign n70591 = pi19 ? n70588 : n70590;
  assign n70592 = pi18 ? n32 : n70591;
  assign n70593 = pi17 ? n32 : n70592;
  assign n70594 = pi16 ? n32 : n70593;
  assign n70595 = pi15 ? n70586 : n70594;
  assign n70596 = pi14 ? n70576 : n70595;
  assign n70597 = pi21 ? n40960 : n40986;
  assign n70598 = pi20 ? n37926 : n70597;
  assign n70599 = pi24 ? n14626 : n316;
  assign n70600 = pi23 ? n14626 : n70599;
  assign n70601 = pi22 ? n70600 : n32;
  assign n70602 = pi21 ? n51564 : n70601;
  assign n70603 = pi20 ? n70602 : n32;
  assign n70604 = pi19 ? n70598 : n70603;
  assign n70605 = pi18 ? n32 : n70604;
  assign n70606 = pi17 ? n32 : n70605;
  assign n70607 = pi16 ? n32 : n70606;
  assign n70608 = pi22 ? n33792 : n37288;
  assign n70609 = pi21 ? n54446 : n70608;
  assign n70610 = pi20 ? n51731 : n70609;
  assign n70611 = pi21 ? n51564 : n59673;
  assign n70612 = pi20 ? n70611 : n32;
  assign n70613 = pi19 ? n70610 : n70612;
  assign n70614 = pi18 ? n32 : n70613;
  assign n70615 = pi17 ? n32 : n70614;
  assign n70616 = pi16 ? n32 : n70615;
  assign n70617 = pi15 ? n70607 : n70616;
  assign n70618 = pi21 ? n51762 : n36659;
  assign n70619 = pi20 ? n51756 : n70618;
  assign n70620 = pi21 ? n59595 : n54564;
  assign n70621 = pi20 ? n70620 : n32;
  assign n70622 = pi19 ? n70619 : n70621;
  assign n70623 = pi18 ? n32 : n70622;
  assign n70624 = pi17 ? n32 : n70623;
  assign n70625 = pi16 ? n32 : n70624;
  assign n70626 = pi21 ? n51270 : n36781;
  assign n70627 = pi20 ? n40054 : n70626;
  assign n70628 = pi23 ? n56620 : n14626;
  assign n70629 = pi22 ? n70628 : n13481;
  assign n70630 = pi21 ? n70629 : n37639;
  assign n70631 = pi20 ? n70630 : n32;
  assign n70632 = pi19 ? n70627 : n70631;
  assign n70633 = pi18 ? n32 : n70632;
  assign n70634 = pi17 ? n32 : n70633;
  assign n70635 = pi16 ? n32 : n70634;
  assign n70636 = pi15 ? n70625 : n70635;
  assign n70637 = pi14 ? n70617 : n70636;
  assign n70638 = pi13 ? n70596 : n70637;
  assign n70639 = pi21 ? n61352 : n36781;
  assign n70640 = pi20 ? n40054 : n70639;
  assign n70641 = pi23 ? n55783 : n14626;
  assign n70642 = pi22 ? n70641 : n59672;
  assign n70643 = pi21 ? n70642 : n32;
  assign n70644 = pi20 ? n70643 : n32;
  assign n70645 = pi19 ? n70640 : n70644;
  assign n70646 = pi18 ? n32 : n70645;
  assign n70647 = pi17 ? n32 : n70646;
  assign n70648 = pi16 ? n32 : n70647;
  assign n70649 = pi20 ? n40054 : n67869;
  assign n70650 = pi22 ? n56607 : n54563;
  assign n70651 = pi21 ? n70650 : n32;
  assign n70652 = pi20 ? n70651 : n32;
  assign n70653 = pi19 ? n70649 : n70652;
  assign n70654 = pi18 ? n32 : n70653;
  assign n70655 = pi17 ? n32 : n70654;
  assign n70656 = pi16 ? n32 : n70655;
  assign n70657 = pi15 ? n70648 : n70656;
  assign n70658 = pi21 ? n62322 : n47397;
  assign n70659 = pi20 ? n40054 : n70658;
  assign n70660 = pi20 ? n67073 : n32;
  assign n70661 = pi19 ? n70659 : n70660;
  assign n70662 = pi18 ? n32 : n70661;
  assign n70663 = pi17 ? n32 : n70662;
  assign n70664 = pi16 ? n32 : n70663;
  assign n70665 = pi21 ? n69710 : n57774;
  assign n70666 = pi20 ? n40054 : n70665;
  assign n70667 = pi19 ? n70666 : n55669;
  assign n70668 = pi18 ? n32 : n70667;
  assign n70669 = pi17 ? n32 : n70668;
  assign n70670 = pi16 ? n32 : n70669;
  assign n70671 = pi15 ? n70664 : n70670;
  assign n70672 = pi14 ? n70657 : n70671;
  assign n70673 = pi21 ? n63401 : n55708;
  assign n70674 = pi20 ? n37926 : n70673;
  assign n70675 = pi20 ? n59466 : n32;
  assign n70676 = pi19 ? n70674 : n70675;
  assign n70677 = pi18 ? n32 : n70676;
  assign n70678 = pi17 ? n32 : n70677;
  assign n70679 = pi16 ? n32 : n70678;
  assign n70680 = pi21 ? n38285 : n68938;
  assign n70681 = pi20 ? n37926 : n70680;
  assign n70682 = pi19 ? n70681 : n70675;
  assign n70683 = pi18 ? n32 : n70682;
  assign n70684 = pi17 ? n32 : n70683;
  assign n70685 = pi16 ? n32 : n70684;
  assign n70686 = pi15 ? n70679 : n70685;
  assign n70687 = pi21 ? n39972 : n51564;
  assign n70688 = pi20 ? n47835 : n70687;
  assign n70689 = pi19 ? n70688 : n37641;
  assign n70690 = pi18 ? n32 : n70689;
  assign n70691 = pi17 ? n32 : n70690;
  assign n70692 = pi16 ? n32 : n70691;
  assign n70693 = pi21 ? n67068 : n51564;
  assign n70694 = pi20 ? n32 : n70693;
  assign n70695 = pi19 ? n70694 : n35482;
  assign n70696 = pi18 ? n32 : n70695;
  assign n70697 = pi17 ? n32 : n70696;
  assign n70698 = pi16 ? n32 : n70697;
  assign n70699 = pi15 ? n70692 : n70698;
  assign n70700 = pi14 ? n70686 : n70699;
  assign n70701 = pi13 ? n70672 : n70700;
  assign n70702 = pi12 ? n70638 : n70701;
  assign n70703 = pi22 ? n56712 : n14626;
  assign n70704 = pi21 ? n70703 : n13481;
  assign n70705 = pi20 ? n32 : n70704;
  assign n70706 = pi19 ? n70705 : n32;
  assign n70707 = pi18 ? n32 : n70706;
  assign n70708 = pi17 ? n32 : n70707;
  assign n70709 = pi16 ? n32 : n70708;
  assign n70710 = pi21 ? n56760 : n61184;
  assign n70711 = pi20 ? n32 : n70710;
  assign n70712 = pi19 ? n70711 : n32;
  assign n70713 = pi18 ? n32 : n70712;
  assign n70714 = pi17 ? n32 : n70713;
  assign n70715 = pi16 ? n32 : n70714;
  assign n70716 = pi15 ? n70709 : n70715;
  assign n70717 = pi22 ? n55799 : n51564;
  assign n70718 = pi21 ? n70717 : n57563;
  assign n70719 = pi20 ? n32 : n70718;
  assign n70720 = pi19 ? n70719 : n32;
  assign n70721 = pi18 ? n32 : n70720;
  assign n70722 = pi17 ? n32 : n70721;
  assign n70723 = pi16 ? n32 : n70722;
  assign n70724 = pi21 ? n55606 : n67964;
  assign n70725 = pi20 ? n32 : n70724;
  assign n70726 = pi19 ? n70725 : n32;
  assign n70727 = pi18 ? n32 : n70726;
  assign n70728 = pi17 ? n32 : n70727;
  assign n70729 = pi16 ? n32 : n70728;
  assign n70730 = pi15 ? n70723 : n70729;
  assign n70731 = pi14 ? n70716 : n70730;
  assign n70732 = pi21 ? n56760 : n37639;
  assign n70733 = pi20 ? n32 : n70732;
  assign n70734 = pi19 ? n70733 : n32;
  assign n70735 = pi18 ? n32 : n70734;
  assign n70736 = pi17 ? n32 : n70735;
  assign n70737 = pi16 ? n32 : n70736;
  assign n70738 = pi20 ? n32 : n62516;
  assign n70739 = pi19 ? n70738 : n32;
  assign n70740 = pi18 ? n32 : n70739;
  assign n70741 = pi17 ? n32 : n70740;
  assign n70742 = pi16 ? n32 : n70741;
  assign n70743 = pi15 ? n70737 : n70742;
  assign n70744 = pi23 ? n32 : n51564;
  assign n70745 = pi22 ? n70744 : n59672;
  assign n70746 = pi21 ? n70745 : n32;
  assign n70747 = pi20 ? n32 : n70746;
  assign n70748 = pi19 ? n70747 : n32;
  assign n70749 = pi18 ? n32 : n70748;
  assign n70750 = pi17 ? n32 : n70749;
  assign n70751 = pi16 ? n32 : n70750;
  assign n70752 = pi22 ? n69890 : n55688;
  assign n70753 = pi21 ? n70752 : n32;
  assign n70754 = pi20 ? n32 : n70753;
  assign n70755 = pi19 ? n70754 : n32;
  assign n70756 = pi18 ? n32 : n70755;
  assign n70757 = pi17 ? n32 : n70756;
  assign n70758 = pi16 ? n32 : n70757;
  assign n70759 = pi15 ? n70751 : n70758;
  assign n70760 = pi14 ? n70743 : n70759;
  assign n70761 = pi13 ? n70731 : n70760;
  assign n70762 = pi12 ? n70761 : n32;
  assign n70763 = pi11 ? n70702 : n70762;
  assign n70764 = pi10 ? n70559 : n70763;
  assign n70765 = pi09 ? n70363 : n70764;
  assign n70766 = pi19 ? n37956 : n70348;
  assign n70767 = pi18 ? n32 : n70766;
  assign n70768 = pi17 ? n32 : n70767;
  assign n70769 = pi16 ? n32 : n70768;
  assign n70770 = pi15 ? n32 : n70769;
  assign n70771 = pi19 ? n37956 : n70354;
  assign n70772 = pi18 ? n32 : n70771;
  assign n70773 = pi17 ? n32 : n70772;
  assign n70774 = pi16 ? n32 : n70773;
  assign n70775 = pi14 ? n70770 : n70774;
  assign n70776 = pi13 ? n32 : n70775;
  assign n70777 = pi12 ? n32 : n70776;
  assign n70778 = pi11 ? n32 : n70777;
  assign n70779 = pi10 ? n32 : n70778;
  assign n70780 = pi19 ? n37956 : n62975;
  assign n70781 = pi18 ? n32 : n70780;
  assign n70782 = pi17 ? n32 : n70781;
  assign n70783 = pi16 ? n32 : n70782;
  assign n70784 = pi19 ? n38998 : n62975;
  assign n70785 = pi18 ? n32 : n70784;
  assign n70786 = pi17 ? n32 : n70785;
  assign n70787 = pi16 ? n32 : n70786;
  assign n70788 = pi15 ? n70783 : n70787;
  assign n70789 = pi15 ? n70787 : n69917;
  assign n70790 = pi14 ? n70788 : n70789;
  assign n70791 = pi19 ? n38377 : n62954;
  assign n70792 = pi18 ? n32 : n70791;
  assign n70793 = pi17 ? n32 : n70792;
  assign n70794 = pi16 ? n32 : n70793;
  assign n70795 = pi14 ? n69927 : n70794;
  assign n70796 = pi13 ? n70790 : n70795;
  assign n70797 = pi19 ? n39454 : n62954;
  assign n70798 = pi18 ? n32 : n70797;
  assign n70799 = pi17 ? n32 : n70798;
  assign n70800 = pi16 ? n32 : n70799;
  assign n70801 = pi19 ? n28158 : n59306;
  assign n70802 = pi18 ? n32 : n70801;
  assign n70803 = pi17 ? n32 : n70802;
  assign n70804 = pi16 ? n32 : n70803;
  assign n70805 = pi22 ? n60210 : n14626;
  assign n70806 = pi21 ? n70805 : n64842;
  assign n70807 = pi20 ? n20563 : n70806;
  assign n70808 = pi19 ? n28158 : n70807;
  assign n70809 = pi18 ? n32 : n70808;
  assign n70810 = pi17 ? n32 : n70809;
  assign n70811 = pi16 ? n32 : n70810;
  assign n70812 = pi15 ? n70804 : n70811;
  assign n70813 = pi19 ? n28158 : n70399;
  assign n70814 = pi18 ? n32 : n70813;
  assign n70815 = pi17 ? n32 : n70814;
  assign n70816 = pi16 ? n32 : n70815;
  assign n70817 = pi19 ? n28158 : n70406;
  assign n70818 = pi18 ? n32 : n70817;
  assign n70819 = pi17 ? n32 : n70818;
  assign n70820 = pi16 ? n32 : n70819;
  assign n70821 = pi15 ? n70816 : n70820;
  assign n70822 = pi14 ? n70812 : n70821;
  assign n70823 = pi13 ? n70800 : n70822;
  assign n70824 = pi12 ? n70796 : n70823;
  assign n70825 = pi19 ? n30118 : n70415;
  assign n70826 = pi18 ? n32 : n70825;
  assign n70827 = pi17 ? n32 : n70826;
  assign n70828 = pi16 ? n32 : n70827;
  assign n70829 = pi19 ? n30118 : n70421;
  assign n70830 = pi18 ? n32 : n70829;
  assign n70831 = pi17 ? n32 : n70830;
  assign n70832 = pi16 ? n32 : n70831;
  assign n70833 = pi15 ? n70828 : n70832;
  assign n70834 = pi22 ? n64140 : n14626;
  assign n70835 = pi21 ? n70834 : n2637;
  assign n70836 = pi20 ? n56539 : n70835;
  assign n70837 = pi19 ? n31264 : n70836;
  assign n70838 = pi18 ? n32 : n70837;
  assign n70839 = pi17 ? n32 : n70838;
  assign n70840 = pi16 ? n32 : n70839;
  assign n70841 = pi19 ? n31264 : n70434;
  assign n70842 = pi18 ? n32 : n70841;
  assign n70843 = pi17 ? n32 : n70842;
  assign n70844 = pi16 ? n32 : n70843;
  assign n70845 = pi15 ? n70840 : n70844;
  assign n70846 = pi14 ? n70833 : n70845;
  assign n70847 = pi19 ? n31264 : n70442;
  assign n70848 = pi18 ? n32 : n70847;
  assign n70849 = pi17 ? n32 : n70848;
  assign n70850 = pi16 ? n32 : n70849;
  assign n70851 = pi20 ? n64913 : n59388;
  assign n70852 = pi19 ? n31264 : n70851;
  assign n70853 = pi18 ? n32 : n70852;
  assign n70854 = pi17 ? n32 : n70853;
  assign n70855 = pi16 ? n32 : n70854;
  assign n70856 = pi15 ? n70850 : n70855;
  assign n70857 = pi22 ? n30868 : n39954;
  assign n70858 = pi21 ? n30868 : n70857;
  assign n70859 = pi20 ? n70858 : n10297;
  assign n70860 = pi19 ? n31264 : n70859;
  assign n70861 = pi18 ? n32 : n70860;
  assign n70862 = pi17 ? n32 : n70861;
  assign n70863 = pi16 ? n32 : n70862;
  assign n70864 = pi21 ? n63179 : n20563;
  assign n70865 = pi20 ? n32 : n70864;
  assign n70866 = pi19 ? n70865 : n70473;
  assign n70867 = pi18 ? n32 : n70866;
  assign n70868 = pi17 ? n32 : n70867;
  assign n70869 = pi16 ? n32 : n70868;
  assign n70870 = pi15 ? n70863 : n70869;
  assign n70871 = pi14 ? n70856 : n70870;
  assign n70872 = pi13 ? n70846 : n70871;
  assign n70873 = pi22 ? n62333 : n45675;
  assign n70874 = pi21 ? n20563 : n70873;
  assign n70875 = pi20 ? n70874 : n70483;
  assign n70876 = pi19 ? n31314 : n70875;
  assign n70877 = pi18 ? n32 : n70876;
  assign n70878 = pi17 ? n32 : n70877;
  assign n70879 = pi16 ? n32 : n70878;
  assign n70880 = pi21 ? n40908 : n36489;
  assign n70881 = pi20 ? n32 : n70880;
  assign n70882 = pi23 ? n30868 : n56064;
  assign n70883 = pi22 ? n70882 : n70491;
  assign n70884 = pi21 ? n20563 : n70883;
  assign n70885 = pi20 ? n70884 : n70495;
  assign n70886 = pi19 ? n70881 : n70885;
  assign n70887 = pi18 ? n32 : n70886;
  assign n70888 = pi17 ? n32 : n70887;
  assign n70889 = pi16 ? n32 : n70888;
  assign n70890 = pi15 ? n70879 : n70889;
  assign n70891 = pi22 ? n41458 : n37173;
  assign n70892 = pi21 ? n70891 : n45016;
  assign n70893 = pi20 ? n32 : n70892;
  assign n70894 = pi23 ? n33792 : n8184;
  assign n70895 = pi22 ? n70894 : n43199;
  assign n70896 = pi21 ? n33792 : n70895;
  assign n70897 = pi20 ? n70896 : n59635;
  assign n70898 = pi19 ? n70893 : n70897;
  assign n70899 = pi18 ? n32 : n70898;
  assign n70900 = pi17 ? n32 : n70899;
  assign n70901 = pi16 ? n32 : n70900;
  assign n70902 = pi22 ? n41481 : n36659;
  assign n70903 = pi21 ? n70902 : n40986;
  assign n70904 = pi20 ? n32 : n70903;
  assign n70905 = pi22 ? n61761 : n69595;
  assign n70906 = pi21 ? n36659 : n70905;
  assign n70907 = pi20 ? n70906 : n4110;
  assign n70908 = pi19 ? n70904 : n70907;
  assign n70909 = pi18 ? n32 : n70908;
  assign n70910 = pi17 ? n32 : n70909;
  assign n70911 = pi16 ? n32 : n70910;
  assign n70912 = pi15 ? n70901 : n70911;
  assign n70913 = pi14 ? n70890 : n70912;
  assign n70914 = pi22 ? n41481 : n37783;
  assign n70915 = pi21 ? n70914 : n40986;
  assign n70916 = pi20 ? n32 : n70915;
  assign n70917 = pi19 ? n70916 : n70527;
  assign n70918 = pi18 ? n32 : n70917;
  assign n70919 = pi17 ? n32 : n70918;
  assign n70920 = pi16 ? n32 : n70919;
  assign n70921 = pi23 ? n37273 : n20563;
  assign n70922 = pi23 ? n20563 : n60408;
  assign n70923 = pi22 ? n70921 : n70922;
  assign n70924 = pi21 ? n70923 : n40986;
  assign n70925 = pi20 ? n32 : n70924;
  assign n70926 = pi23 ? n36659 : n59957;
  assign n70927 = pi22 ? n70926 : n65935;
  assign n70928 = pi21 ? n36659 : n70927;
  assign n70929 = pi20 ? n70928 : n59674;
  assign n70930 = pi19 ? n70925 : n70929;
  assign n70931 = pi18 ? n32 : n70930;
  assign n70932 = pi17 ? n32 : n70931;
  assign n70933 = pi16 ? n32 : n70932;
  assign n70934 = pi15 ? n70920 : n70933;
  assign n70935 = pi23 ? n14626 : n58538;
  assign n70936 = pi22 ? n70935 : n56607;
  assign n70937 = pi21 ? n36659 : n70936;
  assign n70938 = pi20 ? n70937 : n54565;
  assign n70939 = pi19 ? n31314 : n70938;
  assign n70940 = pi18 ? n32 : n70939;
  assign n70941 = pi17 ? n32 : n70940;
  assign n70942 = pi16 ? n32 : n70941;
  assign n70943 = pi22 ? n62283 : n57659;
  assign n70944 = pi21 ? n36659 : n70943;
  assign n70945 = pi20 ? n70944 : n37640;
  assign n70946 = pi19 ? n31264 : n70945;
  assign n70947 = pi18 ? n32 : n70946;
  assign n70948 = pi17 ? n32 : n70947;
  assign n70949 = pi16 ? n32 : n70948;
  assign n70950 = pi15 ? n70942 : n70949;
  assign n70951 = pi14 ? n70934 : n70950;
  assign n70952 = pi13 ? n70913 : n70951;
  assign n70953 = pi12 ? n70872 : n70952;
  assign n70954 = pi11 ? n70824 : n70953;
  assign n70955 = pi23 ? n36782 : n20563;
  assign n70956 = pi22 ? n70955 : n30868;
  assign n70957 = pi21 ? n70956 : n20563;
  assign n70958 = pi20 ? n32 : n70957;
  assign n70959 = pi23 ? n51564 : n57029;
  assign n70960 = pi22 ? n70959 : n65432;
  assign n70961 = pi21 ? n36781 : n70960;
  assign n70962 = pi20 ? n70961 : n32;
  assign n70963 = pi19 ? n70958 : n70962;
  assign n70964 = pi18 ? n32 : n70963;
  assign n70965 = pi17 ? n32 : n70964;
  assign n70966 = pi16 ? n32 : n70965;
  assign n70967 = pi21 ? n68255 : n20563;
  assign n70968 = pi20 ? n32 : n70967;
  assign n70969 = pi22 ? n14626 : n59672;
  assign n70970 = pi21 ? n39972 : n70969;
  assign n70971 = pi20 ? n70970 : n32;
  assign n70972 = pi19 ? n70968 : n70971;
  assign n70973 = pi18 ? n32 : n70972;
  assign n70974 = pi17 ? n32 : n70973;
  assign n70975 = pi16 ? n32 : n70974;
  assign n70976 = pi15 ? n70966 : n70975;
  assign n70977 = pi21 ? n68279 : n36489;
  assign n70978 = pi20 ? n32 : n70977;
  assign n70979 = pi23 ? n43198 : n67465;
  assign n70980 = pi22 ? n70979 : n59672;
  assign n70981 = pi21 ? n39972 : n70980;
  assign n70982 = pi20 ? n70981 : n32;
  assign n70983 = pi19 ? n70978 : n70982;
  assign n70984 = pi18 ? n32 : n70983;
  assign n70985 = pi17 ? n32 : n70984;
  assign n70986 = pi16 ? n32 : n70985;
  assign n70987 = pi22 ? n70921 : n36659;
  assign n70988 = pi21 ? n70987 : n68602;
  assign n70989 = pi20 ? n32 : n70988;
  assign n70990 = pi19 ? n70989 : n70590;
  assign n70991 = pi18 ? n32 : n70990;
  assign n70992 = pi17 ? n32 : n70991;
  assign n70993 = pi16 ? n32 : n70992;
  assign n70994 = pi15 ? n70986 : n70993;
  assign n70995 = pi14 ? n70976 : n70994;
  assign n70996 = pi22 ? n30865 : n30867;
  assign n70997 = pi21 ? n70996 : n40986;
  assign n70998 = pi20 ? n32 : n70997;
  assign n70999 = pi19 ? n70998 : n70603;
  assign n71000 = pi18 ? n32 : n70999;
  assign n71001 = pi17 ? n32 : n71000;
  assign n71002 = pi16 ? n32 : n71001;
  assign n71003 = pi23 ? n34196 : n33792;
  assign n71004 = pi22 ? n71003 : n33792;
  assign n71005 = pi21 ? n71004 : n47360;
  assign n71006 = pi20 ? n32 : n71005;
  assign n71007 = pi19 ? n71006 : n70612;
  assign n71008 = pi18 ? n32 : n71007;
  assign n71009 = pi17 ? n32 : n71008;
  assign n71010 = pi16 ? n32 : n71009;
  assign n71011 = pi15 ? n71002 : n71010;
  assign n71012 = pi22 ? n41097 : n36659;
  assign n71013 = pi21 ? n71012 : n36659;
  assign n71014 = pi20 ? n32 : n71013;
  assign n71015 = pi21 ? n59595 : n58503;
  assign n71016 = pi20 ? n71015 : n32;
  assign n71017 = pi19 ? n71014 : n71016;
  assign n71018 = pi18 ? n32 : n71017;
  assign n71019 = pi17 ? n32 : n71018;
  assign n71020 = pi16 ? n32 : n71019;
  assign n71021 = pi20 ? n32 : n70626;
  assign n71022 = pi21 ? n67426 : n20952;
  assign n71023 = pi20 ? n71022 : n32;
  assign n71024 = pi19 ? n71021 : n71023;
  assign n71025 = pi18 ? n32 : n71024;
  assign n71026 = pi17 ? n32 : n71025;
  assign n71027 = pi16 ? n32 : n71026;
  assign n71028 = pi15 ? n71020 : n71027;
  assign n71029 = pi14 ? n71011 : n71028;
  assign n71030 = pi13 ? n70995 : n71029;
  assign n71031 = pi20 ? n32 : n70639;
  assign n71032 = pi23 ? n64160 : n14626;
  assign n71033 = pi22 ? n71032 : n59672;
  assign n71034 = pi21 ? n71033 : n32;
  assign n71035 = pi20 ? n71034 : n32;
  assign n71036 = pi19 ? n71031 : n71035;
  assign n71037 = pi18 ? n32 : n71036;
  assign n71038 = pi17 ? n32 : n71037;
  assign n71039 = pi16 ? n32 : n71038;
  assign n71040 = pi22 ? n30865 : n36781;
  assign n71041 = pi21 ? n71040 : n36798;
  assign n71042 = pi20 ? n32 : n71041;
  assign n71043 = pi19 ? n71042 : n70652;
  assign n71044 = pi18 ? n32 : n71043;
  assign n71045 = pi17 ? n32 : n71044;
  assign n71046 = pi16 ? n32 : n71045;
  assign n71047 = pi15 ? n71039 : n71046;
  assign n71048 = pi23 ? n20564 : n36798;
  assign n71049 = pi22 ? n71048 : n36798;
  assign n71050 = pi21 ? n71049 : n47397;
  assign n71051 = pi20 ? n32 : n71050;
  assign n71052 = pi19 ? n71051 : n70660;
  assign n71053 = pi18 ? n32 : n71052;
  assign n71054 = pi17 ? n32 : n71053;
  assign n71055 = pi16 ? n32 : n71054;
  assign n71056 = pi23 ? n20564 : n36781;
  assign n71057 = pi22 ? n71056 : n36781;
  assign n71058 = pi21 ? n71057 : n57774;
  assign n71059 = pi20 ? n32 : n71058;
  assign n71060 = pi19 ? n71059 : n56131;
  assign n71061 = pi18 ? n32 : n71060;
  assign n71062 = pi17 ? n32 : n71061;
  assign n71063 = pi16 ? n32 : n71062;
  assign n71064 = pi15 ? n71055 : n71063;
  assign n71065 = pi14 ? n71047 : n71064;
  assign n71066 = pi21 ? n41600 : n55708;
  assign n71067 = pi20 ? n32 : n71066;
  assign n71068 = pi19 ? n71067 : n70675;
  assign n71069 = pi18 ? n32 : n71068;
  assign n71070 = pi17 ? n32 : n71069;
  assign n71071 = pi16 ? n32 : n71070;
  assign n71072 = pi21 ? n45136 : n68938;
  assign n71073 = pi20 ? n32 : n71072;
  assign n71074 = pi19 ? n71073 : n70675;
  assign n71075 = pi18 ? n32 : n71074;
  assign n71076 = pi17 ? n32 : n71075;
  assign n71077 = pi16 ? n32 : n71076;
  assign n71078 = pi15 ? n71071 : n71077;
  assign n71079 = pi22 ? n45135 : n36798;
  assign n71080 = pi21 ? n71079 : n51564;
  assign n71081 = pi20 ? n32 : n71080;
  assign n71082 = pi19 ? n71081 : n37641;
  assign n71083 = pi18 ? n32 : n71082;
  assign n71084 = pi17 ? n32 : n71083;
  assign n71085 = pi16 ? n32 : n71084;
  assign n71086 = pi22 ? n45160 : n14626;
  assign n71087 = pi22 ? n51564 : n62473;
  assign n71088 = pi21 ? n71086 : n71087;
  assign n71089 = pi20 ? n32 : n71088;
  assign n71090 = pi19 ? n71089 : n32;
  assign n71091 = pi18 ? n32 : n71090;
  assign n71092 = pi17 ? n32 : n71091;
  assign n71093 = pi16 ? n32 : n71092;
  assign n71094 = pi15 ? n71085 : n71093;
  assign n71095 = pi14 ? n71078 : n71094;
  assign n71096 = pi13 ? n71065 : n71095;
  assign n71097 = pi12 ? n71030 : n71096;
  assign n71098 = pi22 ? n45652 : n14626;
  assign n71099 = pi21 ? n71098 : n59648;
  assign n71100 = pi20 ? n32 : n71099;
  assign n71101 = pi19 ? n71100 : n32;
  assign n71102 = pi18 ? n32 : n71101;
  assign n71103 = pi17 ? n32 : n71102;
  assign n71104 = pi16 ? n32 : n71103;
  assign n71105 = pi22 ? n46789 : n51564;
  assign n71106 = pi21 ? n71105 : n61184;
  assign n71107 = pi20 ? n32 : n71106;
  assign n71108 = pi19 ? n71107 : n32;
  assign n71109 = pi18 ? n32 : n71108;
  assign n71110 = pi17 ? n32 : n71109;
  assign n71111 = pi16 ? n32 : n71110;
  assign n71112 = pi15 ? n71104 : n71111;
  assign n71113 = pi22 ? n46275 : n51564;
  assign n71114 = pi21 ? n71113 : n57563;
  assign n71115 = pi20 ? n32 : n71114;
  assign n71116 = pi19 ? n71115 : n32;
  assign n71117 = pi18 ? n32 : n71116;
  assign n71118 = pi17 ? n32 : n71117;
  assign n71119 = pi16 ? n32 : n71118;
  assign n71120 = pi22 ? n32 : n13481;
  assign n71121 = pi21 ? n71120 : n67964;
  assign n71122 = pi20 ? n32 : n71121;
  assign n71123 = pi19 ? n71122 : n32;
  assign n71124 = pi18 ? n32 : n71123;
  assign n71125 = pi17 ? n32 : n71124;
  assign n71126 = pi16 ? n32 : n71125;
  assign n71127 = pi15 ? n71119 : n71126;
  assign n71128 = pi14 ? n71112 : n71127;
  assign n71129 = pi22 ? n32 : n51564;
  assign n71130 = pi21 ? n71129 : n37639;
  assign n71131 = pi20 ? n32 : n71130;
  assign n71132 = pi19 ? n71131 : n32;
  assign n71133 = pi18 ? n32 : n71132;
  assign n71134 = pi17 ? n32 : n71133;
  assign n71135 = pi16 ? n32 : n71134;
  assign n71136 = pi21 ? n71120 : n32;
  assign n71137 = pi20 ? n32 : n71136;
  assign n71138 = pi19 ? n71137 : n32;
  assign n71139 = pi18 ? n32 : n71138;
  assign n71140 = pi17 ? n32 : n71139;
  assign n71141 = pi16 ? n32 : n71140;
  assign n71142 = pi15 ? n71135 : n71141;
  assign n71143 = pi24 ? n32 : n51564;
  assign n71144 = pi23 ? n71143 : n51565;
  assign n71145 = pi22 ? n32 : n71144;
  assign n71146 = pi21 ? n71145 : n32;
  assign n71147 = pi20 ? n32 : n71146;
  assign n71148 = pi19 ? n71147 : n32;
  assign n71149 = pi18 ? n32 : n71148;
  assign n71150 = pi17 ? n32 : n71149;
  assign n71151 = pi16 ? n32 : n71150;
  assign n71152 = pi23 ? n69400 : n14362;
  assign n71153 = pi22 ? n32 : n71152;
  assign n71154 = pi21 ? n71153 : n32;
  assign n71155 = pi20 ? n32 : n71154;
  assign n71156 = pi19 ? n71155 : n32;
  assign n71157 = pi18 ? n32 : n71156;
  assign n71158 = pi17 ? n32 : n71157;
  assign n71159 = pi16 ? n32 : n71158;
  assign n71160 = pi15 ? n71151 : n71159;
  assign n71161 = pi14 ? n71142 : n71160;
  assign n71162 = pi13 ? n71128 : n71161;
  assign n71163 = pi12 ? n71162 : n32;
  assign n71164 = pi11 ? n71097 : n71163;
  assign n71165 = pi10 ? n70954 : n71164;
  assign n71166 = pi09 ? n70779 : n71165;
  assign n71167 = pi08 ? n70765 : n71166;
  assign n71168 = pi19 ? n37934 : n70348;
  assign n71169 = pi18 ? n32 : n71168;
  assign n71170 = pi17 ? n32 : n71169;
  assign n71171 = pi16 ? n32 : n71170;
  assign n71172 = pi15 ? n32 : n71171;
  assign n71173 = pi19 ? n37934 : n70354;
  assign n71174 = pi18 ? n32 : n71173;
  assign n71175 = pi17 ? n32 : n71174;
  assign n71176 = pi16 ? n32 : n71175;
  assign n71177 = pi14 ? n71172 : n71176;
  assign n71178 = pi13 ? n32 : n71177;
  assign n71179 = pi12 ? n32 : n71178;
  assign n71180 = pi11 ? n32 : n71179;
  assign n71181 = pi10 ? n32 : n71180;
  assign n71182 = pi19 ? n36868 : n62975;
  assign n71183 = pi18 ? n32 : n71182;
  assign n71184 = pi17 ? n32 : n71183;
  assign n71185 = pi16 ? n32 : n71184;
  assign n71186 = pi15 ? n71185 : n70783;
  assign n71187 = pi14 ? n71186 : n70788;
  assign n71188 = pi19 ? n37321 : n62954;
  assign n71189 = pi18 ? n32 : n71188;
  assign n71190 = pi17 ? n32 : n71189;
  assign n71191 = pi16 ? n32 : n71190;
  assign n71192 = pi14 ? n70367 : n71191;
  assign n71193 = pi13 ? n71187 : n71192;
  assign n71194 = pi19 ? n37334 : n62954;
  assign n71195 = pi18 ? n32 : n71194;
  assign n71196 = pi17 ? n32 : n71195;
  assign n71197 = pi16 ? n32 : n71196;
  assign n71198 = pi19 ? n38377 : n59306;
  assign n71199 = pi18 ? n32 : n71198;
  assign n71200 = pi17 ? n32 : n71199;
  assign n71201 = pi16 ? n32 : n71200;
  assign n71202 = pi19 ? n38377 : n70807;
  assign n71203 = pi18 ? n32 : n71202;
  assign n71204 = pi17 ? n32 : n71203;
  assign n71205 = pi16 ? n32 : n71204;
  assign n71206 = pi15 ? n71201 : n71205;
  assign n71207 = pi19 ? n38377 : n70399;
  assign n71208 = pi18 ? n32 : n71207;
  assign n71209 = pi17 ? n32 : n71208;
  assign n71210 = pi16 ? n32 : n71209;
  assign n71211 = pi21 ? n68565 : n3523;
  assign n71212 = pi20 ? n20563 : n71211;
  assign n71213 = pi19 ? n38377 : n71212;
  assign n71214 = pi18 ? n32 : n71213;
  assign n71215 = pi17 ? n32 : n71214;
  assign n71216 = pi16 ? n32 : n71215;
  assign n71217 = pi15 ? n71210 : n71216;
  assign n71218 = pi14 ? n71206 : n71217;
  assign n71219 = pi13 ? n71197 : n71218;
  assign n71220 = pi12 ? n71193 : n71219;
  assign n71221 = pi19 ? n39454 : n70415;
  assign n71222 = pi18 ? n32 : n71221;
  assign n71223 = pi17 ? n32 : n71222;
  assign n71224 = pi16 ? n32 : n71223;
  assign n71225 = pi19 ? n39454 : n70421;
  assign n71226 = pi18 ? n32 : n71225;
  assign n71227 = pi17 ? n32 : n71226;
  assign n71228 = pi16 ? n32 : n71227;
  assign n71229 = pi15 ? n71224 : n71228;
  assign n71230 = pi19 ? n39454 : n70836;
  assign n71231 = pi18 ? n32 : n71230;
  assign n71232 = pi17 ? n32 : n71231;
  assign n71233 = pi16 ? n32 : n71232;
  assign n71234 = pi20 ? n47158 : n14723;
  assign n71235 = pi19 ? n39454 : n71234;
  assign n71236 = pi18 ? n32 : n71235;
  assign n71237 = pi17 ? n32 : n71236;
  assign n71238 = pi16 ? n32 : n71237;
  assign n71239 = pi15 ? n71233 : n71238;
  assign n71240 = pi14 ? n71229 : n71239;
  assign n71241 = pi20 ? n53367 : n70441;
  assign n71242 = pi19 ? n39454 : n71241;
  assign n71243 = pi18 ? n32 : n71242;
  assign n71244 = pi17 ? n32 : n71243;
  assign n71245 = pi16 ? n32 : n71244;
  assign n71246 = pi22 ? n30867 : n204;
  assign n71247 = pi21 ? n20563 : n71246;
  assign n71248 = pi20 ? n71247 : n59388;
  assign n71249 = pi19 ? n56687 : n71248;
  assign n71250 = pi18 ? n32 : n71249;
  assign n71251 = pi17 ? n32 : n71250;
  assign n71252 = pi16 ? n32 : n71251;
  assign n71253 = pi15 ? n71245 : n71252;
  assign n71254 = pi21 ? n30868 : n53408;
  assign n71255 = pi20 ? n71254 : n68625;
  assign n71256 = pi19 ? n39454 : n71255;
  assign n71257 = pi18 ? n32 : n71256;
  assign n71258 = pi17 ? n32 : n71257;
  assign n71259 = pi16 ? n32 : n71258;
  assign n71260 = pi22 ? n33792 : n14626;
  assign n71261 = pi21 ? n30868 : n71260;
  assign n71262 = pi20 ? n71261 : n67702;
  assign n71263 = pi19 ? n39454 : n71262;
  assign n71264 = pi18 ? n32 : n71263;
  assign n71265 = pi17 ? n32 : n71264;
  assign n71266 = pi16 ? n32 : n71265;
  assign n71267 = pi15 ? n71259 : n71266;
  assign n71268 = pi14 ? n71253 : n71267;
  assign n71269 = pi13 ? n71240 : n71268;
  assign n71270 = pi23 ? n20563 : n56467;
  assign n71271 = pi22 ? n71270 : n204;
  assign n71272 = pi21 ? n20563 : n71271;
  assign n71273 = pi20 ? n71272 : n67719;
  assign n71274 = pi19 ? n28158 : n71273;
  assign n71275 = pi18 ? n32 : n71274;
  assign n71276 = pi17 ? n32 : n71275;
  assign n71277 = pi16 ? n32 : n71276;
  assign n71278 = pi21 ? n28156 : n36489;
  assign n71279 = pi20 ? n32 : n71278;
  assign n71280 = pi22 ? n62742 : n204;
  assign n71281 = pi21 ? n20563 : n71280;
  assign n71282 = pi20 ? n71281 : n6935;
  assign n71283 = pi19 ? n71279 : n71282;
  assign n71284 = pi18 ? n32 : n71283;
  assign n71285 = pi17 ? n32 : n71284;
  assign n71286 = pi16 ? n32 : n71285;
  assign n71287 = pi15 ? n71277 : n71286;
  assign n71288 = pi21 ? n30116 : n45016;
  assign n71289 = pi20 ? n32 : n71288;
  assign n71290 = pi23 ? n139 : n62832;
  assign n71291 = pi22 ? n71290 : n316;
  assign n71292 = pi21 ? n33792 : n71291;
  assign n71293 = pi20 ? n71292 : n59649;
  assign n71294 = pi19 ? n71289 : n71293;
  assign n71295 = pi18 ? n32 : n71294;
  assign n71296 = pi17 ? n32 : n71295;
  assign n71297 = pi16 ? n32 : n71296;
  assign n71298 = pi21 ? n30116 : n40986;
  assign n71299 = pi20 ? n32 : n71298;
  assign n71300 = pi22 ? n61761 : n63317;
  assign n71301 = pi21 ? n36659 : n71300;
  assign n71302 = pi20 ? n71301 : n65434;
  assign n71303 = pi19 ? n71299 : n71302;
  assign n71304 = pi18 ? n32 : n71303;
  assign n71305 = pi17 ? n32 : n71304;
  assign n71306 = pi16 ? n32 : n71305;
  assign n71307 = pi15 ? n71297 : n71306;
  assign n71308 = pi14 ? n71287 : n71307;
  assign n71309 = pi22 ? n40386 : n36659;
  assign n71310 = pi21 ? n30116 : n71309;
  assign n71311 = pi20 ? n32 : n71310;
  assign n71312 = pi22 ? n39976 : n57632;
  assign n71313 = pi21 ? n36659 : n71312;
  assign n71314 = pi20 ? n71313 : n4116;
  assign n71315 = pi19 ? n71311 : n71314;
  assign n71316 = pi18 ? n32 : n71315;
  assign n71317 = pi17 ? n32 : n71316;
  assign n71318 = pi16 ? n32 : n71317;
  assign n71319 = pi21 ? n54400 : n40986;
  assign n71320 = pi20 ? n32 : n71319;
  assign n71321 = pi22 ? n70926 : n2299;
  assign n71322 = pi21 ? n36659 : n71321;
  assign n71323 = pi20 ? n71322 : n51568;
  assign n71324 = pi19 ? n71320 : n71323;
  assign n71325 = pi18 ? n32 : n71324;
  assign n71326 = pi17 ? n32 : n71325;
  assign n71327 = pi16 ? n32 : n71326;
  assign n71328 = pi15 ? n71318 : n71327;
  assign n71329 = pi21 ? n58576 : n40954;
  assign n71330 = pi20 ? n32 : n71329;
  assign n71331 = pi23 ? n157 : n58538;
  assign n71332 = pi22 ? n71331 : n57659;
  assign n71333 = pi21 ? n36659 : n71332;
  assign n71334 = pi20 ? n71333 : n55690;
  assign n71335 = pi19 ? n71330 : n71334;
  assign n71336 = pi18 ? n32 : n71335;
  assign n71337 = pi17 ? n32 : n71336;
  assign n71338 = pi16 ? n32 : n71337;
  assign n71339 = pi21 ? n58576 : n45092;
  assign n71340 = pi20 ? n32 : n71339;
  assign n71341 = pi23 ? n157 : n57517;
  assign n71342 = pi22 ? n71341 : n56678;
  assign n71343 = pi21 ? n36659 : n71342;
  assign n71344 = pi20 ? n71343 : n32;
  assign n71345 = pi19 ? n71340 : n71344;
  assign n71346 = pi18 ? n32 : n71345;
  assign n71347 = pi17 ? n32 : n71346;
  assign n71348 = pi16 ? n32 : n71347;
  assign n71349 = pi15 ? n71338 : n71348;
  assign n71350 = pi14 ? n71328 : n71349;
  assign n71351 = pi13 ? n71308 : n71350;
  assign n71352 = pi12 ? n71269 : n71351;
  assign n71353 = pi11 ? n71220 : n71352;
  assign n71354 = pi22 ? n46757 : n39190;
  assign n71355 = pi22 ? n45106 : n39190;
  assign n71356 = pi21 ? n71354 : n71355;
  assign n71357 = pi20 ? n32 : n71356;
  assign n71358 = pi23 ? n204 : n58566;
  assign n71359 = pi22 ? n71358 : n66784;
  assign n71360 = pi21 ? n36781 : n71359;
  assign n71361 = pi20 ? n71360 : n32;
  assign n71362 = pi19 ? n71357 : n71361;
  assign n71363 = pi18 ? n32 : n71362;
  assign n71364 = pi17 ? n32 : n71363;
  assign n71365 = pi16 ? n32 : n71364;
  assign n71366 = pi23 ? n36781 : n30868;
  assign n71367 = pi22 ? n71366 : n39190;
  assign n71368 = pi21 ? n70144 : n71367;
  assign n71369 = pi20 ? n32 : n71368;
  assign n71370 = pi22 ? n14626 : n51566;
  assign n71371 = pi21 ? n39972 : n71370;
  assign n71372 = pi20 ? n71371 : n32;
  assign n71373 = pi19 ? n71369 : n71372;
  assign n71374 = pi18 ? n32 : n71373;
  assign n71375 = pi17 ? n32 : n71374;
  assign n71376 = pi16 ? n32 : n71375;
  assign n71377 = pi15 ? n71365 : n71376;
  assign n71378 = pi22 ? n45634 : n33792;
  assign n71379 = pi22 ? n38271 : n42109;
  assign n71380 = pi21 ? n71378 : n71379;
  assign n71381 = pi20 ? n32 : n71380;
  assign n71382 = pi23 ? n233 : n65601;
  assign n71383 = pi23 ? n13481 : n51565;
  assign n71384 = pi22 ? n71382 : n71383;
  assign n71385 = pi21 ? n39972 : n71384;
  assign n71386 = pi20 ? n71385 : n32;
  assign n71387 = pi19 ? n71381 : n71386;
  assign n71388 = pi18 ? n32 : n71387;
  assign n71389 = pi17 ? n32 : n71388;
  assign n71390 = pi16 ? n32 : n71389;
  assign n71391 = pi22 ? n45634 : n58710;
  assign n71392 = pi22 ? n36659 : n66336;
  assign n71393 = pi21 ? n71391 : n71392;
  assign n71394 = pi20 ? n32 : n71393;
  assign n71395 = pi21 ? n14626 : n57198;
  assign n71396 = pi20 ? n71395 : n32;
  assign n71397 = pi19 ? n71394 : n71396;
  assign n71398 = pi18 ? n32 : n71397;
  assign n71399 = pi17 ? n32 : n71398;
  assign n71400 = pi16 ? n32 : n71399;
  assign n71401 = pi15 ? n71390 : n71400;
  assign n71402 = pi14 ? n71377 : n71401;
  assign n71403 = pi22 ? n40386 : n58710;
  assign n71404 = pi21 ? n28156 : n71403;
  assign n71405 = pi20 ? n32 : n71404;
  assign n71406 = pi24 ? n51564 : n316;
  assign n71407 = pi23 ? n685 : n71406;
  assign n71408 = pi22 ? n71407 : n32;
  assign n71409 = pi21 ? n51564 : n71408;
  assign n71410 = pi20 ? n71409 : n32;
  assign n71411 = pi19 ? n71405 : n71410;
  assign n71412 = pi18 ? n32 : n71411;
  assign n71413 = pi17 ? n32 : n71412;
  assign n71414 = pi16 ? n32 : n71413;
  assign n71415 = pi22 ? n32 : n37173;
  assign n71416 = pi21 ? n71415 : n67291;
  assign n71417 = pi20 ? n32 : n71416;
  assign n71418 = pi21 ? n51564 : n51567;
  assign n71419 = pi20 ? n71418 : n32;
  assign n71420 = pi19 ? n71417 : n71419;
  assign n71421 = pi18 ? n32 : n71420;
  assign n71422 = pi17 ? n32 : n71421;
  assign n71423 = pi16 ? n32 : n71422;
  assign n71424 = pi15 ? n71414 : n71423;
  assign n71425 = pi22 ? n36659 : n38284;
  assign n71426 = pi21 ? n30155 : n71425;
  assign n71427 = pi20 ? n32 : n71426;
  assign n71428 = pi21 ? n60463 : n928;
  assign n71429 = pi20 ? n71428 : n32;
  assign n71430 = pi19 ? n71427 : n71429;
  assign n71431 = pi18 ? n32 : n71430;
  assign n71432 = pi17 ? n32 : n71431;
  assign n71433 = pi16 ? n32 : n71432;
  assign n71434 = pi21 ? n30155 : n36781;
  assign n71435 = pi20 ? n32 : n71434;
  assign n71436 = pi21 ? n64697 : n32;
  assign n71437 = pi20 ? n71436 : n32;
  assign n71438 = pi19 ? n71435 : n71437;
  assign n71439 = pi18 ? n32 : n71438;
  assign n71440 = pi17 ? n32 : n71439;
  assign n71441 = pi16 ? n32 : n71440;
  assign n71442 = pi15 ? n71433 : n71441;
  assign n71443 = pi14 ? n71424 : n71442;
  assign n71444 = pi13 ? n71402 : n71443;
  assign n71445 = pi22 ? n47380 : n49412;
  assign n71446 = pi21 ? n30116 : n71445;
  assign n71447 = pi20 ? n32 : n71446;
  assign n71448 = pi22 ? n51564 : n71383;
  assign n71449 = pi21 ? n71448 : n32;
  assign n71450 = pi20 ? n71449 : n32;
  assign n71451 = pi19 ? n71447 : n71450;
  assign n71452 = pi18 ? n32 : n71451;
  assign n71453 = pi17 ? n32 : n71452;
  assign n71454 = pi16 ? n32 : n71453;
  assign n71455 = pi22 ? n32 : n54574;
  assign n71456 = pi21 ? n71455 : n53551;
  assign n71457 = pi20 ? n32 : n71456;
  assign n71458 = pi22 ? n61484 : n55688;
  assign n71459 = pi21 ? n71458 : n32;
  assign n71460 = pi20 ? n71459 : n32;
  assign n71461 = pi19 ? n71457 : n71460;
  assign n71462 = pi18 ? n32 : n71461;
  assign n71463 = pi17 ? n32 : n71462;
  assign n71464 = pi16 ? n32 : n71463;
  assign n71465 = pi15 ? n71454 : n71464;
  assign n71466 = pi22 ? n32 : n37276;
  assign n71467 = pi21 ? n71466 : n62511;
  assign n71468 = pi20 ? n32 : n71467;
  assign n71469 = pi20 ? n64354 : n32;
  assign n71470 = pi19 ? n71468 : n71469;
  assign n71471 = pi18 ? n32 : n71470;
  assign n71472 = pi17 ? n32 : n71471;
  assign n71473 = pi16 ? n32 : n71472;
  assign n71474 = pi22 ? n32 : n58736;
  assign n71475 = pi22 ? n62510 : n55641;
  assign n71476 = pi21 ? n71474 : n71475;
  assign n71477 = pi20 ? n32 : n71476;
  assign n71478 = pi19 ? n71477 : n67389;
  assign n71479 = pi18 ? n32 : n71478;
  assign n71480 = pi17 ? n32 : n71479;
  assign n71481 = pi16 ? n32 : n71480;
  assign n71482 = pi15 ? n71473 : n71481;
  assign n71483 = pi14 ? n71465 : n71482;
  assign n71484 = pi22 ? n32 : n37288;
  assign n71485 = pi22 ? n64229 : n14626;
  assign n71486 = pi21 ? n71484 : n71485;
  assign n71487 = pi20 ? n32 : n71486;
  assign n71488 = pi19 ? n71487 : n70675;
  assign n71489 = pi18 ? n32 : n71488;
  assign n71490 = pi17 ? n32 : n71489;
  assign n71491 = pi16 ? n32 : n71490;
  assign n71492 = pi21 ? n65263 : n64307;
  assign n71493 = pi20 ? n32 : n71492;
  assign n71494 = pi19 ? n71493 : n37641;
  assign n71495 = pi18 ? n32 : n71494;
  assign n71496 = pi17 ? n32 : n71495;
  assign n71497 = pi16 ? n32 : n71496;
  assign n71498 = pi15 ? n71491 : n71497;
  assign n71499 = pi21 ? n46727 : n64335;
  assign n71500 = pi20 ? n32 : n71499;
  assign n71501 = pi19 ? n71500 : n37641;
  assign n71502 = pi18 ? n32 : n71501;
  assign n71503 = pi17 ? n32 : n71502;
  assign n71504 = pi16 ? n32 : n71503;
  assign n71505 = pi23 ? n36830 : n51564;
  assign n71506 = pi22 ? n32 : n71505;
  assign n71507 = pi21 ? n71506 : n69293;
  assign n71508 = pi20 ? n32 : n71507;
  assign n71509 = pi19 ? n71508 : n32;
  assign n71510 = pi18 ? n32 : n71509;
  assign n71511 = pi17 ? n32 : n71510;
  assign n71512 = pi16 ? n32 : n71511;
  assign n71513 = pi15 ? n71504 : n71512;
  assign n71514 = pi14 ? n71498 : n71513;
  assign n71515 = pi13 ? n71483 : n71514;
  assign n71516 = pi12 ? n71444 : n71515;
  assign n71517 = pi21 ? n48856 : n59648;
  assign n71518 = pi20 ? n32 : n71517;
  assign n71519 = pi19 ? n71518 : n32;
  assign n71520 = pi18 ? n32 : n71519;
  assign n71521 = pi17 ? n32 : n71520;
  assign n71522 = pi16 ? n32 : n71521;
  assign n71523 = pi23 ? n46274 : n13481;
  assign n71524 = pi22 ? n32 : n71523;
  assign n71525 = pi21 ? n71524 : n61184;
  assign n71526 = pi20 ? n32 : n71525;
  assign n71527 = pi19 ? n71526 : n32;
  assign n71528 = pi18 ? n32 : n71527;
  assign n71529 = pi17 ? n32 : n71528;
  assign n71530 = pi16 ? n32 : n71529;
  assign n71531 = pi15 ? n71522 : n71530;
  assign n71532 = pi23 ? n32 : n60075;
  assign n71533 = pi22 ? n32 : n71532;
  assign n71534 = pi21 ? n71533 : n56129;
  assign n71535 = pi20 ? n32 : n71534;
  assign n71536 = pi19 ? n71535 : n32;
  assign n71537 = pi18 ? n32 : n71536;
  assign n71538 = pi17 ? n32 : n71537;
  assign n71539 = pi16 ? n32 : n71538;
  assign n71540 = pi23 ? n32 : n71143;
  assign n71541 = pi22 ? n32 : n71540;
  assign n71542 = pi21 ? n71541 : n32;
  assign n71543 = pi20 ? n32 : n71542;
  assign n71544 = pi19 ? n71543 : n32;
  assign n71545 = pi18 ? n32 : n71544;
  assign n71546 = pi17 ? n32 : n71545;
  assign n71547 = pi16 ? n32 : n71546;
  assign n71548 = pi15 ? n71539 : n71547;
  assign n71549 = pi14 ? n71531 : n71548;
  assign n71550 = pi21 ? n70313 : n32;
  assign n71551 = pi20 ? n32 : n71550;
  assign n71552 = pi19 ? n71551 : n32;
  assign n71553 = pi18 ? n32 : n71552;
  assign n71554 = pi17 ? n32 : n71553;
  assign n71555 = pi16 ? n32 : n71554;
  assign n71556 = pi15 ? n71547 : n71555;
  assign n71557 = pi23 ? n32 : n51565;
  assign n71558 = pi22 ? n32 : n71557;
  assign n71559 = pi21 ? n71558 : n32;
  assign n71560 = pi20 ? n32 : n71559;
  assign n71561 = pi19 ? n71560 : n32;
  assign n71562 = pi18 ? n32 : n71561;
  assign n71563 = pi17 ? n32 : n71562;
  assign n71564 = pi16 ? n32 : n71563;
  assign n71565 = pi23 ? n32 : n14362;
  assign n71566 = pi22 ? n32 : n71565;
  assign n71567 = pi21 ? n71566 : n32;
  assign n71568 = pi20 ? n32 : n71567;
  assign n71569 = pi19 ? n71568 : n32;
  assign n71570 = pi18 ? n32 : n71569;
  assign n71571 = pi17 ? n32 : n71570;
  assign n71572 = pi16 ? n32 : n71571;
  assign n71573 = pi15 ? n71564 : n71572;
  assign n71574 = pi14 ? n71556 : n71573;
  assign n71575 = pi13 ? n71549 : n71574;
  assign n71576 = pi12 ? n71575 : n32;
  assign n71577 = pi11 ? n71516 : n71576;
  assign n71578 = pi10 ? n71353 : n71577;
  assign n71579 = pi09 ? n71181 : n71578;
  assign n71580 = pi19 ? n38982 : n70348;
  assign n71581 = pi18 ? n32 : n71580;
  assign n71582 = pi17 ? n32 : n71581;
  assign n71583 = pi16 ? n32 : n71582;
  assign n71584 = pi15 ? n32 : n71583;
  assign n71585 = pi19 ? n38982 : n70354;
  assign n71586 = pi18 ? n32 : n71585;
  assign n71587 = pi17 ? n32 : n71586;
  assign n71588 = pi16 ? n32 : n71587;
  assign n71589 = pi14 ? n71584 : n71588;
  assign n71590 = pi13 ? n32 : n71589;
  assign n71591 = pi12 ? n32 : n71590;
  assign n71592 = pi11 ? n32 : n71591;
  assign n71593 = pi10 ? n32 : n71592;
  assign n71594 = pi19 ? n40055 : n62975;
  assign n71595 = pi18 ? n32 : n71594;
  assign n71596 = pi17 ? n32 : n71595;
  assign n71597 = pi16 ? n32 : n71596;
  assign n71598 = pi19 ? n37934 : n62975;
  assign n71599 = pi18 ? n32 : n71598;
  assign n71600 = pi17 ? n32 : n71599;
  assign n71601 = pi16 ? n32 : n71600;
  assign n71602 = pi15 ? n71597 : n71601;
  assign n71603 = pi15 ? n71601 : n70783;
  assign n71604 = pi14 ? n71602 : n71603;
  assign n71605 = pi19 ? n38998 : n62954;
  assign n71606 = pi18 ? n32 : n71605;
  assign n71607 = pi17 ? n32 : n71606;
  assign n71608 = pi16 ? n32 : n71607;
  assign n71609 = pi14 ? n70787 : n71608;
  assign n71610 = pi13 ? n71604 : n71609;
  assign n71611 = pi19 ? n37321 : n59306;
  assign n71612 = pi18 ? n32 : n71611;
  assign n71613 = pi17 ? n32 : n71612;
  assign n71614 = pi16 ? n32 : n71613;
  assign n71615 = pi19 ? n37321 : n70807;
  assign n71616 = pi18 ? n32 : n71615;
  assign n71617 = pi17 ? n32 : n71616;
  assign n71618 = pi16 ? n32 : n71617;
  assign n71619 = pi15 ? n71614 : n71618;
  assign n71620 = pi19 ? n37321 : n70399;
  assign n71621 = pi18 ? n32 : n71620;
  assign n71622 = pi17 ? n32 : n71621;
  assign n71623 = pi16 ? n32 : n71622;
  assign n71624 = pi19 ? n37321 : n71212;
  assign n71625 = pi18 ? n32 : n71624;
  assign n71626 = pi17 ? n32 : n71625;
  assign n71627 = pi16 ? n32 : n71626;
  assign n71628 = pi15 ? n71623 : n71627;
  assign n71629 = pi14 ? n71619 : n71628;
  assign n71630 = pi13 ? n71608 : n71629;
  assign n71631 = pi12 ? n71610 : n71630;
  assign n71632 = pi19 ? n37334 : n70415;
  assign n71633 = pi18 ? n32 : n71632;
  assign n71634 = pi17 ? n32 : n71633;
  assign n71635 = pi16 ? n32 : n71634;
  assign n71636 = pi19 ? n37334 : n70421;
  assign n71637 = pi18 ? n32 : n71636;
  assign n71638 = pi17 ? n32 : n71637;
  assign n71639 = pi16 ? n32 : n71638;
  assign n71640 = pi15 ? n71635 : n71639;
  assign n71641 = pi22 ? n65975 : n14626;
  assign n71642 = pi21 ? n71641 : n2637;
  assign n71643 = pi20 ? n56539 : n71642;
  assign n71644 = pi19 ? n37334 : n71643;
  assign n71645 = pi18 ? n32 : n71644;
  assign n71646 = pi17 ? n32 : n71645;
  assign n71647 = pi16 ? n32 : n71646;
  assign n71648 = pi19 ? n37334 : n71234;
  assign n71649 = pi18 ? n32 : n71648;
  assign n71650 = pi17 ? n32 : n71649;
  assign n71651 = pi16 ? n32 : n71650;
  assign n71652 = pi15 ? n71647 : n71651;
  assign n71653 = pi14 ? n71640 : n71652;
  assign n71654 = pi19 ? n37334 : n71241;
  assign n71655 = pi18 ? n32 : n71654;
  assign n71656 = pi17 ? n32 : n71655;
  assign n71657 = pi16 ? n32 : n71656;
  assign n71658 = pi21 ? n37332 : n46116;
  assign n71659 = pi20 ? n32 : n71658;
  assign n71660 = pi22 ? n112 : n204;
  assign n71661 = pi21 ? n20563 : n71660;
  assign n71662 = pi20 ? n71661 : n59388;
  assign n71663 = pi19 ? n71659 : n71662;
  assign n71664 = pi18 ? n32 : n71663;
  assign n71665 = pi17 ? n32 : n71664;
  assign n71666 = pi16 ? n32 : n71665;
  assign n71667 = pi15 ? n71657 : n71666;
  assign n71668 = pi22 ? n57085 : n20563;
  assign n71669 = pi21 ? n37332 : n71668;
  assign n71670 = pi20 ? n32 : n71669;
  assign n71671 = pi19 ? n71670 : n71255;
  assign n71672 = pi18 ? n32 : n71671;
  assign n71673 = pi17 ? n32 : n71672;
  assign n71674 = pi16 ? n32 : n71673;
  assign n71675 = pi22 ? n62333 : n20563;
  assign n71676 = pi21 ? n37332 : n71675;
  assign n71677 = pi20 ? n32 : n71676;
  assign n71678 = pi19 ? n71677 : n71262;
  assign n71679 = pi18 ? n32 : n71678;
  assign n71680 = pi17 ? n32 : n71679;
  assign n71681 = pi16 ? n32 : n71680;
  assign n71682 = pi15 ? n71674 : n71681;
  assign n71683 = pi14 ? n71667 : n71682;
  assign n71684 = pi13 ? n71653 : n71683;
  assign n71685 = pi22 ? n745 : n204;
  assign n71686 = pi21 ? n20563 : n71685;
  assign n71687 = pi20 ? n71686 : n67719;
  assign n71688 = pi19 ? n38377 : n71687;
  assign n71689 = pi18 ? n32 : n71688;
  assign n71690 = pi17 ? n32 : n71689;
  assign n71691 = pi16 ? n32 : n71690;
  assign n71692 = pi22 ? n63623 : n204;
  assign n71693 = pi21 ? n20563 : n71692;
  assign n71694 = pi20 ? n71693 : n6935;
  assign n71695 = pi19 ? n67802 : n71694;
  assign n71696 = pi18 ? n32 : n71695;
  assign n71697 = pi17 ? n32 : n71696;
  assign n71698 = pi16 ? n32 : n71697;
  assign n71699 = pi15 ? n71691 : n71698;
  assign n71700 = pi23 ? n139 : n55580;
  assign n71701 = pi22 ? n71700 : n316;
  assign n71702 = pi21 ? n33792 : n71701;
  assign n71703 = pi20 ? n71702 : n59649;
  assign n71704 = pi19 ? n67822 : n71703;
  assign n71705 = pi18 ? n32 : n71704;
  assign n71706 = pi17 ? n32 : n71705;
  assign n71707 = pi16 ? n32 : n71706;
  assign n71708 = pi20 ? n32 : n66358;
  assign n71709 = pi23 ? n33792 : n63194;
  assign n71710 = pi23 ? n157 : n14626;
  assign n71711 = pi22 ? n71709 : n71710;
  assign n71712 = pi21 ? n36659 : n71711;
  assign n71713 = pi20 ? n71712 : n65434;
  assign n71714 = pi19 ? n71708 : n71713;
  assign n71715 = pi18 ? n32 : n71714;
  assign n71716 = pi17 ? n32 : n71715;
  assign n71717 = pi16 ? n32 : n71716;
  assign n71718 = pi15 ? n71707 : n71717;
  assign n71719 = pi14 ? n71699 : n71718;
  assign n71720 = pi23 ? n335 : n59957;
  assign n71721 = pi22 ? n71720 : n3762;
  assign n71722 = pi21 ? n36659 : n71721;
  assign n71723 = pi20 ? n71722 : n4116;
  assign n71724 = pi19 ? n71708 : n71723;
  assign n71725 = pi18 ? n32 : n71724;
  assign n71726 = pi17 ? n32 : n71725;
  assign n71727 = pi16 ? n32 : n71726;
  assign n71728 = pi22 ? n60396 : n2299;
  assign n71729 = pi21 ? n36659 : n71728;
  assign n71730 = pi20 ? n71729 : n10011;
  assign n71731 = pi19 ? n71708 : n71730;
  assign n71732 = pi18 ? n32 : n71731;
  assign n71733 = pi17 ? n32 : n71732;
  assign n71734 = pi16 ? n32 : n71733;
  assign n71735 = pi15 ? n71727 : n71734;
  assign n71736 = pi22 ? n71341 : n57659;
  assign n71737 = pi21 ? n36659 : n71736;
  assign n71738 = pi20 ? n71737 : n57716;
  assign n71739 = pi19 ? n39454 : n71738;
  assign n71740 = pi18 ? n32 : n71739;
  assign n71741 = pi17 ? n32 : n71740;
  assign n71742 = pi16 ? n32 : n71741;
  assign n71743 = pi22 ? n18448 : n56678;
  assign n71744 = pi21 ? n36659 : n71743;
  assign n71745 = pi20 ? n71744 : n32;
  assign n71746 = pi19 ? n38377 : n71745;
  assign n71747 = pi18 ? n32 : n71746;
  assign n71748 = pi17 ? n32 : n71747;
  assign n71749 = pi16 ? n32 : n71748;
  assign n71750 = pi15 ? n71742 : n71749;
  assign n71751 = pi14 ? n71735 : n71750;
  assign n71752 = pi13 ? n71719 : n71751;
  assign n71753 = pi12 ? n71684 : n71752;
  assign n71754 = pi11 ? n71631 : n71753;
  assign n71755 = pi21 ? n45620 : n39190;
  assign n71756 = pi20 ? n32 : n71755;
  assign n71757 = pi22 ? n71358 : n54520;
  assign n71758 = pi21 ? n36781 : n71757;
  assign n71759 = pi20 ? n71758 : n32;
  assign n71760 = pi19 ? n71756 : n71759;
  assign n71761 = pi18 ? n32 : n71760;
  assign n71762 = pi17 ? n32 : n71761;
  assign n71763 = pi16 ? n32 : n71762;
  assign n71764 = pi21 ? n45598 : n48173;
  assign n71765 = pi20 ? n32 : n71764;
  assign n71766 = pi22 ? n14626 : n19696;
  assign n71767 = pi21 ? n39972 : n71766;
  assign n71768 = pi20 ? n71767 : n32;
  assign n71769 = pi19 ? n71765 : n71768;
  assign n71770 = pi18 ? n32 : n71769;
  assign n71771 = pi17 ? n32 : n71770;
  assign n71772 = pi16 ? n32 : n71771;
  assign n71773 = pi15 ? n71763 : n71772;
  assign n71774 = pi22 ? n37173 : n42109;
  assign n71775 = pi21 ? n47768 : n71774;
  assign n71776 = pi20 ? n32 : n71775;
  assign n71777 = pi22 ? n71382 : n56665;
  assign n71778 = pi21 ? n39972 : n71777;
  assign n71779 = pi20 ? n71778 : n32;
  assign n71780 = pi19 ? n71776 : n71779;
  assign n71781 = pi18 ? n32 : n71780;
  assign n71782 = pi17 ? n32 : n71781;
  assign n71783 = pi16 ? n32 : n71782;
  assign n71784 = pi22 ? n32 : n37873;
  assign n71785 = pi21 ? n71784 : n67832;
  assign n71786 = pi20 ? n32 : n71785;
  assign n71787 = pi23 ? n14626 : n71406;
  assign n71788 = pi22 ? n71787 : n32;
  assign n71789 = pi21 ? n14626 : n71788;
  assign n71790 = pi20 ? n71789 : n32;
  assign n71791 = pi19 ? n71786 : n71790;
  assign n71792 = pi18 ? n32 : n71791;
  assign n71793 = pi17 ? n32 : n71792;
  assign n71794 = pi16 ? n32 : n71793;
  assign n71795 = pi15 ? n71783 : n71794;
  assign n71796 = pi14 ? n71773 : n71795;
  assign n71797 = pi23 ? n37273 : n60408;
  assign n71798 = pi22 ? n32 : n71797;
  assign n71799 = pi22 ? n46172 : n66956;
  assign n71800 = pi21 ? n71798 : n71799;
  assign n71801 = pi20 ? n32 : n71800;
  assign n71802 = pi21 ? n51564 : n7048;
  assign n71803 = pi20 ? n71802 : n32;
  assign n71804 = pi19 ? n71801 : n71803;
  assign n71805 = pi18 ? n32 : n71804;
  assign n71806 = pi17 ? n32 : n71805;
  assign n71807 = pi16 ? n32 : n71806;
  assign n71808 = pi22 ? n32 : n52391;
  assign n71809 = pi23 ? n55580 : n36659;
  assign n71810 = pi22 ? n52395 : n71809;
  assign n71811 = pi21 ? n71808 : n71810;
  assign n71812 = pi20 ? n32 : n71811;
  assign n71813 = pi21 ? n51564 : n882;
  assign n71814 = pi20 ? n71813 : n32;
  assign n71815 = pi19 ? n71812 : n71814;
  assign n71816 = pi18 ? n32 : n71815;
  assign n71817 = pi17 ? n32 : n71816;
  assign n71818 = pi16 ? n32 : n71817;
  assign n71819 = pi15 ? n71807 : n71818;
  assign n71820 = pi21 ? n39394 : n71425;
  assign n71821 = pi20 ? n32 : n71820;
  assign n71822 = pi19 ? n71821 : n71429;
  assign n71823 = pi18 ? n32 : n71822;
  assign n71824 = pi17 ? n32 : n71823;
  assign n71825 = pi16 ? n32 : n71824;
  assign n71826 = pi21 ? n38375 : n54617;
  assign n71827 = pi20 ? n32 : n71826;
  assign n71828 = pi21 ? n70969 : n32;
  assign n71829 = pi20 ? n71828 : n32;
  assign n71830 = pi19 ? n71827 : n71829;
  assign n71831 = pi18 ? n32 : n71830;
  assign n71832 = pi17 ? n32 : n71831;
  assign n71833 = pi16 ? n32 : n71832;
  assign n71834 = pi15 ? n71825 : n71833;
  assign n71835 = pi14 ? n71819 : n71834;
  assign n71836 = pi13 ? n71796 : n71835;
  assign n71837 = pi23 ? n36830 : n20563;
  assign n71838 = pi22 ? n32 : n71837;
  assign n71839 = pi22 ? n47380 : n36798;
  assign n71840 = pi21 ? n71838 : n71839;
  assign n71841 = pi20 ? n32 : n71840;
  assign n71842 = pi19 ? n71841 : n62367;
  assign n71843 = pi18 ? n32 : n71842;
  assign n71844 = pi17 ? n32 : n71843;
  assign n71845 = pi16 ? n32 : n71844;
  assign n71846 = pi21 ? n46772 : n53551;
  assign n71847 = pi20 ? n32 : n71846;
  assign n71848 = pi22 ? n61484 : n56665;
  assign n71849 = pi21 ? n71848 : n32;
  assign n71850 = pi20 ? n71849 : n32;
  assign n71851 = pi19 ? n71847 : n71850;
  assign n71852 = pi18 ? n32 : n71851;
  assign n71853 = pi17 ? n32 : n71852;
  assign n71854 = pi16 ? n32 : n71853;
  assign n71855 = pi15 ? n71845 : n71854;
  assign n71856 = pi22 ? n62510 : n63717;
  assign n71857 = pi21 ? n46772 : n71856;
  assign n71858 = pi20 ? n32 : n71857;
  assign n71859 = pi19 ? n71858 : n67389;
  assign n71860 = pi18 ? n32 : n71859;
  assign n71861 = pi17 ? n32 : n71860;
  assign n71862 = pi16 ? n32 : n71861;
  assign n71863 = pi22 ? n62510 : n70641;
  assign n71864 = pi21 ? n55516 : n71863;
  assign n71865 = pi20 ? n32 : n71864;
  assign n71866 = pi20 ? n57459 : n32;
  assign n71867 = pi19 ? n71865 : n71866;
  assign n71868 = pi18 ? n32 : n71867;
  assign n71869 = pi17 ? n32 : n71868;
  assign n71870 = pi16 ? n32 : n71869;
  assign n71871 = pi15 ? n71862 : n71870;
  assign n71872 = pi14 ? n71855 : n71871;
  assign n71873 = pi22 ? n64678 : n14626;
  assign n71874 = pi21 ? n46758 : n71873;
  assign n71875 = pi20 ? n32 : n71874;
  assign n71876 = pi19 ? n71875 : n70675;
  assign n71877 = pi18 ? n32 : n71876;
  assign n71878 = pi17 ? n32 : n71877;
  assign n71879 = pi16 ? n32 : n71878;
  assign n71880 = pi23 ? n60075 : n51564;
  assign n71881 = pi22 ? n51564 : n71880;
  assign n71882 = pi21 ? n45635 : n71881;
  assign n71883 = pi20 ? n32 : n71882;
  assign n71884 = pi19 ? n71883 : n37641;
  assign n71885 = pi18 ? n32 : n71884;
  assign n71886 = pi17 ? n32 : n71885;
  assign n71887 = pi16 ? n32 : n71886;
  assign n71888 = pi15 ? n71879 : n71887;
  assign n71889 = pi22 ? n13481 : n69371;
  assign n71890 = pi21 ? n45653 : n71889;
  assign n71891 = pi20 ? n32 : n71890;
  assign n71892 = pi19 ? n71891 : n37641;
  assign n71893 = pi18 ? n32 : n71892;
  assign n71894 = pi17 ? n32 : n71893;
  assign n71895 = pi16 ? n32 : n71894;
  assign n71896 = pi24 ? n14626 : n13481;
  assign n71897 = pi23 ? n71896 : n13481;
  assign n71898 = pi22 ? n51564 : n71897;
  assign n71899 = pi21 ? n70313 : n71898;
  assign n71900 = pi20 ? n32 : n71899;
  assign n71901 = pi19 ? n71900 : n32;
  assign n71902 = pi18 ? n32 : n71901;
  assign n71903 = pi17 ? n32 : n71902;
  assign n71904 = pi16 ? n32 : n71903;
  assign n71905 = pi15 ? n71895 : n71904;
  assign n71906 = pi14 ? n71888 : n71905;
  assign n71907 = pi13 ? n71872 : n71906;
  assign n71908 = pi12 ? n71836 : n71907;
  assign n71909 = pi23 ? n69724 : n32;
  assign n71910 = pi22 ? n13481 : n71909;
  assign n71911 = pi21 ? n46276 : n71910;
  assign n71912 = pi20 ? n32 : n71911;
  assign n71913 = pi19 ? n71912 : n32;
  assign n71914 = pi18 ? n32 : n71913;
  assign n71915 = pi17 ? n32 : n71914;
  assign n71916 = pi16 ? n32 : n71915;
  assign n71917 = pi21 ? n32 : n56129;
  assign n71918 = pi20 ? n32 : n71917;
  assign n71919 = pi19 ? n71918 : n32;
  assign n71920 = pi18 ? n32 : n71919;
  assign n71921 = pi17 ? n32 : n71920;
  assign n71922 = pi16 ? n32 : n71921;
  assign n71923 = pi15 ? n71916 : n71922;
  assign n71924 = pi23 ? n69400 : n13481;
  assign n71925 = pi22 ? n71924 : n14363;
  assign n71926 = pi21 ? n32 : n71925;
  assign n71927 = pi20 ? n32 : n71926;
  assign n71928 = pi19 ? n71927 : n32;
  assign n71929 = pi18 ? n32 : n71928;
  assign n71930 = pi17 ? n32 : n71929;
  assign n71931 = pi16 ? n32 : n71930;
  assign n71932 = pi15 ? n71931 : n32;
  assign n71933 = pi14 ? n71923 : n71932;
  assign n71934 = pi13 ? n71933 : n32;
  assign n71935 = pi12 ? n71934 : n32;
  assign n71936 = pi11 ? n71908 : n71935;
  assign n71937 = pi10 ? n71754 : n71936;
  assign n71938 = pi09 ? n71593 : n71937;
  assign n71939 = pi08 ? n71579 : n71938;
  assign n71940 = pi07 ? n71167 : n71939;
  assign n71941 = pi15 ? n71588 : n71597;
  assign n71942 = pi14 ? n71941 : n71601;
  assign n71943 = pi19 ? n36868 : n62954;
  assign n71944 = pi18 ? n32 : n71943;
  assign n71945 = pi17 ? n32 : n71944;
  assign n71946 = pi16 ? n32 : n71945;
  assign n71947 = pi14 ? n71185 : n71946;
  assign n71948 = pi13 ? n71942 : n71947;
  assign n71949 = pi19 ? n37956 : n67606;
  assign n71950 = pi18 ? n32 : n71949;
  assign n71951 = pi17 ? n32 : n71950;
  assign n71952 = pi16 ? n32 : n71951;
  assign n71953 = pi20 ? n40791 : n61008;
  assign n71954 = pi19 ? n37956 : n71953;
  assign n71955 = pi18 ? n32 : n71954;
  assign n71956 = pi17 ? n32 : n71955;
  assign n71957 = pi16 ? n32 : n71956;
  assign n71958 = pi15 ? n71952 : n71957;
  assign n71959 = pi19 ? n37956 : n62954;
  assign n71960 = pi18 ? n32 : n71959;
  assign n71961 = pi17 ? n32 : n71960;
  assign n71962 = pi16 ? n32 : n71961;
  assign n71963 = pi14 ? n71958 : n71962;
  assign n71964 = pi19 ? n38998 : n59306;
  assign n71965 = pi18 ? n32 : n71964;
  assign n71966 = pi17 ? n32 : n71965;
  assign n71967 = pi16 ? n32 : n71966;
  assign n71968 = pi22 ? n685 : n63009;
  assign n71969 = pi21 ? n61081 : n71968;
  assign n71970 = pi20 ? n20563 : n71969;
  assign n71971 = pi19 ? n38998 : n71970;
  assign n71972 = pi18 ? n32 : n71971;
  assign n71973 = pi17 ? n32 : n71972;
  assign n71974 = pi16 ? n32 : n71973;
  assign n71975 = pi15 ? n71967 : n71974;
  assign n71976 = pi20 ? n47158 : n69484;
  assign n71977 = pi19 ? n38998 : n71976;
  assign n71978 = pi18 ? n32 : n71977;
  assign n71979 = pi17 ? n32 : n71978;
  assign n71980 = pi16 ? n32 : n71979;
  assign n71981 = pi24 ? n36659 : n316;
  assign n71982 = pi23 ? n71981 : n316;
  assign n71983 = pi22 ? n71982 : n316;
  assign n71984 = pi21 ? n71983 : n3523;
  assign n71985 = pi20 ? n40791 : n71984;
  assign n71986 = pi19 ? n38998 : n71985;
  assign n71987 = pi18 ? n32 : n71986;
  assign n71988 = pi17 ? n32 : n71987;
  assign n71989 = pi16 ? n32 : n71988;
  assign n71990 = pi15 ? n71980 : n71989;
  assign n71991 = pi14 ? n71975 : n71990;
  assign n71992 = pi13 ? n71963 : n71991;
  assign n71993 = pi12 ? n71948 : n71992;
  assign n71994 = pi22 ? n71982 : n13481;
  assign n71995 = pi21 ? n71994 : n55560;
  assign n71996 = pi20 ? n59593 : n71995;
  assign n71997 = pi19 ? n38998 : n71996;
  assign n71998 = pi18 ? n32 : n71997;
  assign n71999 = pi17 ? n32 : n71998;
  assign n72000 = pi16 ? n32 : n71999;
  assign n72001 = pi22 ? n65074 : n14626;
  assign n72002 = pi21 ? n72001 : n2637;
  assign n72003 = pi20 ? n53326 : n72002;
  assign n72004 = pi19 ? n38998 : n72003;
  assign n72005 = pi18 ? n32 : n72004;
  assign n72006 = pi17 ? n32 : n72005;
  assign n72007 = pi16 ? n32 : n72006;
  assign n72008 = pi15 ? n72000 : n72007;
  assign n72009 = pi23 ? n65974 : n685;
  assign n72010 = pi22 ? n72009 : n685;
  assign n72011 = pi21 ? n72010 : n2637;
  assign n72012 = pi20 ? n55475 : n72011;
  assign n72013 = pi19 ? n38998 : n72012;
  assign n72014 = pi18 ? n32 : n72013;
  assign n72015 = pi17 ? n32 : n72014;
  assign n72016 = pi16 ? n32 : n72015;
  assign n72017 = pi20 ? n68577 : n59367;
  assign n72018 = pi19 ? n38998 : n72017;
  assign n72019 = pi18 ? n32 : n72018;
  assign n72020 = pi17 ? n32 : n72019;
  assign n72021 = pi16 ? n32 : n72020;
  assign n72022 = pi15 ? n72016 : n72021;
  assign n72023 = pi14 ? n72008 : n72022;
  assign n72024 = pi21 ? n67811 : n51270;
  assign n72025 = pi20 ? n72024 : n70441;
  assign n72026 = pi19 ? n38998 : n72025;
  assign n72027 = pi18 ? n32 : n72026;
  assign n72028 = pi17 ? n32 : n72027;
  assign n72029 = pi16 ? n32 : n72028;
  assign n72030 = pi21 ? n32 : n40908;
  assign n72031 = pi20 ? n32 : n72030;
  assign n72032 = pi21 ? n33792 : n61446;
  assign n72033 = pi20 ? n72032 : n59388;
  assign n72034 = pi19 ? n72031 : n72033;
  assign n72035 = pi18 ? n32 : n72034;
  assign n72036 = pi17 ? n32 : n72035;
  assign n72037 = pi16 ? n32 : n72036;
  assign n72038 = pi15 ? n72029 : n72037;
  assign n72039 = pi21 ? n33792 : n59524;
  assign n72040 = pi21 ? n66824 : n32;
  assign n72041 = pi20 ? n72039 : n72040;
  assign n72042 = pi19 ? n72031 : n72041;
  assign n72043 = pi18 ? n32 : n72042;
  assign n72044 = pi17 ? n32 : n72043;
  assign n72045 = pi16 ? n32 : n72044;
  assign n72046 = pi21 ? n32 : n40950;
  assign n72047 = pi20 ? n32 : n72046;
  assign n72048 = pi22 ? n33792 : n40386;
  assign n72049 = pi21 ? n72048 : n71260;
  assign n72050 = pi22 ? n51564 : n59395;
  assign n72051 = pi21 ? n72050 : n32;
  assign n72052 = pi20 ? n72049 : n72051;
  assign n72053 = pi19 ? n72047 : n72052;
  assign n72054 = pi18 ? n32 : n72053;
  assign n72055 = pi17 ? n32 : n72054;
  assign n72056 = pi16 ? n32 : n72055;
  assign n72057 = pi15 ? n72045 : n72056;
  assign n72058 = pi14 ? n72038 : n72057;
  assign n72059 = pi13 ? n72023 : n72058;
  assign n72060 = pi21 ? n20563 : n53471;
  assign n72061 = pi22 ? n13481 : n396;
  assign n72062 = pi21 ? n72061 : n32;
  assign n72063 = pi20 ? n72060 : n72062;
  assign n72064 = pi19 ? n37321 : n72063;
  assign n72065 = pi18 ? n32 : n72064;
  assign n72066 = pi17 ? n32 : n72065;
  assign n72067 = pi16 ? n32 : n72066;
  assign n72068 = pi20 ? n32 : n66953;
  assign n72069 = pi21 ? n30868 : n64961;
  assign n72070 = pi20 ? n72069 : n72062;
  assign n72071 = pi19 ? n72068 : n72070;
  assign n72072 = pi18 ? n32 : n72071;
  assign n72073 = pi17 ? n32 : n72072;
  assign n72074 = pi16 ? n32 : n72073;
  assign n72075 = pi15 ? n72067 : n72074;
  assign n72076 = pi22 ? n58710 : n685;
  assign n72077 = pi21 ? n33792 : n72076;
  assign n72078 = pi20 ? n72077 : n59649;
  assign n72079 = pi19 ? n72068 : n72078;
  assign n72080 = pi18 ? n32 : n72079;
  assign n72081 = pi17 ? n32 : n72080;
  assign n72082 = pi16 ? n32 : n72081;
  assign n72083 = pi22 ? n37173 : n36659;
  assign n72084 = pi21 ? n32 : n72083;
  assign n72085 = pi20 ? n32 : n72084;
  assign n72086 = pi22 ? n63195 : n51564;
  assign n72087 = pi21 ? n36659 : n72086;
  assign n72088 = pi20 ? n72087 : n65434;
  assign n72089 = pi19 ? n72085 : n72088;
  assign n72090 = pi18 ? n32 : n72089;
  assign n72091 = pi17 ? n32 : n72090;
  assign n72092 = pi16 ? n32 : n72091;
  assign n72093 = pi15 ? n72082 : n72092;
  assign n72094 = pi14 ? n72075 : n72093;
  assign n72095 = pi21 ? n32 : n54446;
  assign n72096 = pi20 ? n32 : n72095;
  assign n72097 = pi21 ? n36659 : n59774;
  assign n72098 = pi20 ? n72097 : n51568;
  assign n72099 = pi19 ? n72096 : n72098;
  assign n72100 = pi18 ? n32 : n72099;
  assign n72101 = pi17 ? n32 : n72100;
  assign n72102 = pi16 ? n32 : n72101;
  assign n72103 = pi21 ? n32 : n51762;
  assign n72104 = pi20 ? n32 : n72103;
  assign n72105 = pi22 ? n36798 : n62880;
  assign n72106 = pi21 ? n36659 : n72105;
  assign n72107 = pi20 ? n72106 : n10011;
  assign n72108 = pi19 ? n72104 : n72107;
  assign n72109 = pi18 ? n32 : n72108;
  assign n72110 = pi17 ? n32 : n72109;
  assign n72111 = pi16 ? n32 : n72110;
  assign n72112 = pi15 ? n72102 : n72111;
  assign n72113 = pi21 ? n32 : n40986;
  assign n72114 = pi20 ? n32 : n72113;
  assign n72115 = pi21 ? n47360 : n63771;
  assign n72116 = pi20 ? n72115 : n57716;
  assign n72117 = pi19 ? n72114 : n72116;
  assign n72118 = pi18 ? n32 : n72117;
  assign n72119 = pi17 ? n32 : n72118;
  assign n72120 = pi16 ? n32 : n72119;
  assign n72121 = pi21 ? n32 : n51270;
  assign n72122 = pi20 ? n32 : n72121;
  assign n72123 = pi21 ? n36781 : n61376;
  assign n72124 = pi20 ? n72123 : n32;
  assign n72125 = pi19 ? n72122 : n72124;
  assign n72126 = pi18 ? n32 : n72125;
  assign n72127 = pi17 ? n32 : n72126;
  assign n72128 = pi16 ? n32 : n72127;
  assign n72129 = pi15 ? n72120 : n72128;
  assign n72130 = pi14 ? n72112 : n72129;
  assign n72131 = pi13 ? n72094 : n72130;
  assign n72132 = pi12 ? n72059 : n72131;
  assign n72133 = pi11 ? n71993 : n72132;
  assign n72134 = pi21 ? n32 : n68713;
  assign n72135 = pi20 ? n32 : n72134;
  assign n72136 = pi21 ? n37878 : n70969;
  assign n72137 = pi20 ? n72136 : n32;
  assign n72138 = pi19 ? n72135 : n72137;
  assign n72139 = pi18 ? n32 : n72138;
  assign n72140 = pi17 ? n32 : n72139;
  assign n72141 = pi16 ? n32 : n72140;
  assign n72142 = pi21 ? n32 : n71309;
  assign n72143 = pi20 ? n32 : n72142;
  assign n72144 = pi21 ? n54617 : n71766;
  assign n72145 = pi20 ? n72144 : n32;
  assign n72146 = pi19 ? n72143 : n72145;
  assign n72147 = pi18 ? n32 : n72146;
  assign n72148 = pi17 ? n32 : n72147;
  assign n72149 = pi16 ? n32 : n72148;
  assign n72150 = pi15 ? n72141 : n72149;
  assign n72151 = pi22 ? n42109 : n36659;
  assign n72152 = pi21 ? n32 : n72151;
  assign n72153 = pi20 ? n32 : n72152;
  assign n72154 = pi21 ? n51564 : n58470;
  assign n72155 = pi20 ? n72154 : n32;
  assign n72156 = pi19 ? n72153 : n72155;
  assign n72157 = pi18 ? n32 : n72156;
  assign n72158 = pi17 ? n32 : n72157;
  assign n72159 = pi16 ? n32 : n72158;
  assign n72160 = pi22 ? n58710 : n36781;
  assign n72161 = pi21 ? n32 : n72160;
  assign n72162 = pi20 ? n32 : n72161;
  assign n72163 = pi21 ? n47397 : n2320;
  assign n72164 = pi20 ? n72163 : n32;
  assign n72165 = pi19 ? n72162 : n72164;
  assign n72166 = pi18 ? n32 : n72165;
  assign n72167 = pi17 ? n32 : n72166;
  assign n72168 = pi16 ? n32 : n72167;
  assign n72169 = pi15 ? n72159 : n72168;
  assign n72170 = pi14 ? n72150 : n72169;
  assign n72171 = pi22 ? n42106 : n68342;
  assign n72172 = pi21 ? n32 : n72171;
  assign n72173 = pi20 ? n32 : n72172;
  assign n72174 = pi20 ? n63405 : n32;
  assign n72175 = pi19 ? n72173 : n72174;
  assign n72176 = pi18 ? n32 : n72175;
  assign n72177 = pi17 ? n32 : n72176;
  assign n72178 = pi16 ? n32 : n72177;
  assign n72179 = pi23 ? n55580 : n14626;
  assign n72180 = pi22 ? n33792 : n72179;
  assign n72181 = pi21 ? n32 : n72180;
  assign n72182 = pi20 ? n32 : n72181;
  assign n72183 = pi21 ? n51564 : n19697;
  assign n72184 = pi20 ? n72183 : n32;
  assign n72185 = pi19 ? n72182 : n72184;
  assign n72186 = pi18 ? n32 : n72185;
  assign n72187 = pi17 ? n32 : n72186;
  assign n72188 = pi16 ? n32 : n72187;
  assign n72189 = pi15 ? n72178 : n72188;
  assign n72190 = pi22 ? n58736 : n72179;
  assign n72191 = pi21 ? n37332 : n72190;
  assign n72192 = pi20 ? n32 : n72191;
  assign n72193 = pi21 ? n63779 : n37639;
  assign n72194 = pi20 ? n72193 : n32;
  assign n72195 = pi19 ? n72192 : n72194;
  assign n72196 = pi18 ? n32 : n72195;
  assign n72197 = pi17 ? n32 : n72196;
  assign n72198 = pi16 ? n32 : n72197;
  assign n72199 = pi21 ? n37332 : n62846;
  assign n72200 = pi20 ? n32 : n72199;
  assign n72201 = pi22 ? n13481 : n59672;
  assign n72202 = pi21 ? n72201 : n32;
  assign n72203 = pi20 ? n72202 : n32;
  assign n72204 = pi19 ? n72200 : n72203;
  assign n72205 = pi18 ? n32 : n72204;
  assign n72206 = pi17 ? n32 : n72205;
  assign n72207 = pi16 ? n32 : n72206;
  assign n72208 = pi15 ? n72198 : n72207;
  assign n72209 = pi14 ? n72189 : n72208;
  assign n72210 = pi13 ? n72170 : n72209;
  assign n72211 = pi23 ? n64110 : n36798;
  assign n72212 = pi22 ? n37288 : n72211;
  assign n72213 = pi21 ? n45653 : n72212;
  assign n72214 = pi20 ? n32 : n72213;
  assign n72215 = pi20 ? n67728 : n32;
  assign n72216 = pi19 ? n72214 : n72215;
  assign n72217 = pi18 ? n32 : n72216;
  assign n72218 = pi17 ? n32 : n72217;
  assign n72219 = pi16 ? n32 : n72218;
  assign n72220 = pi23 ? n56620 : n13481;
  assign n72221 = pi22 ? n56712 : n72220;
  assign n72222 = pi21 ? n45653 : n72221;
  assign n72223 = pi20 ? n32 : n72222;
  assign n72224 = pi19 ? n72223 : n72215;
  assign n72225 = pi18 ? n32 : n72224;
  assign n72226 = pi17 ? n32 : n72225;
  assign n72227 = pi16 ? n32 : n72226;
  assign n72228 = pi15 ? n72219 : n72227;
  assign n72229 = pi23 ? n57517 : n14626;
  assign n72230 = pi22 ? n36798 : n72229;
  assign n72231 = pi21 ? n32 : n72230;
  assign n72232 = pi20 ? n32 : n72231;
  assign n72233 = pi19 ? n72232 : n67389;
  assign n72234 = pi18 ? n32 : n72233;
  assign n72235 = pi17 ? n32 : n72234;
  assign n72236 = pi16 ? n32 : n72235;
  assign n72237 = pi22 ? n36831 : n62411;
  assign n72238 = pi21 ? n32 : n72237;
  assign n72239 = pi20 ? n32 : n72238;
  assign n72240 = pi19 ? n72239 : n54566;
  assign n72241 = pi18 ? n32 : n72240;
  assign n72242 = pi17 ? n32 : n72241;
  assign n72243 = pi16 ? n32 : n72242;
  assign n72244 = pi15 ? n72236 : n72243;
  assign n72245 = pi14 ? n72228 : n72244;
  assign n72246 = pi23 ? n71143 : n43198;
  assign n72247 = pi22 ? n72246 : n13481;
  assign n72248 = pi21 ? n32 : n72247;
  assign n72249 = pi20 ? n32 : n72248;
  assign n72250 = pi19 ? n72249 : n37641;
  assign n72251 = pi18 ? n32 : n72250;
  assign n72252 = pi17 ? n32 : n72251;
  assign n72253 = pi16 ? n32 : n72252;
  assign n72254 = pi22 ? n46789 : n13481;
  assign n72255 = pi21 ? n32 : n72254;
  assign n72256 = pi20 ? n32 : n72255;
  assign n72257 = pi19 ? n72256 : n37641;
  assign n72258 = pi18 ? n32 : n72257;
  assign n72259 = pi17 ? n32 : n72258;
  assign n72260 = pi16 ? n32 : n72259;
  assign n72261 = pi15 ? n72253 : n72260;
  assign n72262 = pi23 ? n69400 : n14626;
  assign n72263 = pi22 ? n72262 : n58452;
  assign n72264 = pi21 ? n32 : n72263;
  assign n72265 = pi20 ? n32 : n72264;
  assign n72266 = pi19 ? n72265 : n32;
  assign n72267 = pi18 ? n32 : n72266;
  assign n72268 = pi17 ? n32 : n72267;
  assign n72269 = pi16 ? n32 : n72268;
  assign n72270 = pi23 ? n63431 : n14626;
  assign n72271 = pi23 ? n70599 : n32;
  assign n72272 = pi22 ? n72270 : n72271;
  assign n72273 = pi21 ? n32 : n72272;
  assign n72274 = pi20 ? n32 : n72273;
  assign n72275 = pi19 ? n72274 : n32;
  assign n72276 = pi18 ? n32 : n72275;
  assign n72277 = pi17 ? n32 : n72276;
  assign n72278 = pi16 ? n32 : n72277;
  assign n72279 = pi15 ? n72269 : n72278;
  assign n72280 = pi14 ? n72261 : n72279;
  assign n72281 = pi13 ? n72245 : n72280;
  assign n72282 = pi12 ? n72210 : n72281;
  assign n72283 = pi22 ? n70744 : n21502;
  assign n72284 = pi21 ? n32 : n72283;
  assign n72285 = pi20 ? n32 : n72284;
  assign n72286 = pi19 ? n72285 : n32;
  assign n72287 = pi18 ? n32 : n72286;
  assign n72288 = pi17 ? n32 : n72287;
  assign n72289 = pi16 ? n32 : n72288;
  assign n72290 = pi22 ? n69890 : n14363;
  assign n72291 = pi21 ? n32 : n72290;
  assign n72292 = pi20 ? n32 : n72291;
  assign n72293 = pi19 ? n72292 : n32;
  assign n72294 = pi18 ? n32 : n72293;
  assign n72295 = pi17 ? n32 : n72294;
  assign n72296 = pi16 ? n32 : n72295;
  assign n72297 = pi15 ? n72289 : n72296;
  assign n72298 = pi15 ? n72296 : n32;
  assign n72299 = pi14 ? n72297 : n72298;
  assign n72300 = pi13 ? n72299 : n32;
  assign n72301 = pi12 ? n72300 : n32;
  assign n72302 = pi11 ? n72282 : n72301;
  assign n72303 = pi10 ? n72133 : n72302;
  assign n72304 = pi09 ? n71593 : n72303;
  assign n72305 = pi19 ? n32 : n70348;
  assign n72306 = pi18 ? n32 : n72305;
  assign n72307 = pi17 ? n32 : n72306;
  assign n72308 = pi16 ? n32 : n72307;
  assign n72309 = pi15 ? n32 : n72308;
  assign n72310 = pi19 ? n32 : n70354;
  assign n72311 = pi18 ? n32 : n72310;
  assign n72312 = pi17 ? n32 : n72311;
  assign n72313 = pi16 ? n32 : n72312;
  assign n72314 = pi14 ? n72309 : n72313;
  assign n72315 = pi13 ? n32 : n72314;
  assign n72316 = pi12 ? n32 : n72315;
  assign n72317 = pi11 ? n32 : n72316;
  assign n72318 = pi10 ? n32 : n72317;
  assign n72319 = pi19 ? n37927 : n70354;
  assign n72320 = pi18 ? n32 : n72319;
  assign n72321 = pi17 ? n32 : n72320;
  assign n72322 = pi16 ? n32 : n72321;
  assign n72323 = pi19 ? n38982 : n62975;
  assign n72324 = pi18 ? n32 : n72323;
  assign n72325 = pi17 ? n32 : n72324;
  assign n72326 = pi16 ? n32 : n72325;
  assign n72327 = pi15 ? n72322 : n72326;
  assign n72328 = pi14 ? n72327 : n71597;
  assign n72329 = pi19 ? n40055 : n62954;
  assign n72330 = pi18 ? n32 : n72329;
  assign n72331 = pi17 ? n32 : n72330;
  assign n72332 = pi16 ? n32 : n72331;
  assign n72333 = pi14 ? n71597 : n72332;
  assign n72334 = pi13 ? n72328 : n72333;
  assign n72335 = pi19 ? n37934 : n67606;
  assign n72336 = pi18 ? n32 : n72335;
  assign n72337 = pi17 ? n32 : n72336;
  assign n72338 = pi16 ? n32 : n72337;
  assign n72339 = pi19 ? n37934 : n71953;
  assign n72340 = pi18 ? n32 : n72339;
  assign n72341 = pi17 ? n32 : n72340;
  assign n72342 = pi16 ? n32 : n72341;
  assign n72343 = pi15 ? n72338 : n72342;
  assign n72344 = pi19 ? n37934 : n62954;
  assign n72345 = pi18 ? n32 : n72344;
  assign n72346 = pi17 ? n32 : n72345;
  assign n72347 = pi16 ? n32 : n72346;
  assign n72348 = pi14 ? n72343 : n72347;
  assign n72349 = pi19 ? n36868 : n59306;
  assign n72350 = pi18 ? n32 : n72349;
  assign n72351 = pi17 ? n32 : n72350;
  assign n72352 = pi16 ? n32 : n72351;
  assign n72353 = pi19 ? n36868 : n58892;
  assign n72354 = pi18 ? n32 : n72353;
  assign n72355 = pi17 ? n32 : n72354;
  assign n72356 = pi16 ? n32 : n72355;
  assign n72357 = pi15 ? n72352 : n72356;
  assign n72358 = pi22 ? n68549 : n685;
  assign n72359 = pi21 ? n72358 : n696;
  assign n72360 = pi20 ? n47158 : n72359;
  assign n72361 = pi19 ? n36868 : n72360;
  assign n72362 = pi18 ? n32 : n72361;
  assign n72363 = pi17 ? n32 : n72362;
  assign n72364 = pi16 ? n32 : n72363;
  assign n72365 = pi19 ? n36868 : n71985;
  assign n72366 = pi18 ? n32 : n72365;
  assign n72367 = pi17 ? n32 : n72366;
  assign n72368 = pi16 ? n32 : n72367;
  assign n72369 = pi15 ? n72364 : n72368;
  assign n72370 = pi14 ? n72357 : n72369;
  assign n72371 = pi13 ? n72348 : n72370;
  assign n72372 = pi12 ? n72334 : n72371;
  assign n72373 = pi19 ? n37956 : n71996;
  assign n72374 = pi18 ? n32 : n72373;
  assign n72375 = pi17 ? n32 : n72374;
  assign n72376 = pi16 ? n32 : n72375;
  assign n72377 = pi19 ? n37956 : n72003;
  assign n72378 = pi18 ? n32 : n72377;
  assign n72379 = pi17 ? n32 : n72378;
  assign n72380 = pi16 ? n32 : n72379;
  assign n72381 = pi15 ? n72376 : n72380;
  assign n72382 = pi23 ? n778 : n685;
  assign n72383 = pi22 ? n72382 : n685;
  assign n72384 = pi21 ? n72383 : n2637;
  assign n72385 = pi20 ? n55475 : n72384;
  assign n72386 = pi19 ? n37956 : n72385;
  assign n72387 = pi18 ? n32 : n72386;
  assign n72388 = pi17 ? n32 : n72387;
  assign n72389 = pi16 ? n32 : n72388;
  assign n72390 = pi19 ? n37956 : n72017;
  assign n72391 = pi18 ? n32 : n72390;
  assign n72392 = pi17 ? n32 : n72391;
  assign n72393 = pi16 ? n32 : n72392;
  assign n72394 = pi15 ? n72389 : n72393;
  assign n72395 = pi14 ? n72381 : n72394;
  assign n72396 = pi19 ? n37956 : n72025;
  assign n72397 = pi18 ? n32 : n72396;
  assign n72398 = pi17 ? n32 : n72397;
  assign n72399 = pi16 ? n32 : n72398;
  assign n72400 = pi19 ? n68257 : n72033;
  assign n72401 = pi18 ? n32 : n72400;
  assign n72402 = pi17 ? n32 : n72401;
  assign n72403 = pi16 ? n32 : n72402;
  assign n72404 = pi15 ? n72399 : n72403;
  assign n72405 = pi19 ? n46189 : n72041;
  assign n72406 = pi18 ? n32 : n72405;
  assign n72407 = pi17 ? n32 : n72406;
  assign n72408 = pi16 ? n32 : n72407;
  assign n72409 = pi22 ? n45597 : n33792;
  assign n72410 = pi21 ? n32 : n72409;
  assign n72411 = pi20 ? n32 : n72410;
  assign n72412 = pi22 ? n33792 : n43571;
  assign n72413 = pi21 ? n72412 : n71260;
  assign n72414 = pi20 ? n72413 : n72051;
  assign n72415 = pi19 ? n72411 : n72414;
  assign n72416 = pi18 ? n32 : n72415;
  assign n72417 = pi17 ? n32 : n72416;
  assign n72418 = pi16 ? n32 : n72417;
  assign n72419 = pi15 ? n72408 : n72418;
  assign n72420 = pi14 ? n72404 : n72419;
  assign n72421 = pi13 ? n72395 : n72420;
  assign n72422 = pi19 ? n37956 : n72063;
  assign n72423 = pi18 ? n32 : n72422;
  assign n72424 = pi17 ? n32 : n72423;
  assign n72425 = pi16 ? n32 : n72424;
  assign n72426 = pi19 ? n46189 : n72070;
  assign n72427 = pi18 ? n32 : n72426;
  assign n72428 = pi17 ? n32 : n72427;
  assign n72429 = pi16 ? n32 : n72428;
  assign n72430 = pi15 ? n72425 : n72429;
  assign n72431 = pi20 ? n72077 : n60045;
  assign n72432 = pi19 ? n46189 : n72431;
  assign n72433 = pi18 ? n32 : n72432;
  assign n72434 = pi17 ? n32 : n72433;
  assign n72435 = pi16 ? n32 : n72434;
  assign n72436 = pi23 ? n37273 : n33792;
  assign n72437 = pi22 ? n72436 : n36659;
  assign n72438 = pi21 ? n32 : n72437;
  assign n72439 = pi20 ? n32 : n72438;
  assign n72440 = pi22 ? n55130 : n51564;
  assign n72441 = pi21 ? n36659 : n72440;
  assign n72442 = pi20 ? n72441 : n65434;
  assign n72443 = pi19 ? n72439 : n72442;
  assign n72444 = pi18 ? n32 : n72443;
  assign n72445 = pi17 ? n32 : n72444;
  assign n72446 = pi16 ? n32 : n72445;
  assign n72447 = pi15 ? n72435 : n72446;
  assign n72448 = pi14 ? n72430 : n72447;
  assign n72449 = pi20 ? n32 : n52743;
  assign n72450 = pi20 ? n72097 : n10011;
  assign n72451 = pi19 ? n72449 : n72450;
  assign n72452 = pi18 ? n32 : n72451;
  assign n72453 = pi17 ? n32 : n72452;
  assign n72454 = pi16 ? n32 : n72453;
  assign n72455 = pi22 ? n51754 : n36659;
  assign n72456 = pi21 ? n32 : n72455;
  assign n72457 = pi20 ? n32 : n72456;
  assign n72458 = pi20 ? n72106 : n32257;
  assign n72459 = pi19 ? n72457 : n72458;
  assign n72460 = pi18 ? n32 : n72459;
  assign n72461 = pi17 ? n32 : n72460;
  assign n72462 = pi16 ? n32 : n72461;
  assign n72463 = pi15 ? n72454 : n72462;
  assign n72464 = pi22 ? n30154 : n36659;
  assign n72465 = pi21 ? n32 : n72464;
  assign n72466 = pi20 ? n32 : n72465;
  assign n72467 = pi20 ? n72115 : n32;
  assign n72468 = pi19 ? n72466 : n72467;
  assign n72469 = pi18 ? n32 : n72468;
  assign n72470 = pi17 ? n32 : n72469;
  assign n72471 = pi16 ? n32 : n72470;
  assign n72472 = pi23 ? n32 : n66385;
  assign n72473 = pi22 ? n72472 : n36781;
  assign n72474 = pi21 ? n32 : n72473;
  assign n72475 = pi20 ? n32 : n72474;
  assign n72476 = pi19 ? n72475 : n72124;
  assign n72477 = pi18 ? n32 : n72476;
  assign n72478 = pi17 ? n32 : n72477;
  assign n72479 = pi16 ? n32 : n72478;
  assign n72480 = pi15 ? n72471 : n72479;
  assign n72481 = pi14 ? n72463 : n72480;
  assign n72482 = pi13 ? n72448 : n72481;
  assign n72483 = pi12 ? n72421 : n72482;
  assign n72484 = pi11 ? n72372 : n72483;
  assign n72485 = pi22 ? n45597 : n36781;
  assign n72486 = pi21 ? n32 : n72485;
  assign n72487 = pi20 ? n32 : n72486;
  assign n72488 = pi21 ? n37878 : n63786;
  assign n72489 = pi20 ? n72488 : n32;
  assign n72490 = pi19 ? n72487 : n72489;
  assign n72491 = pi18 ? n32 : n72490;
  assign n72492 = pi17 ? n32 : n72491;
  assign n72493 = pi16 ? n32 : n72492;
  assign n72494 = pi22 ? n49720 : n36659;
  assign n72495 = pi21 ? n32 : n72494;
  assign n72496 = pi20 ? n32 : n72495;
  assign n72497 = pi21 ? n54617 : n59415;
  assign n72498 = pi20 ? n72497 : n32;
  assign n72499 = pi19 ? n72496 : n72498;
  assign n72500 = pi18 ? n32 : n72499;
  assign n72501 = pi17 ? n32 : n72500;
  assign n72502 = pi16 ? n32 : n72501;
  assign n72503 = pi15 ? n72493 : n72502;
  assign n72504 = pi21 ? n51564 : n60421;
  assign n72505 = pi20 ? n72504 : n32;
  assign n72506 = pi19 ? n72496 : n72505;
  assign n72507 = pi18 ? n32 : n72506;
  assign n72508 = pi17 ? n32 : n72507;
  assign n72509 = pi16 ? n32 : n72508;
  assign n72510 = pi22 ? n51754 : n36781;
  assign n72511 = pi21 ? n32 : n72510;
  assign n72512 = pi20 ? n32 : n72511;
  assign n72513 = pi19 ? n72512 : n72164;
  assign n72514 = pi18 ? n32 : n72513;
  assign n72515 = pi17 ? n32 : n72514;
  assign n72516 = pi16 ? n32 : n72515;
  assign n72517 = pi15 ? n72509 : n72516;
  assign n72518 = pi14 ? n72503 : n72517;
  assign n72519 = pi22 ? n45597 : n52395;
  assign n72520 = pi21 ? n32 : n72519;
  assign n72521 = pi20 ? n32 : n72520;
  assign n72522 = pi19 ? n72521 : n72174;
  assign n72523 = pi18 ? n32 : n72522;
  assign n72524 = pi17 ? n32 : n72523;
  assign n72525 = pi16 ? n32 : n72524;
  assign n72526 = pi22 ? n49720 : n59412;
  assign n72527 = pi21 ? n32 : n72526;
  assign n72528 = pi20 ? n32 : n72527;
  assign n72529 = pi20 ? n59367 : n32;
  assign n72530 = pi19 ? n72528 : n72529;
  assign n72531 = pi18 ? n32 : n72530;
  assign n72532 = pi17 ? n32 : n72531;
  assign n72533 = pi16 ? n32 : n72532;
  assign n72534 = pi15 ? n72525 : n72533;
  assign n72535 = pi22 ? n37251 : n72179;
  assign n72536 = pi21 ? n32 : n72535;
  assign n72537 = pi20 ? n32 : n72536;
  assign n72538 = pi22 ? n14626 : n69725;
  assign n72539 = pi21 ? n72538 : n32;
  assign n72540 = pi20 ? n72539 : n32;
  assign n72541 = pi19 ? n72537 : n72540;
  assign n72542 = pi18 ? n32 : n72541;
  assign n72543 = pi17 ? n32 : n72542;
  assign n72544 = pi16 ? n32 : n72543;
  assign n72545 = pi22 ? n51754 : n62377;
  assign n72546 = pi21 ? n32 : n72545;
  assign n72547 = pi20 ? n32 : n72546;
  assign n72548 = pi22 ? n13481 : n57647;
  assign n72549 = pi21 ? n72548 : n32;
  assign n72550 = pi20 ? n72549 : n32;
  assign n72551 = pi19 ? n72547 : n72550;
  assign n72552 = pi18 ? n32 : n72551;
  assign n72553 = pi17 ? n32 : n72552;
  assign n72554 = pi16 ? n32 : n72553;
  assign n72555 = pi15 ? n72544 : n72554;
  assign n72556 = pi14 ? n72534 : n72555;
  assign n72557 = pi13 ? n72518 : n72556;
  assign n72558 = pi23 ? n59957 : n14626;
  assign n72559 = pi22 ? n37873 : n72558;
  assign n72560 = pi21 ? n32 : n72559;
  assign n72561 = pi20 ? n32 : n72560;
  assign n72562 = pi19 ? n72561 : n72215;
  assign n72563 = pi18 ? n32 : n72562;
  assign n72564 = pi17 ? n32 : n72563;
  assign n72565 = pi16 ? n32 : n72564;
  assign n72566 = pi22 ? n45135 : n62389;
  assign n72567 = pi21 ? n32 : n72566;
  assign n72568 = pi20 ? n32 : n72567;
  assign n72569 = pi19 ? n72568 : n72215;
  assign n72570 = pi18 ? n32 : n72569;
  assign n72571 = pi17 ? n32 : n72570;
  assign n72572 = pi16 ? n32 : n72571;
  assign n72573 = pi15 ? n72565 : n72572;
  assign n72574 = pi22 ? n45160 : n55641;
  assign n72575 = pi21 ? n32 : n72574;
  assign n72576 = pi20 ? n32 : n72575;
  assign n72577 = pi19 ? n72576 : n67389;
  assign n72578 = pi18 ? n32 : n72577;
  assign n72579 = pi17 ? n32 : n72578;
  assign n72580 = pi16 ? n32 : n72579;
  assign n72581 = pi22 ? n45160 : n61484;
  assign n72582 = pi21 ? n32 : n72581;
  assign n72583 = pi20 ? n32 : n72582;
  assign n72584 = pi20 ? n58504 : n32;
  assign n72585 = pi19 ? n72583 : n72584;
  assign n72586 = pi18 ? n32 : n72585;
  assign n72587 = pi17 ? n32 : n72586;
  assign n72588 = pi16 ? n32 : n72587;
  assign n72589 = pi15 ? n72580 : n72588;
  assign n72590 = pi14 ? n72573 : n72589;
  assign n72591 = pi20 ? n32 : n69403;
  assign n72592 = pi19 ? n72591 : n37641;
  assign n72593 = pi18 ? n32 : n72592;
  assign n72594 = pi17 ? n32 : n72593;
  assign n72595 = pi16 ? n32 : n72594;
  assign n72596 = pi21 ? n32 : n71120;
  assign n72597 = pi20 ? n32 : n72596;
  assign n72598 = pi19 ? n72597 : n37641;
  assign n72599 = pi18 ? n32 : n72598;
  assign n72600 = pi17 ? n32 : n72599;
  assign n72601 = pi16 ? n32 : n72600;
  assign n72602 = pi15 ? n72595 : n72601;
  assign n72603 = pi22 ? n32 : n58452;
  assign n72604 = pi21 ? n32 : n72603;
  assign n72605 = pi20 ? n32 : n72604;
  assign n72606 = pi19 ? n72605 : n32;
  assign n72607 = pi18 ? n32 : n72606;
  assign n72608 = pi17 ? n32 : n72607;
  assign n72609 = pi16 ? n32 : n72608;
  assign n72610 = pi22 ? n32 : n21502;
  assign n72611 = pi21 ? n32 : n72610;
  assign n72612 = pi20 ? n32 : n72611;
  assign n72613 = pi19 ? n72612 : n32;
  assign n72614 = pi18 ? n32 : n72613;
  assign n72615 = pi17 ? n32 : n72614;
  assign n72616 = pi16 ? n32 : n72615;
  assign n72617 = pi15 ? n72609 : n72616;
  assign n72618 = pi14 ? n72602 : n72617;
  assign n72619 = pi13 ? n72590 : n72618;
  assign n72620 = pi12 ? n72557 : n72619;
  assign n72621 = pi15 ? n72616 : n32;
  assign n72622 = pi14 ? n72621 : n32;
  assign n72623 = pi13 ? n72622 : n32;
  assign n72624 = pi12 ? n72623 : n32;
  assign n72625 = pi11 ? n72620 : n72624;
  assign n72626 = pi10 ? n72484 : n72625;
  assign n72627 = pi09 ? n72318 : n72626;
  assign n72628 = pi08 ? n72304 : n72627;
  assign n72629 = pi20 ? n31263 : n13040;
  assign n72630 = pi19 ? n32 : n72629;
  assign n72631 = pi18 ? n32 : n72630;
  assign n72632 = pi17 ? n32 : n72631;
  assign n72633 = pi16 ? n32 : n72632;
  assign n72634 = pi15 ? n32 : n72633;
  assign n72635 = pi20 ? n64535 : n1619;
  assign n72636 = pi19 ? n32 : n72635;
  assign n72637 = pi18 ? n32 : n72636;
  assign n72638 = pi17 ? n32 : n72637;
  assign n72639 = pi16 ? n32 : n72638;
  assign n72640 = pi14 ? n72634 : n72639;
  assign n72641 = pi13 ? n32 : n72640;
  assign n72642 = pi12 ? n32 : n72641;
  assign n72643 = pi11 ? n32 : n72642;
  assign n72644 = pi10 ? n32 : n72643;
  assign n72645 = pi22 ? n40342 : n20563;
  assign n72646 = pi21 ? n72645 : n30868;
  assign n72647 = pi20 ? n72646 : n1619;
  assign n72648 = pi19 ? n32 : n72647;
  assign n72649 = pi18 ? n32 : n72648;
  assign n72650 = pi17 ? n32 : n72649;
  assign n72651 = pi16 ? n32 : n72650;
  assign n72652 = pi19 ? n32 : n62975;
  assign n72653 = pi18 ? n32 : n72652;
  assign n72654 = pi17 ? n32 : n72653;
  assign n72655 = pi16 ? n32 : n72654;
  assign n72656 = pi15 ? n72651 : n72655;
  assign n72657 = pi14 ? n72656 : n72326;
  assign n72658 = pi13 ? n72657 : n72333;
  assign n72659 = pi19 ? n40055 : n67606;
  assign n72660 = pi18 ? n32 : n72659;
  assign n72661 = pi17 ? n32 : n72660;
  assign n72662 = pi16 ? n32 : n72661;
  assign n72663 = pi19 ? n40055 : n71953;
  assign n72664 = pi18 ? n32 : n72663;
  assign n72665 = pi17 ? n32 : n72664;
  assign n72666 = pi16 ? n32 : n72665;
  assign n72667 = pi15 ? n72662 : n72666;
  assign n72668 = pi22 ? n32 : n41458;
  assign n72669 = pi21 ? n32 : n72668;
  assign n72670 = pi20 ? n32 : n72669;
  assign n72671 = pi19 ? n72670 : n62954;
  assign n72672 = pi18 ? n32 : n72671;
  assign n72673 = pi17 ? n32 : n72672;
  assign n72674 = pi16 ? n32 : n72673;
  assign n72675 = pi15 ? n72332 : n72674;
  assign n72676 = pi14 ? n72667 : n72675;
  assign n72677 = pi19 ? n40055 : n59306;
  assign n72678 = pi18 ? n32 : n72677;
  assign n72679 = pi17 ? n32 : n72678;
  assign n72680 = pi16 ? n32 : n72679;
  assign n72681 = pi19 ? n40055 : n58892;
  assign n72682 = pi18 ? n32 : n72681;
  assign n72683 = pi17 ? n32 : n72682;
  assign n72684 = pi16 ? n32 : n72683;
  assign n72685 = pi15 ? n72680 : n72684;
  assign n72686 = pi21 ? n63519 : n696;
  assign n72687 = pi20 ? n47158 : n72686;
  assign n72688 = pi19 ? n40055 : n72687;
  assign n72689 = pi18 ? n32 : n72688;
  assign n72690 = pi17 ? n32 : n72689;
  assign n72691 = pi16 ? n32 : n72690;
  assign n72692 = pi22 ? n53175 : n316;
  assign n72693 = pi21 ? n72692 : n3523;
  assign n72694 = pi20 ? n40791 : n72693;
  assign n72695 = pi19 ? n40055 : n72694;
  assign n72696 = pi18 ? n32 : n72695;
  assign n72697 = pi17 ? n32 : n72696;
  assign n72698 = pi16 ? n32 : n72697;
  assign n72699 = pi15 ? n72691 : n72698;
  assign n72700 = pi14 ? n72685 : n72699;
  assign n72701 = pi13 ? n72676 : n72700;
  assign n72702 = pi12 ? n72658 : n72701;
  assign n72703 = pi20 ? n59593 : n69066;
  assign n72704 = pi19 ? n37934 : n72703;
  assign n72705 = pi18 ? n32 : n72704;
  assign n72706 = pi17 ? n32 : n72705;
  assign n72707 = pi16 ? n32 : n72706;
  assign n72708 = pi22 ? n60398 : n14626;
  assign n72709 = pi21 ? n72708 : n2637;
  assign n72710 = pi20 ? n53326 : n72709;
  assign n72711 = pi19 ? n37934 : n72710;
  assign n72712 = pi18 ? n32 : n72711;
  assign n72713 = pi17 ? n32 : n72712;
  assign n72714 = pi16 ? n32 : n72713;
  assign n72715 = pi15 ? n72707 : n72714;
  assign n72716 = pi20 ? n68778 : n72384;
  assign n72717 = pi19 ? n37934 : n72716;
  assign n72718 = pi18 ? n32 : n72717;
  assign n72719 = pi17 ? n32 : n72718;
  assign n72720 = pi16 ? n32 : n72719;
  assign n72721 = pi20 ? n32 : n64225;
  assign n72722 = pi19 ? n72721 : n72017;
  assign n72723 = pi18 ? n32 : n72722;
  assign n72724 = pi17 ? n32 : n72723;
  assign n72725 = pi16 ? n32 : n72724;
  assign n72726 = pi15 ? n72720 : n72725;
  assign n72727 = pi14 ? n72715 : n72726;
  assign n72728 = pi21 ? n32 : n71415;
  assign n72729 = pi20 ? n32 : n72728;
  assign n72730 = pi20 ? n72024 : n61537;
  assign n72731 = pi19 ? n72729 : n72730;
  assign n72732 = pi18 ? n32 : n72731;
  assign n72733 = pi17 ? n32 : n72732;
  assign n72734 = pi16 ? n32 : n72733;
  assign n72735 = pi20 ? n72032 : n58439;
  assign n72736 = pi19 ? n72729 : n72735;
  assign n72737 = pi18 ? n32 : n72736;
  assign n72738 = pi17 ? n32 : n72737;
  assign n72739 = pi16 ? n32 : n72738;
  assign n72740 = pi15 ? n72734 : n72739;
  assign n72741 = pi20 ? n72039 : n11695;
  assign n72742 = pi19 ? n37934 : n72741;
  assign n72743 = pi18 ? n32 : n72742;
  assign n72744 = pi17 ? n32 : n72743;
  assign n72745 = pi16 ? n32 : n72744;
  assign n72746 = pi21 ? n47360 : n71260;
  assign n72747 = pi21 ? n64706 : n32;
  assign n72748 = pi20 ? n72746 : n72747;
  assign n72749 = pi19 ? n37934 : n72748;
  assign n72750 = pi18 ? n32 : n72749;
  assign n72751 = pi17 ? n32 : n72750;
  assign n72752 = pi16 ? n32 : n72751;
  assign n72753 = pi15 ? n72745 : n72752;
  assign n72754 = pi14 ? n72740 : n72753;
  assign n72755 = pi13 ? n72727 : n72754;
  assign n72756 = pi20 ? n72060 : n67728;
  assign n72757 = pi19 ? n36868 : n72756;
  assign n72758 = pi18 ? n32 : n72757;
  assign n72759 = pi17 ? n32 : n72758;
  assign n72760 = pi16 ? n32 : n72759;
  assign n72761 = pi20 ? n72069 : n67728;
  assign n72762 = pi19 ? n36868 : n72761;
  assign n72763 = pi18 ? n32 : n72762;
  assign n72764 = pi17 ? n32 : n72763;
  assign n72765 = pi16 ? n32 : n72764;
  assign n72766 = pi15 ? n72760 : n72765;
  assign n72767 = pi22 ? n52395 : n685;
  assign n72768 = pi21 ? n33792 : n72767;
  assign n72769 = pi20 ? n72768 : n60045;
  assign n72770 = pi19 ? n54402 : n72769;
  assign n72771 = pi18 ? n32 : n72770;
  assign n72772 = pi17 ? n32 : n72771;
  assign n72773 = pi16 ? n32 : n72772;
  assign n72774 = pi21 ? n36659 : n63253;
  assign n72775 = pi20 ? n72774 : n59674;
  assign n72776 = pi19 ? n54402 : n72775;
  assign n72777 = pi18 ? n32 : n72776;
  assign n72778 = pi17 ? n32 : n72777;
  assign n72779 = pi16 ? n32 : n72778;
  assign n72780 = pi15 ? n72773 : n72779;
  assign n72781 = pi14 ? n72766 : n72780;
  assign n72782 = pi20 ? n32 : n58577;
  assign n72783 = pi20 ? n72097 : n57716;
  assign n72784 = pi19 ? n72782 : n72783;
  assign n72785 = pi18 ? n32 : n72784;
  assign n72786 = pi17 ? n32 : n72785;
  assign n72787 = pi16 ? n32 : n72786;
  assign n72788 = pi19 ? n54429 : n72783;
  assign n72789 = pi18 ? n32 : n72788;
  assign n72790 = pi17 ? n32 : n72789;
  assign n72791 = pi16 ? n32 : n72790;
  assign n72792 = pi15 ? n72787 : n72791;
  assign n72793 = pi20 ? n32 : n70145;
  assign n72794 = pi21 ? n39952 : n57733;
  assign n72795 = pi20 ? n72794 : n32;
  assign n72796 = pi19 ? n72793 : n72795;
  assign n72797 = pi18 ? n32 : n72796;
  assign n72798 = pi17 ? n32 : n72797;
  assign n72799 = pi16 ? n32 : n72798;
  assign n72800 = pi21 ? n32 : n71378;
  assign n72801 = pi20 ? n32 : n72800;
  assign n72802 = pi22 ? n43198 : n56186;
  assign n72803 = pi21 ? n36781 : n72802;
  assign n72804 = pi20 ? n72803 : n32;
  assign n72805 = pi19 ? n72801 : n72804;
  assign n72806 = pi18 ? n32 : n72805;
  assign n72807 = pi17 ? n32 : n72806;
  assign n72808 = pi16 ? n32 : n72807;
  assign n72809 = pi15 ? n72799 : n72808;
  assign n72810 = pi14 ? n72792 : n72809;
  assign n72811 = pi13 ? n72781 : n72810;
  assign n72812 = pi12 ? n72755 : n72811;
  assign n72813 = pi11 ? n72702 : n72812;
  assign n72814 = pi21 ? n46260 : n62837;
  assign n72815 = pi20 ? n72814 : n32;
  assign n72816 = pi19 ? n72801 : n72815;
  assign n72817 = pi18 ? n32 : n72816;
  assign n72818 = pi17 ? n32 : n72817;
  assign n72819 = pi16 ? n32 : n72818;
  assign n72820 = pi22 ? n32 : n36659;
  assign n72821 = pi21 ? n32 : n72820;
  assign n72822 = pi20 ? n32 : n72821;
  assign n72823 = pi22 ? n62803 : n21502;
  assign n72824 = pi21 ? n39972 : n72823;
  assign n72825 = pi20 ? n72824 : n32;
  assign n72826 = pi19 ? n72822 : n72825;
  assign n72827 = pi18 ? n32 : n72826;
  assign n72828 = pi17 ? n32 : n72827;
  assign n72829 = pi16 ? n32 : n72828;
  assign n72830 = pi15 ? n72819 : n72829;
  assign n72831 = pi19 ? n65265 : n72505;
  assign n72832 = pi18 ? n32 : n72831;
  assign n72833 = pi17 ? n32 : n72832;
  assign n72834 = pi16 ? n32 : n72833;
  assign n72835 = pi21 ? n55715 : n67964;
  assign n72836 = pi20 ? n72835 : n32;
  assign n72837 = pi19 ? n65265 : n72836;
  assign n72838 = pi18 ? n32 : n72837;
  assign n72839 = pi17 ? n32 : n72838;
  assign n72840 = pi16 ? n32 : n72839;
  assign n72841 = pi15 ? n72834 : n72840;
  assign n72842 = pi14 ? n72830 : n72841;
  assign n72843 = pi22 ? n32 : n37260;
  assign n72844 = pi21 ? n32 : n72843;
  assign n72845 = pi20 ? n32 : n72844;
  assign n72846 = pi22 ? n63317 : n14626;
  assign n72847 = pi21 ? n72846 : n55560;
  assign n72848 = pi20 ? n72847 : n32;
  assign n72849 = pi19 ? n72845 : n72848;
  assign n72850 = pi18 ? n32 : n72849;
  assign n72851 = pi17 ? n32 : n72850;
  assign n72852 = pi16 ? n32 : n72851;
  assign n72853 = pi23 ? n37273 : n51564;
  assign n72854 = pi22 ? n32 : n72853;
  assign n72855 = pi21 ? n32 : n72854;
  assign n72856 = pi20 ? n32 : n72855;
  assign n72857 = pi20 ? n59373 : n32;
  assign n72858 = pi19 ? n72856 : n72857;
  assign n72859 = pi18 ? n32 : n72858;
  assign n72860 = pi17 ? n32 : n72859;
  assign n72861 = pi16 ? n32 : n72860;
  assign n72862 = pi15 ? n72852 : n72861;
  assign n72863 = pi22 ? n32 : n66765;
  assign n72864 = pi21 ? n32 : n72863;
  assign n72865 = pi20 ? n32 : n72864;
  assign n72866 = pi19 ? n72865 : n59605;
  assign n72867 = pi18 ? n32 : n72866;
  assign n72868 = pi17 ? n32 : n72867;
  assign n72869 = pi16 ? n32 : n72868;
  assign n72870 = pi22 ? n32 : n60092;
  assign n72871 = pi21 ? n32 : n72870;
  assign n72872 = pi20 ? n32 : n72871;
  assign n72873 = pi19 ? n72872 : n72215;
  assign n72874 = pi18 ? n32 : n72873;
  assign n72875 = pi17 ? n32 : n72874;
  assign n72876 = pi16 ? n32 : n72875;
  assign n72877 = pi15 ? n72869 : n72876;
  assign n72878 = pi14 ? n72862 : n72877;
  assign n72879 = pi13 ? n72842 : n72878;
  assign n72880 = pi19 ? n65286 : n72215;
  assign n72881 = pi18 ? n32 : n72880;
  assign n72882 = pi17 ? n32 : n72881;
  assign n72883 = pi16 ? n32 : n72882;
  assign n72884 = pi22 ? n32 : n55622;
  assign n72885 = pi21 ? n32 : n72884;
  assign n72886 = pi20 ? n32 : n72885;
  assign n72887 = pi19 ? n72886 : n59675;
  assign n72888 = pi18 ? n32 : n72887;
  assign n72889 = pi17 ? n32 : n72888;
  assign n72890 = pi16 ? n32 : n72889;
  assign n72891 = pi15 ? n72883 : n72890;
  assign n72892 = pi23 ? n46274 : n51564;
  assign n72893 = pi22 ? n32 : n72892;
  assign n72894 = pi21 ? n32 : n72893;
  assign n72895 = pi20 ? n32 : n72894;
  assign n72896 = pi19 ? n72895 : n57717;
  assign n72897 = pi18 ? n32 : n72896;
  assign n72898 = pi17 ? n32 : n72897;
  assign n72899 = pi16 ? n32 : n72898;
  assign n72900 = pi22 ? n32 : n56186;
  assign n72901 = pi21 ? n32 : n72900;
  assign n72902 = pi20 ? n32 : n72901;
  assign n72903 = pi19 ? n72902 : n57717;
  assign n72904 = pi18 ? n32 : n72903;
  assign n72905 = pi17 ? n32 : n72904;
  assign n72906 = pi16 ? n32 : n72905;
  assign n72907 = pi15 ? n72899 : n72906;
  assign n72908 = pi14 ? n72891 : n72907;
  assign n72909 = pi23 ? n71143 : n32;
  assign n72910 = pi22 ? n32 : n72909;
  assign n72911 = pi21 ? n32 : n72910;
  assign n72912 = pi20 ? n32 : n72911;
  assign n72913 = pi19 ? n72912 : n32;
  assign n72914 = pi18 ? n32 : n72913;
  assign n72915 = pi17 ? n32 : n72914;
  assign n72916 = pi16 ? n32 : n72915;
  assign n72917 = pi23 ? n69400 : n32;
  assign n72918 = pi22 ? n32 : n72917;
  assign n72919 = pi21 ? n32 : n72918;
  assign n72920 = pi20 ? n32 : n72919;
  assign n72921 = pi19 ? n72920 : n32;
  assign n72922 = pi18 ? n32 : n72921;
  assign n72923 = pi17 ? n32 : n72922;
  assign n72924 = pi16 ? n32 : n72923;
  assign n72925 = pi15 ? n72916 : n72924;
  assign n72926 = pi14 ? n72601 : n72925;
  assign n72927 = pi13 ? n72908 : n72926;
  assign n72928 = pi12 ? n72879 : n72927;
  assign n72929 = pi15 ? n72924 : n32;
  assign n72930 = pi14 ? n72929 : n32;
  assign n72931 = pi13 ? n72930 : n32;
  assign n72932 = pi12 ? n72931 : n32;
  assign n72933 = pi11 ? n72928 : n72932;
  assign n72934 = pi10 ? n72813 : n72933;
  assign n72935 = pi09 ? n72644 : n72934;
  assign n72936 = pi21 ? n51232 : n30868;
  assign n72937 = pi20 ? n72936 : n1619;
  assign n72938 = pi19 ? n32 : n72937;
  assign n72939 = pi18 ? n32 : n72938;
  assign n72940 = pi17 ? n32 : n72939;
  assign n72941 = pi16 ? n32 : n72940;
  assign n72942 = pi20 ? n31263 : n1619;
  assign n72943 = pi19 ? n32 : n72942;
  assign n72944 = pi18 ? n32 : n72943;
  assign n72945 = pi17 ? n32 : n72944;
  assign n72946 = pi16 ? n32 : n72945;
  assign n72947 = pi15 ? n72941 : n72946;
  assign n72948 = pi14 ? n72947 : n72655;
  assign n72949 = pi19 ? n37927 : n62975;
  assign n72950 = pi18 ? n32 : n72949;
  assign n72951 = pi17 ? n32 : n72950;
  assign n72952 = pi16 ? n32 : n72951;
  assign n72953 = pi19 ? n37927 : n62954;
  assign n72954 = pi18 ? n32 : n72953;
  assign n72955 = pi17 ? n32 : n72954;
  assign n72956 = pi16 ? n32 : n72955;
  assign n72957 = pi14 ? n72952 : n72956;
  assign n72958 = pi13 ? n72948 : n72957;
  assign n72959 = pi22 ? n40386 : n37;
  assign n72960 = pi21 ? n20563 : n72959;
  assign n72961 = pi20 ? n72960 : n61008;
  assign n72962 = pi19 ? n38982 : n72961;
  assign n72963 = pi18 ? n32 : n72962;
  assign n72964 = pi17 ? n32 : n72963;
  assign n72965 = pi16 ? n32 : n72964;
  assign n72966 = pi19 ? n38982 : n71953;
  assign n72967 = pi18 ? n32 : n72966;
  assign n72968 = pi17 ? n32 : n72967;
  assign n72969 = pi16 ? n32 : n72968;
  assign n72970 = pi15 ? n72965 : n72969;
  assign n72971 = pi19 ? n38982 : n62954;
  assign n72972 = pi18 ? n32 : n72971;
  assign n72973 = pi17 ? n32 : n72972;
  assign n72974 = pi16 ? n32 : n72973;
  assign n72975 = pi14 ? n72970 : n72974;
  assign n72976 = pi20 ? n47158 : n67195;
  assign n72977 = pi19 ? n40055 : n72976;
  assign n72978 = pi18 ? n32 : n72977;
  assign n72979 = pi17 ? n32 : n72978;
  assign n72980 = pi16 ? n32 : n72979;
  assign n72981 = pi15 ? n72980 : n72698;
  assign n72982 = pi14 ? n72685 : n72981;
  assign n72983 = pi13 ? n72975 : n72982;
  assign n72984 = pi12 ? n72958 : n72983;
  assign n72985 = pi24 ? n36781 : n13481;
  assign n72986 = pi23 ? n72985 : n13481;
  assign n72987 = pi22 ? n72986 : n13481;
  assign n72988 = pi21 ? n72987 : n55560;
  assign n72989 = pi20 ? n59593 : n72988;
  assign n72990 = pi19 ? n40055 : n72989;
  assign n72991 = pi18 ? n32 : n72990;
  assign n72992 = pi17 ? n32 : n72991;
  assign n72993 = pi16 ? n32 : n72992;
  assign n72994 = pi20 ? n53326 : n71642;
  assign n72995 = pi19 ? n40055 : n72994;
  assign n72996 = pi18 ? n32 : n72995;
  assign n72997 = pi17 ? n32 : n72996;
  assign n72998 = pi16 ? n32 : n72997;
  assign n72999 = pi15 ? n72993 : n72998;
  assign n73000 = pi22 ? n66302 : n685;
  assign n73001 = pi21 ? n73000 : n2637;
  assign n73002 = pi20 ? n68778 : n73001;
  assign n73003 = pi19 ? n72670 : n73002;
  assign n73004 = pi18 ? n32 : n73003;
  assign n73005 = pi17 ? n32 : n73004;
  assign n73006 = pi16 ? n32 : n73005;
  assign n73007 = pi21 ? n40913 : n53385;
  assign n73008 = pi20 ? n73007 : n59367;
  assign n73009 = pi19 ? n51815 : n73008;
  assign n73010 = pi18 ? n32 : n73009;
  assign n73011 = pi17 ? n32 : n73010;
  assign n73012 = pi16 ? n32 : n73011;
  assign n73013 = pi15 ? n73006 : n73012;
  assign n73014 = pi14 ? n72999 : n73013;
  assign n73015 = pi20 ? n32 : n47769;
  assign n73016 = pi21 ? n72048 : n51270;
  assign n73017 = pi20 ? n73016 : n61537;
  assign n73018 = pi19 ? n73015 : n73017;
  assign n73019 = pi18 ? n32 : n73018;
  assign n73020 = pi17 ? n32 : n73019;
  assign n73021 = pi16 ? n32 : n73020;
  assign n73022 = pi21 ? n40955 : n61446;
  assign n73023 = pi20 ? n73022 : n58439;
  assign n73024 = pi19 ? n73015 : n73023;
  assign n73025 = pi18 ? n32 : n73024;
  assign n73026 = pi17 ? n32 : n73025;
  assign n73027 = pi16 ? n32 : n73026;
  assign n73028 = pi15 ? n73021 : n73027;
  assign n73029 = pi19 ? n38982 : n72741;
  assign n73030 = pi18 ? n32 : n73029;
  assign n73031 = pi17 ? n32 : n73030;
  assign n73032 = pi16 ? n32 : n73031;
  assign n73033 = pi20 ? n72413 : n72747;
  assign n73034 = pi19 ? n38982 : n73033;
  assign n73035 = pi18 ? n32 : n73034;
  assign n73036 = pi17 ? n32 : n73035;
  assign n73037 = pi16 ? n32 : n73036;
  assign n73038 = pi15 ? n73032 : n73037;
  assign n73039 = pi14 ? n73028 : n73038;
  assign n73040 = pi13 ? n73014 : n73039;
  assign n73041 = pi19 ? n40055 : n72756;
  assign n73042 = pi18 ? n32 : n73041;
  assign n73043 = pi17 ? n32 : n73042;
  assign n73044 = pi16 ? n32 : n73043;
  assign n73045 = pi19 ? n40055 : n72761;
  assign n73046 = pi18 ? n32 : n73045;
  assign n73047 = pi17 ? n32 : n73046;
  assign n73048 = pi16 ? n32 : n73047;
  assign n73049 = pi15 ? n73044 : n73048;
  assign n73050 = pi22 ? n38284 : n685;
  assign n73051 = pi21 ? n33792 : n73050;
  assign n73052 = pi20 ? n73051 : n60045;
  assign n73053 = pi19 ? n40055 : n73052;
  assign n73054 = pi18 ? n32 : n73053;
  assign n73055 = pi17 ? n32 : n73054;
  assign n73056 = pi16 ? n32 : n73055;
  assign n73057 = pi20 ? n72774 : n58504;
  assign n73058 = pi19 ? n40055 : n73057;
  assign n73059 = pi18 ? n32 : n73058;
  assign n73060 = pi17 ? n32 : n73059;
  assign n73061 = pi16 ? n32 : n73060;
  assign n73062 = pi15 ? n73056 : n73061;
  assign n73063 = pi14 ? n73049 : n73062;
  assign n73064 = pi19 ? n40055 : n72783;
  assign n73065 = pi18 ? n32 : n73064;
  assign n73066 = pi17 ? n32 : n73065;
  assign n73067 = pi16 ? n32 : n73066;
  assign n73068 = pi21 ? n32 : n50666;
  assign n73069 = pi20 ? n32 : n73068;
  assign n73070 = pi20 ? n72097 : n37640;
  assign n73071 = pi19 ? n73069 : n73070;
  assign n73072 = pi18 ? n32 : n73071;
  assign n73073 = pi17 ? n32 : n73072;
  assign n73074 = pi16 ? n32 : n73073;
  assign n73075 = pi15 ? n73067 : n73074;
  assign n73076 = pi19 ? n51815 : n72795;
  assign n73077 = pi18 ? n32 : n73076;
  assign n73078 = pi17 ? n32 : n73077;
  assign n73079 = pi16 ? n32 : n73078;
  assign n73080 = pi22 ? n32 : n71003;
  assign n73081 = pi21 ? n32 : n73080;
  assign n73082 = pi20 ? n32 : n73081;
  assign n73083 = pi19 ? n73082 : n72804;
  assign n73084 = pi18 ? n32 : n73083;
  assign n73085 = pi17 ? n32 : n73084;
  assign n73086 = pi16 ? n32 : n73085;
  assign n73087 = pi15 ? n73079 : n73086;
  assign n73088 = pi14 ? n73075 : n73087;
  assign n73089 = pi13 ? n73063 : n73088;
  assign n73090 = pi12 ? n73040 : n73089;
  assign n73091 = pi11 ? n72984 : n73090;
  assign n73092 = pi19 ? n73015 : n72815;
  assign n73093 = pi18 ? n32 : n73092;
  assign n73094 = pi17 ? n32 : n73093;
  assign n73095 = pi16 ? n32 : n73094;
  assign n73096 = pi22 ? n32 : n41097;
  assign n73097 = pi21 ? n32 : n73096;
  assign n73098 = pi20 ? n32 : n73097;
  assign n73099 = pi19 ? n73098 : n72825;
  assign n73100 = pi18 ? n32 : n73099;
  assign n73101 = pi17 ? n32 : n73100;
  assign n73102 = pi16 ? n32 : n73101;
  assign n73103 = pi15 ? n73095 : n73102;
  assign n73104 = pi22 ? n32 : n39996;
  assign n73105 = pi21 ? n32 : n73104;
  assign n73106 = pi20 ? n32 : n73105;
  assign n73107 = pi19 ? n73106 : n72505;
  assign n73108 = pi18 ? n32 : n73107;
  assign n73109 = pi17 ? n32 : n73108;
  assign n73110 = pi16 ? n32 : n73109;
  assign n73111 = pi21 ? n32 : n45211;
  assign n73112 = pi20 ? n32 : n73111;
  assign n73113 = pi19 ? n73112 : n72836;
  assign n73114 = pi18 ? n32 : n73113;
  assign n73115 = pi17 ? n32 : n73114;
  assign n73116 = pi16 ? n32 : n73115;
  assign n73117 = pi15 ? n73110 : n73116;
  assign n73118 = pi14 ? n73103 : n73117;
  assign n73119 = pi19 ? n73112 : n72848;
  assign n73120 = pi18 ? n32 : n73119;
  assign n73121 = pi17 ? n32 : n73120;
  assign n73122 = pi16 ? n32 : n73121;
  assign n73123 = pi22 ? n32 : n70744;
  assign n73124 = pi21 ? n32 : n73123;
  assign n73125 = pi20 ? n32 : n73124;
  assign n73126 = pi19 ? n73125 : n72857;
  assign n73127 = pi18 ? n32 : n73126;
  assign n73128 = pi17 ? n32 : n73127;
  assign n73129 = pi16 ? n32 : n73128;
  assign n73130 = pi15 ? n73122 : n73129;
  assign n73131 = pi20 ? n32 : n69892;
  assign n73132 = pi19 ? n73131 : n59605;
  assign n73133 = pi18 ? n32 : n73132;
  assign n73134 = pi17 ? n32 : n73133;
  assign n73135 = pi16 ? n32 : n73134;
  assign n73136 = pi23 ? n36782 : n13481;
  assign n73137 = pi22 ? n32 : n73136;
  assign n73138 = pi21 ? n32 : n73137;
  assign n73139 = pi20 ? n32 : n73138;
  assign n73140 = pi19 ? n73139 : n72215;
  assign n73141 = pi18 ? n32 : n73140;
  assign n73142 = pi17 ? n32 : n73141;
  assign n73143 = pi16 ? n32 : n73142;
  assign n73144 = pi15 ? n73135 : n73143;
  assign n73145 = pi14 ? n73130 : n73144;
  assign n73146 = pi13 ? n73118 : n73145;
  assign n73147 = pi23 ? n36830 : n71143;
  assign n73148 = pi22 ? n32 : n73147;
  assign n73149 = pi21 ? n32 : n73148;
  assign n73150 = pi20 ? n32 : n73149;
  assign n73151 = pi19 ? n73150 : n72215;
  assign n73152 = pi18 ? n32 : n73151;
  assign n73153 = pi17 ? n32 : n73152;
  assign n73154 = pi16 ? n32 : n73153;
  assign n73155 = pi19 ? n73150 : n59675;
  assign n73156 = pi18 ? n32 : n73155;
  assign n73157 = pi17 ? n32 : n73156;
  assign n73158 = pi16 ? n32 : n73157;
  assign n73159 = pi15 ? n73154 : n73158;
  assign n73160 = pi20 ? n32 : n70314;
  assign n73161 = pi19 ? n73160 : n57717;
  assign n73162 = pi18 ? n32 : n73161;
  assign n73163 = pi17 ? n32 : n73162;
  assign n73164 = pi16 ? n32 : n73163;
  assign n73165 = pi19 ? n73131 : n57717;
  assign n73166 = pi18 ? n32 : n73165;
  assign n73167 = pi17 ? n32 : n73166;
  assign n73168 = pi16 ? n32 : n73167;
  assign n73169 = pi15 ? n73164 : n73168;
  assign n73170 = pi14 ? n73159 : n73169;
  assign n73171 = pi21 ? n32 : n71566;
  assign n73172 = pi20 ? n32 : n73171;
  assign n73173 = pi19 ? n73172 : n32;
  assign n73174 = pi18 ? n32 : n73173;
  assign n73175 = pi17 ? n32 : n73174;
  assign n73176 = pi16 ? n32 : n73175;
  assign n73177 = pi15 ? n73176 : n32;
  assign n73178 = pi14 ? n73177 : n32;
  assign n73179 = pi13 ? n73170 : n73178;
  assign n73180 = pi12 ? n73146 : n73179;
  assign n73181 = pi11 ? n73180 : n32;
  assign n73182 = pi10 ? n73091 : n73181;
  assign n73183 = pi09 ? n72644 : n73182;
  assign n73184 = pi08 ? n72935 : n73183;
  assign n73185 = pi07 ? n72628 : n73184;
  assign n73186 = pi06 ? n71940 : n73185;
  assign n73187 = pi20 ? n28157 : n13040;
  assign n73188 = pi19 ? n32 : n73187;
  assign n73189 = pi18 ? n32 : n73188;
  assign n73190 = pi17 ? n32 : n73189;
  assign n73191 = pi16 ? n32 : n73190;
  assign n73192 = pi15 ? n32 : n73191;
  assign n73193 = pi20 ? n28157 : n61008;
  assign n73194 = pi19 ? n32 : n73193;
  assign n73195 = pi18 ? n32 : n73194;
  assign n73196 = pi17 ? n32 : n73195;
  assign n73197 = pi16 ? n32 : n73196;
  assign n73198 = pi20 ? n30117 : n61008;
  assign n73199 = pi19 ? n32 : n73198;
  assign n73200 = pi18 ? n32 : n73199;
  assign n73201 = pi17 ? n32 : n73200;
  assign n73202 = pi16 ? n32 : n73201;
  assign n73203 = pi15 ? n73197 : n73202;
  assign n73204 = pi14 ? n73192 : n73203;
  assign n73205 = pi13 ? n32 : n73204;
  assign n73206 = pi12 ? n32 : n73205;
  assign n73207 = pi11 ? n32 : n73206;
  assign n73208 = pi10 ? n32 : n73207;
  assign n73209 = pi20 ? n31263 : n61008;
  assign n73210 = pi19 ? n32 : n73209;
  assign n73211 = pi18 ? n32 : n73210;
  assign n73212 = pi17 ? n32 : n73211;
  assign n73213 = pi16 ? n32 : n73212;
  assign n73214 = pi15 ? n73202 : n73213;
  assign n73215 = pi14 ? n73214 : n72946;
  assign n73216 = pi20 ? n31313 : n1619;
  assign n73217 = pi19 ? n32 : n73216;
  assign n73218 = pi18 ? n32 : n73217;
  assign n73219 = pi17 ? n32 : n73218;
  assign n73220 = pi16 ? n32 : n73219;
  assign n73221 = pi13 ? n73215 : n73220;
  assign n73222 = pi14 ? n72313 : n72655;
  assign n73223 = pi19 ? n37927 : n59306;
  assign n73224 = pi18 ? n32 : n73223;
  assign n73225 = pi17 ? n32 : n73224;
  assign n73226 = pi16 ? n32 : n73225;
  assign n73227 = pi21 ? n46116 : n30868;
  assign n73228 = pi20 ? n73227 : n72686;
  assign n73229 = pi19 ? n37927 : n73228;
  assign n73230 = pi18 ? n32 : n73229;
  assign n73231 = pi17 ? n32 : n73230;
  assign n73232 = pi16 ? n32 : n73231;
  assign n73233 = pi15 ? n73226 : n73232;
  assign n73234 = pi22 ? n64420 : n51564;
  assign n73235 = pi21 ? n73234 : n57433;
  assign n73236 = pi20 ? n40791 : n73235;
  assign n73237 = pi19 ? n37927 : n73236;
  assign n73238 = pi18 ? n32 : n73237;
  assign n73239 = pi17 ? n32 : n73238;
  assign n73240 = pi16 ? n32 : n73239;
  assign n73241 = pi24 ? n30868 : n316;
  assign n73242 = pi23 ? n73241 : n316;
  assign n73243 = pi22 ? n73242 : n316;
  assign n73244 = pi21 ? n73243 : n3523;
  assign n73245 = pi20 ? n54474 : n73244;
  assign n73246 = pi19 ? n37927 : n73245;
  assign n73247 = pi18 ? n32 : n73246;
  assign n73248 = pi17 ? n32 : n73247;
  assign n73249 = pi16 ? n32 : n73248;
  assign n73250 = pi15 ? n73240 : n73249;
  assign n73251 = pi14 ? n73233 : n73250;
  assign n73252 = pi13 ? n73222 : n73251;
  assign n73253 = pi12 ? n73221 : n73252;
  assign n73254 = pi21 ? n39191 : n47360;
  assign n73255 = pi20 ? n73254 : n72988;
  assign n73256 = pi19 ? n38982 : n73255;
  assign n73257 = pi18 ? n32 : n73256;
  assign n73258 = pi17 ? n32 : n73257;
  assign n73259 = pi16 ? n32 : n73258;
  assign n73260 = pi21 ? n36489 : n47360;
  assign n73261 = pi20 ? n73260 : n72384;
  assign n73262 = pi19 ? n38982 : n73261;
  assign n73263 = pi18 ? n32 : n73262;
  assign n73264 = pi17 ? n32 : n73263;
  assign n73265 = pi16 ? n32 : n73264;
  assign n73266 = pi15 ? n73259 : n73265;
  assign n73267 = pi21 ? n52246 : n39952;
  assign n73268 = pi22 ? n66302 : n51564;
  assign n73269 = pi21 ? n73268 : n2637;
  assign n73270 = pi20 ? n73267 : n73269;
  assign n73271 = pi19 ? n38982 : n73270;
  assign n73272 = pi18 ? n32 : n73271;
  assign n73273 = pi17 ? n32 : n73272;
  assign n73274 = pi16 ? n32 : n73273;
  assign n73275 = pi21 ? n64217 : n39952;
  assign n73276 = pi23 ? n65230 : n316;
  assign n73277 = pi22 ? n73276 : n316;
  assign n73278 = pi21 ? n73277 : n928;
  assign n73279 = pi20 ? n73275 : n73278;
  assign n73280 = pi19 ? n38982 : n73279;
  assign n73281 = pi18 ? n32 : n73280;
  assign n73282 = pi17 ? n32 : n73281;
  assign n73283 = pi16 ? n32 : n73282;
  assign n73284 = pi15 ? n73274 : n73283;
  assign n73285 = pi14 ? n73266 : n73284;
  assign n73286 = pi21 ? n37768 : n61352;
  assign n73287 = pi20 ? n73286 : n61537;
  assign n73288 = pi19 ? n38982 : n73287;
  assign n73289 = pi18 ? n32 : n73288;
  assign n73290 = pi17 ? n32 : n73289;
  assign n73291 = pi16 ? n32 : n73290;
  assign n73292 = pi21 ? n37768 : n59524;
  assign n73293 = pi22 ? n685 : n66784;
  assign n73294 = pi21 ? n73293 : n32;
  assign n73295 = pi20 ? n73292 : n73294;
  assign n73296 = pi19 ? n51702 : n73295;
  assign n73297 = pi18 ? n32 : n73296;
  assign n73298 = pi17 ? n32 : n73297;
  assign n73299 = pi16 ? n32 : n73298;
  assign n73300 = pi15 ? n73291 : n73299;
  assign n73301 = pi21 ? n20563 : n61446;
  assign n73302 = pi20 ? n73301 : n70483;
  assign n73303 = pi19 ? n51702 : n73302;
  assign n73304 = pi18 ? n32 : n73303;
  assign n73305 = pi17 ? n32 : n73304;
  assign n73306 = pi16 ? n32 : n73305;
  assign n73307 = pi21 ? n20563 : n71260;
  assign n73308 = pi20 ? n73307 : n68653;
  assign n73309 = pi19 ? n51732 : n73308;
  assign n73310 = pi18 ? n32 : n73309;
  assign n73311 = pi17 ? n32 : n73310;
  assign n73312 = pi16 ? n32 : n73311;
  assign n73313 = pi15 ? n73306 : n73312;
  assign n73314 = pi14 ? n73300 : n73313;
  assign n73315 = pi13 ? n73285 : n73314;
  assign n73316 = pi20 ? n73307 : n67728;
  assign n73317 = pi19 ? n51732 : n73316;
  assign n73318 = pi18 ? n32 : n73317;
  assign n73319 = pi17 ? n32 : n73318;
  assign n73320 = pi16 ? n32 : n73319;
  assign n73321 = pi21 ? n30868 : n69292;
  assign n73322 = pi20 ? n73321 : n62857;
  assign n73323 = pi19 ? n51702 : n73322;
  assign n73324 = pi18 ? n32 : n73323;
  assign n73325 = pi17 ? n32 : n73324;
  assign n73326 = pi16 ? n32 : n73325;
  assign n73327 = pi15 ? n73320 : n73326;
  assign n73328 = pi22 ? n59412 : n51564;
  assign n73329 = pi21 ? n67811 : n73328;
  assign n73330 = pi20 ? n73329 : n3210;
  assign n73331 = pi19 ? n51732 : n73330;
  assign n73332 = pi18 ? n32 : n73331;
  assign n73333 = pi17 ? n32 : n73332;
  assign n73334 = pi16 ? n32 : n73333;
  assign n73335 = pi21 ? n47360 : n69301;
  assign n73336 = pi20 ? n73335 : n32257;
  assign n73337 = pi19 ? n51732 : n73336;
  assign n73338 = pi18 ? n32 : n73337;
  assign n73339 = pi17 ? n32 : n73338;
  assign n73340 = pi16 ? n32 : n73339;
  assign n73341 = pi15 ? n73334 : n73340;
  assign n73342 = pi14 ? n73327 : n73341;
  assign n73343 = pi21 ? n67832 : n59774;
  assign n73344 = pi20 ? n73343 : n37640;
  assign n73345 = pi19 ? n51757 : n73344;
  assign n73346 = pi18 ? n32 : n73345;
  assign n73347 = pi17 ? n32 : n73346;
  assign n73348 = pi16 ? n32 : n73347;
  assign n73349 = pi22 ? n53550 : n51564;
  assign n73350 = pi21 ? n36659 : n73349;
  assign n73351 = pi20 ? n73350 : n32;
  assign n73352 = pi19 ? n49331 : n73351;
  assign n73353 = pi18 ? n32 : n73352;
  assign n73354 = pi17 ? n32 : n73353;
  assign n73355 = pi16 ? n32 : n73354;
  assign n73356 = pi15 ? n73348 : n73355;
  assign n73357 = pi22 ? n32 : n45135;
  assign n73358 = pi21 ? n32 : n73357;
  assign n73359 = pi20 ? n32 : n73358;
  assign n73360 = pi22 ? n55622 : n13481;
  assign n73361 = pi21 ? n36781 : n73360;
  assign n73362 = pi20 ? n73361 : n32;
  assign n73363 = pi19 ? n73359 : n73362;
  assign n73364 = pi18 ? n32 : n73363;
  assign n73365 = pi17 ? n32 : n73364;
  assign n73366 = pi16 ? n32 : n73365;
  assign n73367 = pi21 ? n32 : n55516;
  assign n73368 = pi20 ? n32 : n73367;
  assign n73369 = pi21 ? n36781 : n62438;
  assign n73370 = pi20 ? n73369 : n32;
  assign n73371 = pi19 ? n73368 : n73370;
  assign n73372 = pi18 ? n32 : n73371;
  assign n73373 = pi17 ? n32 : n73372;
  assign n73374 = pi16 ? n32 : n73373;
  assign n73375 = pi15 ? n73366 : n73374;
  assign n73376 = pi14 ? n73356 : n73375;
  assign n73377 = pi13 ? n73342 : n73376;
  assign n73378 = pi12 ? n73315 : n73377;
  assign n73379 = pi11 ? n73253 : n73378;
  assign n73380 = pi21 ? n64961 : n56810;
  assign n73381 = pi20 ? n73380 : n32;
  assign n73382 = pi19 ? n73368 : n73381;
  assign n73383 = pi18 ? n32 : n73382;
  assign n73384 = pi17 ? n32 : n73383;
  assign n73385 = pi16 ? n32 : n73384;
  assign n73386 = pi21 ? n57774 : n57198;
  assign n73387 = pi20 ? n73386 : n32;
  assign n73388 = pi19 ? n48847 : n73387;
  assign n73389 = pi18 ? n32 : n73388;
  assign n73390 = pi17 ? n32 : n73389;
  assign n73391 = pi16 ? n32 : n73390;
  assign n73392 = pi15 ? n73385 : n73391;
  assign n73393 = pi21 ? n63253 : n67964;
  assign n73394 = pi20 ? n73393 : n32;
  assign n73395 = pi19 ? n46202 : n73394;
  assign n73396 = pi18 ? n32 : n73395;
  assign n73397 = pi17 ? n32 : n73396;
  assign n73398 = pi16 ? n32 : n73397;
  assign n73399 = pi22 ? n63328 : n51564;
  assign n73400 = pi21 ? n73399 : n67964;
  assign n73401 = pi20 ? n73400 : n32;
  assign n73402 = pi19 ? n46278 : n73401;
  assign n73403 = pi18 ? n32 : n73402;
  assign n73404 = pi17 ? n32 : n73403;
  assign n73405 = pi16 ? n32 : n73404;
  assign n73406 = pi15 ? n73398 : n73405;
  assign n73407 = pi14 ? n73392 : n73406;
  assign n73408 = pi21 ? n32 : n63433;
  assign n73409 = pi20 ? n32 : n73408;
  assign n73410 = pi21 ? n73399 : n32;
  assign n73411 = pi20 ? n73410 : n32;
  assign n73412 = pi19 ? n73409 : n73411;
  assign n73413 = pi18 ? n32 : n73412;
  assign n73414 = pi17 ? n32 : n73413;
  assign n73415 = pi16 ? n32 : n73414;
  assign n73416 = pi21 ? n32 : n71541;
  assign n73417 = pi20 ? n32 : n73416;
  assign n73418 = pi20 ? n62516 : n32;
  assign n73419 = pi19 ? n73417 : n73418;
  assign n73420 = pi18 ? n32 : n73419;
  assign n73421 = pi17 ? n32 : n73420;
  assign n73422 = pi16 ? n32 : n73421;
  assign n73423 = pi15 ? n73415 : n73422;
  assign n73424 = pi22 ? n61484 : n13481;
  assign n73425 = pi21 ? n73424 : n32;
  assign n73426 = pi20 ? n73425 : n32;
  assign n73427 = pi19 ? n73417 : n73426;
  assign n73428 = pi18 ? n32 : n73427;
  assign n73429 = pi17 ? n32 : n73428;
  assign n73430 = pi16 ? n32 : n73429;
  assign n73431 = pi21 ? n67007 : n32;
  assign n73432 = pi20 ? n73431 : n32;
  assign n73433 = pi19 ? n73160 : n73432;
  assign n73434 = pi18 ? n32 : n73433;
  assign n73435 = pi17 ? n32 : n73434;
  assign n73436 = pi16 ? n32 : n73435;
  assign n73437 = pi15 ? n73430 : n73436;
  assign n73438 = pi14 ? n73423 : n73437;
  assign n73439 = pi13 ? n73407 : n73438;
  assign n73440 = pi22 ? n56186 : n56665;
  assign n73441 = pi21 ? n73440 : n32;
  assign n73442 = pi20 ? n73441 : n32;
  assign n73443 = pi19 ? n73160 : n73442;
  assign n73444 = pi18 ? n32 : n73443;
  assign n73445 = pi17 ? n32 : n73444;
  assign n73446 = pi16 ? n32 : n73445;
  assign n73447 = pi19 ? n32 : n59675;
  assign n73448 = pi18 ? n32 : n73447;
  assign n73449 = pi17 ? n32 : n73448;
  assign n73450 = pi16 ? n32 : n73449;
  assign n73451 = pi15 ? n73446 : n73450;
  assign n73452 = pi19 ? n32 : n57717;
  assign n73453 = pi18 ? n32 : n73452;
  assign n73454 = pi17 ? n32 : n73453;
  assign n73455 = pi16 ? n32 : n73454;
  assign n73456 = pi15 ? n73455 : n73164;
  assign n73457 = pi14 ? n73451 : n73456;
  assign n73458 = pi13 ? n73457 : n32;
  assign n73459 = pi12 ? n73439 : n73458;
  assign n73460 = pi11 ? n73459 : n32;
  assign n73461 = pi10 ? n73379 : n73460;
  assign n73462 = pi09 ? n73208 : n73461;
  assign n73463 = pi20 ? n38376 : n13040;
  assign n73464 = pi19 ? n32 : n73463;
  assign n73465 = pi18 ? n32 : n73464;
  assign n73466 = pi17 ? n32 : n73465;
  assign n73467 = pi16 ? n32 : n73466;
  assign n73468 = pi15 ? n32 : n73467;
  assign n73469 = pi20 ? n38376 : n61008;
  assign n73470 = pi19 ? n32 : n73469;
  assign n73471 = pi18 ? n32 : n73470;
  assign n73472 = pi17 ? n32 : n73471;
  assign n73473 = pi16 ? n32 : n73472;
  assign n73474 = pi14 ? n73468 : n73473;
  assign n73475 = pi13 ? n32 : n73474;
  assign n73476 = pi12 ? n32 : n73475;
  assign n73477 = pi11 ? n32 : n73476;
  assign n73478 = pi10 ? n32 : n73477;
  assign n73479 = pi15 ? n73473 : n73213;
  assign n73480 = pi22 ? n30154 : n60973;
  assign n73481 = pi21 ? n73480 : n20563;
  assign n73482 = pi20 ? n73481 : n1619;
  assign n73483 = pi19 ? n32 : n73482;
  assign n73484 = pi18 ? n32 : n73483;
  assign n73485 = pi17 ? n32 : n73484;
  assign n73486 = pi16 ? n32 : n73485;
  assign n73487 = pi15 ? n72946 : n73486;
  assign n73488 = pi14 ? n73479 : n73487;
  assign n73489 = pi13 ? n73488 : n73220;
  assign n73490 = pi20 ? n59020 : n1619;
  assign n73491 = pi19 ? n32 : n73490;
  assign n73492 = pi18 ? n32 : n73491;
  assign n73493 = pi17 ? n32 : n73492;
  assign n73494 = pi16 ? n32 : n73493;
  assign n73495 = pi22 ? n41458 : n20563;
  assign n73496 = pi21 ? n73495 : n30868;
  assign n73497 = pi20 ? n73496 : n1619;
  assign n73498 = pi19 ? n32 : n73497;
  assign n73499 = pi18 ? n32 : n73498;
  assign n73500 = pi17 ? n32 : n73499;
  assign n73501 = pi16 ? n32 : n73500;
  assign n73502 = pi15 ? n73494 : n73501;
  assign n73503 = pi21 ? n73495 : n20563;
  assign n73504 = pi20 ? n73503 : n1619;
  assign n73505 = pi19 ? n32 : n73504;
  assign n73506 = pi18 ? n32 : n73505;
  assign n73507 = pi17 ? n32 : n73506;
  assign n73508 = pi16 ? n32 : n73507;
  assign n73509 = pi15 ? n73508 : n72946;
  assign n73510 = pi14 ? n73502 : n73509;
  assign n73511 = pi20 ? n31313 : n59305;
  assign n73512 = pi19 ? n32 : n73511;
  assign n73513 = pi18 ? n32 : n73512;
  assign n73514 = pi17 ? n32 : n73513;
  assign n73515 = pi16 ? n32 : n73514;
  assign n73516 = pi20 ? n72646 : n72686;
  assign n73517 = pi19 ? n32 : n73516;
  assign n73518 = pi18 ? n32 : n73517;
  assign n73519 = pi17 ? n32 : n73518;
  assign n73520 = pi16 ? n32 : n73519;
  assign n73521 = pi15 ? n73515 : n73520;
  assign n73522 = pi20 ? n59020 : n73235;
  assign n73523 = pi19 ? n32 : n73522;
  assign n73524 = pi18 ? n32 : n73523;
  assign n73525 = pi17 ? n32 : n73524;
  assign n73526 = pi16 ? n32 : n73525;
  assign n73527 = pi21 ? n37217 : n33792;
  assign n73528 = pi20 ? n73527 : n73244;
  assign n73529 = pi19 ? n32 : n73528;
  assign n73530 = pi18 ? n32 : n73529;
  assign n73531 = pi17 ? n32 : n73530;
  assign n73532 = pi16 ? n32 : n73531;
  assign n73533 = pi15 ? n73526 : n73532;
  assign n73534 = pi14 ? n73521 : n73533;
  assign n73535 = pi13 ? n73510 : n73534;
  assign n73536 = pi12 ? n73489 : n73535;
  assign n73537 = pi24 ? n33792 : n13481;
  assign n73538 = pi23 ? n73537 : n13481;
  assign n73539 = pi22 ? n73538 : n13481;
  assign n73540 = pi21 ? n73539 : n55560;
  assign n73541 = pi20 ? n73254 : n73540;
  assign n73542 = pi19 ? n32 : n73541;
  assign n73543 = pi18 ? n32 : n73542;
  assign n73544 = pi17 ? n32 : n73543;
  assign n73545 = pi16 ? n32 : n73544;
  assign n73546 = pi20 ? n73260 : n73001;
  assign n73547 = pi19 ? n32 : n73546;
  assign n73548 = pi18 ? n32 : n73547;
  assign n73549 = pi17 ? n32 : n73548;
  assign n73550 = pi16 ? n32 : n73549;
  assign n73551 = pi15 ? n73545 : n73550;
  assign n73552 = pi23 ? n1598 : n685;
  assign n73553 = pi22 ? n73552 : n51564;
  assign n73554 = pi21 ? n73553 : n2637;
  assign n73555 = pi20 ? n73267 : n73554;
  assign n73556 = pi19 ? n32 : n73555;
  assign n73557 = pi18 ? n32 : n73556;
  assign n73558 = pi17 ? n32 : n73557;
  assign n73559 = pi16 ? n32 : n73558;
  assign n73560 = pi22 ? n44028 : n316;
  assign n73561 = pi21 ? n73560 : n928;
  assign n73562 = pi20 ? n73275 : n73561;
  assign n73563 = pi19 ? n32 : n73562;
  assign n73564 = pi18 ? n32 : n73563;
  assign n73565 = pi17 ? n32 : n73564;
  assign n73566 = pi16 ? n32 : n73565;
  assign n73567 = pi15 ? n73559 : n73566;
  assign n73568 = pi14 ? n73551 : n73567;
  assign n73569 = pi19 ? n32 : n73287;
  assign n73570 = pi18 ? n32 : n73569;
  assign n73571 = pi17 ? n32 : n73570;
  assign n73572 = pi16 ? n32 : n73571;
  assign n73573 = pi20 ? n73292 : n11695;
  assign n73574 = pi19 ? n32 : n73573;
  assign n73575 = pi18 ? n32 : n73574;
  assign n73576 = pi17 ? n32 : n73575;
  assign n73577 = pi16 ? n32 : n73576;
  assign n73578 = pi15 ? n73572 : n73577;
  assign n73579 = pi21 ? n37784 : n61446;
  assign n73580 = pi20 ? n73579 : n70483;
  assign n73581 = pi19 ? n32 : n73580;
  assign n73582 = pi18 ? n32 : n73581;
  assign n73583 = pi17 ? n32 : n73582;
  assign n73584 = pi16 ? n32 : n73583;
  assign n73585 = pi19 ? n32 : n73308;
  assign n73586 = pi18 ? n32 : n73585;
  assign n73587 = pi17 ? n32 : n73586;
  assign n73588 = pi16 ? n32 : n73587;
  assign n73589 = pi15 ? n73584 : n73588;
  assign n73590 = pi14 ? n73578 : n73589;
  assign n73591 = pi13 ? n73568 : n73590;
  assign n73592 = pi19 ? n37927 : n73316;
  assign n73593 = pi18 ? n32 : n73592;
  assign n73594 = pi17 ? n32 : n73593;
  assign n73595 = pi16 ? n32 : n73594;
  assign n73596 = pi19 ? n49331 : n73322;
  assign n73597 = pi18 ? n32 : n73596;
  assign n73598 = pi17 ? n32 : n73597;
  assign n73599 = pi16 ? n32 : n73598;
  assign n73600 = pi15 ? n73595 : n73599;
  assign n73601 = pi19 ? n49331 : n73330;
  assign n73602 = pi18 ? n32 : n73601;
  assign n73603 = pi17 ? n32 : n73602;
  assign n73604 = pi16 ? n32 : n73603;
  assign n73605 = pi22 ? n52451 : n13481;
  assign n73606 = pi21 ? n47360 : n73605;
  assign n73607 = pi20 ? n73606 : n32257;
  assign n73608 = pi19 ? n73368 : n73607;
  assign n73609 = pi18 ? n32 : n73608;
  assign n73610 = pi17 ? n32 : n73609;
  assign n73611 = pi16 ? n32 : n73610;
  assign n73612 = pi15 ? n73604 : n73611;
  assign n73613 = pi14 ? n73600 : n73612;
  assign n73614 = pi19 ? n73368 : n73344;
  assign n73615 = pi18 ? n32 : n73614;
  assign n73616 = pi17 ? n32 : n73615;
  assign n73617 = pi16 ? n32 : n73616;
  assign n73618 = pi22 ? n59719 : n51564;
  assign n73619 = pi21 ? n36659 : n73618;
  assign n73620 = pi20 ? n73619 : n32;
  assign n73621 = pi19 ? n48847 : n73620;
  assign n73622 = pi18 ? n32 : n73621;
  assign n73623 = pi17 ? n32 : n73622;
  assign n73624 = pi16 ? n32 : n73623;
  assign n73625 = pi15 ? n73617 : n73624;
  assign n73626 = pi22 ? n64606 : n13481;
  assign n73627 = pi21 ? n36781 : n73626;
  assign n73628 = pi20 ? n73627 : n32;
  assign n73629 = pi19 ? n46202 : n73628;
  assign n73630 = pi18 ? n32 : n73629;
  assign n73631 = pi17 ? n32 : n73630;
  assign n73632 = pi16 ? n32 : n73631;
  assign n73633 = pi14 ? n73625 : n73632;
  assign n73634 = pi13 ? n73613 : n73633;
  assign n73635 = pi12 ? n73591 : n73634;
  assign n73636 = pi11 ? n73536 : n73635;
  assign n73637 = pi22 ? n61806 : n21502;
  assign n73638 = pi21 ? n64961 : n73637;
  assign n73639 = pi20 ? n73638 : n32;
  assign n73640 = pi19 ? n32 : n73639;
  assign n73641 = pi18 ? n32 : n73640;
  assign n73642 = pi17 ? n32 : n73641;
  assign n73643 = pi16 ? n32 : n73642;
  assign n73644 = pi22 ? n61806 : n32;
  assign n73645 = pi21 ? n57774 : n73644;
  assign n73646 = pi20 ? n73645 : n32;
  assign n73647 = pi19 ? n32 : n73646;
  assign n73648 = pi18 ? n32 : n73647;
  assign n73649 = pi17 ? n32 : n73648;
  assign n73650 = pi16 ? n32 : n73649;
  assign n73651 = pi15 ? n73643 : n73650;
  assign n73652 = pi21 ? n63253 : n59785;
  assign n73653 = pi20 ? n73652 : n32;
  assign n73654 = pi19 ? n32 : n73653;
  assign n73655 = pi18 ? n32 : n73654;
  assign n73656 = pi17 ? n32 : n73655;
  assign n73657 = pi16 ? n32 : n73656;
  assign n73658 = pi22 ? n71505 : n51564;
  assign n73659 = pi21 ? n73658 : n55560;
  assign n73660 = pi20 ? n73659 : n32;
  assign n73661 = pi19 ? n32 : n73660;
  assign n73662 = pi18 ? n32 : n73661;
  assign n73663 = pi17 ? n32 : n73662;
  assign n73664 = pi16 ? n32 : n73663;
  assign n73665 = pi15 ? n73657 : n73664;
  assign n73666 = pi14 ? n73651 : n73665;
  assign n73667 = pi21 ? n73658 : n32;
  assign n73668 = pi20 ? n73667 : n32;
  assign n73669 = pi19 ? n32 : n73668;
  assign n73670 = pi18 ? n32 : n73669;
  assign n73671 = pi17 ? n32 : n73670;
  assign n73672 = pi16 ? n32 : n73671;
  assign n73673 = pi22 ? n71523 : n13481;
  assign n73674 = pi21 ? n73673 : n32;
  assign n73675 = pi20 ? n73674 : n32;
  assign n73676 = pi19 ? n32 : n73675;
  assign n73677 = pi18 ? n32 : n73676;
  assign n73678 = pi17 ? n32 : n73677;
  assign n73679 = pi16 ? n32 : n73678;
  assign n73680 = pi15 ? n73672 : n73679;
  assign n73681 = pi23 ? n63431 : n13481;
  assign n73682 = pi22 ? n73681 : n13481;
  assign n73683 = pi21 ? n73682 : n32;
  assign n73684 = pi20 ? n73683 : n32;
  assign n73685 = pi19 ? n32 : n73684;
  assign n73686 = pi18 ? n32 : n73685;
  assign n73687 = pi17 ? n32 : n73686;
  assign n73688 = pi16 ? n32 : n73687;
  assign n73689 = pi23 ? n63431 : n71896;
  assign n73690 = pi22 ? n73689 : n32;
  assign n73691 = pi21 ? n73690 : n32;
  assign n73692 = pi20 ? n73691 : n32;
  assign n73693 = pi19 ? n32 : n73692;
  assign n73694 = pi18 ? n32 : n73693;
  assign n73695 = pi17 ? n32 : n73694;
  assign n73696 = pi16 ? n32 : n73695;
  assign n73697 = pi15 ? n73688 : n73696;
  assign n73698 = pi14 ? n73680 : n73697;
  assign n73699 = pi13 ? n73666 : n73698;
  assign n73700 = pi22 ? n71144 : n32;
  assign n73701 = pi21 ? n73700 : n32;
  assign n73702 = pi20 ? n73701 : n32;
  assign n73703 = pi19 ? n32 : n73702;
  assign n73704 = pi18 ? n32 : n73703;
  assign n73705 = pi17 ? n32 : n73704;
  assign n73706 = pi16 ? n32 : n73705;
  assign n73707 = pi22 ? n71152 : n32;
  assign n73708 = pi21 ? n73707 : n32;
  assign n73709 = pi20 ? n73708 : n32;
  assign n73710 = pi19 ? n32 : n73709;
  assign n73711 = pi18 ? n32 : n73710;
  assign n73712 = pi17 ? n32 : n73711;
  assign n73713 = pi16 ? n32 : n73712;
  assign n73714 = pi15 ? n73713 : n73455;
  assign n73715 = pi14 ? n73706 : n73714;
  assign n73716 = pi13 ? n73715 : n32;
  assign n73717 = pi12 ? n73699 : n73716;
  assign n73718 = pi11 ? n73717 : n32;
  assign n73719 = pi10 ? n73636 : n73718;
  assign n73720 = pi09 ? n73478 : n73719;
  assign n73721 = pi08 ? n73462 : n73720;
  assign n73722 = pi20 ? n37333 : n13040;
  assign n73723 = pi19 ? n32 : n73722;
  assign n73724 = pi18 ? n32 : n73723;
  assign n73725 = pi17 ? n32 : n73724;
  assign n73726 = pi16 ? n32 : n73725;
  assign n73727 = pi15 ? n32 : n73726;
  assign n73728 = pi14 ? n73727 : n73473;
  assign n73729 = pi13 ? n32 : n73728;
  assign n73730 = pi12 ? n32 : n73729;
  assign n73731 = pi11 ? n32 : n73730;
  assign n73732 = pi10 ? n32 : n73731;
  assign n73733 = pi20 ? n39395 : n61008;
  assign n73734 = pi19 ? n32 : n73733;
  assign n73735 = pi18 ? n32 : n73734;
  assign n73736 = pi17 ? n32 : n73735;
  assign n73737 = pi16 ? n32 : n73736;
  assign n73738 = pi15 ? n73473 : n73737;
  assign n73739 = pi22 ? n32 : n31993;
  assign n73740 = pi21 ? n73739 : n20563;
  assign n73741 = pi20 ? n73740 : n1619;
  assign n73742 = pi19 ? n32 : n73741;
  assign n73743 = pi18 ? n32 : n73742;
  assign n73744 = pi17 ? n32 : n73743;
  assign n73745 = pi16 ? n32 : n73744;
  assign n73746 = pi21 ? n39394 : n37;
  assign n73747 = pi20 ? n73746 : n1619;
  assign n73748 = pi19 ? n32 : n73747;
  assign n73749 = pi18 ? n32 : n73748;
  assign n73750 = pi17 ? n32 : n73749;
  assign n73751 = pi16 ? n32 : n73750;
  assign n73752 = pi15 ? n73745 : n73751;
  assign n73753 = pi14 ? n73738 : n73752;
  assign n73754 = pi20 ? n28157 : n1619;
  assign n73755 = pi19 ? n32 : n73754;
  assign n73756 = pi18 ? n32 : n73755;
  assign n73757 = pi17 ? n32 : n73756;
  assign n73758 = pi16 ? n32 : n73757;
  assign n73759 = pi20 ? n30117 : n1619;
  assign n73760 = pi19 ? n32 : n73759;
  assign n73761 = pi18 ? n32 : n73760;
  assign n73762 = pi17 ? n32 : n73761;
  assign n73763 = pi16 ? n32 : n73762;
  assign n73764 = pi15 ? n73758 : n73763;
  assign n73765 = pi15 ? n73763 : n72946;
  assign n73766 = pi14 ? n73764 : n73765;
  assign n73767 = pi13 ? n73753 : n73766;
  assign n73768 = pi14 ? n72639 : n73487;
  assign n73769 = pi20 ? n59020 : n67195;
  assign n73770 = pi19 ? n32 : n73769;
  assign n73771 = pi18 ? n32 : n73770;
  assign n73772 = pi17 ? n32 : n73771;
  assign n73773 = pi16 ? n32 : n73772;
  assign n73774 = pi15 ? n73515 : n73773;
  assign n73775 = pi24 ? n99 : n51564;
  assign n73776 = pi23 ? n73775 : n51564;
  assign n73777 = pi22 ? n73776 : n51564;
  assign n73778 = pi21 ? n73777 : n58966;
  assign n73779 = pi20 ? n59020 : n73778;
  assign n73780 = pi19 ? n32 : n73779;
  assign n73781 = pi18 ? n32 : n73780;
  assign n73782 = pi17 ? n32 : n73781;
  assign n73783 = pi16 ? n32 : n73782;
  assign n73784 = pi21 ? n57350 : n33095;
  assign n73785 = pi20 ? n60377 : n73784;
  assign n73786 = pi19 ? n32 : n73785;
  assign n73787 = pi18 ? n32 : n73786;
  assign n73788 = pi17 ? n32 : n73787;
  assign n73789 = pi16 ? n32 : n73788;
  assign n73790 = pi15 ? n73783 : n73789;
  assign n73791 = pi14 ? n73774 : n73790;
  assign n73792 = pi13 ? n73768 : n73791;
  assign n73793 = pi12 ? n73767 : n73792;
  assign n73794 = pi21 ? n30866 : n47360;
  assign n73795 = pi24 ? n335 : n13481;
  assign n73796 = pi23 ? n73795 : n13481;
  assign n73797 = pi22 ? n73796 : n13481;
  assign n73798 = pi21 ? n73797 : n55560;
  assign n73799 = pi20 ? n73794 : n73798;
  assign n73800 = pi19 ? n32 : n73799;
  assign n73801 = pi18 ? n32 : n73800;
  assign n73802 = pi17 ? n32 : n73801;
  assign n73803 = pi16 ? n32 : n73802;
  assign n73804 = pi21 ? n73495 : n47360;
  assign n73805 = pi21 ? n73000 : n59357;
  assign n73806 = pi20 ? n73804 : n73805;
  assign n73807 = pi19 ? n32 : n73806;
  assign n73808 = pi18 ? n32 : n73807;
  assign n73809 = pi17 ? n32 : n73808;
  assign n73810 = pi16 ? n32 : n73809;
  assign n73811 = pi15 ? n73803 : n73810;
  assign n73812 = pi21 ? n73495 : n39952;
  assign n73813 = pi24 ? n204 : n51564;
  assign n73814 = pi23 ? n73813 : n51564;
  assign n73815 = pi22 ? n73814 : n51564;
  assign n73816 = pi21 ? n73815 : n59357;
  assign n73817 = pi20 ? n73812 : n73816;
  assign n73818 = pi19 ? n32 : n73817;
  assign n73819 = pi18 ? n32 : n73818;
  assign n73820 = pi17 ? n32 : n73819;
  assign n73821 = pi16 ? n32 : n73820;
  assign n73822 = pi22 ? n41481 : n30868;
  assign n73823 = pi21 ? n73822 : n39952;
  assign n73824 = pi21 ? n73560 : n37639;
  assign n73825 = pi20 ? n73823 : n73824;
  assign n73826 = pi19 ? n32 : n73825;
  assign n73827 = pi18 ? n32 : n73826;
  assign n73828 = pi17 ? n32 : n73827;
  assign n73829 = pi16 ? n32 : n73828;
  assign n73830 = pi15 ? n73821 : n73829;
  assign n73831 = pi14 ? n73811 : n73830;
  assign n73832 = pi21 ? n63179 : n59524;
  assign n73833 = pi20 ? n73832 : n61537;
  assign n73834 = pi19 ? n32 : n73833;
  assign n73835 = pi18 ? n32 : n73834;
  assign n73836 = pi17 ? n32 : n73835;
  assign n73837 = pi16 ? n32 : n73836;
  assign n73838 = pi22 ? n30154 : n36615;
  assign n73839 = pi21 ? n73838 : n59524;
  assign n73840 = pi20 ? n73839 : n67712;
  assign n73841 = pi19 ? n32 : n73840;
  assign n73842 = pi18 ? n32 : n73841;
  assign n73843 = pi17 ? n32 : n73842;
  assign n73844 = pi16 ? n32 : n73843;
  assign n73845 = pi15 ? n73837 : n73844;
  assign n73846 = pi22 ? n45597 : n39190;
  assign n73847 = pi21 ? n73846 : n53471;
  assign n73848 = pi20 ? n73847 : n67719;
  assign n73849 = pi19 ? n32 : n73848;
  assign n73850 = pi18 ? n32 : n73849;
  assign n73851 = pi17 ? n32 : n73850;
  assign n73852 = pi16 ? n32 : n73851;
  assign n73853 = pi22 ? n45597 : n45106;
  assign n73854 = pi21 ? n73853 : n64961;
  assign n73855 = pi20 ? n73854 : n68653;
  assign n73856 = pi19 ? n32 : n73855;
  assign n73857 = pi18 ? n32 : n73856;
  assign n73858 = pi17 ? n32 : n73857;
  assign n73859 = pi16 ? n32 : n73858;
  assign n73860 = pi15 ? n73852 : n73859;
  assign n73861 = pi14 ? n73845 : n73860;
  assign n73862 = pi13 ? n73831 : n73861;
  assign n73863 = pi22 ? n37216 : n42109;
  assign n73864 = pi21 ? n73863 : n64961;
  assign n73865 = pi20 ? n73864 : n59649;
  assign n73866 = pi19 ? n32 : n73865;
  assign n73867 = pi18 ? n32 : n73866;
  assign n73868 = pi17 ? n32 : n73867;
  assign n73869 = pi16 ? n32 : n73868;
  assign n73870 = pi22 ? n37229 : n66956;
  assign n73871 = pi21 ? n73870 : n59595;
  assign n73872 = pi20 ? n73871 : n62857;
  assign n73873 = pi19 ? n32 : n73872;
  assign n73874 = pi18 ? n32 : n73873;
  assign n73875 = pi17 ? n32 : n73874;
  assign n73876 = pi16 ? n32 : n73875;
  assign n73877 = pi15 ? n73869 : n73876;
  assign n73878 = pi23 ? n55580 : n335;
  assign n73879 = pi22 ? n37229 : n73878;
  assign n73880 = pi21 ? n73879 : n63253;
  assign n73881 = pi20 ? n73880 : n3210;
  assign n73882 = pi19 ? n32 : n73881;
  assign n73883 = pi18 ? n32 : n73882;
  assign n73884 = pi17 ? n32 : n73883;
  assign n73885 = pi16 ? n32 : n73884;
  assign n73886 = pi22 ? n37229 : n36659;
  assign n73887 = pi21 ? n73886 : n59774;
  assign n73888 = pi20 ? n73887 : n32257;
  assign n73889 = pi19 ? n32 : n73888;
  assign n73890 = pi18 ? n32 : n73889;
  assign n73891 = pi17 ? n32 : n73890;
  assign n73892 = pi16 ? n32 : n73891;
  assign n73893 = pi15 ? n73885 : n73892;
  assign n73894 = pi14 ? n73877 : n73893;
  assign n73895 = pi23 ? n56079 : n363;
  assign n73896 = pi22 ? n37804 : n73895;
  assign n73897 = pi21 ? n73896 : n69327;
  assign n73898 = pi20 ? n73897 : n37640;
  assign n73899 = pi19 ? n32 : n73898;
  assign n73900 = pi18 ? n32 : n73899;
  assign n73901 = pi17 ? n32 : n73900;
  assign n73902 = pi16 ? n32 : n73901;
  assign n73903 = pi24 ? n363 : n36781;
  assign n73904 = pi23 ? n73903 : n36781;
  assign n73905 = pi22 ? n37804 : n73904;
  assign n73906 = pi21 ? n73905 : n56760;
  assign n73907 = pi20 ? n73906 : n32;
  assign n73908 = pi19 ? n32 : n73907;
  assign n73909 = pi18 ? n32 : n73908;
  assign n73910 = pi17 ? n32 : n73909;
  assign n73911 = pi16 ? n32 : n73910;
  assign n73912 = pi15 ? n73902 : n73911;
  assign n73913 = pi22 ? n37251 : n57782;
  assign n73914 = pi22 ? n14626 : n62473;
  assign n73915 = pi21 ? n73913 : n73914;
  assign n73916 = pi20 ? n73915 : n32;
  assign n73917 = pi19 ? n32 : n73916;
  assign n73918 = pi18 ? n32 : n73917;
  assign n73919 = pi17 ? n32 : n73918;
  assign n73920 = pi16 ? n32 : n73919;
  assign n73921 = pi21 ? n39968 : n57760;
  assign n73922 = pi20 ? n73921 : n32;
  assign n73923 = pi19 ? n32 : n73922;
  assign n73924 = pi18 ? n32 : n73923;
  assign n73925 = pi17 ? n32 : n73924;
  assign n73926 = pi16 ? n32 : n73925;
  assign n73927 = pi15 ? n73920 : n73926;
  assign n73928 = pi14 ? n73912 : n73927;
  assign n73929 = pi13 ? n73894 : n73928;
  assign n73930 = pi12 ? n73862 : n73929;
  assign n73931 = pi11 ? n73793 : n73930;
  assign n73932 = pi22 ? n37873 : n64678;
  assign n73933 = pi21 ? n73932 : n58470;
  assign n73934 = pi20 ? n73933 : n32;
  assign n73935 = pi19 ? n32 : n73934;
  assign n73936 = pi18 ? n32 : n73935;
  assign n73937 = pi17 ? n32 : n73936;
  assign n73938 = pi16 ? n32 : n73937;
  assign n73939 = pi23 ? n36782 : n14626;
  assign n73940 = pi24 ? n204 : n14626;
  assign n73941 = pi23 ? n73940 : n233;
  assign n73942 = pi22 ? n73939 : n73941;
  assign n73943 = pi21 ? n73942 : n60421;
  assign n73944 = pi20 ? n73943 : n32;
  assign n73945 = pi19 ? n32 : n73944;
  assign n73946 = pi18 ? n32 : n73945;
  assign n73947 = pi17 ? n32 : n73946;
  assign n73948 = pi16 ? n32 : n73947;
  assign n73949 = pi15 ? n73938 : n73948;
  assign n73950 = pi23 ? n14627 : n14626;
  assign n73951 = pi22 ? n36783 : n73950;
  assign n73952 = pi21 ? n73951 : n55560;
  assign n73953 = pi20 ? n73952 : n32;
  assign n73954 = pi19 ? n32 : n73953;
  assign n73955 = pi18 ? n32 : n73954;
  assign n73956 = pi17 ? n32 : n73955;
  assign n73957 = pi16 ? n32 : n73956;
  assign n73958 = pi23 ? n71143 : n51564;
  assign n73959 = pi24 ? n233 : n51564;
  assign n73960 = pi23 ? n73959 : n51564;
  assign n73961 = pi22 ? n73958 : n73960;
  assign n73962 = pi21 ? n73961 : n55560;
  assign n73963 = pi20 ? n73962 : n32;
  assign n73964 = pi19 ? n32 : n73963;
  assign n73965 = pi18 ? n32 : n73964;
  assign n73966 = pi17 ? n32 : n73965;
  assign n73967 = pi16 ? n32 : n73966;
  assign n73968 = pi15 ? n73957 : n73967;
  assign n73969 = pi14 ? n73949 : n73968;
  assign n73970 = pi22 ? n70744 : n51564;
  assign n73971 = pi21 ? n73970 : n32;
  assign n73972 = pi20 ? n73971 : n32;
  assign n73973 = pi19 ? n32 : n73972;
  assign n73974 = pi18 ? n32 : n73973;
  assign n73975 = pi17 ? n32 : n73974;
  assign n73976 = pi16 ? n32 : n73975;
  assign n73977 = pi23 ? n69724 : n13481;
  assign n73978 = pi22 ? n71924 : n73977;
  assign n73979 = pi21 ? n73978 : n32;
  assign n73980 = pi20 ? n73979 : n32;
  assign n73981 = pi19 ? n32 : n73980;
  assign n73982 = pi18 ? n32 : n73981;
  assign n73983 = pi17 ? n32 : n73982;
  assign n73984 = pi16 ? n32 : n73983;
  assign n73985 = pi15 ? n73976 : n73984;
  assign n73986 = pi22 ? n69890 : n13481;
  assign n73987 = pi21 ? n73986 : n32;
  assign n73988 = pi20 ? n73987 : n32;
  assign n73989 = pi19 ? n32 : n73988;
  assign n73990 = pi18 ? n32 : n73989;
  assign n73991 = pi17 ? n32 : n73990;
  assign n73992 = pi16 ? n32 : n73991;
  assign n73993 = pi22 ? n69401 : n32;
  assign n73994 = pi21 ? n73993 : n32;
  assign n73995 = pi20 ? n73994 : n32;
  assign n73996 = pi19 ? n32 : n73995;
  assign n73997 = pi18 ? n32 : n73996;
  assign n73998 = pi17 ? n32 : n73997;
  assign n73999 = pi16 ? n32 : n73998;
  assign n74000 = pi15 ? n73992 : n73999;
  assign n74001 = pi14 ? n73985 : n74000;
  assign n74002 = pi13 ? n73969 : n74001;
  assign n74003 = pi12 ? n74002 : n32;
  assign n74004 = pi11 ? n74003 : n32;
  assign n74005 = pi10 ? n73931 : n74004;
  assign n74006 = pi09 ? n73732 : n74005;
  assign n74007 = pi20 ? n37320 : n13040;
  assign n74008 = pi19 ? n32 : n74007;
  assign n74009 = pi18 ? n32 : n74008;
  assign n74010 = pi17 ? n32 : n74009;
  assign n74011 = pi16 ? n32 : n74010;
  assign n74012 = pi15 ? n32 : n74011;
  assign n74013 = pi20 ? n37320 : n61008;
  assign n74014 = pi19 ? n32 : n74013;
  assign n74015 = pi18 ? n32 : n74014;
  assign n74016 = pi17 ? n32 : n74015;
  assign n74017 = pi16 ? n32 : n74016;
  assign n74018 = pi14 ? n74012 : n74017;
  assign n74019 = pi13 ? n32 : n74018;
  assign n74020 = pi12 ? n32 : n74019;
  assign n74021 = pi11 ? n32 : n74020;
  assign n74022 = pi10 ? n32 : n74021;
  assign n74023 = pi15 ? n74017 : n73737;
  assign n74024 = pi20 ? n39395 : n1619;
  assign n74025 = pi19 ? n32 : n74024;
  assign n74026 = pi18 ? n32 : n74025;
  assign n74027 = pi17 ? n32 : n74026;
  assign n74028 = pi16 ? n32 : n74027;
  assign n74029 = pi21 ? n28156 : n35230;
  assign n74030 = pi20 ? n74029 : n1619;
  assign n74031 = pi19 ? n32 : n74030;
  assign n74032 = pi18 ? n32 : n74031;
  assign n74033 = pi17 ? n32 : n74032;
  assign n74034 = pi16 ? n32 : n74033;
  assign n74035 = pi15 ? n74028 : n74034;
  assign n74036 = pi14 ? n74023 : n74035;
  assign n74037 = pi15 ? n73758 : n74028;
  assign n74038 = pi14 ? n74037 : n74028;
  assign n74039 = pi13 ? n74036 : n74038;
  assign n74040 = pi20 ? n50676 : n1619;
  assign n74041 = pi19 ? n32 : n74040;
  assign n74042 = pi18 ? n32 : n74041;
  assign n74043 = pi17 ? n32 : n74042;
  assign n74044 = pi16 ? n32 : n74043;
  assign n74045 = pi14 ? n74044 : n74028;
  assign n74046 = pi20 ? n28157 : n59305;
  assign n74047 = pi19 ? n32 : n74046;
  assign n74048 = pi18 ? n32 : n74047;
  assign n74049 = pi17 ? n32 : n74048;
  assign n74050 = pi16 ? n32 : n74049;
  assign n74051 = pi20 ? n63353 : n67195;
  assign n74052 = pi19 ? n32 : n74051;
  assign n74053 = pi18 ? n32 : n74052;
  assign n74054 = pi17 ? n32 : n74053;
  assign n74055 = pi16 ? n32 : n74054;
  assign n74056 = pi15 ? n74050 : n74055;
  assign n74057 = pi20 ? n63353 : n73778;
  assign n74058 = pi19 ? n32 : n74057;
  assign n74059 = pi18 ? n32 : n74058;
  assign n74060 = pi17 ? n32 : n74059;
  assign n74061 = pi16 ? n32 : n74060;
  assign n74062 = pi21 ? n30155 : n33792;
  assign n74063 = pi20 ? n74062 : n73784;
  assign n74064 = pi19 ? n32 : n74063;
  assign n74065 = pi18 ? n32 : n74064;
  assign n74066 = pi17 ? n32 : n74065;
  assign n74067 = pi16 ? n32 : n74066;
  assign n74068 = pi15 ? n74061 : n74067;
  assign n74069 = pi14 ? n74056 : n74068;
  assign n74070 = pi13 ? n74045 : n74069;
  assign n74071 = pi12 ? n74039 : n74070;
  assign n74072 = pi21 ? n30155 : n47360;
  assign n74073 = pi23 ? n6960 : n13481;
  assign n74074 = pi22 ? n74073 : n13481;
  assign n74075 = pi21 ? n74074 : n37639;
  assign n74076 = pi20 ? n74072 : n74075;
  assign n74077 = pi19 ? n32 : n74076;
  assign n74078 = pi18 ? n32 : n74077;
  assign n74079 = pi17 ? n32 : n74078;
  assign n74080 = pi16 ? n32 : n74079;
  assign n74081 = pi20 ? n74072 : n73805;
  assign n74082 = pi19 ? n32 : n74081;
  assign n74083 = pi18 ? n32 : n74082;
  assign n74084 = pi17 ? n32 : n74083;
  assign n74085 = pi16 ? n32 : n74084;
  assign n74086 = pi15 ? n74080 : n74085;
  assign n74087 = pi21 ? n30155 : n39952;
  assign n74088 = pi20 ? n74087 : n73816;
  assign n74089 = pi19 ? n32 : n74088;
  assign n74090 = pi18 ? n32 : n74089;
  assign n74091 = pi17 ? n32 : n74090;
  assign n74092 = pi16 ? n32 : n74091;
  assign n74093 = pi21 ? n68255 : n39952;
  assign n74094 = pi20 ? n74093 : n73824;
  assign n74095 = pi19 ? n32 : n74094;
  assign n74096 = pi18 ? n32 : n74095;
  assign n74097 = pi17 ? n32 : n74096;
  assign n74098 = pi16 ? n32 : n74097;
  assign n74099 = pi15 ? n74092 : n74098;
  assign n74100 = pi14 ? n74086 : n74099;
  assign n74101 = pi22 ? n13481 : n61712;
  assign n74102 = pi21 ? n74101 : n32;
  assign n74103 = pi20 ? n73832 : n74102;
  assign n74104 = pi19 ? n32 : n74103;
  assign n74105 = pi18 ? n32 : n74104;
  assign n74106 = pi17 ? n32 : n74105;
  assign n74107 = pi16 ? n32 : n74106;
  assign n74108 = pi15 ? n74107 : n73844;
  assign n74109 = pi20 ? n73854 : n5667;
  assign n74110 = pi19 ? n32 : n74109;
  assign n74111 = pi18 ? n32 : n74110;
  assign n74112 = pi17 ? n32 : n74111;
  assign n74113 = pi16 ? n32 : n74112;
  assign n74114 = pi15 ? n73852 : n74113;
  assign n74115 = pi14 ? n74108 : n74114;
  assign n74116 = pi13 ? n74100 : n74115;
  assign n74117 = pi22 ? n49720 : n42109;
  assign n74118 = pi21 ? n74117 : n64961;
  assign n74119 = pi20 ? n74118 : n60045;
  assign n74120 = pi19 ? n32 : n74119;
  assign n74121 = pi18 ? n32 : n74120;
  assign n74122 = pi17 ? n32 : n74121;
  assign n74123 = pi16 ? n32 : n74122;
  assign n74124 = pi24 ? n99 : n36781;
  assign n74125 = pi23 ? n74124 : n33792;
  assign n74126 = pi22 ? n51754 : n74125;
  assign n74127 = pi21 ? n74126 : n59595;
  assign n74128 = pi20 ? n74127 : n62857;
  assign n74129 = pi19 ? n32 : n74128;
  assign n74130 = pi18 ? n32 : n74129;
  assign n74131 = pi17 ? n32 : n74130;
  assign n74132 = pi16 ? n32 : n74131;
  assign n74133 = pi15 ? n74123 : n74132;
  assign n74134 = pi23 ? n8184 : n335;
  assign n74135 = pi22 ? n51754 : n74134;
  assign n74136 = pi21 ? n74135 : n63253;
  assign n74137 = pi20 ? n74136 : n3210;
  assign n74138 = pi19 ? n32 : n74137;
  assign n74139 = pi18 ? n32 : n74138;
  assign n74140 = pi17 ? n32 : n74139;
  assign n74141 = pi16 ? n32 : n74140;
  assign n74142 = pi21 ? n72455 : n59774;
  assign n74143 = pi20 ? n74142 : n2653;
  assign n74144 = pi19 ? n32 : n74143;
  assign n74145 = pi18 ? n32 : n74144;
  assign n74146 = pi17 ? n32 : n74145;
  assign n74147 = pi16 ? n32 : n74146;
  assign n74148 = pi15 ? n74141 : n74147;
  assign n74149 = pi14 ? n74133 : n74148;
  assign n74150 = pi23 ? n19714 : n363;
  assign n74151 = pi22 ? n45516 : n74150;
  assign n74152 = pi21 ? n74151 : n69327;
  assign n74153 = pi20 ? n74152 : n32;
  assign n74154 = pi19 ? n32 : n74153;
  assign n74155 = pi18 ? n32 : n74154;
  assign n74156 = pi17 ? n32 : n74155;
  assign n74157 = pi16 ? n32 : n74156;
  assign n74158 = pi22 ? n46757 : n36781;
  assign n74159 = pi21 ? n74158 : n56760;
  assign n74160 = pi20 ? n74159 : n32;
  assign n74161 = pi19 ? n32 : n74160;
  assign n74162 = pi18 ? n32 : n74161;
  assign n74163 = pi17 ? n32 : n74162;
  assign n74164 = pi16 ? n32 : n74163;
  assign n74165 = pi15 ? n74157 : n74164;
  assign n74166 = pi22 ? n46757 : n62510;
  assign n74167 = pi21 ? n74166 : n73914;
  assign n74168 = pi20 ? n74167 : n32;
  assign n74169 = pi19 ? n32 : n74168;
  assign n74170 = pi18 ? n32 : n74169;
  assign n74171 = pi17 ? n32 : n74170;
  assign n74172 = pi16 ? n32 : n74171;
  assign n74173 = pi21 ? n59129 : n60421;
  assign n74174 = pi20 ? n74173 : n32;
  assign n74175 = pi19 ? n32 : n74174;
  assign n74176 = pi18 ? n32 : n74175;
  assign n74177 = pi17 ? n32 : n74176;
  assign n74178 = pi16 ? n32 : n74177;
  assign n74179 = pi15 ? n74172 : n74178;
  assign n74180 = pi14 ? n74165 : n74179;
  assign n74181 = pi13 ? n74149 : n74180;
  assign n74182 = pi12 ? n74116 : n74181;
  assign n74183 = pi11 ? n74071 : n74182;
  assign n74184 = pi22 ? n45634 : n64678;
  assign n74185 = pi21 ? n74184 : n60421;
  assign n74186 = pi20 ? n74185 : n32;
  assign n74187 = pi19 ? n32 : n74186;
  assign n74188 = pi18 ? n32 : n74187;
  assign n74189 = pi17 ? n32 : n74188;
  assign n74190 = pi16 ? n32 : n74189;
  assign n74191 = pi23 ? n58566 : n14626;
  assign n74192 = pi22 ? n45652 : n74191;
  assign n74193 = pi21 ? n74192 : n60421;
  assign n74194 = pi20 ? n74193 : n32;
  assign n74195 = pi19 ? n32 : n74194;
  assign n74196 = pi18 ? n32 : n74195;
  assign n74197 = pi17 ? n32 : n74196;
  assign n74198 = pi16 ? n32 : n74197;
  assign n74199 = pi15 ? n74190 : n74198;
  assign n74200 = pi21 ? n71098 : n1009;
  assign n74201 = pi20 ? n74200 : n32;
  assign n74202 = pi19 ? n32 : n74201;
  assign n74203 = pi18 ? n32 : n74202;
  assign n74204 = pi17 ? n32 : n74203;
  assign n74205 = pi16 ? n32 : n74204;
  assign n74206 = pi23 ? n63306 : n51564;
  assign n74207 = pi22 ? n46275 : n74206;
  assign n74208 = pi21 ? n74207 : n32;
  assign n74209 = pi20 ? n74208 : n32;
  assign n74210 = pi19 ? n32 : n74209;
  assign n74211 = pi18 ? n32 : n74210;
  assign n74212 = pi17 ? n32 : n74211;
  assign n74213 = pi16 ? n32 : n74212;
  assign n74214 = pi15 ? n74205 : n74213;
  assign n74215 = pi14 ? n74199 : n74214;
  assign n74216 = pi22 ? n63432 : n51564;
  assign n74217 = pi21 ? n74216 : n32;
  assign n74218 = pi20 ? n74217 : n32;
  assign n74219 = pi19 ? n32 : n74218;
  assign n74220 = pi18 ? n32 : n74219;
  assign n74221 = pi17 ? n32 : n74220;
  assign n74222 = pi16 ? n32 : n74221;
  assign n74223 = pi22 ? n71540 : n73977;
  assign n74224 = pi21 ? n74223 : n32;
  assign n74225 = pi20 ? n74224 : n32;
  assign n74226 = pi19 ? n32 : n74225;
  assign n74227 = pi18 ? n32 : n74226;
  assign n74228 = pi17 ? n32 : n74227;
  assign n74229 = pi16 ? n32 : n74228;
  assign n74230 = pi15 ? n74222 : n74229;
  assign n74231 = pi21 ? n69402 : n32;
  assign n74232 = pi20 ? n74231 : n32;
  assign n74233 = pi19 ? n32 : n74232;
  assign n74234 = pi18 ? n32 : n74233;
  assign n74235 = pi17 ? n32 : n74234;
  assign n74236 = pi16 ? n32 : n74235;
  assign n74237 = pi15 ? n74236 : n73999;
  assign n74238 = pi14 ? n74230 : n74237;
  assign n74239 = pi13 ? n74215 : n74238;
  assign n74240 = pi12 ? n74239 : n32;
  assign n74241 = pi11 ? n74240 : n32;
  assign n74242 = pi10 ? n74183 : n74241;
  assign n74243 = pi09 ? n74022 : n74242;
  assign n74244 = pi08 ? n74006 : n74243;
  assign n74245 = pi07 ? n73721 : n74244;
  assign n74246 = pi21 ? n20563 : n13039;
  assign n74247 = pi20 ? n38997 : n74246;
  assign n74248 = pi19 ? n32 : n74247;
  assign n74249 = pi18 ? n32 : n74248;
  assign n74250 = pi17 ? n32 : n74249;
  assign n74251 = pi16 ? n32 : n74250;
  assign n74252 = pi15 ? n32 : n74251;
  assign n74253 = pi21 ? n32 : n31293;
  assign n74254 = pi20 ? n74253 : n61008;
  assign n74255 = pi19 ? n32 : n74254;
  assign n74256 = pi18 ? n32 : n74255;
  assign n74257 = pi17 ? n32 : n74256;
  assign n74258 = pi16 ? n32 : n74257;
  assign n74259 = pi14 ? n74252 : n74258;
  assign n74260 = pi13 ? n32 : n74259;
  assign n74261 = pi12 ? n32 : n74260;
  assign n74262 = pi11 ? n32 : n74261;
  assign n74263 = pi10 ? n32 : n74262;
  assign n74264 = pi20 ? n37333 : n61008;
  assign n74265 = pi19 ? n32 : n74264;
  assign n74266 = pi18 ? n32 : n74265;
  assign n74267 = pi17 ? n32 : n74266;
  assign n74268 = pi16 ? n32 : n74267;
  assign n74269 = pi15 ? n74258 : n74268;
  assign n74270 = pi20 ? n38376 : n1619;
  assign n74271 = pi19 ? n32 : n74270;
  assign n74272 = pi18 ? n32 : n74271;
  assign n74273 = pi17 ? n32 : n74272;
  assign n74274 = pi16 ? n32 : n74273;
  assign n74275 = pi14 ? n74269 : n74274;
  assign n74276 = pi14 ? n74274 : n74028;
  assign n74277 = pi13 ? n74275 : n74276;
  assign n74278 = pi22 ? n59303 : n14626;
  assign n74279 = pi21 ? n74278 : n65115;
  assign n74280 = pi20 ? n28157 : n74279;
  assign n74281 = pi19 ? n32 : n74280;
  assign n74282 = pi18 ? n32 : n74281;
  assign n74283 = pi17 ? n32 : n74282;
  assign n74284 = pi16 ? n32 : n74283;
  assign n74285 = pi20 ? n48254 : n67195;
  assign n74286 = pi19 ? n32 : n74285;
  assign n74287 = pi18 ? n32 : n74286;
  assign n74288 = pi17 ? n32 : n74287;
  assign n74289 = pi16 ? n32 : n74288;
  assign n74290 = pi15 ? n74284 : n74289;
  assign n74291 = pi21 ? n46060 : n33792;
  assign n74292 = pi22 ? n63921 : n316;
  assign n74293 = pi21 ? n74292 : n54546;
  assign n74294 = pi20 ? n74291 : n74293;
  assign n74295 = pi19 ? n32 : n74294;
  assign n74296 = pi18 ? n32 : n74295;
  assign n74297 = pi17 ? n32 : n74296;
  assign n74298 = pi16 ? n32 : n74297;
  assign n74299 = pi23 ? n33792 : n56458;
  assign n74300 = pi22 ? n32 : n74299;
  assign n74301 = pi21 ? n74300 : n33792;
  assign n74302 = pi20 ? n74301 : n73784;
  assign n74303 = pi19 ? n32 : n74302;
  assign n74304 = pi18 ? n32 : n74303;
  assign n74305 = pi17 ? n32 : n74304;
  assign n74306 = pi16 ? n32 : n74305;
  assign n74307 = pi15 ? n74298 : n74306;
  assign n74308 = pi14 ? n74290 : n74307;
  assign n74309 = pi13 ? n74045 : n74308;
  assign n74310 = pi12 ? n74277 : n74309;
  assign n74311 = pi23 ? n20564 : n62332;
  assign n74312 = pi22 ? n32 : n74311;
  assign n74313 = pi21 ? n74312 : n36781;
  assign n74314 = pi22 ? n16717 : n14626;
  assign n74315 = pi21 ? n74314 : n2637;
  assign n74316 = pi20 ? n74313 : n74315;
  assign n74317 = pi19 ? n32 : n74316;
  assign n74318 = pi18 ? n32 : n74317;
  assign n74319 = pi17 ? n32 : n74318;
  assign n74320 = pi16 ? n32 : n74319;
  assign n74321 = pi21 ? n39394 : n36781;
  assign n74322 = pi22 ? n73552 : n685;
  assign n74323 = pi21 ? n74322 : n59357;
  assign n74324 = pi20 ? n74321 : n74323;
  assign n74325 = pi19 ? n32 : n74324;
  assign n74326 = pi18 ? n32 : n74325;
  assign n74327 = pi17 ? n32 : n74326;
  assign n74328 = pi16 ? n32 : n74327;
  assign n74329 = pi15 ? n74320 : n74328;
  assign n74330 = pi21 ? n28156 : n36798;
  assign n74331 = pi22 ? n73814 : n316;
  assign n74332 = pi21 ? n74331 : n928;
  assign n74333 = pi20 ? n74330 : n74332;
  assign n74334 = pi19 ? n32 : n74333;
  assign n74335 = pi18 ? n32 : n74334;
  assign n74336 = pi17 ? n32 : n74335;
  assign n74337 = pi16 ? n32 : n74336;
  assign n74338 = pi21 ? n72668 : n36798;
  assign n74339 = pi20 ? n74338 : n73824;
  assign n74340 = pi19 ? n32 : n74339;
  assign n74341 = pi18 ? n32 : n74340;
  assign n74342 = pi17 ? n32 : n74341;
  assign n74343 = pi16 ? n32 : n74342;
  assign n74344 = pi15 ? n74337 : n74343;
  assign n74345 = pi14 ? n74329 : n74344;
  assign n74346 = pi21 ? n56529 : n43198;
  assign n74347 = pi20 ? n74346 : n70472;
  assign n74348 = pi19 ? n32 : n74347;
  assign n74349 = pi18 ? n32 : n74348;
  assign n74350 = pi17 ? n32 : n74349;
  assign n74351 = pi16 ? n32 : n74350;
  assign n74352 = pi22 ? n32 : n41481;
  assign n74353 = pi21 ? n74352 : n43198;
  assign n74354 = pi20 ? n74353 : n70483;
  assign n74355 = pi19 ? n32 : n74354;
  assign n74356 = pi18 ? n32 : n74355;
  assign n74357 = pi17 ? n32 : n74356;
  assign n74358 = pi16 ? n32 : n74357;
  assign n74359 = pi15 ? n74351 : n74358;
  assign n74360 = pi21 ? n64224 : n14626;
  assign n74361 = pi20 ? n74360 : n70495;
  assign n74362 = pi19 ? n32 : n74361;
  assign n74363 = pi18 ? n32 : n74362;
  assign n74364 = pi17 ? n32 : n74363;
  assign n74365 = pi16 ? n32 : n74364;
  assign n74366 = pi22 ? n32 : n70123;
  assign n74367 = pi21 ? n74366 : n14626;
  assign n74368 = pi20 ? n74367 : n59635;
  assign n74369 = pi19 ? n32 : n74368;
  assign n74370 = pi18 ? n32 : n74369;
  assign n74371 = pi17 ? n32 : n74370;
  assign n74372 = pi16 ? n32 : n74371;
  assign n74373 = pi15 ? n74365 : n74372;
  assign n74374 = pi14 ? n74359 : n74373;
  assign n74375 = pi13 ? n74345 : n74374;
  assign n74376 = pi22 ? n30115 : n42109;
  assign n74377 = pi21 ? n74376 : n14626;
  assign n74378 = pi20 ? n74377 : n7724;
  assign n74379 = pi19 ? n32 : n74378;
  assign n74380 = pi18 ? n32 : n74379;
  assign n74381 = pi17 ? n32 : n74380;
  assign n74382 = pi16 ? n32 : n74381;
  assign n74383 = pi24 ? n30868 : n36781;
  assign n74384 = pi23 ? n74383 : n33792;
  assign n74385 = pi22 ? n30115 : n74384;
  assign n74386 = pi21 ? n74385 : n13481;
  assign n74387 = pi20 ? n74386 : n3210;
  assign n74388 = pi19 ? n32 : n74387;
  assign n74389 = pi18 ? n32 : n74388;
  assign n74390 = pi17 ? n32 : n74389;
  assign n74391 = pi16 ? n32 : n74390;
  assign n74392 = pi15 ? n74382 : n74391;
  assign n74393 = pi24 ? n335 : n36659;
  assign n74394 = pi23 ? n62832 : n74393;
  assign n74395 = pi22 ? n46165 : n74394;
  assign n74396 = pi21 ? n74395 : n59691;
  assign n74397 = pi20 ? n74396 : n60045;
  assign n74398 = pi19 ? n32 : n74397;
  assign n74399 = pi18 ? n32 : n74398;
  assign n74400 = pi17 ? n32 : n74399;
  assign n74401 = pi16 ? n32 : n74400;
  assign n74402 = pi22 ? n46165 : n36659;
  assign n74403 = pi21 ? n74402 : n63771;
  assign n74404 = pi20 ? n74403 : n37640;
  assign n74405 = pi19 ? n32 : n74404;
  assign n74406 = pi18 ? n32 : n74405;
  assign n74407 = pi17 ? n32 : n74406;
  assign n74408 = pi16 ? n32 : n74407;
  assign n74409 = pi15 ? n74401 : n74408;
  assign n74410 = pi14 ? n74392 : n74409;
  assign n74411 = pi22 ? n45516 : n69207;
  assign n74412 = pi21 ? n74411 : n59595;
  assign n74413 = pi20 ? n74412 : n32;
  assign n74414 = pi19 ? n32 : n74413;
  assign n74415 = pi18 ? n32 : n74414;
  assign n74416 = pi17 ? n32 : n74415;
  assign n74417 = pi16 ? n32 : n74416;
  assign n74418 = pi23 ? n4882 : n233;
  assign n74419 = pi22 ? n74418 : n51564;
  assign n74420 = pi21 ? n74158 : n74419;
  assign n74421 = pi20 ? n74420 : n32;
  assign n74422 = pi19 ? n32 : n74421;
  assign n74423 = pi18 ? n32 : n74422;
  assign n74424 = pi17 ? n32 : n74423;
  assign n74425 = pi16 ? n32 : n74424;
  assign n74426 = pi15 ? n74417 : n74425;
  assign n74427 = pi22 ? n46757 : n67348;
  assign n74428 = pi21 ? n74427 : n57746;
  assign n74429 = pi20 ? n74428 : n32;
  assign n74430 = pi19 ? n32 : n74429;
  assign n74431 = pi18 ? n32 : n74430;
  assign n74432 = pi17 ? n32 : n74431;
  assign n74433 = pi16 ? n32 : n74432;
  assign n74434 = pi22 ? n45634 : n63717;
  assign n74435 = pi21 ? n74434 : n60421;
  assign n74436 = pi20 ? n74435 : n32;
  assign n74437 = pi19 ? n32 : n74436;
  assign n74438 = pi18 ? n32 : n74437;
  assign n74439 = pi17 ? n32 : n74438;
  assign n74440 = pi16 ? n32 : n74439;
  assign n74441 = pi15 ? n74433 : n74440;
  assign n74442 = pi14 ? n74426 : n74441;
  assign n74443 = pi13 ? n74410 : n74442;
  assign n74444 = pi12 ? n74375 : n74443;
  assign n74445 = pi11 ? n74310 : n74444;
  assign n74446 = pi23 ? n51564 : n14627;
  assign n74447 = pi22 ? n45634 : n74446;
  assign n74448 = pi21 ? n74447 : n60421;
  assign n74449 = pi20 ? n74448 : n32;
  assign n74450 = pi19 ? n32 : n74449;
  assign n74451 = pi18 ? n32 : n74450;
  assign n74452 = pi17 ? n32 : n74451;
  assign n74453 = pi16 ? n32 : n74452;
  assign n74454 = pi22 ? n32 : n67362;
  assign n74455 = pi21 ? n74454 : n55560;
  assign n74456 = pi20 ? n74455 : n32;
  assign n74457 = pi19 ? n32 : n74456;
  assign n74458 = pi18 ? n32 : n74457;
  assign n74459 = pi17 ? n32 : n74458;
  assign n74460 = pi16 ? n32 : n74459;
  assign n74461 = pi15 ? n74453 : n74460;
  assign n74462 = pi22 ? n32 : n73958;
  assign n74463 = pi21 ? n74462 : n1009;
  assign n74464 = pi20 ? n74463 : n32;
  assign n74465 = pi19 ? n32 : n74464;
  assign n74466 = pi18 ? n32 : n74465;
  assign n74467 = pi17 ? n32 : n74466;
  assign n74468 = pi16 ? n32 : n74467;
  assign n74469 = pi22 ? n32 : n74206;
  assign n74470 = pi21 ? n74469 : n32;
  assign n74471 = pi20 ? n74470 : n32;
  assign n74472 = pi19 ? n32 : n74471;
  assign n74473 = pi18 ? n32 : n74472;
  assign n74474 = pi17 ? n32 : n74473;
  assign n74475 = pi16 ? n32 : n74474;
  assign n74476 = pi15 ? n74468 : n74475;
  assign n74477 = pi14 ? n74461 : n74476;
  assign n74478 = pi22 ? n32 : n73977;
  assign n74479 = pi21 ? n74478 : n32;
  assign n74480 = pi20 ? n74479 : n32;
  assign n74481 = pi19 ? n32 : n74480;
  assign n74482 = pi18 ? n32 : n74481;
  assign n74483 = pi17 ? n32 : n74482;
  assign n74484 = pi16 ? n32 : n74483;
  assign n74485 = pi22 ? n32 : n53982;
  assign n74486 = pi21 ? n74485 : n32;
  assign n74487 = pi20 ? n74486 : n32;
  assign n74488 = pi19 ? n32 : n74487;
  assign n74489 = pi18 ? n32 : n74488;
  assign n74490 = pi17 ? n32 : n74489;
  assign n74491 = pi16 ? n32 : n74490;
  assign n74492 = pi15 ? n74484 : n74491;
  assign n74493 = pi22 ? n32 : n14363;
  assign n74494 = pi21 ? n74493 : n32;
  assign n74495 = pi20 ? n74494 : n32;
  assign n74496 = pi19 ? n32 : n74495;
  assign n74497 = pi18 ? n32 : n74496;
  assign n74498 = pi17 ? n32 : n74497;
  assign n74499 = pi16 ? n32 : n74498;
  assign n74500 = pi15 ? n74499 : n32;
  assign n74501 = pi14 ? n74492 : n74500;
  assign n74502 = pi13 ? n74477 : n74501;
  assign n74503 = pi12 ? n74502 : n32;
  assign n74504 = pi11 ? n74503 : n32;
  assign n74505 = pi10 ? n74445 : n74504;
  assign n74506 = pi09 ? n74263 : n74505;
  assign n74507 = pi20 ? n38997 : n61008;
  assign n74508 = pi19 ? n32 : n74507;
  assign n74509 = pi18 ? n32 : n74508;
  assign n74510 = pi17 ? n32 : n74509;
  assign n74511 = pi16 ? n32 : n74510;
  assign n74512 = pi14 ? n74252 : n74511;
  assign n74513 = pi13 ? n32 : n74512;
  assign n74514 = pi12 ? n32 : n74513;
  assign n74515 = pi11 ? n32 : n74514;
  assign n74516 = pi10 ? n32 : n74515;
  assign n74517 = pi15 ? n74511 : n74017;
  assign n74518 = pi20 ? n37333 : n1619;
  assign n74519 = pi19 ? n32 : n74518;
  assign n74520 = pi18 ? n32 : n74519;
  assign n74521 = pi17 ? n32 : n74520;
  assign n74522 = pi16 ? n32 : n74521;
  assign n74523 = pi14 ? n74517 : n74522;
  assign n74524 = pi13 ? n74523 : n74522;
  assign n74525 = pi20 ? n45502 : n1619;
  assign n74526 = pi19 ? n32 : n74525;
  assign n74527 = pi18 ? n32 : n74526;
  assign n74528 = pi17 ? n32 : n74527;
  assign n74529 = pi16 ? n32 : n74528;
  assign n74530 = pi15 ? n74522 : n74274;
  assign n74531 = pi14 ? n74529 : n74530;
  assign n74532 = pi20 ? n38376 : n74279;
  assign n74533 = pi19 ? n32 : n74532;
  assign n74534 = pi18 ? n32 : n74533;
  assign n74535 = pi17 ? n32 : n74534;
  assign n74536 = pi16 ? n32 : n74535;
  assign n74537 = pi20 ? n45599 : n67195;
  assign n74538 = pi19 ? n32 : n74537;
  assign n74539 = pi18 ? n32 : n74538;
  assign n74540 = pi17 ? n32 : n74539;
  assign n74541 = pi16 ? n32 : n74540;
  assign n74542 = pi15 ? n74536 : n74541;
  assign n74543 = pi21 ? n45598 : n33792;
  assign n74544 = pi21 ? n64858 : n54546;
  assign n74545 = pi20 ? n74543 : n74544;
  assign n74546 = pi19 ? n32 : n74545;
  assign n74547 = pi18 ? n32 : n74546;
  assign n74548 = pi17 ? n32 : n74547;
  assign n74549 = pi16 ? n32 : n74548;
  assign n74550 = pi21 ? n39394 : n33792;
  assign n74551 = pi20 ? n74550 : n73784;
  assign n74552 = pi19 ? n32 : n74551;
  assign n74553 = pi18 ? n32 : n74552;
  assign n74554 = pi17 ? n32 : n74553;
  assign n74555 = pi16 ? n32 : n74554;
  assign n74556 = pi15 ? n74549 : n74555;
  assign n74557 = pi14 ? n74542 : n74556;
  assign n74558 = pi13 ? n74531 : n74557;
  assign n74559 = pi12 ? n74524 : n74558;
  assign n74560 = pi22 ? n59525 : n14626;
  assign n74561 = pi21 ? n74560 : n2637;
  assign n74562 = pi20 ? n74321 : n74561;
  assign n74563 = pi19 ? n32 : n74562;
  assign n74564 = pi18 ? n32 : n74563;
  assign n74565 = pi17 ? n32 : n74564;
  assign n74566 = pi16 ? n32 : n74565;
  assign n74567 = pi15 ? n74566 : n74328;
  assign n74568 = pi21 ? n39394 : n36798;
  assign n74569 = pi20 ? n74568 : n74332;
  assign n74570 = pi19 ? n32 : n74569;
  assign n74571 = pi18 ? n32 : n74570;
  assign n74572 = pi17 ? n32 : n74571;
  assign n74573 = pi16 ? n32 : n74572;
  assign n74574 = pi21 ? n73560 : n1009;
  assign n74575 = pi20 ? n74338 : n74574;
  assign n74576 = pi19 ? n32 : n74575;
  assign n74577 = pi18 ? n32 : n74576;
  assign n74578 = pi17 ? n32 : n74577;
  assign n74579 = pi16 ? n32 : n74578;
  assign n74580 = pi15 ? n74573 : n74579;
  assign n74581 = pi14 ? n74567 : n74580;
  assign n74582 = pi20 ? n74353 : n70472;
  assign n74583 = pi19 ? n32 : n74582;
  assign n74584 = pi18 ? n32 : n74583;
  assign n74585 = pi17 ? n32 : n74584;
  assign n74586 = pi16 ? n32 : n74585;
  assign n74587 = pi15 ? n74586 : n74358;
  assign n74588 = pi23 ? n37273 : n30868;
  assign n74589 = pi22 ? n32 : n74588;
  assign n74590 = pi21 ? n74589 : n14626;
  assign n74591 = pi20 ? n74590 : n70495;
  assign n74592 = pi19 ? n32 : n74591;
  assign n74593 = pi18 ? n32 : n74592;
  assign n74594 = pi17 ? n32 : n74593;
  assign n74595 = pi16 ? n32 : n74594;
  assign n74596 = pi22 ? n32 : n72436;
  assign n74597 = pi21 ? n74596 : n14626;
  assign n74598 = pi20 ? n74597 : n59635;
  assign n74599 = pi19 ? n32 : n74598;
  assign n74600 = pi18 ? n32 : n74599;
  assign n74601 = pi17 ? n32 : n74600;
  assign n74602 = pi16 ? n32 : n74601;
  assign n74603 = pi15 ? n74595 : n74602;
  assign n74604 = pi14 ? n74587 : n74603;
  assign n74605 = pi13 ? n74581 : n74604;
  assign n74606 = pi21 ? n49721 : n14626;
  assign n74607 = pi20 ? n74606 : n7724;
  assign n74608 = pi19 ? n32 : n74607;
  assign n74609 = pi18 ? n32 : n74608;
  assign n74610 = pi17 ? n32 : n74609;
  assign n74611 = pi16 ? n32 : n74610;
  assign n74612 = pi24 ? n36659 : n335;
  assign n74613 = pi23 ? n32 : n74612;
  assign n74614 = pi22 ? n32 : n74613;
  assign n74615 = pi21 ? n74614 : n13481;
  assign n74616 = pi20 ? n74615 : n3210;
  assign n74617 = pi19 ? n32 : n74616;
  assign n74618 = pi18 ? n32 : n74617;
  assign n74619 = pi17 ? n32 : n74618;
  assign n74620 = pi16 ? n32 : n74619;
  assign n74621 = pi15 ? n74611 : n74620;
  assign n74622 = pi24 ? n33792 : n32;
  assign n74623 = pi23 ? n74622 : n74393;
  assign n74624 = pi22 ? n32 : n74623;
  assign n74625 = pi21 ? n74624 : n59691;
  assign n74626 = pi20 ? n74625 : n60045;
  assign n74627 = pi19 ? n32 : n74626;
  assign n74628 = pi18 ? n32 : n74627;
  assign n74629 = pi17 ? n32 : n74628;
  assign n74630 = pi16 ? n32 : n74629;
  assign n74631 = pi23 ? n36782 : n363;
  assign n74632 = pi22 ? n32 : n74631;
  assign n74633 = pi21 ? n74632 : n63771;
  assign n74634 = pi20 ? n74633 : n37640;
  assign n74635 = pi19 ? n32 : n74634;
  assign n74636 = pi18 ? n32 : n74635;
  assign n74637 = pi17 ? n32 : n74636;
  assign n74638 = pi16 ? n32 : n74637;
  assign n74639 = pi15 ? n74630 : n74638;
  assign n74640 = pi14 ? n74621 : n74639;
  assign n74641 = pi23 ? n56079 : n36781;
  assign n74642 = pi22 ? n32 : n74641;
  assign n74643 = pi21 ? n74642 : n59595;
  assign n74644 = pi20 ? n74643 : n32;
  assign n74645 = pi19 ? n32 : n74644;
  assign n74646 = pi18 ? n32 : n74645;
  assign n74647 = pi17 ? n32 : n74646;
  assign n74648 = pi16 ? n32 : n74647;
  assign n74649 = pi22 ? n32 : n57782;
  assign n74650 = pi23 ? n60075 : n233;
  assign n74651 = pi22 ? n74650 : n51564;
  assign n74652 = pi21 ? n74649 : n74651;
  assign n74653 = pi20 ? n74652 : n32;
  assign n74654 = pi19 ? n32 : n74653;
  assign n74655 = pi18 ? n32 : n74654;
  assign n74656 = pi17 ? n32 : n74655;
  assign n74657 = pi16 ? n32 : n74656;
  assign n74658 = pi15 ? n74648 : n74657;
  assign n74659 = pi24 ? n36781 : n32;
  assign n74660 = pi23 ? n74659 : n43198;
  assign n74661 = pi22 ? n32 : n74660;
  assign n74662 = pi21 ? n74661 : n57746;
  assign n74663 = pi20 ? n74662 : n32;
  assign n74664 = pi19 ? n32 : n74663;
  assign n74665 = pi18 ? n32 : n74664;
  assign n74666 = pi17 ? n32 : n74665;
  assign n74667 = pi16 ? n32 : n74666;
  assign n74668 = pi21 ? n50786 : n60421;
  assign n74669 = pi20 ? n74668 : n32;
  assign n74670 = pi19 ? n32 : n74669;
  assign n74671 = pi18 ? n32 : n74670;
  assign n74672 = pi17 ? n32 : n74671;
  assign n74673 = pi16 ? n32 : n74672;
  assign n74674 = pi15 ? n74667 : n74673;
  assign n74675 = pi14 ? n74658 : n74674;
  assign n74676 = pi13 ? n74640 : n74675;
  assign n74677 = pi12 ? n74605 : n74676;
  assign n74678 = pi11 ? n74559 : n74677;
  assign n74679 = pi22 ? n32 : n72270;
  assign n74680 = pi21 ? n74679 : n60421;
  assign n74681 = pi20 ? n74680 : n32;
  assign n74682 = pi19 ? n32 : n74681;
  assign n74683 = pi18 ? n32 : n74682;
  assign n74684 = pi17 ? n32 : n74683;
  assign n74685 = pi16 ? n32 : n74684;
  assign n74686 = pi21 ? n74679 : n55560;
  assign n74687 = pi20 ? n74686 : n32;
  assign n74688 = pi19 ? n32 : n74687;
  assign n74689 = pi18 ? n32 : n74688;
  assign n74690 = pi17 ? n32 : n74689;
  assign n74691 = pi16 ? n32 : n74690;
  assign n74692 = pi15 ? n74685 : n74691;
  assign n74693 = pi21 ? n74462 : n20952;
  assign n74694 = pi20 ? n74693 : n32;
  assign n74695 = pi19 ? n32 : n74694;
  assign n74696 = pi18 ? n32 : n74695;
  assign n74697 = pi17 ? n32 : n74696;
  assign n74698 = pi16 ? n32 : n74697;
  assign n74699 = pi21 ? n74462 : n32;
  assign n74700 = pi20 ? n74699 : n32;
  assign n74701 = pi19 ? n32 : n74700;
  assign n74702 = pi18 ? n32 : n74701;
  assign n74703 = pi17 ? n32 : n74702;
  assign n74704 = pi16 ? n32 : n74703;
  assign n74705 = pi15 ? n74698 : n74704;
  assign n74706 = pi14 ? n74692 : n74705;
  assign n74707 = pi22 ? n32 : n71924;
  assign n74708 = pi21 ? n74707 : n32;
  assign n74709 = pi20 ? n74708 : n32;
  assign n74710 = pi19 ? n32 : n74709;
  assign n74711 = pi18 ? n32 : n74710;
  assign n74712 = pi17 ? n32 : n74711;
  assign n74713 = pi16 ? n32 : n74712;
  assign n74714 = pi15 ? n74713 : n32;
  assign n74715 = pi14 ? n74714 : n32;
  assign n74716 = pi13 ? n74706 : n74715;
  assign n74717 = pi12 ? n74716 : n32;
  assign n74718 = pi11 ? n74717 : n32;
  assign n74719 = pi10 ? n74678 : n74718;
  assign n74720 = pi09 ? n74516 : n74719;
  assign n74721 = pi08 ? n74506 : n74720;
  assign n74722 = pi20 ? n37955 : n74246;
  assign n74723 = pi19 ? n32 : n74722;
  assign n74724 = pi18 ? n32 : n74723;
  assign n74725 = pi17 ? n32 : n74724;
  assign n74726 = pi16 ? n32 : n74725;
  assign n74727 = pi15 ? n32 : n74726;
  assign n74728 = pi20 ? n37955 : n61008;
  assign n74729 = pi19 ? n32 : n74728;
  assign n74730 = pi18 ? n32 : n74729;
  assign n74731 = pi17 ? n32 : n74730;
  assign n74732 = pi16 ? n32 : n74731;
  assign n74733 = pi14 ? n74727 : n74732;
  assign n74734 = pi13 ? n32 : n74733;
  assign n74735 = pi12 ? n32 : n74734;
  assign n74736 = pi11 ? n32 : n74735;
  assign n74737 = pi10 ? n32 : n74736;
  assign n74738 = pi20 ? n37320 : n1619;
  assign n74739 = pi19 ? n32 : n74738;
  assign n74740 = pi18 ? n32 : n74739;
  assign n74741 = pi17 ? n32 : n74740;
  assign n74742 = pi16 ? n32 : n74741;
  assign n74743 = pi15 ? n74742 : n74522;
  assign n74744 = pi14 ? n74517 : n74743;
  assign n74745 = pi20 ? n37320 : n66577;
  assign n74746 = pi19 ? n32 : n74745;
  assign n74747 = pi18 ? n32 : n74746;
  assign n74748 = pi17 ? n32 : n74747;
  assign n74749 = pi16 ? n32 : n74748;
  assign n74750 = pi15 ? n74742 : n74749;
  assign n74751 = pi14 ? n74522 : n74750;
  assign n74752 = pi13 ? n74744 : n74751;
  assign n74753 = pi20 ? n47192 : n1619;
  assign n74754 = pi19 ? n32 : n74753;
  assign n74755 = pi18 ? n32 : n74754;
  assign n74756 = pi17 ? n32 : n74755;
  assign n74757 = pi16 ? n32 : n74756;
  assign n74758 = pi14 ? n74757 : n74743;
  assign n74759 = pi24 ? n20563 : n14626;
  assign n74760 = pi23 ? n74759 : n14626;
  assign n74761 = pi22 ? n74760 : n14626;
  assign n74762 = pi21 ? n74761 : n64842;
  assign n74763 = pi20 ? n37333 : n74762;
  assign n74764 = pi19 ? n32 : n74763;
  assign n74765 = pi18 ? n32 : n74764;
  assign n74766 = pi17 ? n32 : n74765;
  assign n74767 = pi16 ? n32 : n74766;
  assign n74768 = pi20 ? n45502 : n68542;
  assign n74769 = pi19 ? n32 : n74768;
  assign n74770 = pi18 ? n32 : n74769;
  assign n74771 = pi17 ? n32 : n74770;
  assign n74772 = pi16 ? n32 : n74771;
  assign n74773 = pi15 ? n74767 : n74772;
  assign n74774 = pi21 ? n37332 : n33792;
  assign n74775 = pi21 ? n57350 : n3523;
  assign n74776 = pi20 ? n74774 : n74775;
  assign n74777 = pi19 ? n32 : n74776;
  assign n74778 = pi18 ? n32 : n74777;
  assign n74779 = pi17 ? n32 : n74778;
  assign n74780 = pi16 ? n32 : n74779;
  assign n74781 = pi21 ? n67642 : n33095;
  assign n74782 = pi20 ? n60777 : n74781;
  assign n74783 = pi19 ? n32 : n74782;
  assign n74784 = pi18 ? n32 : n74783;
  assign n74785 = pi17 ? n32 : n74784;
  assign n74786 = pi16 ? n32 : n74785;
  assign n74787 = pi15 ? n74780 : n74786;
  assign n74788 = pi14 ? n74773 : n74787;
  assign n74789 = pi13 ? n74758 : n74788;
  assign n74790 = pi12 ? n74752 : n74789;
  assign n74791 = pi21 ? n37332 : n36781;
  assign n74792 = pi20 ? n74791 : n71642;
  assign n74793 = pi19 ? n32 : n74792;
  assign n74794 = pi18 ? n32 : n74793;
  assign n74795 = pi17 ? n32 : n74794;
  assign n74796 = pi16 ? n32 : n74795;
  assign n74797 = pi21 ? n74322 : n928;
  assign n74798 = pi20 ? n74791 : n74797;
  assign n74799 = pi19 ? n32 : n74798;
  assign n74800 = pi18 ? n32 : n74799;
  assign n74801 = pi17 ? n32 : n74800;
  assign n74802 = pi16 ? n32 : n74801;
  assign n74803 = pi15 ? n74796 : n74802;
  assign n74804 = pi21 ? n37332 : n36798;
  assign n74805 = pi23 ? n8133 : n316;
  assign n74806 = pi22 ? n74805 : n316;
  assign n74807 = pi21 ? n74806 : n928;
  assign n74808 = pi20 ? n74804 : n74807;
  assign n74809 = pi19 ? n32 : n74808;
  assign n74810 = pi18 ? n32 : n74809;
  assign n74811 = pi17 ? n32 : n74810;
  assign n74812 = pi16 ? n32 : n74811;
  assign n74813 = pi20 ? n74804 : n74574;
  assign n74814 = pi19 ? n32 : n74813;
  assign n74815 = pi18 ? n32 : n74814;
  assign n74816 = pi17 ? n32 : n74815;
  assign n74817 = pi16 ? n32 : n74816;
  assign n74818 = pi15 ? n74812 : n74817;
  assign n74819 = pi14 ? n74803 : n74818;
  assign n74820 = pi21 ? n38375 : n43198;
  assign n74821 = pi20 ? n74820 : n67702;
  assign n74822 = pi19 ? n32 : n74821;
  assign n74823 = pi18 ? n32 : n74822;
  assign n74824 = pi17 ? n32 : n74823;
  assign n74825 = pi16 ? n32 : n74824;
  assign n74826 = pi20 ? n74820 : n67719;
  assign n74827 = pi19 ? n32 : n74826;
  assign n74828 = pi18 ? n32 : n74827;
  assign n74829 = pi17 ? n32 : n74828;
  assign n74830 = pi16 ? n32 : n74829;
  assign n74831 = pi15 ? n74825 : n74830;
  assign n74832 = pi21 ? n45598 : n14626;
  assign n74833 = pi20 ? n74832 : n6935;
  assign n74834 = pi19 ? n32 : n74833;
  assign n74835 = pi18 ? n32 : n74834;
  assign n74836 = pi17 ? n32 : n74835;
  assign n74837 = pi16 ? n32 : n74836;
  assign n74838 = pi21 ? n55516 : n14626;
  assign n74839 = pi20 ? n74838 : n59649;
  assign n74840 = pi19 ? n32 : n74839;
  assign n74841 = pi18 ? n32 : n74840;
  assign n74842 = pi17 ? n32 : n74841;
  assign n74843 = pi16 ? n32 : n74842;
  assign n74844 = pi15 ? n74837 : n74843;
  assign n74845 = pi14 ? n74831 : n74844;
  assign n74846 = pi13 ? n74819 : n74845;
  assign n74847 = pi21 ? n49721 : n57746;
  assign n74848 = pi20 ? n74847 : n7724;
  assign n74849 = pi19 ? n32 : n74848;
  assign n74850 = pi18 ? n32 : n74849;
  assign n74851 = pi17 ? n32 : n74850;
  assign n74852 = pi16 ? n32 : n74851;
  assign n74853 = pi21 ? n51755 : n13481;
  assign n74854 = pi20 ? n74853 : n3210;
  assign n74855 = pi19 ? n32 : n74854;
  assign n74856 = pi18 ? n32 : n74855;
  assign n74857 = pi17 ? n32 : n74856;
  assign n74858 = pi16 ? n32 : n74857;
  assign n74859 = pi15 ? n74852 : n74858;
  assign n74860 = pi21 ? n51755 : n63771;
  assign n74861 = pi20 ? n74860 : n60045;
  assign n74862 = pi19 ? n32 : n74861;
  assign n74863 = pi18 ? n32 : n74862;
  assign n74864 = pi17 ? n32 : n74863;
  assign n74865 = pi16 ? n32 : n74864;
  assign n74866 = pi21 ? n73357 : n56760;
  assign n74867 = pi20 ? n74866 : n32;
  assign n74868 = pi19 ? n32 : n74867;
  assign n74869 = pi18 ? n32 : n74868;
  assign n74870 = pi17 ? n32 : n74869;
  assign n74871 = pi16 ? n32 : n74870;
  assign n74872 = pi15 ? n74865 : n74871;
  assign n74873 = pi14 ? n74859 : n74872;
  assign n74874 = pi21 ? n73357 : n57746;
  assign n74875 = pi20 ? n74874 : n32;
  assign n74876 = pi19 ? n32 : n74875;
  assign n74877 = pi18 ? n32 : n74876;
  assign n74878 = pi17 ? n32 : n74877;
  assign n74879 = pi16 ? n32 : n74878;
  assign n74880 = pi22 ? n67362 : n13481;
  assign n74881 = pi21 ? n46772 : n74880;
  assign n74882 = pi20 ? n74881 : n32;
  assign n74883 = pi19 ? n32 : n74882;
  assign n74884 = pi18 ? n32 : n74883;
  assign n74885 = pi17 ? n32 : n74884;
  assign n74886 = pi16 ? n32 : n74885;
  assign n74887 = pi15 ? n74879 : n74886;
  assign n74888 = pi21 ? n46276 : n60795;
  assign n74889 = pi20 ? n74888 : n32;
  assign n74890 = pi19 ? n32 : n74889;
  assign n74891 = pi18 ? n32 : n74890;
  assign n74892 = pi17 ? n32 : n74891;
  assign n74893 = pi16 ? n32 : n74892;
  assign n74894 = pi21 ? n46790 : n60421;
  assign n74895 = pi20 ? n74894 : n32;
  assign n74896 = pi19 ? n32 : n74895;
  assign n74897 = pi18 ? n32 : n74896;
  assign n74898 = pi17 ? n32 : n74897;
  assign n74899 = pi16 ? n32 : n74898;
  assign n74900 = pi15 ? n74893 : n74899;
  assign n74901 = pi14 ? n74887 : n74900;
  assign n74902 = pi13 ? n74873 : n74901;
  assign n74903 = pi12 ? n74846 : n74902;
  assign n74904 = pi11 ? n74790 : n74903;
  assign n74905 = pi23 ? n32 : n14626;
  assign n74906 = pi22 ? n32 : n74905;
  assign n74907 = pi22 ? n62473 : n32;
  assign n74908 = pi21 ? n74906 : n74907;
  assign n74909 = pi20 ? n74908 : n32;
  assign n74910 = pi19 ? n32 : n74909;
  assign n74911 = pi18 ? n32 : n74910;
  assign n74912 = pi17 ? n32 : n74911;
  assign n74913 = pi16 ? n32 : n74912;
  assign n74914 = pi21 ? n74906 : n53983;
  assign n74915 = pi20 ? n74914 : n32;
  assign n74916 = pi19 ? n32 : n74915;
  assign n74917 = pi18 ? n32 : n74916;
  assign n74918 = pi17 ? n32 : n74917;
  assign n74919 = pi16 ? n32 : n74918;
  assign n74920 = pi15 ? n74913 : n74919;
  assign n74921 = pi21 ? n73123 : n1009;
  assign n74922 = pi20 ? n74921 : n32;
  assign n74923 = pi19 ? n32 : n74922;
  assign n74924 = pi18 ? n32 : n74923;
  assign n74925 = pi17 ? n32 : n74924;
  assign n74926 = pi16 ? n32 : n74925;
  assign n74927 = pi21 ? n73123 : n32;
  assign n74928 = pi20 ? n74927 : n32;
  assign n74929 = pi19 ? n32 : n74928;
  assign n74930 = pi18 ? n32 : n74929;
  assign n74931 = pi17 ? n32 : n74930;
  assign n74932 = pi16 ? n32 : n74931;
  assign n74933 = pi15 ? n74926 : n74932;
  assign n74934 = pi14 ? n74920 : n74933;
  assign n74935 = pi21 ? n69891 : n32;
  assign n74936 = pi20 ? n74935 : n32;
  assign n74937 = pi19 ? n32 : n74936;
  assign n74938 = pi18 ? n32 : n74937;
  assign n74939 = pi17 ? n32 : n74938;
  assign n74940 = pi16 ? n32 : n74939;
  assign n74941 = pi15 ? n74940 : n32;
  assign n74942 = pi14 ? n74941 : n32;
  assign n74943 = pi13 ? n74934 : n74942;
  assign n74944 = pi12 ? n74943 : n32;
  assign n74945 = pi11 ? n74944 : n32;
  assign n74946 = pi10 ? n74904 : n74945;
  assign n74947 = pi09 ? n74737 : n74946;
  assign n74948 = pi15 ? n74732 : n74511;
  assign n74949 = pi20 ? n38997 : n1619;
  assign n74950 = pi19 ? n32 : n74949;
  assign n74951 = pi18 ? n32 : n74950;
  assign n74952 = pi17 ? n32 : n74951;
  assign n74953 = pi16 ? n32 : n74952;
  assign n74954 = pi15 ? n74953 : n74742;
  assign n74955 = pi14 ? n74948 : n74954;
  assign n74956 = pi14 ? n74742 : n74750;
  assign n74957 = pi13 ? n74955 : n74956;
  assign n74958 = pi14 ? n74757 : n74742;
  assign n74959 = pi21 ? n47321 : n33792;
  assign n74960 = pi20 ? n74959 : n74775;
  assign n74961 = pi19 ? n32 : n74960;
  assign n74962 = pi18 ? n32 : n74961;
  assign n74963 = pi17 ? n32 : n74962;
  assign n74964 = pi16 ? n32 : n74963;
  assign n74965 = pi20 ? n59715 : n74781;
  assign n74966 = pi19 ? n32 : n74965;
  assign n74967 = pi18 ? n32 : n74966;
  assign n74968 = pi17 ? n32 : n74967;
  assign n74969 = pi16 ? n32 : n74968;
  assign n74970 = pi15 ? n74964 : n74969;
  assign n74971 = pi14 ? n74773 : n74970;
  assign n74972 = pi13 ? n74958 : n74971;
  assign n74973 = pi12 ? n74957 : n74972;
  assign n74974 = pi21 ? n55516 : n36781;
  assign n74975 = pi20 ? n74974 : n71642;
  assign n74976 = pi19 ? n32 : n74975;
  assign n74977 = pi18 ? n32 : n74976;
  assign n74978 = pi17 ? n32 : n74977;
  assign n74979 = pi16 ? n32 : n74978;
  assign n74980 = pi21 ? n32 : n36781;
  assign n74981 = pi20 ? n74980 : n74797;
  assign n74982 = pi19 ? n32 : n74981;
  assign n74983 = pi18 ? n32 : n74982;
  assign n74984 = pi17 ? n32 : n74983;
  assign n74985 = pi16 ? n32 : n74984;
  assign n74986 = pi15 ? n74979 : n74985;
  assign n74987 = pi21 ? n32 : n36798;
  assign n74988 = pi20 ? n74987 : n74807;
  assign n74989 = pi19 ? n32 : n74988;
  assign n74990 = pi18 ? n32 : n74989;
  assign n74991 = pi17 ? n32 : n74990;
  assign n74992 = pi16 ? n32 : n74991;
  assign n74993 = pi20 ? n74987 : n74574;
  assign n74994 = pi19 ? n32 : n74993;
  assign n74995 = pi18 ? n32 : n74994;
  assign n74996 = pi17 ? n32 : n74995;
  assign n74997 = pi16 ? n32 : n74996;
  assign n74998 = pi15 ? n74992 : n74997;
  assign n74999 = pi14 ? n74986 : n74998;
  assign n75000 = pi21 ? n37332 : n43198;
  assign n75001 = pi20 ? n75000 : n67702;
  assign n75002 = pi19 ? n32 : n75001;
  assign n75003 = pi18 ? n32 : n75002;
  assign n75004 = pi17 ? n32 : n75003;
  assign n75005 = pi16 ? n32 : n75004;
  assign n75006 = pi20 ? n75000 : n67719;
  assign n75007 = pi19 ? n32 : n75006;
  assign n75008 = pi18 ? n32 : n75007;
  assign n75009 = pi17 ? n32 : n75008;
  assign n75010 = pi16 ? n32 : n75009;
  assign n75011 = pi15 ? n75005 : n75010;
  assign n75012 = pi21 ? n47321 : n14626;
  assign n75013 = pi20 ? n75012 : n6935;
  assign n75014 = pi19 ? n32 : n75013;
  assign n75015 = pi18 ? n32 : n75014;
  assign n75016 = pi17 ? n32 : n75015;
  assign n75017 = pi16 ? n32 : n75016;
  assign n75018 = pi20 ? n66541 : n59649;
  assign n75019 = pi19 ? n32 : n75018;
  assign n75020 = pi18 ? n32 : n75019;
  assign n75021 = pi17 ? n32 : n75020;
  assign n75022 = pi16 ? n32 : n75021;
  assign n75023 = pi15 ? n75017 : n75022;
  assign n75024 = pi14 ? n75011 : n75023;
  assign n75025 = pi13 ? n74999 : n75024;
  assign n75026 = pi21 ? n55516 : n57746;
  assign n75027 = pi20 ? n75026 : n7724;
  assign n75028 = pi19 ? n32 : n75027;
  assign n75029 = pi18 ? n32 : n75028;
  assign n75030 = pi17 ? n32 : n75029;
  assign n75031 = pi16 ? n32 : n75030;
  assign n75032 = pi21 ? n46758 : n13481;
  assign n75033 = pi20 ? n75032 : n3210;
  assign n75034 = pi19 ? n32 : n75033;
  assign n75035 = pi18 ? n32 : n75034;
  assign n75036 = pi17 ? n32 : n75035;
  assign n75037 = pi16 ? n32 : n75036;
  assign n75038 = pi15 ? n75031 : n75037;
  assign n75039 = pi23 ? n14626 : n71896;
  assign n75040 = pi22 ? n43198 : n75039;
  assign n75041 = pi21 ? n51755 : n75040;
  assign n75042 = pi20 ? n75041 : n60045;
  assign n75043 = pi19 ? n32 : n75042;
  assign n75044 = pi18 ? n32 : n75043;
  assign n75045 = pi17 ? n32 : n75044;
  assign n75046 = pi16 ? n32 : n75045;
  assign n75047 = pi21 ? n32 : n56760;
  assign n75048 = pi20 ? n75047 : n32;
  assign n75049 = pi19 ? n32 : n75048;
  assign n75050 = pi18 ? n32 : n75049;
  assign n75051 = pi17 ? n32 : n75050;
  assign n75052 = pi16 ? n32 : n75051;
  assign n75053 = pi15 ? n75046 : n75052;
  assign n75054 = pi14 ? n75038 : n75053;
  assign n75055 = pi21 ? n32 : n57746;
  assign n75056 = pi20 ? n75055 : n32;
  assign n75057 = pi19 ? n32 : n75056;
  assign n75058 = pi18 ? n32 : n75057;
  assign n75059 = pi17 ? n32 : n75058;
  assign n75060 = pi16 ? n32 : n75059;
  assign n75061 = pi21 ? n46276 : n74880;
  assign n75062 = pi20 ? n75061 : n32;
  assign n75063 = pi19 ? n32 : n75062;
  assign n75064 = pi18 ? n32 : n75063;
  assign n75065 = pi17 ? n32 : n75064;
  assign n75066 = pi16 ? n32 : n75065;
  assign n75067 = pi15 ? n75060 : n75066;
  assign n75068 = pi23 ? n65601 : n51564;
  assign n75069 = pi22 ? n75068 : n706;
  assign n75070 = pi21 ? n63433 : n75069;
  assign n75071 = pi20 ? n75070 : n32;
  assign n75072 = pi19 ? n32 : n75071;
  assign n75073 = pi18 ? n32 : n75072;
  assign n75074 = pi17 ? n32 : n75073;
  assign n75075 = pi16 ? n32 : n75074;
  assign n75076 = pi22 ? n71897 : n32;
  assign n75077 = pi21 ? n63433 : n75076;
  assign n75078 = pi20 ? n75077 : n32;
  assign n75079 = pi19 ? n32 : n75078;
  assign n75080 = pi18 ? n32 : n75079;
  assign n75081 = pi17 ? n32 : n75080;
  assign n75082 = pi16 ? n32 : n75081;
  assign n75083 = pi15 ? n75075 : n75082;
  assign n75084 = pi14 ? n75067 : n75083;
  assign n75085 = pi13 ? n75054 : n75084;
  assign n75086 = pi12 ? n75025 : n75085;
  assign n75087 = pi11 ? n74973 : n75086;
  assign n75088 = pi23 ? n13481 : n316;
  assign n75089 = pi22 ? n75088 : n32;
  assign n75090 = pi21 ? n71541 : n75089;
  assign n75091 = pi20 ? n75090 : n32;
  assign n75092 = pi19 ? n32 : n75091;
  assign n75093 = pi18 ? n32 : n75092;
  assign n75094 = pi17 ? n32 : n75093;
  assign n75095 = pi16 ? n32 : n75094;
  assign n75096 = pi21 ? n32 : n1009;
  assign n75097 = pi20 ? n75096 : n32;
  assign n75098 = pi19 ? n32 : n75097;
  assign n75099 = pi18 ? n32 : n75098;
  assign n75100 = pi17 ? n32 : n75099;
  assign n75101 = pi16 ? n32 : n75100;
  assign n75102 = pi15 ? n75095 : n75101;
  assign n75103 = pi21 ? n32 : n20952;
  assign n75104 = pi20 ? n75103 : n32;
  assign n75105 = pi19 ? n32 : n75104;
  assign n75106 = pi18 ? n32 : n75105;
  assign n75107 = pi17 ? n32 : n75106;
  assign n75108 = pi16 ? n32 : n75107;
  assign n75109 = pi15 ? n75108 : n32;
  assign n75110 = pi14 ? n75102 : n75109;
  assign n75111 = pi13 ? n75110 : n32;
  assign n75112 = pi12 ? n75111 : n32;
  assign n75113 = pi11 ? n75112 : n32;
  assign n75114 = pi10 ? n75087 : n75113;
  assign n75115 = pi09 ? n74737 : n75114;
  assign n75116 = pi08 ? n74947 : n75115;
  assign n75117 = pi07 ? n74721 : n75116;
  assign n75118 = pi06 ? n74245 : n75117;
  assign n75119 = pi05 ? n73186 : n75118;
  assign n75120 = pi22 ? n39 : n30868;
  assign n75121 = pi21 ? n32 : n75120;
  assign n75122 = pi20 ? n75121 : n13040;
  assign n75123 = pi19 ? n32 : n75122;
  assign n75124 = pi18 ? n32 : n75123;
  assign n75125 = pi17 ? n32 : n75124;
  assign n75126 = pi16 ? n32 : n75125;
  assign n75127 = pi15 ? n32 : n75126;
  assign n75128 = pi22 ? n39 : n33792;
  assign n75129 = pi21 ? n32 : n75128;
  assign n75130 = pi20 ? n75129 : n61008;
  assign n75131 = pi19 ? n32 : n75130;
  assign n75132 = pi18 ? n32 : n75131;
  assign n75133 = pi17 ? n32 : n75132;
  assign n75134 = pi16 ? n32 : n75133;
  assign n75135 = pi22 ? n30115 : n33792;
  assign n75136 = pi21 ? n32 : n75135;
  assign n75137 = pi20 ? n75136 : n61008;
  assign n75138 = pi19 ? n32 : n75137;
  assign n75139 = pi18 ? n32 : n75138;
  assign n75140 = pi17 ? n32 : n75139;
  assign n75141 = pi16 ? n32 : n75140;
  assign n75142 = pi15 ? n75134 : n75141;
  assign n75143 = pi14 ? n75127 : n75142;
  assign n75144 = pi13 ? n32 : n75143;
  assign n75145 = pi12 ? n32 : n75144;
  assign n75146 = pi11 ? n32 : n75145;
  assign n75147 = pi10 ? n32 : n75146;
  assign n75148 = pi20 ? n38997 : n66577;
  assign n75149 = pi19 ? n32 : n75148;
  assign n75150 = pi18 ? n32 : n75149;
  assign n75151 = pi17 ? n32 : n75150;
  assign n75152 = pi16 ? n32 : n75151;
  assign n75153 = pi15 ? n75152 : n74953;
  assign n75154 = pi14 ? n74511 : n75153;
  assign n75155 = pi13 ? n74511 : n75154;
  assign n75156 = pi21 ? n30868 : n1618;
  assign n75157 = pi20 ? n72030 : n75156;
  assign n75158 = pi19 ? n32 : n75157;
  assign n75159 = pi18 ? n32 : n75158;
  assign n75160 = pi17 ? n32 : n75159;
  assign n75161 = pi16 ? n32 : n75160;
  assign n75162 = pi14 ? n74511 : n75161;
  assign n75163 = pi22 ? n65354 : n685;
  assign n75164 = pi21 ? n75163 : n71968;
  assign n75165 = pi20 ? n37320 : n75164;
  assign n75166 = pi19 ? n32 : n75165;
  assign n75167 = pi18 ? n32 : n75166;
  assign n75168 = pi17 ? n32 : n75167;
  assign n75169 = pi16 ? n32 : n75168;
  assign n75170 = pi20 ? n65200 : n69484;
  assign n75171 = pi19 ? n32 : n75170;
  assign n75172 = pi18 ? n32 : n75171;
  assign n75173 = pi17 ? n32 : n75172;
  assign n75174 = pi16 ? n32 : n75173;
  assign n75175 = pi15 ? n75169 : n75174;
  assign n75176 = pi20 ? n62445 : n74775;
  assign n75177 = pi19 ? n32 : n75176;
  assign n75178 = pi18 ? n32 : n75177;
  assign n75179 = pi17 ? n32 : n75178;
  assign n75180 = pi16 ? n32 : n75179;
  assign n75181 = pi22 ? n68564 : n13481;
  assign n75182 = pi21 ? n75181 : n55560;
  assign n75183 = pi20 ? n72113 : n75182;
  assign n75184 = pi19 ? n32 : n75183;
  assign n75185 = pi18 ? n32 : n75184;
  assign n75186 = pi17 ? n32 : n75185;
  assign n75187 = pi16 ? n32 : n75186;
  assign n75188 = pi15 ? n75180 : n75187;
  assign n75189 = pi14 ? n75175 : n75188;
  assign n75190 = pi13 ? n75162 : n75189;
  assign n75191 = pi12 ? n75155 : n75190;
  assign n75192 = pi24 ? n36659 : n14626;
  assign n75193 = pi23 ? n75192 : n14626;
  assign n75194 = pi22 ? n75193 : n685;
  assign n75195 = pi21 ? n75194 : n2637;
  assign n75196 = pi20 ? n72121 : n75195;
  assign n75197 = pi19 ? n32 : n75196;
  assign n75198 = pi18 ? n32 : n75197;
  assign n75199 = pi17 ? n32 : n75198;
  assign n75200 = pi16 ? n32 : n75199;
  assign n75201 = pi21 ? n32 : n61373;
  assign n75202 = pi21 ? n73553 : n928;
  assign n75203 = pi20 ? n75201 : n75202;
  assign n75204 = pi19 ? n32 : n75203;
  assign n75205 = pi18 ? n32 : n75204;
  assign n75206 = pi17 ? n32 : n75205;
  assign n75207 = pi16 ? n32 : n75206;
  assign n75208 = pi15 ? n75200 : n75207;
  assign n75209 = pi22 ? n73276 : n13481;
  assign n75210 = pi21 ? n75209 : n928;
  assign n75211 = pi20 ? n75201 : n75210;
  assign n75212 = pi19 ? n32 : n75211;
  assign n75213 = pi18 ? n32 : n75212;
  assign n75214 = pi17 ? n32 : n75213;
  assign n75215 = pi16 ? n32 : n75214;
  assign n75216 = pi21 ? n32 : n68724;
  assign n75217 = pi23 ? n70599 : n316;
  assign n75218 = pi22 ? n75217 : n13481;
  assign n75219 = pi21 ? n75218 : n1009;
  assign n75220 = pi20 ? n75216 : n75219;
  assign n75221 = pi19 ? n32 : n75220;
  assign n75222 = pi18 ? n32 : n75221;
  assign n75223 = pi17 ? n32 : n75222;
  assign n75224 = pi16 ? n32 : n75223;
  assign n75225 = pi15 ? n75215 : n75224;
  assign n75226 = pi14 ? n75208 : n75225;
  assign n75227 = pi21 ? n32 : n53471;
  assign n75228 = pi20 ? n75227 : n72051;
  assign n75229 = pi19 ? n32 : n75228;
  assign n75230 = pi18 ? n32 : n75229;
  assign n75231 = pi17 ? n32 : n75230;
  assign n75232 = pi16 ? n32 : n75231;
  assign n75233 = pi21 ? n32 : n64961;
  assign n75234 = pi20 ? n75233 : n72062;
  assign n75235 = pi19 ? n32 : n75234;
  assign n75236 = pi18 ? n32 : n75235;
  assign n75237 = pi17 ? n32 : n75236;
  assign n75238 = pi16 ? n32 : n75237;
  assign n75239 = pi15 ? n75232 : n75238;
  assign n75240 = pi22 ? n64325 : n14626;
  assign n75241 = pi21 ? n32 : n75240;
  assign n75242 = pi20 ? n75241 : n59649;
  assign n75243 = pi19 ? n32 : n75242;
  assign n75244 = pi18 ? n32 : n75243;
  assign n75245 = pi17 ? n32 : n75244;
  assign n75246 = pi16 ? n32 : n75245;
  assign n75247 = pi15 ? n75238 : n75246;
  assign n75248 = pi14 ? n75239 : n75247;
  assign n75249 = pi13 ? n75226 : n75248;
  assign n75250 = pi22 ? n72211 : n13481;
  assign n75251 = pi21 ? n32 : n75250;
  assign n75252 = pi20 ? n75251 : n60045;
  assign n75253 = pi19 ? n32 : n75252;
  assign n75254 = pi18 ? n32 : n75253;
  assign n75255 = pi17 ? n32 : n75254;
  assign n75256 = pi16 ? n32 : n75255;
  assign n75257 = pi22 ? n36831 : n13481;
  assign n75258 = pi21 ? n32 : n75257;
  assign n75259 = pi20 ? n75258 : n60045;
  assign n75260 = pi19 ? n32 : n75259;
  assign n75261 = pi18 ? n32 : n75260;
  assign n75262 = pi17 ? n32 : n75261;
  assign n75263 = pi16 ? n32 : n75262;
  assign n75264 = pi15 ? n75256 : n75263;
  assign n75265 = pi22 ? n49843 : n13481;
  assign n75266 = pi21 ? n32 : n75265;
  assign n75267 = pi20 ? n75266 : n60045;
  assign n75268 = pi19 ? n32 : n75267;
  assign n75269 = pi18 ? n32 : n75268;
  assign n75270 = pi17 ? n32 : n75269;
  assign n75271 = pi16 ? n32 : n75270;
  assign n75272 = pi20 ? n75266 : n32;
  assign n75273 = pi19 ? n32 : n75272;
  assign n75274 = pi18 ? n32 : n75273;
  assign n75275 = pi17 ? n32 : n75274;
  assign n75276 = pi16 ? n32 : n75275;
  assign n75277 = pi15 ? n75271 : n75276;
  assign n75278 = pi14 ? n75264 : n75277;
  assign n75279 = pi22 ? n72270 : n13481;
  assign n75280 = pi21 ? n32 : n75279;
  assign n75281 = pi20 ? n75280 : n32;
  assign n75282 = pi19 ? n32 : n75281;
  assign n75283 = pi18 ? n32 : n75282;
  assign n75284 = pi17 ? n32 : n75283;
  assign n75285 = pi16 ? n32 : n75284;
  assign n75286 = pi21 ? n32 : n74880;
  assign n75287 = pi20 ? n75286 : n32;
  assign n75288 = pi19 ? n32 : n75287;
  assign n75289 = pi18 ? n32 : n75288;
  assign n75290 = pi17 ? n32 : n75289;
  assign n75291 = pi16 ? n32 : n75290;
  assign n75292 = pi15 ? n75285 : n75291;
  assign n75293 = pi22 ? n74206 : n706;
  assign n75294 = pi21 ? n32 : n75293;
  assign n75295 = pi20 ? n75294 : n32;
  assign n75296 = pi19 ? n32 : n75295;
  assign n75297 = pi18 ? n32 : n75296;
  assign n75298 = pi17 ? n32 : n75297;
  assign n75299 = pi16 ? n32 : n75298;
  assign n75300 = pi21 ? n32 : n75076;
  assign n75301 = pi20 ? n75300 : n32;
  assign n75302 = pi19 ? n32 : n75301;
  assign n75303 = pi18 ? n32 : n75302;
  assign n75304 = pi17 ? n32 : n75303;
  assign n75305 = pi16 ? n32 : n75304;
  assign n75306 = pi15 ? n75299 : n75305;
  assign n75307 = pi14 ? n75292 : n75306;
  assign n75308 = pi13 ? n75278 : n75307;
  assign n75309 = pi12 ? n75249 : n75308;
  assign n75310 = pi11 ? n75191 : n75309;
  assign n75311 = pi21 ? n32 : n55560;
  assign n75312 = pi20 ? n75311 : n32;
  assign n75313 = pi19 ? n32 : n75312;
  assign n75314 = pi18 ? n32 : n75313;
  assign n75315 = pi17 ? n32 : n75314;
  assign n75316 = pi16 ? n32 : n75315;
  assign n75317 = pi15 ? n75316 : n75108;
  assign n75318 = pi14 ? n75317 : n32;
  assign n75319 = pi13 ? n75318 : n32;
  assign n75320 = pi12 ? n75319 : n32;
  assign n75321 = pi11 ? n75320 : n32;
  assign n75322 = pi10 ? n75310 : n75321;
  assign n75323 = pi09 ? n75147 : n75322;
  assign n75324 = pi20 ? n60055 : n13040;
  assign n75325 = pi19 ? n32 : n75324;
  assign n75326 = pi18 ? n32 : n75325;
  assign n75327 = pi17 ? n32 : n75326;
  assign n75328 = pi16 ? n32 : n75327;
  assign n75329 = pi15 ? n32 : n75328;
  assign n75330 = pi20 ? n70117 : n61008;
  assign n75331 = pi19 ? n32 : n75330;
  assign n75332 = pi18 ? n32 : n75331;
  assign n75333 = pi17 ? n32 : n75332;
  assign n75334 = pi16 ? n32 : n75333;
  assign n75335 = pi15 ? n75141 : n75334;
  assign n75336 = pi14 ? n75329 : n75335;
  assign n75337 = pi13 ? n32 : n75336;
  assign n75338 = pi12 ? n32 : n75337;
  assign n75339 = pi11 ? n32 : n75338;
  assign n75340 = pi10 ? n32 : n75339;
  assign n75341 = pi14 ? n74732 : n74948;
  assign n75342 = pi13 ? n75341 : n75154;
  assign n75343 = pi21 ? n32 : n41459;
  assign n75344 = pi20 ? n75343 : n75156;
  assign n75345 = pi19 ? n32 : n75344;
  assign n75346 = pi18 ? n32 : n75345;
  assign n75347 = pi17 ? n32 : n75346;
  assign n75348 = pi16 ? n32 : n75347;
  assign n75349 = pi15 ? n75161 : n75348;
  assign n75350 = pi14 ? n74511 : n75349;
  assign n75351 = pi24 ? n30868 : n14626;
  assign n75352 = pi23 ? n75351 : n14626;
  assign n75353 = pi22 ? n75352 : n685;
  assign n75354 = pi21 ? n75353 : n71968;
  assign n75355 = pi20 ? n38997 : n75354;
  assign n75356 = pi19 ? n32 : n75355;
  assign n75357 = pi18 ? n32 : n75356;
  assign n75358 = pi17 ? n32 : n75357;
  assign n75359 = pi16 ? n32 : n75358;
  assign n75360 = pi20 ? n72030 : n69484;
  assign n75361 = pi19 ? n32 : n75360;
  assign n75362 = pi18 ? n32 : n75361;
  assign n75363 = pi17 ? n32 : n75362;
  assign n75364 = pi16 ? n32 : n75363;
  assign n75365 = pi15 ? n75359 : n75364;
  assign n75366 = pi21 ? n67642 : n3523;
  assign n75367 = pi20 ? n62445 : n75366;
  assign n75368 = pi19 ? n32 : n75367;
  assign n75369 = pi18 ? n32 : n75368;
  assign n75370 = pi17 ? n32 : n75369;
  assign n75371 = pi16 ? n32 : n75370;
  assign n75372 = pi22 ? n30865 : n36659;
  assign n75373 = pi21 ? n32 : n75372;
  assign n75374 = pi20 ? n75373 : n71995;
  assign n75375 = pi19 ? n32 : n75374;
  assign n75376 = pi18 ? n32 : n75375;
  assign n75377 = pi17 ? n32 : n75376;
  assign n75378 = pi16 ? n32 : n75377;
  assign n75379 = pi15 ? n75371 : n75378;
  assign n75380 = pi14 ? n75365 : n75379;
  assign n75381 = pi13 ? n75350 : n75380;
  assign n75382 = pi12 ? n75342 : n75381;
  assign n75383 = pi21 ? n32 : n71040;
  assign n75384 = pi22 ? n66891 : n685;
  assign n75385 = pi21 ? n75384 : n2637;
  assign n75386 = pi20 ? n75383 : n75385;
  assign n75387 = pi19 ? n32 : n75386;
  assign n75388 = pi18 ? n32 : n75387;
  assign n75389 = pi17 ? n32 : n75388;
  assign n75390 = pi16 ? n32 : n75389;
  assign n75391 = pi22 ? n40342 : n36798;
  assign n75392 = pi21 ? n32 : n75391;
  assign n75393 = pi23 ? n67465 : n685;
  assign n75394 = pi22 ? n75393 : n51564;
  assign n75395 = pi21 ? n75394 : n928;
  assign n75396 = pi20 ? n75392 : n75395;
  assign n75397 = pi19 ? n32 : n75396;
  assign n75398 = pi18 ? n32 : n75397;
  assign n75399 = pi17 ? n32 : n75398;
  assign n75400 = pi16 ? n32 : n75399;
  assign n75401 = pi15 ? n75390 : n75400;
  assign n75402 = pi20 ? n75392 : n75210;
  assign n75403 = pi19 ? n32 : n75402;
  assign n75404 = pi18 ? n32 : n75403;
  assign n75405 = pi17 ? n32 : n75404;
  assign n75406 = pi16 ? n32 : n75405;
  assign n75407 = pi22 ? n71003 : n43198;
  assign n75408 = pi21 ? n32 : n75407;
  assign n75409 = pi20 ? n75408 : n75219;
  assign n75410 = pi19 ? n32 : n75409;
  assign n75411 = pi18 ? n32 : n75410;
  assign n75412 = pi17 ? n32 : n75411;
  assign n75413 = pi16 ? n32 : n75412;
  assign n75414 = pi15 ? n75406 : n75413;
  assign n75415 = pi14 ? n75401 : n75414;
  assign n75416 = pi22 ? n37251 : n43198;
  assign n75417 = pi21 ? n32 : n75416;
  assign n75418 = pi20 ? n75417 : n72051;
  assign n75419 = pi19 ? n32 : n75418;
  assign n75420 = pi18 ? n32 : n75419;
  assign n75421 = pi17 ? n32 : n75420;
  assign n75422 = pi16 ? n32 : n75421;
  assign n75423 = pi22 ? n37873 : n14626;
  assign n75424 = pi21 ? n32 : n75423;
  assign n75425 = pi20 ? n75424 : n72062;
  assign n75426 = pi19 ? n32 : n75425;
  assign n75427 = pi18 ? n32 : n75426;
  assign n75428 = pi17 ? n32 : n75427;
  assign n75429 = pi16 ? n32 : n75428;
  assign n75430 = pi15 ? n75422 : n75429;
  assign n75431 = pi22 ? n36783 : n14626;
  assign n75432 = pi21 ? n32 : n75431;
  assign n75433 = pi20 ? n75432 : n60045;
  assign n75434 = pi19 ? n32 : n75433;
  assign n75435 = pi18 ? n32 : n75434;
  assign n75436 = pi17 ? n32 : n75435;
  assign n75437 = pi16 ? n32 : n75436;
  assign n75438 = pi15 ? n75429 : n75437;
  assign n75439 = pi14 ? n75430 : n75438;
  assign n75440 = pi13 ? n75415 : n75439;
  assign n75441 = pi20 ? n75266 : n1822;
  assign n75442 = pi19 ? n32 : n75441;
  assign n75443 = pi18 ? n32 : n75442;
  assign n75444 = pi17 ? n32 : n75443;
  assign n75445 = pi16 ? n32 : n75444;
  assign n75446 = pi15 ? n75445 : n75276;
  assign n75447 = pi14 ? n75263 : n75446;
  assign n75448 = pi22 ? n72270 : n706;
  assign n75449 = pi21 ? n32 : n75448;
  assign n75450 = pi20 ? n75449 : n32;
  assign n75451 = pi19 ? n32 : n75450;
  assign n75452 = pi18 ? n32 : n75451;
  assign n75453 = pi17 ? n32 : n75452;
  assign n75454 = pi16 ? n32 : n75453;
  assign n75455 = pi15 ? n75285 : n75454;
  assign n75456 = pi22 ? n74206 : n14363;
  assign n75457 = pi21 ? n32 : n75456;
  assign n75458 = pi20 ? n75457 : n32;
  assign n75459 = pi19 ? n32 : n75458;
  assign n75460 = pi18 ? n32 : n75459;
  assign n75461 = pi17 ? n32 : n75460;
  assign n75462 = pi16 ? n32 : n75461;
  assign n75463 = pi23 ? n51565 : n13481;
  assign n75464 = pi22 ? n75463 : n32;
  assign n75465 = pi21 ? n32 : n75464;
  assign n75466 = pi20 ? n75465 : n32;
  assign n75467 = pi19 ? n32 : n75466;
  assign n75468 = pi18 ? n32 : n75467;
  assign n75469 = pi17 ? n32 : n75468;
  assign n75470 = pi16 ? n32 : n75469;
  assign n75471 = pi15 ? n75462 : n75470;
  assign n75472 = pi14 ? n75455 : n75471;
  assign n75473 = pi13 ? n75447 : n75472;
  assign n75474 = pi12 ? n75440 : n75473;
  assign n75475 = pi11 ? n75382 : n75474;
  assign n75476 = pi10 ? n75475 : n32;
  assign n75477 = pi09 ? n75340 : n75476;
  assign n75478 = pi08 ? n75323 : n75477;
  assign n75479 = pi20 ? n46061 : n13040;
  assign n75480 = pi19 ? n32 : n75479;
  assign n75481 = pi18 ? n32 : n75480;
  assign n75482 = pi17 ? n32 : n75481;
  assign n75483 = pi16 ? n32 : n75482;
  assign n75484 = pi15 ? n32 : n75483;
  assign n75485 = pi20 ? n54444 : n61008;
  assign n75486 = pi19 ? n32 : n75485;
  assign n75487 = pi18 ? n32 : n75486;
  assign n75488 = pi17 ? n32 : n75487;
  assign n75489 = pi16 ? n32 : n75488;
  assign n75490 = pi14 ? n75484 : n75489;
  assign n75491 = pi13 ? n32 : n75490;
  assign n75492 = pi12 ? n32 : n75491;
  assign n75493 = pi11 ? n32 : n75492;
  assign n75494 = pi10 ? n32 : n75493;
  assign n75495 = pi20 ? n36867 : n61008;
  assign n75496 = pi19 ? n32 : n75495;
  assign n75497 = pi18 ? n32 : n75496;
  assign n75498 = pi17 ? n32 : n75497;
  assign n75499 = pi16 ? n32 : n75498;
  assign n75500 = pi15 ? n75499 : n74732;
  assign n75501 = pi14 ? n75499 : n75500;
  assign n75502 = pi20 ? n37955 : n1619;
  assign n75503 = pi19 ? n32 : n75502;
  assign n75504 = pi18 ? n32 : n75503;
  assign n75505 = pi17 ? n32 : n75504;
  assign n75506 = pi16 ? n32 : n75505;
  assign n75507 = pi14 ? n74732 : n75506;
  assign n75508 = pi13 ? n75501 : n75507;
  assign n75509 = pi20 ? n51233 : n61008;
  assign n75510 = pi19 ? n32 : n75509;
  assign n75511 = pi18 ? n32 : n75510;
  assign n75512 = pi17 ? n32 : n75511;
  assign n75513 = pi16 ? n32 : n75512;
  assign n75514 = pi15 ? n74732 : n75513;
  assign n75515 = pi20 ? n46188 : n75156;
  assign n75516 = pi19 ? n32 : n75515;
  assign n75517 = pi18 ? n32 : n75516;
  assign n75518 = pi17 ? n32 : n75517;
  assign n75519 = pi16 ? n32 : n75518;
  assign n75520 = pi20 ? n68256 : n75156;
  assign n75521 = pi19 ? n32 : n75520;
  assign n75522 = pi18 ? n32 : n75521;
  assign n75523 = pi17 ? n32 : n75522;
  assign n75524 = pi16 ? n32 : n75523;
  assign n75525 = pi15 ? n75519 : n75524;
  assign n75526 = pi14 ? n75514 : n75525;
  assign n75527 = pi20 ? n38997 : n68542;
  assign n75528 = pi19 ? n32 : n75527;
  assign n75529 = pi18 ? n32 : n75528;
  assign n75530 = pi17 ? n32 : n75529;
  assign n75531 = pi16 ? n32 : n75530;
  assign n75532 = pi15 ? n75531 : n75364;
  assign n75533 = pi20 ? n72046 : n75366;
  assign n75534 = pi19 ? n32 : n75533;
  assign n75535 = pi18 ? n32 : n75534;
  assign n75536 = pi17 ? n32 : n75535;
  assign n75537 = pi16 ? n32 : n75536;
  assign n75538 = pi20 ? n75373 : n68156;
  assign n75539 = pi19 ? n32 : n75538;
  assign n75540 = pi18 ? n32 : n75539;
  assign n75541 = pi17 ? n32 : n75540;
  assign n75542 = pi16 ? n32 : n75541;
  assign n75543 = pi15 ? n75537 : n75542;
  assign n75544 = pi14 ? n75532 : n75543;
  assign n75545 = pi13 ? n75526 : n75544;
  assign n75546 = pi12 ? n75508 : n75545;
  assign n75547 = pi22 ? n40342 : n36781;
  assign n75548 = pi21 ? n32 : n75547;
  assign n75549 = pi21 ? n59324 : n2637;
  assign n75550 = pi20 ? n75548 : n75549;
  assign n75551 = pi19 ? n32 : n75550;
  assign n75552 = pi18 ? n32 : n75551;
  assign n75553 = pi17 ? n32 : n75552;
  assign n75554 = pi16 ? n32 : n75553;
  assign n75555 = pi22 ? n65218 : n51564;
  assign n75556 = pi21 ? n75555 : n928;
  assign n75557 = pi20 ? n75392 : n75556;
  assign n75558 = pi19 ? n32 : n75557;
  assign n75559 = pi18 ? n32 : n75558;
  assign n75560 = pi17 ? n32 : n75559;
  assign n75561 = pi16 ? n32 : n75560;
  assign n75562 = pi15 ? n75554 : n75561;
  assign n75563 = pi22 ? n71003 : n36798;
  assign n75564 = pi21 ? n32 : n75563;
  assign n75565 = pi23 ? n21112 : n13481;
  assign n75566 = pi22 ? n75565 : n13481;
  assign n75567 = pi21 ? n75566 : n37639;
  assign n75568 = pi20 ? n75564 : n75567;
  assign n75569 = pi19 ? n32 : n75568;
  assign n75570 = pi18 ? n32 : n75569;
  assign n75571 = pi17 ? n32 : n75570;
  assign n75572 = pi16 ? n32 : n75571;
  assign n75573 = pi23 ? n13482 : n13481;
  assign n75574 = pi22 ? n75573 : n13481;
  assign n75575 = pi21 ? n75574 : n20952;
  assign n75576 = pi20 ? n75408 : n75575;
  assign n75577 = pi19 ? n32 : n75576;
  assign n75578 = pi18 ? n32 : n75577;
  assign n75579 = pi17 ? n32 : n75578;
  assign n75580 = pi16 ? n32 : n75579;
  assign n75581 = pi15 ? n75572 : n75580;
  assign n75582 = pi14 ? n75562 : n75581;
  assign n75583 = pi22 ? n41097 : n43198;
  assign n75584 = pi21 ? n32 : n75583;
  assign n75585 = pi20 ? n75584 : n72747;
  assign n75586 = pi19 ? n32 : n75585;
  assign n75587 = pi18 ? n32 : n75586;
  assign n75588 = pi17 ? n32 : n75587;
  assign n75589 = pi16 ? n32 : n75588;
  assign n75590 = pi22 ? n39996 : n14626;
  assign n75591 = pi21 ? n32 : n75590;
  assign n75592 = pi20 ? n75591 : n67728;
  assign n75593 = pi19 ? n32 : n75592;
  assign n75594 = pi18 ? n32 : n75593;
  assign n75595 = pi17 ? n32 : n75594;
  assign n75596 = pi16 ? n32 : n75595;
  assign n75597 = pi15 ? n75589 : n75596;
  assign n75598 = pi22 ? n45160 : n57632;
  assign n75599 = pi21 ? n32 : n75598;
  assign n75600 = pi20 ? n75599 : n60045;
  assign n75601 = pi19 ? n32 : n75600;
  assign n75602 = pi18 ? n32 : n75601;
  assign n75603 = pi17 ? n32 : n75602;
  assign n75604 = pi16 ? n32 : n75603;
  assign n75605 = pi15 ? n75596 : n75604;
  assign n75606 = pi14 ? n75597 : n75605;
  assign n75607 = pi13 ? n75582 : n75606;
  assign n75608 = pi22 ? n45160 : n13481;
  assign n75609 = pi21 ? n32 : n75608;
  assign n75610 = pi20 ? n75609 : n60045;
  assign n75611 = pi19 ? n32 : n75610;
  assign n75612 = pi18 ? n32 : n75611;
  assign n75613 = pi17 ? n32 : n75612;
  assign n75614 = pi16 ? n32 : n75613;
  assign n75615 = pi20 ? n72255 : n60045;
  assign n75616 = pi19 ? n32 : n75615;
  assign n75617 = pi18 ? n32 : n75616;
  assign n75618 = pi17 ? n32 : n75617;
  assign n75619 = pi16 ? n32 : n75618;
  assign n75620 = pi15 ? n75614 : n75619;
  assign n75621 = pi20 ? n72255 : n1822;
  assign n75622 = pi19 ? n32 : n75621;
  assign n75623 = pi18 ? n32 : n75622;
  assign n75624 = pi17 ? n32 : n75623;
  assign n75625 = pi16 ? n32 : n75624;
  assign n75626 = pi22 ? n74905 : n13481;
  assign n75627 = pi21 ? n32 : n75626;
  assign n75628 = pi20 ? n75627 : n32;
  assign n75629 = pi19 ? n32 : n75628;
  assign n75630 = pi18 ? n32 : n75629;
  assign n75631 = pi17 ? n32 : n75630;
  assign n75632 = pi16 ? n32 : n75631;
  assign n75633 = pi15 ? n75625 : n75632;
  assign n75634 = pi14 ? n75620 : n75633;
  assign n75635 = pi22 ? n70744 : n13481;
  assign n75636 = pi21 ? n32 : n75635;
  assign n75637 = pi20 ? n75636 : n32;
  assign n75638 = pi19 ? n32 : n75637;
  assign n75639 = pi18 ? n32 : n75638;
  assign n75640 = pi17 ? n32 : n75639;
  assign n75641 = pi16 ? n32 : n75640;
  assign n75642 = pi22 ? n70744 : n14363;
  assign n75643 = pi21 ? n32 : n75642;
  assign n75644 = pi20 ? n75643 : n32;
  assign n75645 = pi19 ? n32 : n75644;
  assign n75646 = pi18 ? n32 : n75645;
  assign n75647 = pi17 ? n32 : n75646;
  assign n75648 = pi16 ? n32 : n75647;
  assign n75649 = pi15 ? n75641 : n75648;
  assign n75650 = pi20 ? n72291 : n32;
  assign n75651 = pi19 ? n32 : n75650;
  assign n75652 = pi18 ? n32 : n75651;
  assign n75653 = pi17 ? n32 : n75652;
  assign n75654 = pi16 ? n32 : n75653;
  assign n75655 = pi22 ? n69890 : n32;
  assign n75656 = pi21 ? n32 : n75655;
  assign n75657 = pi20 ? n75656 : n32;
  assign n75658 = pi19 ? n32 : n75657;
  assign n75659 = pi18 ? n32 : n75658;
  assign n75660 = pi17 ? n32 : n75659;
  assign n75661 = pi16 ? n32 : n75660;
  assign n75662 = pi15 ? n75654 : n75661;
  assign n75663 = pi14 ? n75649 : n75662;
  assign n75664 = pi13 ? n75634 : n75663;
  assign n75665 = pi12 ? n75607 : n75664;
  assign n75666 = pi11 ? n75546 : n75665;
  assign n75667 = pi10 ? n75666 : n32;
  assign n75668 = pi09 ? n75494 : n75667;
  assign n75669 = pi20 ? n60055 : n75156;
  assign n75670 = pi19 ? n32 : n75669;
  assign n75671 = pi18 ? n32 : n75670;
  assign n75672 = pi17 ? n32 : n75671;
  assign n75673 = pi16 ? n32 : n75672;
  assign n75674 = pi15 ? n75519 : n75673;
  assign n75675 = pi14 ? n75514 : n75674;
  assign n75676 = pi20 ? n37955 : n58879;
  assign n75677 = pi19 ? n32 : n75676;
  assign n75678 = pi18 ? n32 : n75677;
  assign n75679 = pi17 ? n32 : n75678;
  assign n75680 = pi16 ? n32 : n75679;
  assign n75681 = pi20 ? n68256 : n69484;
  assign n75682 = pi19 ? n32 : n75681;
  assign n75683 = pi18 ? n32 : n75682;
  assign n75684 = pi17 ? n32 : n75683;
  assign n75685 = pi16 ? n32 : n75684;
  assign n75686 = pi15 ? n75680 : n75685;
  assign n75687 = pi20 ? n68280 : n72693;
  assign n75688 = pi19 ? n32 : n75687;
  assign n75689 = pi18 ? n32 : n75688;
  assign n75690 = pi17 ? n32 : n75689;
  assign n75691 = pi16 ? n32 : n75690;
  assign n75692 = pi24 ? n139 : n13481;
  assign n75693 = pi23 ? n75692 : n13481;
  assign n75694 = pi22 ? n75693 : n13481;
  assign n75695 = pi21 ? n75694 : n55560;
  assign n75696 = pi20 ? n72465 : n75695;
  assign n75697 = pi19 ? n32 : n75696;
  assign n75698 = pi18 ? n32 : n75697;
  assign n75699 = pi17 ? n32 : n75698;
  assign n75700 = pi16 ? n32 : n75699;
  assign n75701 = pi15 ? n75691 : n75700;
  assign n75702 = pi14 ? n75686 : n75701;
  assign n75703 = pi13 ? n75675 : n75702;
  assign n75704 = pi12 ? n75508 : n75703;
  assign n75705 = pi21 ? n62630 : n2637;
  assign n75706 = pi20 ? n72486 : n75705;
  assign n75707 = pi19 ? n32 : n75706;
  assign n75708 = pi18 ? n32 : n75707;
  assign n75709 = pi17 ? n32 : n75708;
  assign n75710 = pi16 ? n32 : n75709;
  assign n75711 = pi22 ? n45597 : n36798;
  assign n75712 = pi21 ? n32 : n75711;
  assign n75713 = pi20 ? n75712 : n75556;
  assign n75714 = pi19 ? n32 : n75713;
  assign n75715 = pi18 ? n32 : n75714;
  assign n75716 = pi17 ? n32 : n75715;
  assign n75717 = pi16 ? n32 : n75716;
  assign n75718 = pi15 ? n75710 : n75717;
  assign n75719 = pi22 ? n49720 : n36798;
  assign n75720 = pi21 ? n32 : n75719;
  assign n75721 = pi22 ? n71897 : n13481;
  assign n75722 = pi21 ? n75721 : n37639;
  assign n75723 = pi20 ? n75720 : n75722;
  assign n75724 = pi19 ? n32 : n75723;
  assign n75725 = pi18 ? n32 : n75724;
  assign n75726 = pi17 ? n32 : n75725;
  assign n75727 = pi16 ? n32 : n75726;
  assign n75728 = pi21 ? n32 : n59137;
  assign n75729 = pi20 ? n75728 : n75575;
  assign n75730 = pi19 ? n32 : n75729;
  assign n75731 = pi18 ? n32 : n75730;
  assign n75732 = pi17 ? n32 : n75731;
  assign n75733 = pi16 ? n32 : n75732;
  assign n75734 = pi15 ? n75727 : n75733;
  assign n75735 = pi14 ? n75718 : n75734;
  assign n75736 = pi22 ? n51754 : n43198;
  assign n75737 = pi21 ? n32 : n75736;
  assign n75738 = pi20 ? n75737 : n72747;
  assign n75739 = pi19 ? n32 : n75738;
  assign n75740 = pi18 ? n32 : n75739;
  assign n75741 = pi17 ? n32 : n75740;
  assign n75742 = pi16 ? n32 : n75741;
  assign n75743 = pi22 ? n45135 : n14626;
  assign n75744 = pi21 ? n32 : n75743;
  assign n75745 = pi20 ? n75744 : n67728;
  assign n75746 = pi19 ? n32 : n75745;
  assign n75747 = pi18 ? n32 : n75746;
  assign n75748 = pi17 ? n32 : n75747;
  assign n75749 = pi16 ? n32 : n75748;
  assign n75750 = pi15 ? n75742 : n75749;
  assign n75751 = pi15 ? n75749 : n75604;
  assign n75752 = pi14 ? n75750 : n75751;
  assign n75753 = pi13 ? n75735 : n75752;
  assign n75754 = pi22 ? n69401 : n14363;
  assign n75755 = pi21 ? n32 : n75754;
  assign n75756 = pi20 ? n75755 : n32;
  assign n75757 = pi19 ? n32 : n75756;
  assign n75758 = pi18 ? n32 : n75757;
  assign n75759 = pi17 ? n32 : n75758;
  assign n75760 = pi16 ? n32 : n75759;
  assign n75761 = pi15 ? n75760 : n32;
  assign n75762 = pi14 ? n75649 : n75761;
  assign n75763 = pi13 ? n75634 : n75762;
  assign n75764 = pi12 ? n75753 : n75763;
  assign n75765 = pi11 ? n75704 : n75764;
  assign n75766 = pi10 ? n75765 : n32;
  assign n75767 = pi09 ? n75494 : n75766;
  assign n75768 = pi08 ? n75668 : n75767;
  assign n75769 = pi07 ? n75478 : n75768;
  assign n75770 = pi20 ? n40054 : n74246;
  assign n75771 = pi19 ? n32 : n75770;
  assign n75772 = pi18 ? n32 : n75771;
  assign n75773 = pi17 ? n32 : n75772;
  assign n75774 = pi16 ? n32 : n75773;
  assign n75775 = pi15 ? n32 : n75774;
  assign n75776 = pi20 ? n40054 : n61008;
  assign n75777 = pi19 ? n32 : n75776;
  assign n75778 = pi18 ? n32 : n75777;
  assign n75779 = pi17 ? n32 : n75778;
  assign n75780 = pi16 ? n32 : n75779;
  assign n75781 = pi14 ? n75775 : n75780;
  assign n75782 = pi13 ? n32 : n75781;
  assign n75783 = pi12 ? n32 : n75782;
  assign n75784 = pi11 ? n32 : n75783;
  assign n75785 = pi10 ? n32 : n75784;
  assign n75786 = pi20 ? n37933 : n61008;
  assign n75787 = pi19 ? n32 : n75786;
  assign n75788 = pi18 ? n32 : n75787;
  assign n75789 = pi17 ? n32 : n75788;
  assign n75790 = pi16 ? n32 : n75789;
  assign n75791 = pi15 ? n75790 : n75499;
  assign n75792 = pi14 ? n75790 : n75791;
  assign n75793 = pi20 ? n60055 : n1619;
  assign n75794 = pi19 ? n32 : n75793;
  assign n75795 = pi18 ? n32 : n75794;
  assign n75796 = pi17 ? n32 : n75795;
  assign n75797 = pi16 ? n32 : n75796;
  assign n75798 = pi20 ? n60055 : n61008;
  assign n75799 = pi19 ? n32 : n75798;
  assign n75800 = pi18 ? n32 : n75799;
  assign n75801 = pi17 ? n32 : n75800;
  assign n75802 = pi16 ? n32 : n75801;
  assign n75803 = pi15 ? n75797 : n75802;
  assign n75804 = pi14 ? n75499 : n75803;
  assign n75805 = pi13 ? n75792 : n75804;
  assign n75806 = pi20 ? n36867 : n75156;
  assign n75807 = pi19 ? n32 : n75806;
  assign n75808 = pi18 ? n32 : n75807;
  assign n75809 = pi17 ? n32 : n75808;
  assign n75810 = pi16 ? n32 : n75809;
  assign n75811 = pi14 ? n75499 : n75810;
  assign n75812 = pi20 ? n37955 : n72686;
  assign n75813 = pi19 ? n32 : n75812;
  assign n75814 = pi18 ? n32 : n75813;
  assign n75815 = pi17 ? n32 : n75814;
  assign n75816 = pi16 ? n32 : n75815;
  assign n75817 = pi21 ? n68550 : n57433;
  assign n75818 = pi20 ? n68256 : n75817;
  assign n75819 = pi19 ? n32 : n75818;
  assign n75820 = pi18 ? n32 : n75819;
  assign n75821 = pi17 ? n32 : n75820;
  assign n75822 = pi16 ? n32 : n75821;
  assign n75823 = pi15 ? n75816 : n75822;
  assign n75824 = pi20 ? n68280 : n73244;
  assign n75825 = pi19 ? n32 : n75824;
  assign n75826 = pi18 ? n32 : n75825;
  assign n75827 = pi17 ? n32 : n75826;
  assign n75828 = pi16 ? n32 : n75827;
  assign n75829 = pi20 ? n68280 : n69066;
  assign n75830 = pi19 ? n32 : n75829;
  assign n75831 = pi18 ? n32 : n75830;
  assign n75832 = pi17 ? n32 : n75831;
  assign n75833 = pi16 ? n32 : n75832;
  assign n75834 = pi15 ? n75828 : n75833;
  assign n75835 = pi14 ? n75823 : n75834;
  assign n75836 = pi13 ? n75811 : n75835;
  assign n75837 = pi12 ? n75805 : n75836;
  assign n75838 = pi21 ? n63026 : n2637;
  assign n75839 = pi20 ? n72410 : n75838;
  assign n75840 = pi19 ? n32 : n75839;
  assign n75841 = pi18 ? n32 : n75840;
  assign n75842 = pi17 ? n32 : n75841;
  assign n75843 = pi16 ? n32 : n75842;
  assign n75844 = pi22 ? n45597 : n70065;
  assign n75845 = pi21 ? n32 : n75844;
  assign n75846 = pi20 ? n75845 : n73278;
  assign n75847 = pi19 ? n32 : n75846;
  assign n75848 = pi18 ? n32 : n75847;
  assign n75849 = pi17 ? n32 : n75848;
  assign n75850 = pi16 ? n32 : n75849;
  assign n75851 = pi15 ? n75843 : n75850;
  assign n75852 = pi21 ? n65025 : n32;
  assign n75853 = pi20 ? n75720 : n75852;
  assign n75854 = pi19 ? n32 : n75853;
  assign n75855 = pi18 ? n32 : n75854;
  assign n75856 = pi17 ? n32 : n75855;
  assign n75857 = pi16 ? n32 : n75856;
  assign n75858 = pi15 ? n75727 : n75857;
  assign n75859 = pi14 ? n75851 : n75858;
  assign n75860 = pi20 ? n75737 : n6935;
  assign n75861 = pi19 ? n32 : n75860;
  assign n75862 = pi18 ? n32 : n75861;
  assign n75863 = pi17 ? n32 : n75862;
  assign n75864 = pi16 ? n32 : n75863;
  assign n75865 = pi22 ? n45634 : n14626;
  assign n75866 = pi21 ? n32 : n75865;
  assign n75867 = pi20 ? n75866 : n67728;
  assign n75868 = pi19 ? n32 : n75867;
  assign n75869 = pi18 ? n32 : n75868;
  assign n75870 = pi17 ? n32 : n75869;
  assign n75871 = pi16 ? n32 : n75870;
  assign n75872 = pi15 ? n75864 : n75871;
  assign n75873 = pi21 ? n32 : n71098;
  assign n75874 = pi20 ? n75873 : n62857;
  assign n75875 = pi19 ? n32 : n75874;
  assign n75876 = pi18 ? n32 : n75875;
  assign n75877 = pi17 ? n32 : n75876;
  assign n75878 = pi16 ? n32 : n75877;
  assign n75879 = pi20 ? n75873 : n60045;
  assign n75880 = pi19 ? n32 : n75879;
  assign n75881 = pi18 ? n32 : n75880;
  assign n75882 = pi17 ? n32 : n75881;
  assign n75883 = pi16 ? n32 : n75882;
  assign n75884 = pi15 ? n75878 : n75883;
  assign n75885 = pi14 ? n75872 : n75884;
  assign n75886 = pi13 ? n75859 : n75885;
  assign n75887 = pi22 ? n46275 : n62803;
  assign n75888 = pi21 ? n32 : n75887;
  assign n75889 = pi20 ? n75888 : n60045;
  assign n75890 = pi19 ? n32 : n75889;
  assign n75891 = pi18 ? n32 : n75890;
  assign n75892 = pi17 ? n32 : n75891;
  assign n75893 = pi16 ? n32 : n75892;
  assign n75894 = pi21 ? n32 : n71113;
  assign n75895 = pi20 ? n75894 : n2701;
  assign n75896 = pi19 ? n32 : n75895;
  assign n75897 = pi18 ? n32 : n75896;
  assign n75898 = pi17 ? n32 : n75897;
  assign n75899 = pi16 ? n32 : n75898;
  assign n75900 = pi15 ? n75893 : n75899;
  assign n75901 = pi22 ? n63432 : n56186;
  assign n75902 = pi21 ? n32 : n75901;
  assign n75903 = pi20 ? n75902 : n20953;
  assign n75904 = pi19 ? n32 : n75903;
  assign n75905 = pi18 ? n32 : n75904;
  assign n75906 = pi17 ? n32 : n75905;
  assign n75907 = pi16 ? n32 : n75906;
  assign n75908 = pi21 ? n32 : n74223;
  assign n75909 = pi20 ? n75908 : n32;
  assign n75910 = pi19 ? n32 : n75909;
  assign n75911 = pi18 ? n32 : n75910;
  assign n75912 = pi17 ? n32 : n75911;
  assign n75913 = pi16 ? n32 : n75912;
  assign n75914 = pi15 ? n75907 : n75913;
  assign n75915 = pi14 ? n75900 : n75914;
  assign n75916 = pi22 ? n71540 : n53982;
  assign n75917 = pi21 ? n32 : n75916;
  assign n75918 = pi20 ? n75917 : n32;
  assign n75919 = pi19 ? n32 : n75918;
  assign n75920 = pi18 ? n32 : n75919;
  assign n75921 = pi17 ? n32 : n75920;
  assign n75922 = pi16 ? n32 : n75921;
  assign n75923 = pi15 ? n75922 : n75760;
  assign n75924 = pi14 ? n75923 : n32;
  assign n75925 = pi13 ? n75915 : n75924;
  assign n75926 = pi12 ? n75886 : n75925;
  assign n75927 = pi11 ? n75837 : n75926;
  assign n75928 = pi10 ? n75927 : n32;
  assign n75929 = pi09 ? n75785 : n75928;
  assign n75930 = pi20 ? n38981 : n74246;
  assign n75931 = pi19 ? n32 : n75930;
  assign n75932 = pi18 ? n32 : n75931;
  assign n75933 = pi17 ? n32 : n75932;
  assign n75934 = pi16 ? n32 : n75933;
  assign n75935 = pi15 ? n32 : n75934;
  assign n75936 = pi20 ? n38981 : n61008;
  assign n75937 = pi19 ? n32 : n75936;
  assign n75938 = pi18 ? n32 : n75937;
  assign n75939 = pi17 ? n32 : n75938;
  assign n75940 = pi16 ? n32 : n75939;
  assign n75941 = pi15 ? n75940 : n75780;
  assign n75942 = pi14 ? n75935 : n75941;
  assign n75943 = pi13 ? n32 : n75942;
  assign n75944 = pi12 ? n32 : n75943;
  assign n75945 = pi11 ? n32 : n75944;
  assign n75946 = pi10 ? n32 : n75945;
  assign n75947 = pi20 ? n54401 : n61008;
  assign n75948 = pi19 ? n32 : n75947;
  assign n75949 = pi18 ? n32 : n75948;
  assign n75950 = pi17 ? n32 : n75949;
  assign n75951 = pi16 ? n32 : n75950;
  assign n75952 = pi20 ? n37933 : n75156;
  assign n75953 = pi19 ? n32 : n75952;
  assign n75954 = pi18 ? n32 : n75953;
  assign n75955 = pi17 ? n32 : n75954;
  assign n75956 = pi16 ? n32 : n75955;
  assign n75957 = pi14 ? n75951 : n75956;
  assign n75958 = pi20 ? n36867 : n72686;
  assign n75959 = pi19 ? n32 : n75958;
  assign n75960 = pi18 ? n32 : n75959;
  assign n75961 = pi17 ? n32 : n75960;
  assign n75962 = pi16 ? n32 : n75961;
  assign n75963 = pi20 ? n60055 : n75817;
  assign n75964 = pi19 ? n32 : n75963;
  assign n75965 = pi18 ? n32 : n75964;
  assign n75966 = pi17 ? n32 : n75965;
  assign n75967 = pi16 ? n32 : n75966;
  assign n75968 = pi15 ? n75962 : n75967;
  assign n75969 = pi20 ? n75136 : n73244;
  assign n75970 = pi19 ? n32 : n75969;
  assign n75971 = pi18 ? n32 : n75970;
  assign n75972 = pi17 ? n32 : n75971;
  assign n75973 = pi16 ? n32 : n75972;
  assign n75974 = pi20 ? n70117 : n69066;
  assign n75975 = pi19 ? n32 : n75974;
  assign n75976 = pi18 ? n32 : n75975;
  assign n75977 = pi17 ? n32 : n75976;
  assign n75978 = pi16 ? n32 : n75977;
  assign n75979 = pi15 ? n75973 : n75978;
  assign n75980 = pi14 ? n75968 : n75979;
  assign n75981 = pi13 ? n75957 : n75980;
  assign n75982 = pi12 ? n75805 : n75981;
  assign n75983 = pi22 ? n72382 : n51564;
  assign n75984 = pi21 ? n75983 : n2637;
  assign n75985 = pi20 ? n70117 : n75984;
  assign n75986 = pi19 ? n32 : n75985;
  assign n75987 = pi18 ? n32 : n75986;
  assign n75988 = pi17 ? n32 : n75987;
  assign n75989 = pi16 ? n32 : n75988;
  assign n75990 = pi22 ? n45516 : n70065;
  assign n75991 = pi21 ? n32 : n75990;
  assign n75992 = pi21 ? n62639 : n928;
  assign n75993 = pi20 ? n75991 : n75992;
  assign n75994 = pi19 ? n32 : n75993;
  assign n75995 = pi18 ? n32 : n75994;
  assign n75996 = pi17 ? n32 : n75995;
  assign n75997 = pi16 ? n32 : n75996;
  assign n75998 = pi15 ? n75989 : n75997;
  assign n75999 = pi22 ? n45516 : n36798;
  assign n76000 = pi21 ? n32 : n75999;
  assign n76001 = pi21 ? n63544 : n37639;
  assign n76002 = pi20 ? n76000 : n76001;
  assign n76003 = pi19 ? n32 : n76002;
  assign n76004 = pi18 ? n32 : n76003;
  assign n76005 = pi17 ? n32 : n76004;
  assign n76006 = pi16 ? n32 : n76005;
  assign n76007 = pi22 ? n46757 : n36798;
  assign n76008 = pi21 ? n32 : n76007;
  assign n76009 = pi20 ? n76008 : n75852;
  assign n76010 = pi19 ? n32 : n76009;
  assign n76011 = pi18 ? n32 : n76010;
  assign n76012 = pi17 ? n32 : n76011;
  assign n76013 = pi16 ? n32 : n76012;
  assign n76014 = pi15 ? n76006 : n76013;
  assign n76015 = pi14 ? n75998 : n76014;
  assign n76016 = pi22 ? n45634 : n43198;
  assign n76017 = pi21 ? n32 : n76016;
  assign n76018 = pi20 ? n76017 : n6935;
  assign n76019 = pi19 ? n32 : n76018;
  assign n76020 = pi18 ? n32 : n76019;
  assign n76021 = pi17 ? n32 : n76020;
  assign n76022 = pi16 ? n32 : n76021;
  assign n76023 = pi15 ? n76022 : n75871;
  assign n76024 = pi14 ? n76023 : n75884;
  assign n76025 = pi13 ? n76015 : n76024;
  assign n76026 = pi21 ? n32 : n74216;
  assign n76027 = pi20 ? n76026 : n53984;
  assign n76028 = pi19 ? n32 : n76027;
  assign n76029 = pi18 ? n32 : n76028;
  assign n76030 = pi17 ? n32 : n76029;
  assign n76031 = pi16 ? n32 : n76030;
  assign n76032 = pi15 ? n75893 : n76031;
  assign n76033 = pi22 ? n71540 : n13481;
  assign n76034 = pi21 ? n32 : n76033;
  assign n76035 = pi20 ? n76034 : n20953;
  assign n76036 = pi19 ? n32 : n76035;
  assign n76037 = pi18 ? n32 : n76036;
  assign n76038 = pi17 ? n32 : n76037;
  assign n76039 = pi16 ? n32 : n76038;
  assign n76040 = pi20 ? n76034 : n32;
  assign n76041 = pi19 ? n32 : n76040;
  assign n76042 = pi18 ? n32 : n76041;
  assign n76043 = pi17 ? n32 : n76042;
  assign n76044 = pi16 ? n32 : n76043;
  assign n76045 = pi15 ? n76039 : n76044;
  assign n76046 = pi14 ? n76032 : n76045;
  assign n76047 = pi21 ? n32 : n74493;
  assign n76048 = pi20 ? n76047 : n32;
  assign n76049 = pi19 ? n32 : n76048;
  assign n76050 = pi18 ? n32 : n76049;
  assign n76051 = pi17 ? n32 : n76050;
  assign n76052 = pi16 ? n32 : n76051;
  assign n76053 = pi14 ? n76052 : n32;
  assign n76054 = pi13 ? n76046 : n76053;
  assign n76055 = pi12 ? n76025 : n76054;
  assign n76056 = pi11 ? n75982 : n76055;
  assign n76057 = pi10 ? n76056 : n32;
  assign n76058 = pi09 ? n75946 : n76057;
  assign n76059 = pi08 ? n75929 : n76058;
  assign n76060 = pi21 ? n20563 : n13049;
  assign n76061 = pi20 ? n38981 : n76060;
  assign n76062 = pi19 ? n32 : n76061;
  assign n76063 = pi18 ? n32 : n76062;
  assign n76064 = pi17 ? n32 : n76063;
  assign n76065 = pi16 ? n32 : n76064;
  assign n76066 = pi15 ? n32 : n76065;
  assign n76067 = pi14 ? n76066 : n75940;
  assign n76068 = pi13 ? n32 : n76067;
  assign n76069 = pi12 ? n32 : n76068;
  assign n76070 = pi11 ? n32 : n76069;
  assign n76071 = pi10 ? n32 : n76070;
  assign n76072 = pi15 ? n75780 : n75790;
  assign n76073 = pi14 ? n75780 : n76072;
  assign n76074 = pi20 ? n46061 : n61008;
  assign n76075 = pi19 ? n32 : n76074;
  assign n76076 = pi18 ? n32 : n76075;
  assign n76077 = pi17 ? n32 : n76076;
  assign n76078 = pi16 ? n32 : n76077;
  assign n76079 = pi15 ? n75790 : n76078;
  assign n76080 = pi20 ? n37933 : n66577;
  assign n76081 = pi19 ? n32 : n76080;
  assign n76082 = pi18 ? n32 : n76081;
  assign n76083 = pi17 ? n32 : n76082;
  assign n76084 = pi16 ? n32 : n76083;
  assign n76085 = pi15 ? n76084 : n75790;
  assign n76086 = pi14 ? n76079 : n76085;
  assign n76087 = pi13 ? n76073 : n76086;
  assign n76088 = pi14 ? n75790 : n75956;
  assign n76089 = pi22 ? n30115 : n39190;
  assign n76090 = pi21 ? n32 : n76089;
  assign n76091 = pi20 ? n76090 : n67195;
  assign n76092 = pi19 ? n32 : n76091;
  assign n76093 = pi18 ? n32 : n76092;
  assign n76094 = pi17 ? n32 : n76093;
  assign n76095 = pi16 ? n32 : n76094;
  assign n76096 = pi21 ? n63922 : n58966;
  assign n76097 = pi20 ? n60055 : n76096;
  assign n76098 = pi19 ? n32 : n76097;
  assign n76099 = pi18 ? n32 : n76098;
  assign n76100 = pi17 ? n32 : n76099;
  assign n76101 = pi16 ? n32 : n76100;
  assign n76102 = pi15 ? n76095 : n76101;
  assign n76103 = pi20 ? n75136 : n75366;
  assign n76104 = pi19 ? n32 : n76103;
  assign n76105 = pi18 ? n32 : n76104;
  assign n76106 = pi17 ? n32 : n76105;
  assign n76107 = pi16 ? n32 : n76106;
  assign n76108 = pi22 ? n46165 : n58710;
  assign n76109 = pi21 ? n32 : n76108;
  assign n76110 = pi20 ? n76109 : n69066;
  assign n76111 = pi19 ? n32 : n76110;
  assign n76112 = pi18 ? n32 : n76111;
  assign n76113 = pi17 ? n32 : n76112;
  assign n76114 = pi16 ? n32 : n76113;
  assign n76115 = pi15 ? n76107 : n76114;
  assign n76116 = pi14 ? n76102 : n76115;
  assign n76117 = pi13 ? n76088 : n76116;
  assign n76118 = pi12 ? n76087 : n76117;
  assign n76119 = pi22 ? n46165 : n36781;
  assign n76120 = pi21 ? n32 : n76119;
  assign n76121 = pi23 ? n59885 : n51564;
  assign n76122 = pi22 ? n76121 : n51564;
  assign n76123 = pi21 ? n76122 : n59357;
  assign n76124 = pi20 ? n76120 : n76123;
  assign n76125 = pi19 ? n32 : n76124;
  assign n76126 = pi18 ? n32 : n76125;
  assign n76127 = pi17 ? n32 : n76126;
  assign n76128 = pi16 ? n32 : n76127;
  assign n76129 = pi22 ? n45516 : n36781;
  assign n76130 = pi21 ? n32 : n76129;
  assign n76131 = pi20 ? n76130 : n75992;
  assign n76132 = pi19 ? n32 : n76131;
  assign n76133 = pi18 ? n32 : n76132;
  assign n76134 = pi17 ? n32 : n76133;
  assign n76135 = pi16 ? n32 : n76134;
  assign n76136 = pi15 ? n76128 : n76135;
  assign n76137 = pi20 ? n76008 : n72747;
  assign n76138 = pi19 ? n32 : n76137;
  assign n76139 = pi18 ? n32 : n76138;
  assign n76140 = pi17 ? n32 : n76139;
  assign n76141 = pi16 ? n32 : n76140;
  assign n76142 = pi15 ? n76006 : n76141;
  assign n76143 = pi14 ? n76136 : n76142;
  assign n76144 = pi20 ? n48857 : n6935;
  assign n76145 = pi19 ? n32 : n76144;
  assign n76146 = pi18 ? n32 : n76145;
  assign n76147 = pi17 ? n32 : n76146;
  assign n76148 = pi16 ? n32 : n76147;
  assign n76149 = pi20 ? n63830 : n67728;
  assign n76150 = pi19 ? n32 : n76149;
  assign n76151 = pi18 ? n32 : n76150;
  assign n76152 = pi17 ? n32 : n76151;
  assign n76153 = pi16 ? n32 : n76152;
  assign n76154 = pi15 ? n76148 : n76153;
  assign n76155 = pi20 ? n63830 : n62857;
  assign n76156 = pi19 ? n32 : n76155;
  assign n76157 = pi18 ? n32 : n76156;
  assign n76158 = pi17 ? n32 : n76157;
  assign n76159 = pi16 ? n32 : n76158;
  assign n76160 = pi22 ? n32 : n57197;
  assign n76161 = pi21 ? n32 : n76160;
  assign n76162 = pi20 ? n76161 : n60045;
  assign n76163 = pi19 ? n32 : n76162;
  assign n76164 = pi18 ? n32 : n76163;
  assign n76165 = pi17 ? n32 : n76164;
  assign n76166 = pi16 ? n32 : n76165;
  assign n76167 = pi15 ? n76159 : n76166;
  assign n76168 = pi14 ? n76154 : n76167;
  assign n76169 = pi13 ? n76143 : n76168;
  assign n76170 = pi21 ? n32 : n71129;
  assign n76171 = pi20 ? n76170 : n60045;
  assign n76172 = pi19 ? n32 : n76171;
  assign n76173 = pi18 ? n32 : n76172;
  assign n76174 = pi17 ? n32 : n76173;
  assign n76175 = pi16 ? n32 : n76174;
  assign n76176 = pi20 ? n72901 : n53984;
  assign n76177 = pi19 ? n32 : n76176;
  assign n76178 = pi18 ? n32 : n76177;
  assign n76179 = pi17 ? n32 : n76178;
  assign n76180 = pi16 ? n32 : n76179;
  assign n76181 = pi15 ? n76175 : n76180;
  assign n76182 = pi20 ? n72596 : n20953;
  assign n76183 = pi19 ? n32 : n76182;
  assign n76184 = pi18 ? n32 : n76183;
  assign n76185 = pi17 ? n32 : n76184;
  assign n76186 = pi16 ? n32 : n76185;
  assign n76187 = pi20 ? n72611 : n32;
  assign n76188 = pi19 ? n32 : n76187;
  assign n76189 = pi18 ? n32 : n76188;
  assign n76190 = pi17 ? n32 : n76189;
  assign n76191 = pi16 ? n32 : n76190;
  assign n76192 = pi15 ? n76186 : n76191;
  assign n76193 = pi14 ? n76181 : n76192;
  assign n76194 = pi15 ? n76052 : n32;
  assign n76195 = pi14 ? n76194 : n32;
  assign n76196 = pi13 ? n76193 : n76195;
  assign n76197 = pi12 ? n76169 : n76196;
  assign n76198 = pi11 ? n76118 : n76197;
  assign n76199 = pi10 ? n76198 : n32;
  assign n76200 = pi09 ? n76071 : n76199;
  assign n76201 = pi20 ? n6783 : n76060;
  assign n76202 = pi19 ? n32 : n76201;
  assign n76203 = pi18 ? n32 : n76202;
  assign n76204 = pi17 ? n32 : n76203;
  assign n76205 = pi16 ? n32 : n76204;
  assign n76206 = pi15 ? n32 : n76205;
  assign n76207 = pi20 ? n6783 : n61008;
  assign n76208 = pi19 ? n32 : n76207;
  assign n76209 = pi18 ? n32 : n76208;
  assign n76210 = pi17 ? n32 : n76209;
  assign n76211 = pi16 ? n32 : n76210;
  assign n76212 = pi15 ? n76211 : n75940;
  assign n76213 = pi14 ? n76206 : n76212;
  assign n76214 = pi13 ? n32 : n76213;
  assign n76215 = pi12 ? n32 : n76214;
  assign n76216 = pi11 ? n32 : n76215;
  assign n76217 = pi10 ? n32 : n76216;
  assign n76218 = pi15 ? n75780 : n76078;
  assign n76219 = pi20 ? n40054 : n66577;
  assign n76220 = pi19 ? n32 : n76219;
  assign n76221 = pi18 ? n32 : n76220;
  assign n76222 = pi17 ? n32 : n76221;
  assign n76223 = pi16 ? n32 : n76222;
  assign n76224 = pi15 ? n76223 : n75780;
  assign n76225 = pi14 ? n76218 : n76224;
  assign n76226 = pi13 ? n76073 : n76225;
  assign n76227 = pi20 ? n40054 : n75156;
  assign n76228 = pi19 ? n32 : n76227;
  assign n76229 = pi18 ? n32 : n76228;
  assign n76230 = pi17 ? n32 : n76229;
  assign n76231 = pi16 ? n32 : n76230;
  assign n76232 = pi14 ? n75780 : n76231;
  assign n76233 = pi20 ? n64225 : n67195;
  assign n76234 = pi19 ? n32 : n76233;
  assign n76235 = pi18 ? n32 : n76234;
  assign n76236 = pi17 ? n32 : n76235;
  assign n76237 = pi16 ? n32 : n76236;
  assign n76238 = pi20 ? n46061 : n76096;
  assign n76239 = pi19 ? n32 : n76238;
  assign n76240 = pi18 ? n32 : n76239;
  assign n76241 = pi17 ? n32 : n76240;
  assign n76242 = pi16 ? n32 : n76241;
  assign n76243 = pi15 ? n76237 : n76242;
  assign n76244 = pi20 ? n54444 : n75366;
  assign n76245 = pi19 ? n32 : n76244;
  assign n76246 = pi18 ? n32 : n76245;
  assign n76247 = pi17 ? n32 : n76246;
  assign n76248 = pi16 ? n32 : n76247;
  assign n76249 = pi22 ? n32 : n58710;
  assign n76250 = pi21 ? n32 : n76249;
  assign n76251 = pi23 ? n7420 : n13481;
  assign n76252 = pi22 ? n76251 : n13481;
  assign n76253 = pi21 ? n76252 : n37639;
  assign n76254 = pi20 ? n76250 : n76253;
  assign n76255 = pi19 ? n32 : n76254;
  assign n76256 = pi18 ? n32 : n76255;
  assign n76257 = pi17 ? n32 : n76256;
  assign n76258 = pi16 ? n32 : n76257;
  assign n76259 = pi15 ? n76248 : n76258;
  assign n76260 = pi14 ? n76243 : n76259;
  assign n76261 = pi13 ? n76232 : n76260;
  assign n76262 = pi12 ? n76226 : n76261;
  assign n76263 = pi20 ? n65264 : n76123;
  assign n76264 = pi19 ? n32 : n76263;
  assign n76265 = pi18 ? n32 : n76264;
  assign n76266 = pi17 ? n32 : n76265;
  assign n76267 = pi16 ? n32 : n76266;
  assign n76268 = pi20 ? n65264 : n75992;
  assign n76269 = pi19 ? n32 : n76268;
  assign n76270 = pi18 ? n32 : n76269;
  assign n76271 = pi17 ? n32 : n76270;
  assign n76272 = pi16 ? n32 : n76271;
  assign n76273 = pi15 ? n76267 : n76272;
  assign n76274 = pi23 ? n1598 : n13481;
  assign n76275 = pi22 ? n76274 : n61712;
  assign n76276 = pi21 ? n76275 : n32;
  assign n76277 = pi20 ? n48822 : n76276;
  assign n76278 = pi19 ? n32 : n76277;
  assign n76279 = pi18 ? n32 : n76278;
  assign n76280 = pi17 ? n32 : n76279;
  assign n76281 = pi16 ? n32 : n76280;
  assign n76282 = pi20 ? n48822 : n72747;
  assign n76283 = pi19 ? n32 : n76282;
  assign n76284 = pi18 ? n32 : n76283;
  assign n76285 = pi17 ? n32 : n76284;
  assign n76286 = pi16 ? n32 : n76285;
  assign n76287 = pi15 ? n76281 : n76286;
  assign n76288 = pi14 ? n76273 : n76287;
  assign n76289 = pi20 ? n63830 : n60045;
  assign n76290 = pi19 ? n32 : n76289;
  assign n76291 = pi18 ? n32 : n76290;
  assign n76292 = pi17 ? n32 : n76291;
  assign n76293 = pi16 ? n32 : n76292;
  assign n76294 = pi15 ? n76148 : n76293;
  assign n76295 = pi14 ? n76294 : n76167;
  assign n76296 = pi13 ? n76288 : n76295;
  assign n76297 = pi20 ? n76170 : n53984;
  assign n76298 = pi19 ? n32 : n76297;
  assign n76299 = pi18 ? n32 : n76298;
  assign n76300 = pi17 ? n32 : n76299;
  assign n76301 = pi16 ? n32 : n76300;
  assign n76302 = pi20 ? n72901 : n20953;
  assign n76303 = pi19 ? n32 : n76302;
  assign n76304 = pi18 ? n32 : n76303;
  assign n76305 = pi17 ? n32 : n76304;
  assign n76306 = pi16 ? n32 : n76305;
  assign n76307 = pi15 ? n76301 : n76306;
  assign n76308 = pi23 ? n69724 : n14362;
  assign n76309 = pi22 ? n32 : n76308;
  assign n76310 = pi21 ? n32 : n76309;
  assign n76311 = pi20 ? n76310 : n32;
  assign n76312 = pi19 ? n32 : n76311;
  assign n76313 = pi18 ? n32 : n76312;
  assign n76314 = pi17 ? n32 : n76313;
  assign n76315 = pi16 ? n32 : n76314;
  assign n76316 = pi15 ? n76315 : n32;
  assign n76317 = pi14 ? n76307 : n76316;
  assign n76318 = pi13 ? n76317 : n32;
  assign n76319 = pi12 ? n76296 : n76318;
  assign n76320 = pi11 ? n76262 : n76319;
  assign n76321 = pi10 ? n76320 : n32;
  assign n76322 = pi09 ? n76217 : n76321;
  assign n76323 = pi08 ? n76200 : n76322;
  assign n76324 = pi07 ? n76059 : n76323;
  assign n76325 = pi06 ? n75769 : n76324;
  assign n76326 = pi20 ? n37926 : n13050;
  assign n76327 = pi19 ? n32 : n76326;
  assign n76328 = pi18 ? n32 : n76327;
  assign n76329 = pi17 ? n32 : n76328;
  assign n76330 = pi16 ? n32 : n76329;
  assign n76331 = pi15 ? n32 : n76330;
  assign n76332 = pi20 ? n37926 : n61008;
  assign n76333 = pi19 ? n32 : n76332;
  assign n76334 = pi18 ? n32 : n76333;
  assign n76335 = pi17 ? n32 : n76334;
  assign n76336 = pi16 ? n32 : n76335;
  assign n76337 = pi14 ? n76331 : n76336;
  assign n76338 = pi13 ? n32 : n76337;
  assign n76339 = pi12 ? n32 : n76338;
  assign n76340 = pi11 ? n32 : n76339;
  assign n76341 = pi10 ? n32 : n76340;
  assign n76342 = pi14 ? n75940 : n75941;
  assign n76343 = pi21 ? n32 : n73739;
  assign n76344 = pi20 ? n76343 : n61008;
  assign n76345 = pi19 ? n32 : n76344;
  assign n76346 = pi18 ? n32 : n76345;
  assign n76347 = pi17 ? n32 : n76346;
  assign n76348 = pi16 ? n32 : n76347;
  assign n76349 = pi15 ? n75780 : n76348;
  assign n76350 = pi14 ? n76349 : n75780;
  assign n76351 = pi13 ? n76342 : n76350;
  assign n76352 = pi21 ? n33792 : n1618;
  assign n76353 = pi20 ? n73068 : n76352;
  assign n76354 = pi19 ? n32 : n76353;
  assign n76355 = pi18 ? n32 : n76354;
  assign n76356 = pi17 ? n32 : n76355;
  assign n76357 = pi16 ? n32 : n76356;
  assign n76358 = pi15 ? n76231 : n76357;
  assign n76359 = pi14 ? n75780 : n76358;
  assign n76360 = pi22 ? n32 : n64662;
  assign n76361 = pi21 ? n32 : n76360;
  assign n76362 = pi20 ? n76361 : n74544;
  assign n76363 = pi19 ? n32 : n76362;
  assign n76364 = pi18 ? n32 : n76363;
  assign n76365 = pi17 ? n32 : n76364;
  assign n76366 = pi16 ? n32 : n76365;
  assign n76367 = pi15 ? n76237 : n76366;
  assign n76368 = pi23 ? n30868 : n55580;
  assign n76369 = pi22 ? n32 : n76368;
  assign n76370 = pi21 ? n32 : n76369;
  assign n76371 = pi20 ? n76370 : n71211;
  assign n76372 = pi19 ? n32 : n76371;
  assign n76373 = pi18 ? n32 : n76372;
  assign n76374 = pi17 ? n32 : n76373;
  assign n76375 = pi16 ? n32 : n76374;
  assign n76376 = pi20 ? n76250 : n75705;
  assign n76377 = pi19 ? n32 : n76376;
  assign n76378 = pi18 ? n32 : n76377;
  assign n76379 = pi17 ? n32 : n76378;
  assign n76380 = pi16 ? n32 : n76379;
  assign n76381 = pi15 ? n76375 : n76380;
  assign n76382 = pi14 ? n76367 : n76381;
  assign n76383 = pi13 ? n76359 : n76382;
  assign n76384 = pi12 ? n76351 : n76383;
  assign n76385 = pi22 ? n64161 : n316;
  assign n76386 = pi21 ? n76385 : n59357;
  assign n76387 = pi20 ? n73105 : n76386;
  assign n76388 = pi19 ? n32 : n76387;
  assign n76389 = pi18 ? n32 : n76388;
  assign n76390 = pi17 ? n32 : n76389;
  assign n76391 = pi16 ? n32 : n76390;
  assign n76392 = pi20 ? n73105 : n75992;
  assign n76393 = pi19 ? n32 : n76392;
  assign n76394 = pi18 ? n32 : n76393;
  assign n76395 = pi17 ? n32 : n76394;
  assign n76396 = pi16 ? n32 : n76395;
  assign n76397 = pi15 ? n76391 : n76396;
  assign n76398 = pi22 ? n32 : n43191;
  assign n76399 = pi21 ? n32 : n76398;
  assign n76400 = pi22 ? n75393 : n759;
  assign n76401 = pi21 ? n76400 : n32;
  assign n76402 = pi20 ? n76399 : n76401;
  assign n76403 = pi19 ? n32 : n76402;
  assign n76404 = pi18 ? n32 : n76403;
  assign n76405 = pi17 ? n32 : n76404;
  assign n76406 = pi16 ? n32 : n76405;
  assign n76407 = pi23 ? n36782 : n43198;
  assign n76408 = pi22 ? n32 : n76407;
  assign n76409 = pi21 ? n32 : n76408;
  assign n76410 = pi20 ? n76409 : n72747;
  assign n76411 = pi19 ? n32 : n76410;
  assign n76412 = pi18 ? n32 : n76411;
  assign n76413 = pi17 ? n32 : n76412;
  assign n76414 = pi16 ? n32 : n76413;
  assign n76415 = pi15 ? n76406 : n76414;
  assign n76416 = pi14 ? n76397 : n76415;
  assign n76417 = pi23 ? n36830 : n43198;
  assign n76418 = pi22 ? n32 : n76417;
  assign n76419 = pi21 ? n32 : n76418;
  assign n76420 = pi20 ? n76419 : n72062;
  assign n76421 = pi19 ? n32 : n76420;
  assign n76422 = pi18 ? n32 : n76421;
  assign n76423 = pi17 ? n32 : n76422;
  assign n76424 = pi16 ? n32 : n76423;
  assign n76425 = pi23 ? n36830 : n14626;
  assign n76426 = pi22 ? n32 : n76425;
  assign n76427 = pi21 ? n32 : n76426;
  assign n76428 = pi20 ? n76427 : n3210;
  assign n76429 = pi19 ? n32 : n76428;
  assign n76430 = pi18 ? n32 : n76429;
  assign n76431 = pi17 ? n32 : n76430;
  assign n76432 = pi16 ? n32 : n76431;
  assign n76433 = pi15 ? n76424 : n76432;
  assign n76434 = pi23 ? n46274 : n14626;
  assign n76435 = pi22 ? n32 : n76434;
  assign n76436 = pi21 ? n32 : n76435;
  assign n76437 = pi20 ? n76436 : n60045;
  assign n76438 = pi19 ? n32 : n76437;
  assign n76439 = pi18 ? n32 : n76438;
  assign n76440 = pi17 ? n32 : n76439;
  assign n76441 = pi16 ? n32 : n76440;
  assign n76442 = pi23 ? n63431 : n51564;
  assign n76443 = pi22 ? n32 : n76442;
  assign n76444 = pi21 ? n32 : n76443;
  assign n76445 = pi20 ? n76444 : n60045;
  assign n76446 = pi19 ? n32 : n76445;
  assign n76447 = pi18 ? n32 : n76446;
  assign n76448 = pi17 ? n32 : n76447;
  assign n76449 = pi16 ? n32 : n76448;
  assign n76450 = pi15 ? n76441 : n76449;
  assign n76451 = pi14 ? n76433 : n76450;
  assign n76452 = pi13 ? n76416 : n76451;
  assign n76453 = pi20 ? n76444 : n53984;
  assign n76454 = pi19 ? n32 : n76453;
  assign n76455 = pi18 ? n32 : n76454;
  assign n76456 = pi17 ? n32 : n76455;
  assign n76457 = pi16 ? n32 : n76456;
  assign n76458 = pi23 ? n71143 : n13481;
  assign n76459 = pi22 ? n32 : n76458;
  assign n76460 = pi21 ? n32 : n76459;
  assign n76461 = pi20 ? n76460 : n20953;
  assign n76462 = pi19 ? n32 : n76461;
  assign n76463 = pi18 ? n32 : n76462;
  assign n76464 = pi17 ? n32 : n76463;
  assign n76465 = pi16 ? n32 : n76464;
  assign n76466 = pi15 ? n76457 : n76465;
  assign n76467 = pi20 ? n73171 : n32;
  assign n76468 = pi19 ? n32 : n76467;
  assign n76469 = pi18 ? n32 : n76468;
  assign n76470 = pi17 ? n32 : n76469;
  assign n76471 = pi16 ? n32 : n76470;
  assign n76472 = pi15 ? n76471 : n32;
  assign n76473 = pi14 ? n76466 : n76472;
  assign n76474 = pi13 ? n76473 : n32;
  assign n76475 = pi12 ? n76452 : n76474;
  assign n76476 = pi11 ? n76384 : n76475;
  assign n76477 = pi10 ? n76476 : n32;
  assign n76478 = pi09 ? n76341 : n76477;
  assign n76479 = pi21 ? n30843 : n13049;
  assign n76480 = pi20 ? n32 : n76479;
  assign n76481 = pi19 ? n32 : n76480;
  assign n76482 = pi18 ? n32 : n76481;
  assign n76483 = pi17 ? n32 : n76482;
  assign n76484 = pi16 ? n32 : n76483;
  assign n76485 = pi15 ? n32 : n76484;
  assign n76486 = pi14 ? n76485 : n76336;
  assign n76487 = pi13 ? n32 : n76486;
  assign n76488 = pi12 ? n32 : n76487;
  assign n76489 = pi11 ? n32 : n76488;
  assign n76490 = pi10 ? n32 : n76489;
  assign n76491 = pi20 ? n38981 : n75156;
  assign n76492 = pi19 ? n32 : n76491;
  assign n76493 = pi18 ? n32 : n76492;
  assign n76494 = pi17 ? n32 : n76493;
  assign n76495 = pi16 ? n32 : n76494;
  assign n76496 = pi20 ? n47848 : n76352;
  assign n76497 = pi19 ? n32 : n76496;
  assign n76498 = pi18 ? n32 : n76497;
  assign n76499 = pi17 ? n32 : n76498;
  assign n76500 = pi16 ? n32 : n76499;
  assign n76501 = pi15 ? n76495 : n76500;
  assign n76502 = pi14 ? n75940 : n76501;
  assign n76503 = pi20 ? n73068 : n68542;
  assign n76504 = pi19 ? n32 : n76503;
  assign n76505 = pi18 ? n32 : n76504;
  assign n76506 = pi17 ? n32 : n76505;
  assign n76507 = pi16 ? n32 : n76506;
  assign n76508 = pi23 ? n34196 : n55567;
  assign n76509 = pi22 ? n32 : n76508;
  assign n76510 = pi21 ? n32 : n76509;
  assign n76511 = pi24 ? n33792 : n51564;
  assign n76512 = pi23 ? n76511 : n51564;
  assign n76513 = pi22 ? n76512 : n316;
  assign n76514 = pi21 ? n76513 : n54546;
  assign n76515 = pi20 ? n76510 : n76514;
  assign n76516 = pi19 ? n32 : n76515;
  assign n76517 = pi18 ? n32 : n76516;
  assign n76518 = pi17 ? n32 : n76517;
  assign n76519 = pi16 ? n32 : n76518;
  assign n76520 = pi15 ? n76507 : n76519;
  assign n76521 = pi23 ? n34196 : n62832;
  assign n76522 = pi22 ? n32 : n76521;
  assign n76523 = pi21 ? n32 : n76522;
  assign n76524 = pi20 ? n76523 : n71211;
  assign n76525 = pi19 ? n32 : n76524;
  assign n76526 = pi18 ? n32 : n76525;
  assign n76527 = pi17 ? n32 : n76526;
  assign n76528 = pi16 ? n32 : n76527;
  assign n76529 = pi20 ? n73097 : n75705;
  assign n76530 = pi19 ? n32 : n76529;
  assign n76531 = pi18 ? n32 : n76530;
  assign n76532 = pi17 ? n32 : n76531;
  assign n76533 = pi16 ? n32 : n76532;
  assign n76534 = pi15 ? n76528 : n76533;
  assign n76535 = pi14 ? n76520 : n76534;
  assign n76536 = pi13 ? n76502 : n76535;
  assign n76537 = pi12 ? n75940 : n76536;
  assign n76538 = pi20 ? n73111 : n76386;
  assign n76539 = pi19 ? n32 : n76538;
  assign n76540 = pi18 ? n32 : n76539;
  assign n76541 = pi17 ? n32 : n76540;
  assign n76542 = pi16 ? n32 : n76541;
  assign n76543 = pi20 ? n73111 : n74807;
  assign n76544 = pi19 ? n32 : n76543;
  assign n76545 = pi18 ? n32 : n76544;
  assign n76546 = pi17 ? n32 : n76545;
  assign n76547 = pi16 ? n32 : n76546;
  assign n76548 = pi15 ? n76542 : n76547;
  assign n76549 = pi20 ? n52863 : n76401;
  assign n76550 = pi19 ? n32 : n76549;
  assign n76551 = pi18 ? n32 : n76550;
  assign n76552 = pi17 ? n32 : n76551;
  assign n76553 = pi16 ? n32 : n76552;
  assign n76554 = pi20 ? n52872 : n72747;
  assign n76555 = pi19 ? n32 : n76554;
  assign n76556 = pi18 ? n32 : n76555;
  assign n76557 = pi17 ? n32 : n76556;
  assign n76558 = pi16 ? n32 : n76557;
  assign n76559 = pi15 ? n76553 : n76558;
  assign n76560 = pi14 ? n76548 : n76559;
  assign n76561 = pi20 ? n52872 : n72062;
  assign n76562 = pi19 ? n32 : n76561;
  assign n76563 = pi18 ? n32 : n76562;
  assign n76564 = pi17 ? n32 : n76563;
  assign n76565 = pi16 ? n32 : n76564;
  assign n76566 = pi21 ? n32 : n74679;
  assign n76567 = pi20 ? n76566 : n3210;
  assign n76568 = pi19 ? n32 : n76567;
  assign n76569 = pi18 ? n32 : n76568;
  assign n76570 = pi17 ? n32 : n76569;
  assign n76571 = pi16 ? n32 : n76570;
  assign n76572 = pi15 ? n76565 : n76571;
  assign n76573 = pi20 ? n76566 : n60045;
  assign n76574 = pi19 ? n32 : n76573;
  assign n76575 = pi18 ? n32 : n76574;
  assign n76576 = pi17 ? n32 : n76575;
  assign n76577 = pi16 ? n32 : n76576;
  assign n76578 = pi21 ? n32 : n74462;
  assign n76579 = pi20 ? n76578 : n37640;
  assign n76580 = pi19 ? n32 : n76579;
  assign n76581 = pi18 ? n32 : n76580;
  assign n76582 = pi17 ? n32 : n76581;
  assign n76583 = pi16 ? n32 : n76582;
  assign n76584 = pi15 ? n76577 : n76583;
  assign n76585 = pi14 ? n76572 : n76584;
  assign n76586 = pi13 ? n76560 : n76585;
  assign n76587 = pi20 ? n76578 : n53984;
  assign n76588 = pi19 ? n32 : n76587;
  assign n76589 = pi18 ? n32 : n76588;
  assign n76590 = pi17 ? n32 : n76589;
  assign n76591 = pi16 ? n32 : n76590;
  assign n76592 = pi21 ? n32 : n71558;
  assign n76593 = pi20 ? n76592 : n32;
  assign n76594 = pi19 ? n32 : n76593;
  assign n76595 = pi18 ? n32 : n76594;
  assign n76596 = pi17 ? n32 : n76595;
  assign n76597 = pi16 ? n32 : n76596;
  assign n76598 = pi15 ? n76591 : n76597;
  assign n76599 = pi14 ? n76598 : n32;
  assign n76600 = pi13 ? n76599 : n32;
  assign n76601 = pi12 ? n76586 : n76600;
  assign n76602 = pi11 ? n76537 : n76601;
  assign n76603 = pi10 ? n76602 : n32;
  assign n76604 = pi09 ? n76490 : n76603;
  assign n76605 = pi08 ? n76478 : n76604;
  assign n76606 = pi20 ? n32 : n61008;
  assign n76607 = pi19 ? n32 : n76606;
  assign n76608 = pi18 ? n32 : n76607;
  assign n76609 = pi17 ? n32 : n76608;
  assign n76610 = pi16 ? n32 : n76609;
  assign n76611 = pi14 ? n76485 : n76610;
  assign n76612 = pi13 ? n32 : n76611;
  assign n76613 = pi12 ? n32 : n76612;
  assign n76614 = pi11 ? n32 : n76613;
  assign n76615 = pi10 ? n32 : n76614;
  assign n76616 = pi15 ? n76336 : n75940;
  assign n76617 = pi20 ? n47848 : n61008;
  assign n76618 = pi19 ? n32 : n76617;
  assign n76619 = pi18 ? n32 : n76618;
  assign n76620 = pi17 ? n32 : n76619;
  assign n76621 = pi16 ? n32 : n76620;
  assign n76622 = pi15 ? n75940 : n76621;
  assign n76623 = pi14 ? n76616 : n76622;
  assign n76624 = pi13 ? n76336 : n76623;
  assign n76625 = pi20 ? n47848 : n68542;
  assign n76626 = pi19 ? n32 : n76625;
  assign n76627 = pi18 ? n32 : n76626;
  assign n76628 = pi17 ? n32 : n76627;
  assign n76629 = pi16 ? n32 : n76628;
  assign n76630 = pi23 ? n32 : n55567;
  assign n76631 = pi22 ? n32 : n76630;
  assign n76632 = pi21 ? n32 : n76631;
  assign n76633 = pi20 ? n76632 : n75366;
  assign n76634 = pi19 ? n32 : n76633;
  assign n76635 = pi18 ? n32 : n76634;
  assign n76636 = pi17 ? n32 : n76635;
  assign n76637 = pi16 ? n32 : n76636;
  assign n76638 = pi15 ? n76629 : n76637;
  assign n76639 = pi23 ? n32 : n55580;
  assign n76640 = pi22 ? n32 : n76639;
  assign n76641 = pi21 ? n32 : n76640;
  assign n76642 = pi20 ? n76641 : n71211;
  assign n76643 = pi19 ? n32 : n76642;
  assign n76644 = pi18 ? n32 : n76643;
  assign n76645 = pi17 ? n32 : n76644;
  assign n76646 = pi16 ? n32 : n76645;
  assign n76647 = pi20 ? n73358 : n75549;
  assign n76648 = pi19 ? n32 : n76647;
  assign n76649 = pi18 ? n32 : n76648;
  assign n76650 = pi17 ? n32 : n76649;
  assign n76651 = pi16 ? n32 : n76650;
  assign n76652 = pi15 ? n76646 : n76651;
  assign n76653 = pi14 ? n76638 : n76652;
  assign n76654 = pi13 ? n76502 : n76653;
  assign n76655 = pi12 ? n76624 : n76654;
  assign n76656 = pi21 ? n58913 : n928;
  assign n76657 = pi20 ? n73358 : n76656;
  assign n76658 = pi19 ? n32 : n76657;
  assign n76659 = pi18 ? n32 : n76658;
  assign n76660 = pi17 ? n32 : n76659;
  assign n76661 = pi16 ? n32 : n76660;
  assign n76662 = pi20 ? n70297 : n74807;
  assign n76663 = pi19 ? n32 : n76662;
  assign n76664 = pi18 ? n32 : n76663;
  assign n76665 = pi17 ? n32 : n76664;
  assign n76666 = pi16 ? n32 : n76665;
  assign n76667 = pi15 ? n76661 : n76666;
  assign n76668 = pi22 ? n73960 : n59672;
  assign n76669 = pi21 ? n76668 : n32;
  assign n76670 = pi20 ? n52918 : n76669;
  assign n76671 = pi19 ? n32 : n76670;
  assign n76672 = pi18 ? n32 : n76671;
  assign n76673 = pi17 ? n32 : n76672;
  assign n76674 = pi16 ? n32 : n76673;
  assign n76675 = pi23 ? n63431 : n43198;
  assign n76676 = pi22 ? n32 : n76675;
  assign n76677 = pi21 ? n32 : n76676;
  assign n76678 = pi22 ? n75217 : n396;
  assign n76679 = pi21 ? n76678 : n32;
  assign n76680 = pi20 ? n76677 : n76679;
  assign n76681 = pi19 ? n32 : n76680;
  assign n76682 = pi18 ? n32 : n76681;
  assign n76683 = pi17 ? n32 : n76682;
  assign n76684 = pi16 ? n32 : n76683;
  assign n76685 = pi15 ? n76674 : n76684;
  assign n76686 = pi14 ? n76667 : n76685;
  assign n76687 = pi21 ? n32 : n74906;
  assign n76688 = pi20 ? n76687 : n67728;
  assign n76689 = pi19 ? n32 : n76688;
  assign n76690 = pi18 ? n32 : n76689;
  assign n76691 = pi17 ? n32 : n76690;
  assign n76692 = pi16 ? n32 : n76691;
  assign n76693 = pi20 ? n76687 : n3210;
  assign n76694 = pi19 ? n32 : n76693;
  assign n76695 = pi18 ? n32 : n76694;
  assign n76696 = pi17 ? n32 : n76695;
  assign n76697 = pi16 ? n32 : n76696;
  assign n76698 = pi15 ? n76692 : n76697;
  assign n76699 = pi20 ? n73124 : n60045;
  assign n76700 = pi19 ? n32 : n76699;
  assign n76701 = pi18 ? n32 : n76700;
  assign n76702 = pi17 ? n32 : n76701;
  assign n76703 = pi16 ? n32 : n76702;
  assign n76704 = pi20 ? n69892 : n37640;
  assign n76705 = pi19 ? n32 : n76704;
  assign n76706 = pi18 ? n32 : n76705;
  assign n76707 = pi17 ? n32 : n76706;
  assign n76708 = pi16 ? n32 : n76707;
  assign n76709 = pi15 ? n76703 : n76708;
  assign n76710 = pi14 ? n76698 : n76709;
  assign n76711 = pi13 ? n76686 : n76710;
  assign n76712 = pi19 ? n32 : n69893;
  assign n76713 = pi18 ? n32 : n76712;
  assign n76714 = pi17 ? n32 : n76713;
  assign n76715 = pi16 ? n32 : n76714;
  assign n76716 = pi15 ? n76715 : n32;
  assign n76717 = pi14 ? n76716 : n32;
  assign n76718 = pi13 ? n76717 : n32;
  assign n76719 = pi12 ? n76711 : n76718;
  assign n76720 = pi11 ? n76655 : n76719;
  assign n76721 = pi10 ? n76720 : n32;
  assign n76722 = pi09 ? n76615 : n76721;
  assign n76723 = pi21 ? n180 : n13049;
  assign n76724 = pi20 ? n32 : n76723;
  assign n76725 = pi19 ? n32 : n76724;
  assign n76726 = pi18 ? n32 : n76725;
  assign n76727 = pi17 ? n32 : n76726;
  assign n76728 = pi16 ? n32 : n76727;
  assign n76729 = pi15 ? n32 : n76728;
  assign n76730 = pi14 ? n76729 : n76610;
  assign n76731 = pi13 ? n32 : n76730;
  assign n76732 = pi12 ? n32 : n76731;
  assign n76733 = pi11 ? n32 : n76732;
  assign n76734 = pi10 ? n32 : n76733;
  assign n76735 = pi14 ? n76336 : n76610;
  assign n76736 = pi15 ? n76610 : n76336;
  assign n76737 = pi14 ? n76736 : n76212;
  assign n76738 = pi13 ? n76735 : n76737;
  assign n76739 = pi20 ? n47835 : n75156;
  assign n76740 = pi19 ? n32 : n76739;
  assign n76741 = pi18 ? n32 : n76740;
  assign n76742 = pi17 ? n32 : n76741;
  assign n76743 = pi16 ? n32 : n76742;
  assign n76744 = pi20 ? n73367 : n76352;
  assign n76745 = pi19 ? n32 : n76744;
  assign n76746 = pi18 ? n32 : n76745;
  assign n76747 = pi17 ? n32 : n76746;
  assign n76748 = pi16 ? n32 : n76747;
  assign n76749 = pi15 ? n76743 : n76748;
  assign n76750 = pi14 ? n76336 : n76749;
  assign n76751 = pi20 ? n73367 : n72359;
  assign n76752 = pi19 ? n32 : n76751;
  assign n76753 = pi18 ? n32 : n76752;
  assign n76754 = pi17 ? n32 : n76753;
  assign n76755 = pi16 ? n32 : n76754;
  assign n76756 = pi20 ? n48846 : n71984;
  assign n76757 = pi19 ? n32 : n76756;
  assign n76758 = pi18 ? n32 : n76757;
  assign n76759 = pi17 ? n32 : n76758;
  assign n76760 = pi16 ? n32 : n76759;
  assign n76761 = pi15 ? n76755 : n76760;
  assign n76762 = pi20 ? n73358 : n75705;
  assign n76763 = pi19 ? n32 : n76762;
  assign n76764 = pi18 ? n32 : n76763;
  assign n76765 = pi17 ? n32 : n76764;
  assign n76766 = pi16 ? n32 : n76765;
  assign n76767 = pi15 ? n76760 : n76766;
  assign n76768 = pi14 ? n76761 : n76767;
  assign n76769 = pi13 ? n76750 : n76768;
  assign n76770 = pi12 ? n76738 : n76769;
  assign n76771 = pi20 ? n70297 : n73278;
  assign n76772 = pi19 ? n32 : n76771;
  assign n76773 = pi18 ? n32 : n76772;
  assign n76774 = pi17 ? n32 : n76773;
  assign n76775 = pi16 ? n32 : n76774;
  assign n76776 = pi15 ? n76661 : n76775;
  assign n76777 = pi22 ? n74206 : n59672;
  assign n76778 = pi21 ? n76777 : n32;
  assign n76779 = pi20 ? n52918 : n76778;
  assign n76780 = pi19 ? n32 : n76779;
  assign n76781 = pi18 ? n32 : n76780;
  assign n76782 = pi17 ? n32 : n76781;
  assign n76783 = pi16 ? n32 : n76782;
  assign n76784 = pi20 ? n52918 : n76679;
  assign n76785 = pi19 ? n32 : n76784;
  assign n76786 = pi18 ? n32 : n76785;
  assign n76787 = pi17 ? n32 : n76786;
  assign n76788 = pi16 ? n32 : n76787;
  assign n76789 = pi15 ? n76783 : n76788;
  assign n76790 = pi14 ? n76776 : n76789;
  assign n76791 = pi20 ? n69892 : n60045;
  assign n76792 = pi19 ? n32 : n76791;
  assign n76793 = pi18 ? n32 : n76792;
  assign n76794 = pi17 ? n32 : n76793;
  assign n76795 = pi16 ? n32 : n76794;
  assign n76796 = pi23 ? n32 : n3690;
  assign n76797 = pi22 ? n32 : n76796;
  assign n76798 = pi21 ? n32 : n76797;
  assign n76799 = pi20 ? n76798 : n37640;
  assign n76800 = pi19 ? n32 : n76799;
  assign n76801 = pi18 ? n32 : n76800;
  assign n76802 = pi17 ? n32 : n76801;
  assign n76803 = pi16 ? n32 : n76802;
  assign n76804 = pi15 ? n76795 : n76803;
  assign n76805 = pi14 ? n76698 : n76804;
  assign n76806 = pi13 ? n76790 : n76805;
  assign n76807 = pi20 ? n70314 : n20953;
  assign n76808 = pi19 ? n32 : n76807;
  assign n76809 = pi18 ? n32 : n76808;
  assign n76810 = pi17 ? n32 : n76809;
  assign n76811 = pi16 ? n32 : n76810;
  assign n76812 = pi15 ? n76811 : n32;
  assign n76813 = pi14 ? n76812 : n32;
  assign n76814 = pi13 ? n76813 : n32;
  assign n76815 = pi12 ? n76806 : n76814;
  assign n76816 = pi11 ? n76770 : n76815;
  assign n76817 = pi10 ? n76816 : n32;
  assign n76818 = pi09 ? n76734 : n76817;
  assign n76819 = pi08 ? n76722 : n76818;
  assign n76820 = pi07 ? n76605 : n76819;
  assign n76821 = pi21 ? n34011 : n13049;
  assign n76822 = pi20 ? n32 : n76821;
  assign n76823 = pi19 ? n32 : n76822;
  assign n76824 = pi18 ? n32 : n76823;
  assign n76825 = pi17 ? n32 : n76824;
  assign n76826 = pi16 ? n32 : n76825;
  assign n76827 = pi15 ? n32 : n76826;
  assign n76828 = pi21 ? n180 : n1618;
  assign n76829 = pi20 ? n32 : n76828;
  assign n76830 = pi19 ? n32 : n76829;
  assign n76831 = pi18 ? n32 : n76830;
  assign n76832 = pi17 ? n32 : n76831;
  assign n76833 = pi16 ? n32 : n76832;
  assign n76834 = pi14 ? n76827 : n76833;
  assign n76835 = pi13 ? n32 : n76834;
  assign n76836 = pi12 ? n32 : n76835;
  assign n76837 = pi11 ? n32 : n76836;
  assign n76838 = pi10 ? n32 : n76837;
  assign n76839 = pi20 ? n32 : n66577;
  assign n76840 = pi19 ? n32 : n76839;
  assign n76841 = pi18 ? n32 : n76840;
  assign n76842 = pi17 ? n32 : n76841;
  assign n76843 = pi16 ? n32 : n76842;
  assign n76844 = pi21 ? n30843 : n1618;
  assign n76845 = pi20 ? n32 : n76844;
  assign n76846 = pi19 ? n32 : n76845;
  assign n76847 = pi18 ? n32 : n76846;
  assign n76848 = pi17 ? n32 : n76847;
  assign n76849 = pi16 ? n32 : n76848;
  assign n76850 = pi15 ? n76843 : n76849;
  assign n76851 = pi14 ? n76843 : n76850;
  assign n76852 = pi21 ? n37231 : n1618;
  assign n76853 = pi20 ? n32 : n76852;
  assign n76854 = pi19 ? n32 : n76853;
  assign n76855 = pi18 ? n32 : n76854;
  assign n76856 = pi17 ? n32 : n76855;
  assign n76857 = pi16 ? n32 : n76856;
  assign n76858 = pi15 ? n76857 : n76849;
  assign n76859 = pi20 ? n37926 : n66577;
  assign n76860 = pi19 ? n32 : n76859;
  assign n76861 = pi18 ? n32 : n76860;
  assign n76862 = pi17 ? n32 : n76861;
  assign n76863 = pi16 ? n32 : n76862;
  assign n76864 = pi15 ? n76863 : n76336;
  assign n76865 = pi14 ? n76858 : n76864;
  assign n76866 = pi13 ? n76851 : n76865;
  assign n76867 = pi21 ? n36516 : n1618;
  assign n76868 = pi20 ? n47835 : n76867;
  assign n76869 = pi19 ? n32 : n76868;
  assign n76870 = pi18 ? n32 : n76869;
  assign n76871 = pi17 ? n32 : n76870;
  assign n76872 = pi16 ? n32 : n76871;
  assign n76873 = pi15 ? n76872 : n76748;
  assign n76874 = pi14 ? n76863 : n76873;
  assign n76875 = pi20 ? n46201 : n71211;
  assign n76876 = pi19 ? n32 : n76875;
  assign n76877 = pi18 ? n32 : n76876;
  assign n76878 = pi17 ? n32 : n76877;
  assign n76879 = pi16 ? n32 : n76878;
  assign n76880 = pi15 ? n76755 : n76879;
  assign n76881 = pi23 ? n71981 : n13481;
  assign n76882 = pi22 ? n76881 : n13481;
  assign n76883 = pi21 ? n76882 : n55667;
  assign n76884 = pi20 ? n32 : n76883;
  assign n76885 = pi19 ? n32 : n76884;
  assign n76886 = pi18 ? n32 : n76885;
  assign n76887 = pi17 ? n32 : n76886;
  assign n76888 = pi16 ? n32 : n76887;
  assign n76889 = pi23 ? n62628 : n51564;
  assign n76890 = pi22 ? n76889 : n316;
  assign n76891 = pi21 ? n76890 : n59357;
  assign n76892 = pi20 ? n46201 : n76891;
  assign n76893 = pi19 ? n32 : n76892;
  assign n76894 = pi18 ? n32 : n76893;
  assign n76895 = pi17 ? n32 : n76894;
  assign n76896 = pi16 ? n32 : n76895;
  assign n76897 = pi15 ? n76888 : n76896;
  assign n76898 = pi14 ? n76880 : n76897;
  assign n76899 = pi13 ? n76874 : n76898;
  assign n76900 = pi12 ? n76866 : n76899;
  assign n76901 = pi23 ? n32 : n4262;
  assign n76902 = pi22 ? n32 : n76901;
  assign n76903 = pi21 ? n32 : n76902;
  assign n76904 = pi21 ? n62079 : n37639;
  assign n76905 = pi20 ? n76903 : n76904;
  assign n76906 = pi19 ? n32 : n76905;
  assign n76907 = pi18 ? n32 : n76906;
  assign n76908 = pi17 ? n32 : n76907;
  assign n76909 = pi16 ? n32 : n76908;
  assign n76910 = pi22 ? n65231 : n13481;
  assign n76911 = pi21 ? n76910 : n37639;
  assign n76912 = pi20 ? n52918 : n76911;
  assign n76913 = pi19 ? n32 : n76912;
  assign n76914 = pi18 ? n32 : n76913;
  assign n76915 = pi17 ? n32 : n76914;
  assign n76916 = pi16 ? n32 : n76915;
  assign n76917 = pi15 ? n76909 : n76916;
  assign n76918 = pi23 ? n70599 : n13481;
  assign n76919 = pi22 ? n76918 : n55688;
  assign n76920 = pi21 ? n76919 : n32;
  assign n76921 = pi20 ? n76687 : n76920;
  assign n76922 = pi19 ? n32 : n76921;
  assign n76923 = pi18 ? n32 : n76922;
  assign n76924 = pi17 ? n32 : n76923;
  assign n76925 = pi16 ? n32 : n76924;
  assign n76926 = pi14 ? n76917 : n76925;
  assign n76927 = pi20 ? n73408 : n55668;
  assign n76928 = pi19 ? n32 : n76927;
  assign n76929 = pi18 ? n32 : n76928;
  assign n76930 = pi17 ? n32 : n76929;
  assign n76931 = pi16 ? n32 : n76930;
  assign n76932 = pi20 ? n73408 : n60045;
  assign n76933 = pi19 ? n32 : n76932;
  assign n76934 = pi18 ? n32 : n76933;
  assign n76935 = pi17 ? n32 : n76934;
  assign n76936 = pi16 ? n32 : n76935;
  assign n76937 = pi15 ? n76931 : n76936;
  assign n76938 = pi20 ? n73416 : n37640;
  assign n76939 = pi19 ? n32 : n76938;
  assign n76940 = pi18 ? n32 : n76939;
  assign n76941 = pi17 ? n32 : n76940;
  assign n76942 = pi16 ? n32 : n76941;
  assign n76943 = pi20 ? n76798 : n1822;
  assign n76944 = pi19 ? n32 : n76943;
  assign n76945 = pi18 ? n32 : n76944;
  assign n76946 = pi17 ? n32 : n76945;
  assign n76947 = pi16 ? n32 : n76946;
  assign n76948 = pi15 ? n76942 : n76947;
  assign n76949 = pi14 ? n76937 : n76948;
  assign n76950 = pi13 ? n76926 : n76949;
  assign n76951 = pi12 ? n76950 : n32;
  assign n76952 = pi11 ? n76900 : n76951;
  assign n76953 = pi10 ? n76952 : n32;
  assign n76954 = pi09 ? n76838 : n76953;
  assign n76955 = pi15 ? n76843 : n76833;
  assign n76956 = pi14 ? n76843 : n76955;
  assign n76957 = pi15 ? n76857 : n76833;
  assign n76958 = pi14 ? n76957 : n76864;
  assign n76959 = pi13 ? n76956 : n76958;
  assign n76960 = pi20 ? n47835 : n66577;
  assign n76961 = pi19 ? n32 : n76960;
  assign n76962 = pi18 ? n32 : n76961;
  assign n76963 = pi17 ? n32 : n76962;
  assign n76964 = pi16 ? n32 : n76963;
  assign n76965 = pi15 ? n76964 : n76843;
  assign n76966 = pi20 ? n32 : n76867;
  assign n76967 = pi19 ? n32 : n76966;
  assign n76968 = pi18 ? n32 : n76967;
  assign n76969 = pi17 ? n32 : n76968;
  assign n76970 = pi16 ? n32 : n76969;
  assign n76971 = pi20 ? n32 : n76352;
  assign n76972 = pi19 ? n32 : n76971;
  assign n76973 = pi18 ? n32 : n76972;
  assign n76974 = pi17 ? n32 : n76973;
  assign n76975 = pi16 ? n32 : n76974;
  assign n76976 = pi15 ? n76970 : n76975;
  assign n76977 = pi14 ? n76965 : n76976;
  assign n76978 = pi20 ? n32 : n72359;
  assign n76979 = pi19 ? n32 : n76978;
  assign n76980 = pi18 ? n32 : n76979;
  assign n76981 = pi17 ? n32 : n76980;
  assign n76982 = pi16 ? n32 : n76981;
  assign n76983 = pi20 ? n32 : n71211;
  assign n76984 = pi19 ? n32 : n76983;
  assign n76985 = pi18 ? n32 : n76984;
  assign n76986 = pi17 ? n32 : n76985;
  assign n76987 = pi16 ? n32 : n76986;
  assign n76988 = pi15 ? n76982 : n76987;
  assign n76989 = pi21 ? n72987 : n56129;
  assign n76990 = pi20 ? n32 : n76989;
  assign n76991 = pi19 ? n32 : n76990;
  assign n76992 = pi18 ? n32 : n76991;
  assign n76993 = pi17 ? n32 : n76992;
  assign n76994 = pi16 ? n32 : n76993;
  assign n76995 = pi20 ? n32 : n76386;
  assign n76996 = pi19 ? n32 : n76995;
  assign n76997 = pi18 ? n32 : n76996;
  assign n76998 = pi17 ? n32 : n76997;
  assign n76999 = pi16 ? n32 : n76998;
  assign n77000 = pi15 ? n76994 : n76999;
  assign n77001 = pi14 ? n76988 : n77000;
  assign n77002 = pi13 ? n76977 : n77001;
  assign n77003 = pi12 ? n76959 : n77002;
  assign n77004 = pi24 ? n157 : n13481;
  assign n77005 = pi23 ? n77004 : n13481;
  assign n77006 = pi22 ? n77005 : n13481;
  assign n77007 = pi21 ? n77006 : n37639;
  assign n77008 = pi20 ? n76903 : n77007;
  assign n77009 = pi19 ? n32 : n77008;
  assign n77010 = pi18 ? n32 : n77009;
  assign n77011 = pi17 ? n32 : n77010;
  assign n77012 = pi16 ? n32 : n77011;
  assign n77013 = pi20 ? n46277 : n76001;
  assign n77014 = pi19 ? n32 : n77013;
  assign n77015 = pi18 ? n32 : n77014;
  assign n77016 = pi17 ? n32 : n77015;
  assign n77017 = pi16 ? n32 : n77016;
  assign n77018 = pi15 ? n77012 : n77017;
  assign n77019 = pi23 ? n32 : n3719;
  assign n77020 = pi22 ? n32 : n77019;
  assign n77021 = pi21 ? n32 : n77020;
  assign n77022 = pi22 ? n71897 : n56665;
  assign n77023 = pi21 ? n77022 : n32;
  assign n77024 = pi20 ? n77021 : n77023;
  assign n77025 = pi19 ? n32 : n77024;
  assign n77026 = pi18 ? n32 : n77025;
  assign n77027 = pi17 ? n32 : n77026;
  assign n77028 = pi16 ? n32 : n77027;
  assign n77029 = pi22 ? n75573 : n56665;
  assign n77030 = pi21 ? n77029 : n32;
  assign n77031 = pi20 ? n73408 : n77030;
  assign n77032 = pi19 ? n32 : n77031;
  assign n77033 = pi18 ? n32 : n77032;
  assign n77034 = pi17 ? n32 : n77033;
  assign n77035 = pi16 ? n32 : n77034;
  assign n77036 = pi15 ? n77028 : n77035;
  assign n77037 = pi14 ? n77018 : n77036;
  assign n77038 = pi20 ? n73408 : n56130;
  assign n77039 = pi19 ? n32 : n77038;
  assign n77040 = pi18 ? n32 : n77039;
  assign n77041 = pi17 ? n32 : n77040;
  assign n77042 = pi16 ? n32 : n77041;
  assign n77043 = pi24 ? n32 : n685;
  assign n77044 = pi23 ? n32 : n77043;
  assign n77045 = pi22 ? n32 : n77044;
  assign n77046 = pi21 ? n32 : n77045;
  assign n77047 = pi20 ? n77046 : n60045;
  assign n77048 = pi19 ? n32 : n77047;
  assign n77049 = pi18 ? n32 : n77048;
  assign n77050 = pi17 ? n32 : n77049;
  assign n77051 = pi16 ? n32 : n77050;
  assign n77052 = pi15 ? n77042 : n77051;
  assign n77053 = pi19 ? n32 : n70331;
  assign n77054 = pi18 ? n32 : n77053;
  assign n77055 = pi17 ? n32 : n77054;
  assign n77056 = pi16 ? n32 : n77055;
  assign n77057 = pi15 ? n77056 : n76811;
  assign n77058 = pi14 ? n77052 : n77057;
  assign n77059 = pi13 ? n77037 : n77058;
  assign n77060 = pi12 ? n77059 : n32;
  assign n77061 = pi11 ? n77003 : n77060;
  assign n77062 = pi10 ? n77061 : n32;
  assign n77063 = pi09 ? n76838 : n77062;
  assign n77064 = pi08 ? n76954 : n77063;
  assign n77065 = pi21 ? n65 : n13049;
  assign n77066 = pi20 ? n32 : n77065;
  assign n77067 = pi19 ? n32 : n77066;
  assign n77068 = pi18 ? n32 : n77067;
  assign n77069 = pi17 ? n32 : n77068;
  assign n77070 = pi16 ? n32 : n77069;
  assign n77071 = pi15 ? n32 : n77070;
  assign n77072 = pi14 ? n77071 : n76833;
  assign n77073 = pi13 ? n32 : n77072;
  assign n77074 = pi12 ? n32 : n77073;
  assign n77075 = pi11 ? n32 : n77074;
  assign n77076 = pi10 ? n32 : n77075;
  assign n77077 = pi15 ? n76849 : n76610;
  assign n77078 = pi14 ? n76833 : n77077;
  assign n77079 = pi13 ? n76833 : n77078;
  assign n77080 = pi15 ? n76849 : n76970;
  assign n77081 = pi21 ? n48221 : n1618;
  assign n77082 = pi20 ? n32 : n77081;
  assign n77083 = pi19 ? n32 : n77082;
  assign n77084 = pi18 ? n32 : n77083;
  assign n77085 = pi17 ? n32 : n77084;
  assign n77086 = pi16 ? n32 : n77085;
  assign n77087 = pi15 ? n77086 : n76975;
  assign n77088 = pi14 ? n77080 : n77087;
  assign n77089 = pi24 ? n36659 : n685;
  assign n77090 = pi23 ? n77089 : n685;
  assign n77091 = pi22 ? n77090 : n685;
  assign n77092 = pi21 ? n77091 : n696;
  assign n77093 = pi20 ? n32 : n77092;
  assign n77094 = pi19 ? n32 : n77093;
  assign n77095 = pi18 ? n32 : n77094;
  assign n77096 = pi17 ? n32 : n77095;
  assign n77097 = pi16 ? n32 : n77096;
  assign n77098 = pi20 ? n32 : n71984;
  assign n77099 = pi19 ? n32 : n77098;
  assign n77100 = pi18 ? n32 : n77099;
  assign n77101 = pi17 ? n32 : n77100;
  assign n77102 = pi16 ? n32 : n77101;
  assign n77103 = pi15 ? n77097 : n77102;
  assign n77104 = pi23 ? n71143 : n316;
  assign n77105 = pi22 ? n77104 : n316;
  assign n77106 = pi21 ? n77105 : n928;
  assign n77107 = pi20 ? n32 : n77106;
  assign n77108 = pi19 ? n32 : n77107;
  assign n77109 = pi18 ? n32 : n77108;
  assign n77110 = pi17 ? n32 : n77109;
  assign n77111 = pi16 ? n32 : n77110;
  assign n77112 = pi15 ? n76994 : n77111;
  assign n77113 = pi14 ? n77103 : n77112;
  assign n77114 = pi13 ? n77088 : n77113;
  assign n77115 = pi12 ? n77079 : n77114;
  assign n77116 = pi21 ? n62647 : n37639;
  assign n77117 = pi20 ? n46225 : n77116;
  assign n77118 = pi19 ? n32 : n77117;
  assign n77119 = pi18 ? n32 : n77118;
  assign n77120 = pi17 ? n32 : n77119;
  assign n77121 = pi16 ? n32 : n77120;
  assign n77122 = pi22 ? n62427 : n13481;
  assign n77123 = pi21 ? n77122 : n37639;
  assign n77124 = pi20 ? n46277 : n77123;
  assign n77125 = pi19 ? n32 : n77124;
  assign n77126 = pi18 ? n32 : n77125;
  assign n77127 = pi17 ? n32 : n77126;
  assign n77128 = pi16 ? n32 : n77127;
  assign n77129 = pi15 ? n77121 : n77128;
  assign n77130 = pi22 ? n62427 : n56665;
  assign n77131 = pi21 ? n77130 : n32;
  assign n77132 = pi20 ? n46277 : n77131;
  assign n77133 = pi19 ? n32 : n77132;
  assign n77134 = pi18 ? n32 : n77133;
  assign n77135 = pi17 ? n32 : n77134;
  assign n77136 = pi16 ? n32 : n77135;
  assign n77137 = pi22 ? n73977 : n56665;
  assign n77138 = pi21 ? n77137 : n32;
  assign n77139 = pi20 ? n73408 : n77138;
  assign n77140 = pi19 ? n32 : n77139;
  assign n77141 = pi18 ? n32 : n77140;
  assign n77142 = pi17 ? n32 : n77141;
  assign n77143 = pi16 ? n32 : n77142;
  assign n77144 = pi15 ? n77136 : n77143;
  assign n77145 = pi14 ? n77129 : n77144;
  assign n77146 = pi20 ? n32 : n56130;
  assign n77147 = pi19 ? n32 : n77146;
  assign n77148 = pi18 ? n32 : n77147;
  assign n77149 = pi17 ? n32 : n77148;
  assign n77150 = pi16 ? n32 : n77149;
  assign n77151 = pi19 ? n32 : n70326;
  assign n77152 = pi18 ? n32 : n77151;
  assign n77153 = pi17 ? n32 : n77152;
  assign n77154 = pi16 ? n32 : n77153;
  assign n77155 = pi15 ? n77150 : n77154;
  assign n77156 = pi14 ? n77155 : n77057;
  assign n77157 = pi13 ? n77145 : n77156;
  assign n77158 = pi12 ? n77157 : n32;
  assign n77159 = pi11 ? n77115 : n77158;
  assign n77160 = pi10 ? n77159 : n32;
  assign n77161 = pi09 ? n77076 : n77160;
  assign n77162 = pi15 ? n76833 : n76610;
  assign n77163 = pi14 ? n76833 : n77162;
  assign n77164 = pi13 ? n76833 : n77163;
  assign n77165 = pi15 ? n76833 : n76970;
  assign n77166 = pi14 ? n77165 : n77087;
  assign n77167 = pi23 ? n77043 : n685;
  assign n77168 = pi22 ? n77167 : n685;
  assign n77169 = pi21 ? n77168 : n696;
  assign n77170 = pi20 ? n32 : n77169;
  assign n77171 = pi19 ? n32 : n77170;
  assign n77172 = pi18 ? n32 : n77171;
  assign n77173 = pi17 ? n32 : n77172;
  assign n77174 = pi16 ? n32 : n77173;
  assign n77175 = pi15 ? n77174 : n77102;
  assign n77176 = pi22 ? n71924 : n13481;
  assign n77177 = pi21 ? n77176 : n56129;
  assign n77178 = pi20 ? n32 : n77177;
  assign n77179 = pi19 ? n32 : n77178;
  assign n77180 = pi18 ? n32 : n77179;
  assign n77181 = pi17 ? n32 : n77180;
  assign n77182 = pi16 ? n32 : n77181;
  assign n77183 = pi21 ? n8440 : n928;
  assign n77184 = pi20 ? n32 : n77183;
  assign n77185 = pi19 ? n32 : n77184;
  assign n77186 = pi18 ? n32 : n77185;
  assign n77187 = pi17 ? n32 : n77186;
  assign n77188 = pi16 ? n32 : n77187;
  assign n77189 = pi15 ? n77182 : n77188;
  assign n77190 = pi14 ? n77175 : n77189;
  assign n77191 = pi13 ? n77166 : n77190;
  assign n77192 = pi12 ? n77164 : n77191;
  assign n77193 = pi20 ? n32 : n77116;
  assign n77194 = pi19 ? n32 : n77193;
  assign n77195 = pi18 ? n32 : n77194;
  assign n77196 = pi17 ? n32 : n77195;
  assign n77197 = pi16 ? n32 : n77196;
  assign n77198 = pi21 ? n76910 : n32;
  assign n77199 = pi20 ? n32 : n77198;
  assign n77200 = pi19 ? n32 : n77199;
  assign n77201 = pi18 ? n32 : n77200;
  assign n77202 = pi17 ? n32 : n77201;
  assign n77203 = pi16 ? n32 : n77202;
  assign n77204 = pi15 ? n77197 : n77203;
  assign n77205 = pi22 ? n59784 : n14363;
  assign n77206 = pi21 ? n77205 : n32;
  assign n77207 = pi20 ? n32 : n77206;
  assign n77208 = pi19 ? n32 : n77207;
  assign n77209 = pi18 ? n32 : n77208;
  assign n77210 = pi17 ? n32 : n77209;
  assign n77211 = pi16 ? n32 : n77210;
  assign n77212 = pi15 ? n77136 : n77211;
  assign n77213 = pi14 ? n77204 : n77212;
  assign n77214 = pi15 ? n77154 : n77056;
  assign n77215 = pi20 ? n32 : n20953;
  assign n77216 = pi19 ? n32 : n77215;
  assign n77217 = pi18 ? n32 : n77216;
  assign n77218 = pi17 ? n32 : n77217;
  assign n77219 = pi16 ? n32 : n77218;
  assign n77220 = pi15 ? n77219 : n32;
  assign n77221 = pi14 ? n77214 : n77220;
  assign n77222 = pi13 ? n77213 : n77221;
  assign n77223 = pi12 ? n77222 : n32;
  assign n77224 = pi11 ? n77192 : n77223;
  assign n77225 = pi10 ? n77224 : n32;
  assign n77226 = pi09 ? n77076 : n77225;
  assign n77227 = pi08 ? n77161 : n77226;
  assign n77228 = pi07 ? n77064 : n77227;
  assign n77229 = pi06 ? n76820 : n77228;
  assign n77230 = pi05 ? n76325 : n77229;
  assign n77231 = pi04 ? n75119 : n77230;
  assign n77232 = pi03 ? n70347 : n77231;
  assign n77233 = pi22 ? n39291 : n37;
  assign n77234 = pi21 ? n77233 : n1618;
  assign n77235 = pi20 ? n32 : n77234;
  assign n77236 = pi19 ? n32 : n77235;
  assign n77237 = pi18 ? n32 : n77236;
  assign n77238 = pi17 ? n32 : n77237;
  assign n77239 = pi16 ? n32 : n77238;
  assign n77240 = pi15 ? n76833 : n77239;
  assign n77241 = pi14 ? n76833 : n77240;
  assign n77242 = pi23 ? n77043 : n51564;
  assign n77243 = pi22 ? n77242 : n51564;
  assign n77244 = pi21 ? n77243 : n57433;
  assign n77245 = pi20 ? n32 : n77244;
  assign n77246 = pi19 ? n32 : n77245;
  assign n77247 = pi18 ? n32 : n77246;
  assign n77248 = pi17 ? n32 : n77247;
  assign n77249 = pi16 ? n32 : n77248;
  assign n77250 = pi21 ? n8440 : n3523;
  assign n77251 = pi20 ? n32 : n77250;
  assign n77252 = pi19 ? n32 : n77251;
  assign n77253 = pi18 ? n32 : n77252;
  assign n77254 = pi17 ? n32 : n77253;
  assign n77255 = pi16 ? n32 : n77254;
  assign n77256 = pi15 ? n77249 : n77255;
  assign n77257 = pi14 ? n77256 : n77189;
  assign n77258 = pi13 ? n77241 : n77257;
  assign n77259 = pi12 ? n76833 : n77258;
  assign n77260 = pi21 ? n77176 : n37639;
  assign n77261 = pi20 ? n32 : n77260;
  assign n77262 = pi19 ? n32 : n77261;
  assign n77263 = pi18 ? n32 : n77262;
  assign n77264 = pi17 ? n32 : n77263;
  assign n77265 = pi16 ? n32 : n77264;
  assign n77266 = pi21 ? n75209 : n32;
  assign n77267 = pi20 ? n32 : n77266;
  assign n77268 = pi19 ? n32 : n77267;
  assign n77269 = pi18 ? n32 : n77268;
  assign n77270 = pi17 ? n32 : n77269;
  assign n77271 = pi16 ? n32 : n77270;
  assign n77272 = pi15 ? n77265 : n77271;
  assign n77273 = pi22 ? n75565 : n56665;
  assign n77274 = pi21 ? n77273 : n32;
  assign n77275 = pi20 ? n32 : n77274;
  assign n77276 = pi19 ? n32 : n77275;
  assign n77277 = pi18 ? n32 : n77276;
  assign n77278 = pi17 ? n32 : n77277;
  assign n77279 = pi16 ? n32 : n77278;
  assign n77280 = pi21 ? n33095 : n32;
  assign n77281 = pi20 ? n32 : n77280;
  assign n77282 = pi19 ? n32 : n77281;
  assign n77283 = pi18 ? n32 : n77282;
  assign n77284 = pi17 ? n32 : n77283;
  assign n77285 = pi16 ? n32 : n77284;
  assign n77286 = pi15 ? n77279 : n77285;
  assign n77287 = pi14 ? n77272 : n77286;
  assign n77288 = pi13 ? n77287 : n77221;
  assign n77289 = pi12 ? n77288 : n32;
  assign n77290 = pi11 ? n77259 : n77289;
  assign n77291 = pi10 ? n77290 : n32;
  assign n77292 = pi09 ? n77076 : n77291;
  assign n77293 = pi22 ? n73958 : n51564;
  assign n77294 = pi21 ? n77293 : n58966;
  assign n77295 = pi20 ? n32 : n77294;
  assign n77296 = pi19 ? n32 : n77295;
  assign n77297 = pi18 ? n32 : n77296;
  assign n77298 = pi17 ? n32 : n77297;
  assign n77299 = pi16 ? n32 : n77298;
  assign n77300 = pi15 ? n77299 : n77255;
  assign n77301 = pi14 ? n77300 : n77189;
  assign n77302 = pi13 ? n76833 : n77301;
  assign n77303 = pi12 ? n76833 : n77302;
  assign n77304 = pi22 ? n8439 : n13481;
  assign n77305 = pi21 ? n77304 : n32;
  assign n77306 = pi20 ? n32 : n77305;
  assign n77307 = pi19 ? n32 : n77306;
  assign n77308 = pi18 ? n32 : n77307;
  assign n77309 = pi17 ? n32 : n77308;
  assign n77310 = pi16 ? n32 : n77309;
  assign n77311 = pi15 ? n77265 : n77310;
  assign n77312 = pi14 ? n77311 : n77286;
  assign n77313 = pi13 ? n77312 : n77221;
  assign n77314 = pi12 ? n77313 : n32;
  assign n77315 = pi11 ? n77303 : n77314;
  assign n77316 = pi10 ? n77315 : n32;
  assign n77317 = pi09 ? n77076 : n77316;
  assign n77318 = pi08 ? n77292 : n77317;
  assign n77319 = pi22 ? n73958 : n13481;
  assign n77320 = pi21 ? n77319 : n54564;
  assign n77321 = pi20 ? n32 : n77320;
  assign n77322 = pi19 ? n32 : n77321;
  assign n77323 = pi18 ? n32 : n77322;
  assign n77324 = pi17 ? n32 : n77323;
  assign n77325 = pi16 ? n32 : n77324;
  assign n77326 = pi15 ? n77325 : n77188;
  assign n77327 = pi14 ? n77300 : n77326;
  assign n77328 = pi13 ? n76833 : n77327;
  assign n77329 = pi12 ? n76833 : n77328;
  assign n77330 = pi21 ? n77319 : n32;
  assign n77331 = pi20 ? n32 : n77330;
  assign n77332 = pi19 ? n32 : n77331;
  assign n77333 = pi18 ? n32 : n77332;
  assign n77334 = pi17 ? n32 : n77333;
  assign n77335 = pi16 ? n32 : n77334;
  assign n77336 = pi22 ? n8439 : n396;
  assign n77337 = pi21 ? n77336 : n32;
  assign n77338 = pi20 ? n32 : n77337;
  assign n77339 = pi19 ? n32 : n77338;
  assign n77340 = pi18 ? n32 : n77339;
  assign n77341 = pi17 ? n32 : n77340;
  assign n77342 = pi16 ? n32 : n77341;
  assign n77343 = pi15 ? n77335 : n77342;
  assign n77344 = pi22 ? n73960 : n706;
  assign n77345 = pi21 ? n77344 : n32;
  assign n77346 = pi20 ? n32 : n77345;
  assign n77347 = pi19 ? n32 : n77346;
  assign n77348 = pi18 ? n32 : n77347;
  assign n77349 = pi17 ? n32 : n77348;
  assign n77350 = pi16 ? n32 : n77349;
  assign n77351 = pi20 ? n32 : n3210;
  assign n77352 = pi19 ? n32 : n77351;
  assign n77353 = pi18 ? n32 : n77352;
  assign n77354 = pi17 ? n32 : n77353;
  assign n77355 = pi16 ? n32 : n77354;
  assign n77356 = pi15 ? n77350 : n77355;
  assign n77357 = pi14 ? n77343 : n77356;
  assign n77358 = pi20 ? n32 : n2653;
  assign n77359 = pi19 ? n32 : n77358;
  assign n77360 = pi18 ? n32 : n77359;
  assign n77361 = pi17 ? n32 : n77360;
  assign n77362 = pi16 ? n32 : n77361;
  assign n77363 = pi20 ? n32 : n1822;
  assign n77364 = pi19 ? n32 : n77363;
  assign n77365 = pi18 ? n32 : n77364;
  assign n77366 = pi17 ? n32 : n77365;
  assign n77367 = pi16 ? n32 : n77366;
  assign n77368 = pi15 ? n77362 : n77367;
  assign n77369 = pi14 ? n77368 : n32;
  assign n77370 = pi13 ? n77357 : n77369;
  assign n77371 = pi12 ? n77370 : n32;
  assign n77372 = pi11 ? n77329 : n77371;
  assign n77373 = pi10 ? n77372 : n32;
  assign n77374 = pi09 ? n77076 : n77373;
  assign n77375 = pi15 ? n77362 : n77219;
  assign n77376 = pi14 ? n77375 : n32;
  assign n77377 = pi13 ? n77357 : n77376;
  assign n77378 = pi12 ? n77377 : n32;
  assign n77379 = pi11 ? n77329 : n77378;
  assign n77380 = pi10 ? n77379 : n32;
  assign n77381 = pi09 ? n77076 : n77380;
  assign n77382 = pi08 ? n77374 : n77381;
  assign n77383 = pi07 ? n77318 : n77382;
  assign n77384 = pi22 ? n73958 : n316;
  assign n77385 = pi21 ? n77384 : n54546;
  assign n77386 = pi20 ? n32 : n77385;
  assign n77387 = pi19 ? n32 : n77386;
  assign n77388 = pi18 ? n32 : n77387;
  assign n77389 = pi17 ? n32 : n77388;
  assign n77390 = pi16 ? n32 : n77389;
  assign n77391 = pi15 ? n77390 : n77255;
  assign n77392 = pi21 ? n77384 : n54564;
  assign n77393 = pi20 ? n32 : n77392;
  assign n77394 = pi19 ? n32 : n77393;
  assign n77395 = pi18 ? n32 : n77394;
  assign n77396 = pi17 ? n32 : n77395;
  assign n77397 = pi16 ? n32 : n77396;
  assign n77398 = pi15 ? n77397 : n77188;
  assign n77399 = pi14 ? n77391 : n77398;
  assign n77400 = pi13 ? n76833 : n77399;
  assign n77401 = pi12 ? n76833 : n77400;
  assign n77402 = pi21 ? n77384 : n32;
  assign n77403 = pi20 ? n32 : n77402;
  assign n77404 = pi19 ? n32 : n77403;
  assign n77405 = pi18 ? n32 : n77404;
  assign n77406 = pi17 ? n32 : n77405;
  assign n77407 = pi16 ? n32 : n77406;
  assign n77408 = pi15 ? n77407 : n77342;
  assign n77409 = pi21 ? n75293 : n32;
  assign n77410 = pi20 ? n32 : n77409;
  assign n77411 = pi19 ? n32 : n77410;
  assign n77412 = pi18 ? n32 : n77411;
  assign n77413 = pi17 ? n32 : n77412;
  assign n77414 = pi16 ? n32 : n77413;
  assign n77415 = pi15 ? n77414 : n77355;
  assign n77416 = pi14 ? n77408 : n77415;
  assign n77417 = pi13 ? n77416 : n77376;
  assign n77418 = pi12 ? n77417 : n32;
  assign n77419 = pi11 ? n77401 : n77418;
  assign n77420 = pi10 ? n77419 : n32;
  assign n77421 = pi09 ? n77076 : n77420;
  assign n77422 = pi15 ? n77362 : n32;
  assign n77423 = pi14 ? n77422 : n32;
  assign n77424 = pi13 ? n77416 : n77423;
  assign n77425 = pi12 ? n77424 : n32;
  assign n77426 = pi11 ? n77401 : n77425;
  assign n77427 = pi10 ? n77426 : n32;
  assign n77428 = pi09 ? n77076 : n77427;
  assign n77429 = pi08 ? n77421 : n77428;
  assign n77430 = pi21 ? n8440 : n882;
  assign n77431 = pi20 ? n32 : n77430;
  assign n77432 = pi19 ? n32 : n77431;
  assign n77433 = pi18 ? n32 : n77432;
  assign n77434 = pi17 ? n32 : n77433;
  assign n77435 = pi16 ? n32 : n77434;
  assign n77436 = pi15 ? n77435 : n77188;
  assign n77437 = pi14 ? n77255 : n77436;
  assign n77438 = pi13 ? n76833 : n77437;
  assign n77439 = pi12 ? n76833 : n77438;
  assign n77440 = pi21 ? n8440 : n32;
  assign n77441 = pi20 ? n32 : n77440;
  assign n77442 = pi19 ? n32 : n77441;
  assign n77443 = pi18 ? n32 : n77442;
  assign n77444 = pi17 ? n32 : n77443;
  assign n77445 = pi16 ? n32 : n77444;
  assign n77446 = pi15 ? n77445 : n77342;
  assign n77447 = pi22 ? n11681 : n706;
  assign n77448 = pi21 ? n77447 : n32;
  assign n77449 = pi20 ? n32 : n77448;
  assign n77450 = pi19 ? n32 : n77449;
  assign n77451 = pi18 ? n32 : n77450;
  assign n77452 = pi17 ? n32 : n77451;
  assign n77453 = pi16 ? n32 : n77452;
  assign n77454 = pi15 ? n77453 : n77154;
  assign n77455 = pi14 ? n77446 : n77454;
  assign n77456 = pi15 ? n77056 : n32;
  assign n77457 = pi14 ? n77456 : n32;
  assign n77458 = pi13 ? n77455 : n77457;
  assign n77459 = pi12 ? n77458 : n32;
  assign n77460 = pi11 ? n77439 : n77459;
  assign n77461 = pi10 ? n77460 : n32;
  assign n77462 = pi09 ? n77076 : n77461;
  assign n77463 = pi22 ? n8439 : n706;
  assign n77464 = pi21 ? n77463 : n32;
  assign n77465 = pi20 ? n32 : n77464;
  assign n77466 = pi19 ? n32 : n77465;
  assign n77467 = pi18 ? n32 : n77466;
  assign n77468 = pi17 ? n32 : n77467;
  assign n77469 = pi16 ? n32 : n77468;
  assign n77470 = pi15 ? n77469 : n77154;
  assign n77471 = pi14 ? n77446 : n77470;
  assign n77472 = pi13 ? n77471 : n77457;
  assign n77473 = pi12 ? n77472 : n32;
  assign n77474 = pi11 ? n77439 : n77473;
  assign n77475 = pi10 ? n77474 : n32;
  assign n77476 = pi09 ? n77076 : n77475;
  assign n77477 = pi08 ? n77462 : n77476;
  assign n77478 = pi07 ? n77429 : n77477;
  assign n77479 = pi06 ? n77383 : n77478;
  assign n77480 = pi23 ? n3690 : n13481;
  assign n77481 = pi22 ? n77480 : n13481;
  assign n77482 = pi21 ? n77481 : n55667;
  assign n77483 = pi20 ? n32 : n77482;
  assign n77484 = pi19 ? n32 : n77483;
  assign n77485 = pi18 ? n32 : n77484;
  assign n77486 = pi17 ? n32 : n77485;
  assign n77487 = pi16 ? n32 : n77486;
  assign n77488 = pi15 ? n77255 : n77487;
  assign n77489 = pi21 ? n77481 : n37639;
  assign n77490 = pi20 ? n32 : n77489;
  assign n77491 = pi19 ? n32 : n77490;
  assign n77492 = pi18 ? n32 : n77491;
  assign n77493 = pi17 ? n32 : n77492;
  assign n77494 = pi16 ? n32 : n77493;
  assign n77495 = pi15 ? n77435 : n77494;
  assign n77496 = pi14 ? n77488 : n77495;
  assign n77497 = pi13 ? n76833 : n77496;
  assign n77498 = pi12 ? n76833 : n77497;
  assign n77499 = pi21 ? n77481 : n32;
  assign n77500 = pi20 ? n32 : n77499;
  assign n77501 = pi19 ? n32 : n77500;
  assign n77502 = pi18 ? n32 : n77501;
  assign n77503 = pi17 ? n32 : n77502;
  assign n77504 = pi16 ? n32 : n77503;
  assign n77505 = pi22 ? n77480 : n55688;
  assign n77506 = pi21 ? n77505 : n32;
  assign n77507 = pi20 ? n32 : n77506;
  assign n77508 = pi19 ? n32 : n77507;
  assign n77509 = pi18 ? n32 : n77508;
  assign n77510 = pi17 ? n32 : n77509;
  assign n77511 = pi16 ? n32 : n77510;
  assign n77512 = pi15 ? n77504 : n77511;
  assign n77513 = pi22 ? n77480 : n706;
  assign n77514 = pi21 ? n77513 : n32;
  assign n77515 = pi20 ? n32 : n77514;
  assign n77516 = pi19 ? n32 : n77515;
  assign n77517 = pi18 ? n32 : n77516;
  assign n77518 = pi17 ? n32 : n77517;
  assign n77519 = pi16 ? n32 : n77518;
  assign n77520 = pi15 ? n77519 : n77056;
  assign n77521 = pi14 ? n77512 : n77520;
  assign n77522 = pi13 ? n77521 : n32;
  assign n77523 = pi12 ? n77522 : n32;
  assign n77524 = pi11 ? n77498 : n77523;
  assign n77525 = pi10 ? n77524 : n32;
  assign n77526 = pi09 ? n77076 : n77525;
  assign n77527 = pi15 ? n77255 : n77182;
  assign n77528 = pi15 ? n77435 : n77265;
  assign n77529 = pi14 ? n77527 : n77528;
  assign n77530 = pi13 ? n76833 : n77529;
  assign n77531 = pi12 ? n76833 : n77530;
  assign n77532 = pi21 ? n77176 : n32;
  assign n77533 = pi20 ? n32 : n77532;
  assign n77534 = pi19 ? n32 : n77533;
  assign n77535 = pi18 ? n32 : n77534;
  assign n77536 = pi17 ? n32 : n77535;
  assign n77537 = pi16 ? n32 : n77536;
  assign n77538 = pi22 ? n71924 : n56665;
  assign n77539 = pi21 ? n77538 : n32;
  assign n77540 = pi20 ? n32 : n77539;
  assign n77541 = pi19 ? n32 : n77540;
  assign n77542 = pi18 ? n32 : n77541;
  assign n77543 = pi17 ? n32 : n77542;
  assign n77544 = pi16 ? n32 : n77543;
  assign n77545 = pi15 ? n77537 : n77544;
  assign n77546 = pi21 ? n71925 : n32;
  assign n77547 = pi20 ? n32 : n77546;
  assign n77548 = pi19 ? n32 : n77547;
  assign n77549 = pi18 ? n32 : n77548;
  assign n77550 = pi17 ? n32 : n77549;
  assign n77551 = pi16 ? n32 : n77550;
  assign n77552 = pi15 ? n77551 : n77056;
  assign n77553 = pi14 ? n77545 : n77552;
  assign n77554 = pi13 ? n77553 : n32;
  assign n77555 = pi12 ? n77554 : n32;
  assign n77556 = pi11 ? n77531 : n77555;
  assign n77557 = pi10 ? n77556 : n32;
  assign n77558 = pi09 ? n77076 : n77557;
  assign n77559 = pi08 ? n77526 : n77558;
  assign n77560 = pi22 ? n77167 : n316;
  assign n77561 = pi21 ? n77560 : n3494;
  assign n77562 = pi20 ? n32 : n77561;
  assign n77563 = pi19 ? n32 : n77562;
  assign n77564 = pi18 ? n32 : n77563;
  assign n77565 = pi17 ? n32 : n77564;
  assign n77566 = pi16 ? n32 : n77565;
  assign n77567 = pi21 ? n77304 : n55667;
  assign n77568 = pi20 ? n32 : n77567;
  assign n77569 = pi19 ? n32 : n77568;
  assign n77570 = pi18 ? n32 : n77569;
  assign n77571 = pi17 ? n32 : n77570;
  assign n77572 = pi16 ? n32 : n77571;
  assign n77573 = pi15 ? n77566 : n77572;
  assign n77574 = pi14 ? n77573 : n77528;
  assign n77575 = pi13 ? n76833 : n77574;
  assign n77576 = pi12 ? n76833 : n77575;
  assign n77577 = pi15 ? n77551 : n77219;
  assign n77578 = pi14 ? n77545 : n77577;
  assign n77579 = pi13 ? n77578 : n32;
  assign n77580 = pi12 ? n77579 : n32;
  assign n77581 = pi11 ? n77576 : n77580;
  assign n77582 = pi10 ? n77581 : n32;
  assign n77583 = pi09 ? n77076 : n77582;
  assign n77584 = pi15 ? n77537 : n77551;
  assign n77585 = pi14 ? n77584 : n32;
  assign n77586 = pi13 ? n77585 : n32;
  assign n77587 = pi12 ? n77586 : n32;
  assign n77588 = pi11 ? n77576 : n77587;
  assign n77589 = pi10 ? n77588 : n32;
  assign n77590 = pi09 ? n77076 : n77589;
  assign n77591 = pi08 ? n77583 : n77590;
  assign n77592 = pi07 ? n77559 : n77591;
  assign n77593 = pi23 ? n36659 : n32;
  assign n77594 = pi22 ? n37 : n77593;
  assign n77595 = pi21 ? n65 : n77594;
  assign n77596 = pi20 ? n32 : n77595;
  assign n77597 = pi19 ? n32 : n77596;
  assign n77598 = pi18 ? n32 : n77597;
  assign n77599 = pi17 ? n32 : n77598;
  assign n77600 = pi16 ? n32 : n77599;
  assign n77601 = pi15 ? n32 : n77600;
  assign n77602 = pi14 ? n77601 : n76833;
  assign n77603 = pi13 ? n32 : n77602;
  assign n77604 = pi12 ? n32 : n77603;
  assign n77605 = pi11 ? n32 : n77604;
  assign n77606 = pi10 ? n32 : n77605;
  assign n77607 = pi15 ? n76833 : n77255;
  assign n77608 = pi15 ? n77182 : n77265;
  assign n77609 = pi14 ? n77607 : n77608;
  assign n77610 = pi13 ? n76833 : n77609;
  assign n77611 = pi12 ? n76833 : n77610;
  assign n77612 = pi11 ? n77611 : n77587;
  assign n77613 = pi10 ? n77612 : n32;
  assign n77614 = pi09 ? n77606 : n77613;
  assign n77615 = pi22 ? n71924 : n32;
  assign n77616 = pi21 ? n77615 : n32;
  assign n77617 = pi20 ? n32 : n77616;
  assign n77618 = pi19 ? n32 : n77617;
  assign n77619 = pi18 ? n32 : n77618;
  assign n77620 = pi17 ? n32 : n77619;
  assign n77621 = pi16 ? n32 : n77620;
  assign n77622 = pi15 ? n77537 : n77621;
  assign n77623 = pi14 ? n77622 : n32;
  assign n77624 = pi13 ? n77623 : n32;
  assign n77625 = pi12 ? n77624 : n32;
  assign n77626 = pi11 ? n77611 : n77625;
  assign n77627 = pi10 ? n77626 : n32;
  assign n77628 = pi09 ? n77606 : n77627;
  assign n77629 = pi08 ? n77614 : n77628;
  assign n77630 = pi21 ? n77304 : n19697;
  assign n77631 = pi20 ? n32 : n77630;
  assign n77632 = pi19 ? n32 : n77631;
  assign n77633 = pi18 ? n32 : n77632;
  assign n77634 = pi17 ? n32 : n77633;
  assign n77635 = pi16 ? n32 : n77634;
  assign n77636 = pi15 ? n77635 : n77310;
  assign n77637 = pi14 ? n77607 : n77636;
  assign n77638 = pi13 ? n76833 : n77637;
  assign n77639 = pi12 ? n76833 : n77638;
  assign n77640 = pi15 ? n77621 : n32;
  assign n77641 = pi14 ? n77640 : n32;
  assign n77642 = pi13 ? n77641 : n32;
  assign n77643 = pi12 ? n77642 : n32;
  assign n77644 = pi11 ? n77639 : n77643;
  assign n77645 = pi10 ? n77644 : n32;
  assign n77646 = pi09 ? n77606 : n77645;
  assign n77647 = pi07 ? n77629 : n77646;
  assign n77648 = pi06 ? n77592 : n77647;
  assign n77649 = pi05 ? n77479 : n77648;
  assign n77650 = pi21 ? n65 : n19793;
  assign n77651 = pi20 ? n32 : n77650;
  assign n77652 = pi19 ? n32 : n77651;
  assign n77653 = pi18 ? n32 : n77652;
  assign n77654 = pi17 ? n32 : n77653;
  assign n77655 = pi16 ? n32 : n77654;
  assign n77656 = pi15 ? n32 : n77655;
  assign n77657 = pi14 ? n77656 : n76833;
  assign n77658 = pi13 ? n32 : n77657;
  assign n77659 = pi12 ? n32 : n77658;
  assign n77660 = pi11 ? n32 : n77659;
  assign n77661 = pi10 ? n32 : n77660;
  assign n77662 = pi21 ? n8440 : n19697;
  assign n77663 = pi20 ? n32 : n77662;
  assign n77664 = pi19 ? n32 : n77663;
  assign n77665 = pi18 ? n32 : n77664;
  assign n77666 = pi17 ? n32 : n77665;
  assign n77667 = pi16 ? n32 : n77666;
  assign n77668 = pi15 ? n77667 : n77511;
  assign n77669 = pi14 ? n77607 : n77668;
  assign n77670 = pi13 ? n76833 : n77669;
  assign n77671 = pi12 ? n76833 : n77670;
  assign n77672 = pi11 ? n77671 : n32;
  assign n77673 = pi10 ? n77672 : n32;
  assign n77674 = pi09 ? n77661 : n77673;
  assign n77675 = pi15 ? n77667 : n77544;
  assign n77676 = pi14 ? n77607 : n77675;
  assign n77677 = pi13 ? n76833 : n77676;
  assign n77678 = pi12 ? n76833 : n77677;
  assign n77679 = pi11 ? n77678 : n32;
  assign n77680 = pi10 ? n77679 : n32;
  assign n77681 = pi09 ? n77661 : n77680;
  assign n77682 = pi08 ? n77674 : n77681;
  assign n77683 = pi15 ? n77188 : n32;
  assign n77684 = pi14 ? n77607 : n77683;
  assign n77685 = pi13 ? n76833 : n77684;
  assign n77686 = pi12 ? n76833 : n77685;
  assign n77687 = pi11 ? n77686 : n32;
  assign n77688 = pi10 ? n77687 : n32;
  assign n77689 = pi09 ? n77661 : n77688;
  assign n77690 = pi08 ? n77681 : n77689;
  assign n77691 = pi07 ? n77682 : n77690;
  assign n77692 = pi15 ? n76833 : n77182;
  assign n77693 = pi15 ? n77265 : n32;
  assign n77694 = pi14 ? n77692 : n77693;
  assign n77695 = pi13 ? n76833 : n77694;
  assign n77696 = pi12 ? n76833 : n77695;
  assign n77697 = pi11 ? n77696 : n32;
  assign n77698 = pi10 ? n77697 : n32;
  assign n77699 = pi09 ? n77661 : n77698;
  assign n77700 = pi14 ? n77692 : n32;
  assign n77701 = pi13 ? n76833 : n77700;
  assign n77702 = pi12 ? n76833 : n77701;
  assign n77703 = pi11 ? n77702 : n32;
  assign n77704 = pi10 ? n77703 : n32;
  assign n77705 = pi09 ? n77661 : n77704;
  assign n77706 = pi07 ? n77699 : n77705;
  assign n77707 = pi06 ? n77691 : n77706;
  assign n77708 = pi15 ? n76833 : n32;
  assign n77709 = pi14 ? n77708 : n32;
  assign n77710 = pi13 ? n76833 : n77709;
  assign n77711 = pi12 ? n76833 : n77710;
  assign n77712 = pi11 ? n77711 : n32;
  assign n77713 = pi10 ? n77712 : n32;
  assign n77714 = pi09 ? n77661 : n77713;
  assign n77715 = pi08 ? n77705 : n77714;
  assign n77716 = pi07 ? n77715 : n77714;
  assign n77717 = pi06 ? n77716 : n77714;
  assign n77718 = pi05 ? n77707 : n77717;
  assign n77719 = pi04 ? n77649 : n77718;
  assign n77720 = pi23 ? n36781 : n32;
  assign n77721 = pi22 ? n99 : n77720;
  assign n77722 = pi21 ? n127 : n77721;
  assign n77723 = pi20 ? n32 : n77722;
  assign n77724 = pi19 ? n32 : n77723;
  assign n77725 = pi18 ? n32 : n77724;
  assign n77726 = pi17 ? n32 : n77725;
  assign n77727 = pi16 ? n32 : n77726;
  assign n77728 = pi15 ? n32 : n77727;
  assign n77729 = pi14 ? n77728 : n76833;
  assign n77730 = pi13 ? n32 : n77729;
  assign n77731 = pi12 ? n32 : n77730;
  assign n77732 = pi11 ? n32 : n77731;
  assign n77733 = pi10 ? n32 : n77732;
  assign n77734 = pi09 ? n77733 : n77713;
  assign n77735 = pi21 ? n149 : n5482;
  assign n77736 = pi20 ? n32 : n77735;
  assign n77737 = pi19 ? n32 : n77736;
  assign n77738 = pi18 ? n32 : n77737;
  assign n77739 = pi17 ? n32 : n77738;
  assign n77740 = pi16 ? n32 : n77739;
  assign n77741 = pi15 ? n32 : n77740;
  assign n77742 = pi14 ? n77741 : n76833;
  assign n77743 = pi13 ? n32 : n77742;
  assign n77744 = pi12 ? n32 : n77743;
  assign n77745 = pi11 ? n32 : n77744;
  assign n77746 = pi10 ? n32 : n77745;
  assign n77747 = pi09 ? n77746 : n77713;
  assign n77748 = pi07 ? n77734 : n77747;
  assign n77749 = pi06 ? n77714 : n77748;
  assign n77750 = pi05 ? n77749 : n77747;
  assign n77751 = pi22 ? n148 : n139;
  assign n77752 = pi23 ? n36798 : n32;
  assign n77753 = pi22 ? n139 : n77752;
  assign n77754 = pi21 ? n77751 : n77753;
  assign n77755 = pi20 ? n32 : n77754;
  assign n77756 = pi19 ? n32 : n77755;
  assign n77757 = pi18 ? n32 : n77756;
  assign n77758 = pi17 ? n32 : n77757;
  assign n77759 = pi16 ? n32 : n77758;
  assign n77760 = pi15 ? n32 : n77759;
  assign n77761 = pi14 ? n77760 : n76833;
  assign n77762 = pi13 ? n32 : n77761;
  assign n77763 = pi12 ? n32 : n77762;
  assign n77764 = pi11 ? n32 : n77763;
  assign n77765 = pi10 ? n32 : n77764;
  assign n77766 = pi09 ? n77765 : n77713;
  assign n77767 = pi23 ? n32 : n139;
  assign n77768 = pi22 ? n77767 : n139;
  assign n77769 = pi21 ? n77768 : n6184;
  assign n77770 = pi20 ? n32 : n77769;
  assign n77771 = pi19 ? n32 : n77770;
  assign n77772 = pi18 ? n32 : n77771;
  assign n77773 = pi17 ? n32 : n77772;
  assign n77774 = pi16 ? n32 : n77773;
  assign n77775 = pi15 ? n32 : n77774;
  assign n77776 = pi14 ? n77775 : n76833;
  assign n77777 = pi13 ? n32 : n77776;
  assign n77778 = pi12 ? n32 : n77777;
  assign n77779 = pi11 ? n32 : n77778;
  assign n77780 = pi10 ? n32 : n77779;
  assign n77781 = pi09 ? n77780 : n77713;
  assign n77782 = pi07 ? n77766 : n77781;
  assign n77783 = pi06 ? n77782 : n77781;
  assign n77784 = pi05 ? n77747 : n77783;
  assign n77785 = pi04 ? n77750 : n77784;
  assign n77786 = pi03 ? n77719 : n77785;
  assign n77787 = pi02 ? n77232 : n77786;
  assign n77788 = pi14 ? n76833 : n32;
  assign n77789 = pi13 ? n76833 : n77788;
  assign n77790 = pi12 ? n76833 : n77789;
  assign n77791 = pi11 ? n77790 : n32;
  assign n77792 = pi10 ? n77791 : n32;
  assign n77793 = pi09 ? n77780 : n77792;
  assign n77794 = pi07 ? n77781 : n77793;
  assign n77795 = pi23 ? n43198 : n32;
  assign n77796 = pi22 ? n139 : n77795;
  assign n77797 = pi21 ? n77768 : n77796;
  assign n77798 = pi20 ? n32 : n77797;
  assign n77799 = pi19 ? n32 : n77798;
  assign n77800 = pi18 ? n32 : n77799;
  assign n77801 = pi17 ? n32 : n77800;
  assign n77802 = pi16 ? n32 : n77801;
  assign n77803 = pi15 ? n32 : n77802;
  assign n77804 = pi14 ? n77803 : n76833;
  assign n77805 = pi13 ? n32 : n77804;
  assign n77806 = pi12 ? n32 : n77805;
  assign n77807 = pi11 ? n32 : n77806;
  assign n77808 = pi10 ? n32 : n77807;
  assign n77809 = pi09 ? n77808 : n77792;
  assign n77810 = pi21 ? n77768 : n13102;
  assign n77811 = pi20 ? n32 : n77810;
  assign n77812 = pi19 ? n32 : n77811;
  assign n77813 = pi18 ? n32 : n77812;
  assign n77814 = pi17 ? n32 : n77813;
  assign n77815 = pi16 ? n32 : n77814;
  assign n77816 = pi15 ? n32 : n77815;
  assign n77817 = pi14 ? n77816 : n76833;
  assign n77818 = pi13 ? n32 : n77817;
  assign n77819 = pi12 ? n32 : n77818;
  assign n77820 = pi11 ? n32 : n77819;
  assign n77821 = pi10 ? n32 : n77820;
  assign n77822 = pi09 ? n77821 : n77792;
  assign n77823 = pi07 ? n77809 : n77822;
  assign n77824 = pi06 ? n77794 : n77823;
  assign n77825 = pi05 ? n77781 : n77824;
  assign n77826 = pi22 ? n49720 : n335;
  assign n77827 = pi21 ? n77826 : n20800;
  assign n77828 = pi20 ? n32 : n77827;
  assign n77829 = pi19 ? n32 : n77828;
  assign n77830 = pi18 ? n32 : n77829;
  assign n77831 = pi17 ? n32 : n77830;
  assign n77832 = pi16 ? n32 : n77831;
  assign n77833 = pi15 ? n32 : n77832;
  assign n77834 = pi14 ? n77833 : n76833;
  assign n77835 = pi13 ? n32 : n77834;
  assign n77836 = pi12 ? n32 : n77835;
  assign n77837 = pi11 ? n32 : n77836;
  assign n77838 = pi10 ? n32 : n77837;
  assign n77839 = pi09 ? n77838 : n77792;
  assign n77840 = pi23 ? n32 : n335;
  assign n77841 = pi22 ? n77840 : n335;
  assign n77842 = pi21 ? n77841 : n20800;
  assign n77843 = pi20 ? n32 : n77842;
  assign n77844 = pi19 ? n32 : n77843;
  assign n77845 = pi18 ? n32 : n77844;
  assign n77846 = pi17 ? n32 : n77845;
  assign n77847 = pi16 ? n32 : n77846;
  assign n77848 = pi15 ? n32 : n77847;
  assign n77849 = pi14 ? n77848 : n76833;
  assign n77850 = pi13 ? n32 : n77849;
  assign n77851 = pi12 ? n32 : n77850;
  assign n77852 = pi11 ? n32 : n77851;
  assign n77853 = pi10 ? n32 : n77852;
  assign n77854 = pi09 ? n77853 : n77792;
  assign n77855 = pi07 ? n77839 : n77854;
  assign n77856 = pi22 ? n335 : n59341;
  assign n77857 = pi21 ? n77841 : n77856;
  assign n77858 = pi20 ? n32 : n77857;
  assign n77859 = pi19 ? n32 : n77858;
  assign n77860 = pi18 ? n32 : n77859;
  assign n77861 = pi17 ? n32 : n77860;
  assign n77862 = pi16 ? n32 : n77861;
  assign n77863 = pi15 ? n32 : n77862;
  assign n77864 = pi14 ? n77863 : n76833;
  assign n77865 = pi13 ? n32 : n77864;
  assign n77866 = pi12 ? n32 : n77865;
  assign n77867 = pi11 ? n32 : n77866;
  assign n77868 = pi10 ? n32 : n77867;
  assign n77869 = pi09 ? n77868 : n77792;
  assign n77870 = pi07 ? n77854 : n77869;
  assign n77871 = pi06 ? n77855 : n77870;
  assign n77872 = pi05 ? n77822 : n77871;
  assign n77873 = pi04 ? n77825 : n77872;
  assign n77874 = pi21 ? n77841 : n8260;
  assign n77875 = pi20 ? n32 : n77874;
  assign n77876 = pi19 ? n32 : n77875;
  assign n77877 = pi18 ? n32 : n77876;
  assign n77878 = pi17 ? n32 : n77877;
  assign n77879 = pi16 ? n32 : n77878;
  assign n77880 = pi15 ? n32 : n77879;
  assign n77881 = pi14 ? n77880 : n76833;
  assign n77882 = pi13 ? n32 : n77881;
  assign n77883 = pi12 ? n32 : n77882;
  assign n77884 = pi11 ? n32 : n77883;
  assign n77885 = pi10 ? n32 : n77884;
  assign n77886 = pi09 ? n77885 : n77792;
  assign n77887 = pi07 ? n77869 : n77886;
  assign n77888 = pi06 ? n77887 : n77886;
  assign n77889 = pi22 ? n77840 : n36659;
  assign n77890 = pi22 ? n36659 : n1407;
  assign n77891 = pi21 ? n77889 : n77890;
  assign n77892 = pi20 ? n32 : n77891;
  assign n77893 = pi19 ? n32 : n77892;
  assign n77894 = pi18 ? n32 : n77893;
  assign n77895 = pi17 ? n32 : n77894;
  assign n77896 = pi16 ? n32 : n77895;
  assign n77897 = pi15 ? n32 : n77896;
  assign n77898 = pi14 ? n77897 : n76833;
  assign n77899 = pi13 ? n32 : n77898;
  assign n77900 = pi12 ? n32 : n77899;
  assign n77901 = pi11 ? n32 : n77900;
  assign n77902 = pi10 ? n32 : n77901;
  assign n77903 = pi09 ? n77902 : n77792;
  assign n77904 = pi21 ? n72455 : n77890;
  assign n77905 = pi20 ? n32 : n77904;
  assign n77906 = pi19 ? n32 : n77905;
  assign n77907 = pi18 ? n32 : n77906;
  assign n77908 = pi17 ? n32 : n77907;
  assign n77909 = pi16 ? n32 : n77908;
  assign n77910 = pi15 ? n32 : n77909;
  assign n77911 = pi14 ? n77910 : n76833;
  assign n77912 = pi13 ? n32 : n77911;
  assign n77913 = pi12 ? n32 : n77912;
  assign n77914 = pi11 ? n32 : n77913;
  assign n77915 = pi10 ? n32 : n77914;
  assign n77916 = pi09 ? n77915 : n77792;
  assign n77917 = pi07 ? n77903 : n77916;
  assign n77918 = pi23 ? n32 : n363;
  assign n77919 = pi22 ? n77918 : n363;
  assign n77920 = pi21 ? n77919 : n1408;
  assign n77921 = pi20 ? n32 : n77920;
  assign n77922 = pi19 ? n32 : n77921;
  assign n77923 = pi18 ? n32 : n77922;
  assign n77924 = pi17 ? n32 : n77923;
  assign n77925 = pi16 ? n32 : n77924;
  assign n77926 = pi15 ? n32 : n77925;
  assign n77927 = pi14 ? n77926 : n76833;
  assign n77928 = pi13 ? n32 : n77927;
  assign n77929 = pi12 ? n32 : n77928;
  assign n77930 = pi11 ? n32 : n77929;
  assign n77931 = pi10 ? n32 : n77930;
  assign n77932 = pi09 ? n77931 : n77792;
  assign n77933 = pi06 ? n77917 : n77932;
  assign n77934 = pi05 ? n77888 : n77933;
  assign n77935 = pi22 ? n363 : n58452;
  assign n77936 = pi21 ? n77919 : n77935;
  assign n77937 = pi20 ? n32 : n77936;
  assign n77938 = pi19 ? n32 : n77937;
  assign n77939 = pi18 ? n32 : n77938;
  assign n77940 = pi17 ? n32 : n77939;
  assign n77941 = pi16 ? n32 : n77940;
  assign n77942 = pi15 ? n32 : n77941;
  assign n77943 = pi14 ? n77942 : n76833;
  assign n77944 = pi13 ? n32 : n77943;
  assign n77945 = pi12 ? n32 : n77944;
  assign n77946 = pi11 ? n32 : n77945;
  assign n77947 = pi10 ? n32 : n77946;
  assign n77948 = pi09 ? n77947 : n77792;
  assign n77949 = pi22 ? n36781 : n21502;
  assign n77950 = pi21 ? n45136 : n77949;
  assign n77951 = pi20 ? n32 : n77950;
  assign n77952 = pi19 ? n32 : n77951;
  assign n77953 = pi18 ? n32 : n77952;
  assign n77954 = pi17 ? n32 : n77953;
  assign n77955 = pi16 ? n32 : n77954;
  assign n77956 = pi15 ? n32 : n77955;
  assign n77957 = pi14 ? n77956 : n76833;
  assign n77958 = pi13 ? n32 : n77957;
  assign n77959 = pi12 ? n32 : n77958;
  assign n77960 = pi11 ? n32 : n77959;
  assign n77961 = pi10 ? n32 : n77960;
  assign n77962 = pi09 ? n77961 : n77792;
  assign n77963 = pi23 ? n74659 : n32;
  assign n77964 = pi22 ? n36781 : n77963;
  assign n77965 = pi21 ? n45136 : n77964;
  assign n77966 = pi20 ? n32 : n77965;
  assign n77967 = pi19 ? n32 : n77966;
  assign n77968 = pi18 ? n32 : n77967;
  assign n77969 = pi17 ? n32 : n77968;
  assign n77970 = pi16 ? n32 : n77969;
  assign n77971 = pi15 ? n32 : n77970;
  assign n77972 = pi14 ? n77971 : n76833;
  assign n77973 = pi13 ? n32 : n77972;
  assign n77974 = pi12 ? n32 : n77973;
  assign n77975 = pi11 ? n32 : n77974;
  assign n77976 = pi10 ? n32 : n77975;
  assign n77977 = pi09 ? n77976 : n77792;
  assign n77978 = pi08 ? n77962 : n77977;
  assign n77979 = pi14 ? n32 : n76833;
  assign n77980 = pi13 ? n32 : n77979;
  assign n77981 = pi12 ? n32 : n77980;
  assign n77982 = pi11 ? n32 : n77981;
  assign n77983 = pi10 ? n32 : n77982;
  assign n77984 = pi09 ? n77983 : n77792;
  assign n77985 = pi08 ? n77984 : n32;
  assign n77986 = pi07 ? n77978 : n77985;
  assign n77987 = pi06 ? n77948 : n77986;
  assign n77988 = pi05 ? n77987 : n32;
  assign n77989 = pi04 ? n77934 : n77988;
  assign n77990 = pi03 ? n77873 : n77989;
  assign n77991 = pi02 ? n77990 : n32;
  assign n77992 = pi01 ? n77787 : n77991;
  assign n77993 = pi00 ? n55176 : n77992;
  assign po0 = ~n77993;
endmodule


