// Benchmark "DD" written by ABC on Wed Jun 26 12:37:42 2019

module DD ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17,
    po0, po1, po2, po3, po4, po5, po6  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
    n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
    n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
    n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
    n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
    n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
    n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
    n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
    n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
    n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
    n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
    n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
    n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
    n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
    n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
    n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
    n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
    n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
    n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
    n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
    n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
    n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
    n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
    n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
    n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
    n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
    n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
    n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
    n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
    n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
    n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
    n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
    n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
    n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
    n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
    n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
    n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
    n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
    n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
    n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
    n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
    n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
    n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
    n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
    n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
    n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
    n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
    n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
    n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
    n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
    n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
    n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
    n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
    n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
    n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
    n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
    n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
    n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
    n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
    n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
    n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
    n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
    n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
    n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
    n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
    n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
    n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
    n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
    n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
    n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
    n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
    n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
    n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
    n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
    n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
    n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
    n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
    n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
    n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
    n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
    n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
    n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
    n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
    n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
    n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
    n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
    n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
    n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
    n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
    n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
    n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
    n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
    n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
    n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
    n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
    n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
    n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
    n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
    n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
    n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
    n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417;
  assign n26 = 1'b1;
  assign n27 = pi17 ? n26 : ~n26;
  assign n28 = pi16 ? n26 : n27;
  assign n29 = pi15 ? n28 : ~n26;
  assign n30 = pi14 ? n29 : ~n26;
  assign n31 = pi13 ? n26 : n30;
  assign n32 = pi12 ? n26 : n31;
  assign n33 = pi11 ? n26 : n32;
  assign n34 = pi10 ? n33 : n32;
  assign n35 = pi09 ? n26 : n34;
  assign n36 = pi08 ? n26 : n35;
  assign n37 = pi15 ? n26 : ~n26;
  assign n38 = pi14 ? n37 : ~n26;
  assign n39 = pi13 ? n26 : n38;
  assign n40 = pi12 ? n26 : n39;
  assign n41 = pi11 ? n32 : n40;
  assign n42 = pi10 ? n41 : n40;
  assign n43 = pi09 ? n32 : n42;
  assign n44 = pi16 ? n26 : ~n26;
  assign n45 = pi15 ? n26 : n44;
  assign n46 = pi14 ? n26 : ~n45;
  assign n47 = pi13 ? n26 : n46;
  assign n48 = pi12 ? n26 : n47;
  assign n49 = pi11 ? n48 : n26;
  assign n50 = pi10 ? n49 : n26;
  assign n51 = pi09 ? n50 : n34;
  assign n52 = pi08 ? n43 : n51;
  assign n53 = pi07 ? n36 : n52;
  assign n54 = pi09 ? n42 : n50;
  assign n55 = pi09 ? n34 : n42;
  assign n56 = pi08 ? n54 : n55;
  assign n57 = pi14 ? n26 : ~n26;
  assign n58 = pi13 ? n26 : n57;
  assign n59 = pi12 ? n26 : n58;
  assign n60 = pi16 ? n27 : n26;
  assign n61 = pi15 ? n60 : n26;
  assign n62 = pi14 ? n61 : n26;
  assign n63 = pi15 ? n26 : n28;
  assign n64 = pi14 ? n26 : ~n63;
  assign n65 = pi13 ? n62 : n64;
  assign n66 = pi12 ? n26 : n65;
  assign n67 = pi11 ? n59 : n66;
  assign n68 = pi14 ? n26 : n45;
  assign n69 = pi13 ? n26 : n68;
  assign n70 = pi16 ? n27 : ~n26;
  assign n71 = pi15 ? n26 : n70;
  assign n72 = pi14 ? n71 : ~n26;
  assign n73 = pi15 ? n28 : n26;
  assign n74 = pi14 ? n26 : n73;
  assign n75 = pi13 ? n72 : ~n74;
  assign n76 = pi12 ? n69 : ~n75;
  assign n77 = pi14 ? n26 : n71;
  assign n78 = pi13 ? n26 : n77;
  assign n79 = pi14 ? n45 : ~n26;
  assign n80 = pi13 ? n79 : ~n26;
  assign n81 = pi12 ? n78 : ~n80;
  assign n82 = pi11 ? n76 : n81;
  assign n83 = pi10 ? n67 : n82;
  assign n84 = pi09 ? n40 : n83;
  assign n85 = pi08 ? n51 : n84;
  assign n86 = pi07 ? n56 : n85;
  assign n87 = pi06 ? n53 : n86;
  assign n88 = pi05 ? n26 : n87;
  assign n89 = pi13 ? n26 : ~n26;
  assign n90 = pi12 ? n26 : n89;
  assign n91 = pi11 ? n26 : n90;
  assign n92 = pi10 ? n91 : n90;
  assign n93 = pi09 ? n26 : n92;
  assign n94 = pi08 ? n26 : n93;
  assign n95 = pi13 ? n68 : ~n26;
  assign n96 = pi12 ? n26 : n95;
  assign n97 = pi14 ? n26 : n63;
  assign n98 = pi13 ? n68 : ~n97;
  assign n99 = pi12 ? n26 : n98;
  assign n100 = pi11 ? n96 : n99;
  assign n101 = pi10 ? n96 : n100;
  assign n102 = pi11 ? n99 : n90;
  assign n103 = pi10 ? n99 : n102;
  assign n104 = pi09 ? n101 : n103;
  assign n105 = pi14 ? n45 : ~n63;
  assign n106 = pi13 ? n26 : n105;
  assign n107 = pi12 ? n26 : n106;
  assign n108 = pi13 ? n26 : n74;
  assign n109 = pi12 ? n26 : n108;
  assign n110 = pi11 ? n107 : n109;
  assign n111 = pi10 ? n110 : n26;
  assign n112 = pi10 ? n91 : n100;
  assign n113 = pi09 ? n111 : n112;
  assign n114 = pi08 ? n104 : n113;
  assign n115 = pi07 ? n94 : n114;
  assign n116 = pi09 ? n103 : n111;
  assign n117 = pi09 ? n112 : n103;
  assign n118 = pi08 ? n116 : n117;
  assign n119 = pi10 ? n91 : n32;
  assign n120 = pi09 ? n111 : n119;
  assign n121 = pi10 ? n32 : n40;
  assign n122 = pi13 ? n26 : n79;
  assign n123 = pi12 ? n26 : n122;
  assign n124 = pi13 ? n26 : n97;
  assign n125 = pi15 ? n44 : ~n26;
  assign n126 = pi14 ? n125 : ~n26;
  assign n127 = pi13 ? n126 : ~n57;
  assign n128 = pi12 ? n124 : ~n127;
  assign n129 = pi11 ? n123 : n128;
  assign n130 = pi14 ? n26 : n125;
  assign n131 = pi15 ? n28 : ~n44;
  assign n132 = pi14 ? n26 : n131;
  assign n133 = pi13 ? n130 : ~n132;
  assign n134 = pi12 ? n78 : ~n133;
  assign n135 = pi13 ? n130 : ~n26;
  assign n136 = pi12 ? n78 : ~n135;
  assign n137 = pi11 ? n134 : n136;
  assign n138 = pi10 ? n129 : n137;
  assign n139 = pi09 ? n121 : n138;
  assign n140 = pi08 ? n120 : n139;
  assign n141 = pi07 ? n118 : n140;
  assign n142 = pi06 ? n115 : n141;
  assign n143 = pi14 ? n26 : n37;
  assign n144 = pi13 ? n143 : ~n143;
  assign n145 = pi12 ? n26 : n144;
  assign n146 = pi11 ? n26 : n145;
  assign n147 = pi15 ? n44 : ~n44;
  assign n148 = pi14 ? n63 : ~n147;
  assign n149 = pi14 ? n26 : n147;
  assign n150 = pi13 ? n148 : ~n149;
  assign n151 = pi12 ? n26 : n150;
  assign n152 = pi15 ? n70 : ~n44;
  assign n153 = pi14 ? n26 : ~n152;
  assign n154 = pi13 ? n153 : ~n149;
  assign n155 = pi12 ? n26 : n154;
  assign n156 = pi11 ? n151 : n155;
  assign n157 = pi10 ? n146 : n156;
  assign n158 = pi09 ? n26 : n157;
  assign n159 = pi08 ? n26 : n158;
  assign n160 = pi14 ? n26 : ~n147;
  assign n161 = pi13 ? n160 : ~n149;
  assign n162 = pi12 ? n26 : n161;
  assign n163 = pi15 ? n60 : n44;
  assign n164 = pi14 ? n26 : n163;
  assign n165 = pi13 ? n164 : ~n149;
  assign n166 = pi12 ? n26 : n165;
  assign n167 = pi11 ? n162 : n166;
  assign n168 = pi15 ? n70 : ~n26;
  assign n169 = pi14 ? n26 : n168;
  assign n170 = pi13 ? n169 : ~n130;
  assign n171 = pi12 ? n26 : n170;
  assign n172 = pi13 ? n130 : ~n130;
  assign n173 = pi12 ? n26 : n172;
  assign n174 = pi11 ? n171 : n173;
  assign n175 = pi10 ? n167 : n174;
  assign n176 = pi14 ? n26 : n29;
  assign n177 = pi13 ? n176 : ~n130;
  assign n178 = pi12 ? n26 : n177;
  assign n179 = pi11 ? n173 : n178;
  assign n180 = pi13 ? n143 : ~n68;
  assign n181 = pi12 ? n26 : n180;
  assign n182 = pi11 ? n181 : n90;
  assign n183 = pi10 ? n179 : n182;
  assign n184 = pi09 ? n175 : n183;
  assign n185 = pi13 ? n26 : n132;
  assign n186 = pi12 ? n26 : n185;
  assign n187 = pi11 ? n123 : n186;
  assign n188 = pi10 ? n187 : n26;
  assign n189 = pi10 ? n146 : n174;
  assign n190 = pi09 ? n188 : n189;
  assign n191 = pi08 ? n184 : n190;
  assign n192 = pi07 ? n159 : n191;
  assign n193 = pi09 ? n183 : n188;
  assign n194 = pi09 ? n189 : n183;
  assign n195 = pi08 ? n193 : n194;
  assign n196 = pi10 ? n91 : n41;
  assign n197 = pi09 ? n188 : n196;
  assign n198 = pi14 ? n63 : n26;
  assign n199 = pi13 ? n198 : n38;
  assign n200 = pi12 ? n26 : n199;
  assign n201 = pi11 ? n200 : n40;
  assign n202 = pi14 ? n37 : ~n63;
  assign n203 = pi13 ? n26 : n202;
  assign n204 = pi12 ? n26 : n203;
  assign n205 = pi11 ? n40 : n204;
  assign n206 = pi10 ? n201 : n205;
  assign n207 = pi13 ? n38 : ~n57;
  assign n208 = pi12 ? n69 : ~n207;
  assign n209 = pi11 ? n107 : n208;
  assign n210 = pi13 ? n130 : ~n64;
  assign n211 = pi12 ? n78 : ~n210;
  assign n212 = pi13 ? n77 : ~n26;
  assign n213 = pi12 ? n69 : ~n212;
  assign n214 = pi11 ? n211 : n213;
  assign n215 = pi10 ? n209 : n214;
  assign n216 = pi09 ? n206 : n215;
  assign n217 = pi08 ? n197 : n216;
  assign n218 = pi07 ? n195 : n217;
  assign n219 = pi06 ? n192 : n218;
  assign n220 = pi05 ? n142 : n219;
  assign n221 = pi04 ? n88 : n220;
  assign n222 = pi03 ? n26 : n221;
  assign n223 = pi02 ? n26 : n222;
  assign n224 = pi14 ? n63 : n37;
  assign n225 = pi13 ? n224 : ~n169;
  assign n226 = pi12 ? n26 : n225;
  assign n227 = pi13 ? n224 : ~n57;
  assign n228 = pi12 ? n26 : n227;
  assign n229 = pi11 ? n226 : n228;
  assign n230 = pi10 ? n146 : n229;
  assign n231 = pi09 ? n26 : n230;
  assign n232 = pi08 ? n26 : n231;
  assign n233 = pi15 ? n44 : n26;
  assign n234 = pi14 ? n63 : ~n233;
  assign n235 = pi13 ? n234 : ~n57;
  assign n236 = pi12 ? n26 : n235;
  assign n237 = pi13 ? n57 : ~n57;
  assign n238 = pi12 ? n26 : n237;
  assign n239 = pi11 ? n236 : n238;
  assign n240 = pi14 ? n63 : ~n26;
  assign n241 = pi13 ? n169 : ~n240;
  assign n242 = pi12 ? n26 : n241;
  assign n243 = pi13 ? n130 : ~n79;
  assign n244 = pi12 ? n26 : n243;
  assign n245 = pi11 ? n242 : n244;
  assign n246 = pi10 ? n239 : n245;
  assign n247 = pi10 ? n26 : n91;
  assign n248 = pi09 ? n246 : n247;
  assign n249 = pi15 ? n28 : ~n28;
  assign n250 = pi14 ? n26 : n249;
  assign n251 = pi13 ? n26 : n250;
  assign n252 = pi12 ? n26 : n251;
  assign n253 = pi11 ? n123 : n252;
  assign n254 = pi10 ? n253 : n26;
  assign n255 = pi10 ? n146 : n245;
  assign n256 = pi09 ? n254 : n255;
  assign n257 = pi08 ? n248 : n256;
  assign n258 = pi07 ? n232 : n257;
  assign n259 = pi09 ? n247 : n254;
  assign n260 = pi09 ? n255 : n247;
  assign n261 = pi08 ? n259 : n260;
  assign n262 = pi13 ? n26 : ~n68;
  assign n263 = pi12 ? n26 : n262;
  assign n264 = pi11 ? n26 : n263;
  assign n265 = pi10 ? n264 : n263;
  assign n266 = pi09 ? n254 : n265;
  assign n267 = pi11 ? n90 : n263;
  assign n268 = pi10 ? n263 : n267;
  assign n269 = pi14 ? n147 : n45;
  assign n270 = pi13 ? n26 : ~n269;
  assign n271 = pi12 ? n26 : n270;
  assign n272 = pi11 ? n263 : n271;
  assign n273 = pi13 ? n143 : ~n26;
  assign n274 = pi12 ? n26 : ~n273;
  assign n275 = pi12 ? n78 : ~n212;
  assign n276 = pi11 ? n274 : n275;
  assign n277 = pi10 ? n272 : n276;
  assign n278 = pi09 ? n268 : n277;
  assign n279 = pi08 ? n266 : n278;
  assign n280 = pi07 ? n261 : n279;
  assign n281 = pi06 ? n258 : n280;
  assign n282 = pi13 ? n143 : ~n57;
  assign n283 = pi12 ? n26 : n282;
  assign n284 = pi14 ? n45 : n37;
  assign n285 = pi13 ? n284 : ~n57;
  assign n286 = pi12 ? n26 : n285;
  assign n287 = pi11 ? n283 : n286;
  assign n288 = pi10 ? n146 : n287;
  assign n289 = pi09 ? n26 : n288;
  assign n290 = pi08 ? n26 : n289;
  assign n291 = pi16 ? n26 : ~n27;
  assign n292 = pi15 ? n291 : n26;
  assign n293 = pi14 ? n45 : ~n292;
  assign n294 = pi13 ? n293 : ~n240;
  assign n295 = pi12 ? n26 : n294;
  assign n296 = pi13 ? n240 : ~n79;
  assign n297 = pi12 ? n26 : n296;
  assign n298 = pi11 ? n295 : n297;
  assign n299 = pi13 ? n57 : ~n72;
  assign n300 = pi12 ? n26 : n299;
  assign n301 = pi13 ? n169 : ~n126;
  assign n302 = pi12 ? n26 : n301;
  assign n303 = pi11 ? n300 : n302;
  assign n304 = pi10 ? n298 : n303;
  assign n305 = pi09 ? n304 : n247;
  assign n306 = pi13 ? n26 : n240;
  assign n307 = pi12 ? n26 : n306;
  assign n308 = pi11 ? n123 : n307;
  assign n309 = pi10 ? n308 : n26;
  assign n310 = pi13 ? n57 : ~n240;
  assign n311 = pi12 ? n26 : n310;
  assign n312 = pi11 ? n311 : n302;
  assign n313 = pi10 ? n146 : n312;
  assign n314 = pi09 ? n309 : n313;
  assign n315 = pi08 ? n305 : n314;
  assign n316 = pi07 ? n290 : n315;
  assign n317 = pi09 ? n247 : n309;
  assign n318 = pi09 ? n313 : n247;
  assign n319 = pi08 ? n317 : n318;
  assign n320 = pi15 ? n26 : ~n44;
  assign n321 = pi14 ? n26 : n320;
  assign n322 = pi13 ? n321 : ~n143;
  assign n323 = pi12 ? n26 : n322;
  assign n324 = pi11 ? n26 : n323;
  assign n325 = pi13 ? n68 : ~n143;
  assign n326 = pi12 ? n26 : n325;
  assign n327 = pi15 ? n26 : n60;
  assign n328 = pi14 ? n327 : n45;
  assign n329 = pi13 ? n328 : ~n143;
  assign n330 = pi12 ? n26 : n329;
  assign n331 = pi11 ? n326 : n330;
  assign n332 = pi10 ? n324 : n331;
  assign n333 = pi09 ? n309 : n332;
  assign n334 = pi13 ? n68 : ~n68;
  assign n335 = pi12 ? n26 : n334;
  assign n336 = pi14 ? n26 : n44;
  assign n337 = pi13 ? n26 : ~n336;
  assign n338 = pi12 ? n26 : n337;
  assign n339 = pi11 ? n335 : n338;
  assign n340 = pi14 ? n233 : n37;
  assign n341 = pi13 ? n340 : ~n26;
  assign n342 = pi12 ? n26 : ~n341;
  assign n343 = pi12 ? n26 : ~n212;
  assign n344 = pi11 ? n342 : n343;
  assign n345 = pi10 ? n339 : n344;
  assign n346 = pi09 ? n326 : n345;
  assign n347 = pi08 ? n333 : n346;
  assign n348 = pi07 ? n319 : n347;
  assign n349 = pi06 ? n316 : n348;
  assign n350 = pi05 ? n281 : n349;
  assign n351 = pi14 ? n26 : ~n233;
  assign n352 = pi13 ? n351 : ~n130;
  assign n353 = pi12 ? n26 : n352;
  assign n354 = pi13 ? n72 : ~n240;
  assign n355 = pi12 ? n26 : n354;
  assign n356 = pi11 ? n353 : n355;
  assign n357 = pi10 ? n146 : n356;
  assign n358 = pi09 ? n26 : n357;
  assign n359 = pi08 ? n26 : n358;
  assign n360 = pi13 ? n72 : ~n79;
  assign n361 = pi12 ? n26 : n360;
  assign n362 = pi13 ? n72 : ~n72;
  assign n363 = pi12 ? n26 : n362;
  assign n364 = pi11 ? n361 : n363;
  assign n365 = pi13 ? n79 : ~n38;
  assign n366 = pi12 ? n26 : n365;
  assign n367 = pi13 ? n240 : ~n126;
  assign n368 = pi12 ? n26 : n367;
  assign n369 = pi11 ? n366 : n368;
  assign n370 = pi10 ? n364 : n369;
  assign n371 = pi10 ? n26 : n264;
  assign n372 = pi09 ? n370 : n371;
  assign n373 = pi13 ? n97 : ~n26;
  assign n374 = pi12 ? n26 : n373;
  assign n375 = pi13 ? n176 : ~n143;
  assign n376 = pi12 ? n26 : n375;
  assign n377 = pi11 ? n374 : n376;
  assign n378 = pi10 ? n377 : n312;
  assign n379 = pi09 ? n32 : n378;
  assign n380 = pi08 ? n372 : n379;
  assign n381 = pi07 ? n359 : n380;
  assign n382 = pi09 ? n371 : n32;
  assign n383 = pi09 ? n378 : n371;
  assign n384 = pi08 ? n382 : n383;
  assign n385 = pi11 ? n374 : n326;
  assign n386 = pi13 ? n143 : ~n169;
  assign n387 = pi12 ? n26 : n386;
  assign n388 = pi11 ? n387 : n283;
  assign n389 = pi10 ? n385 : n388;
  assign n390 = pi09 ? n32 : n389;
  assign n391 = pi13 ? n79 : ~n57;
  assign n392 = pi12 ? n26 : n391;
  assign n393 = pi11 ? n283 : n392;
  assign n394 = pi13 ? n38 : ~n72;
  assign n395 = pi12 ? n26 : n394;
  assign n396 = pi14 ? n168 : ~n45;
  assign n397 = pi13 ? n396 : n26;
  assign n398 = pi12 ? n26 : n397;
  assign n399 = pi11 ? n395 : n398;
  assign n400 = pi10 ? n393 : n399;
  assign n401 = pi09 ? n283 : n400;
  assign n402 = pi08 ? n390 : n401;
  assign n403 = pi07 ? n384 : n402;
  assign n404 = pi06 ? n381 : n403;
  assign n405 = pi11 ? n26 : n376;
  assign n406 = pi14 ? n26 : ~n292;
  assign n407 = pi13 ? n406 : ~n240;
  assign n408 = pi12 ? n26 : n407;
  assign n409 = pi13 ? n57 : ~n79;
  assign n410 = pi12 ? n26 : n409;
  assign n411 = pi11 ? n408 : n410;
  assign n412 = pi10 ? n405 : n411;
  assign n413 = pi09 ? n26 : n412;
  assign n414 = pi08 ? n26 : n413;
  assign n415 = pi14 ? n320 : ~n26;
  assign n416 = pi13 ? n415 : ~n72;
  assign n417 = pi12 ? n26 : n416;
  assign n418 = pi13 ? n38 : ~n38;
  assign n419 = pi12 ? n26 : n418;
  assign n420 = pi11 ? n417 : n419;
  assign n421 = pi13 ? n30 : ~n38;
  assign n422 = pi12 ? n26 : n421;
  assign n423 = pi13 ? n30 : ~n126;
  assign n424 = pi12 ? n26 : n423;
  assign n425 = pi11 ? n422 : n424;
  assign n426 = pi10 ? n420 : n425;
  assign n427 = pi13 ? n176 : ~n77;
  assign n428 = pi12 ? n26 : n427;
  assign n429 = pi11 ? n26 : n428;
  assign n430 = pi10 ? n26 : n429;
  assign n431 = pi09 ? n426 : n430;
  assign n432 = pi15 ? n28 : n44;
  assign n433 = pi14 ? n26 : n432;
  assign n434 = pi13 ? n433 : ~n77;
  assign n435 = pi12 ? n26 : n434;
  assign n436 = pi11 ? n435 : n99;
  assign n437 = pi10 ? n436 : n99;
  assign n438 = pi14 ? n63 : n29;
  assign n439 = pi13 ? n438 : ~n143;
  assign n440 = pi12 ? n26 : n439;
  assign n441 = pi11 ? n99 : n440;
  assign n442 = pi15 ? n26 : n27;
  assign n443 = pi14 ? n442 : ~n26;
  assign n444 = pi13 ? n240 : ~n443;
  assign n445 = pi12 ? n26 : n444;
  assign n446 = pi13 ? n57 : ~n126;
  assign n447 = pi12 ? n26 : n446;
  assign n448 = pi11 ? n445 : n447;
  assign n449 = pi10 ? n441 : n448;
  assign n450 = pi09 ? n437 : n449;
  assign n451 = pi08 ? n431 : n450;
  assign n452 = pi07 ? n414 : n451;
  assign n453 = pi09 ? n430 : n437;
  assign n454 = pi09 ? n449 : n430;
  assign n455 = pi08 ? n453 : n454;
  assign n456 = pi13 ? n433 : ~n143;
  assign n457 = pi12 ? n26 : n456;
  assign n458 = pi11 ? n99 : n457;
  assign n459 = pi14 ? n73 : n29;
  assign n460 = pi13 ? n459 : ~n130;
  assign n461 = pi12 ? n26 : n460;
  assign n462 = pi11 ? n178 : n461;
  assign n463 = pi10 ? n458 : n462;
  assign n464 = pi09 ? n437 : n463;
  assign n465 = pi14 ? n292 : n29;
  assign n466 = pi13 ? n465 : ~n169;
  assign n467 = pi12 ? n26 : n466;
  assign n468 = pi11 ? n461 : n467;
  assign n469 = pi13 ? n465 : ~n57;
  assign n470 = pi12 ? n26 : n469;
  assign n471 = pi13 ? n176 : ~n57;
  assign n472 = pi12 ? n26 : n471;
  assign n473 = pi11 ? n470 : n472;
  assign n474 = pi10 ? n468 : n473;
  assign n475 = pi13 ? n406 : ~n57;
  assign n476 = pi12 ? n26 : n475;
  assign n477 = pi11 ? n476 : n238;
  assign n478 = pi14 ? n233 : n26;
  assign n479 = pi13 ? n478 : n72;
  assign n480 = pi12 ? n26 : ~n479;
  assign n481 = pi14 ? n168 : ~n63;
  assign n482 = pi13 ? n481 : ~n126;
  assign n483 = pi12 ? n26 : n482;
  assign n484 = pi11 ? n480 : n483;
  assign n485 = pi10 ? n477 : n484;
  assign n486 = pi09 ? n474 : n485;
  assign n487 = pi08 ? n464 : n486;
  assign n488 = pi07 ? n455 : n487;
  assign n489 = pi06 ? n452 : n488;
  assign n490 = pi05 ? n404 : n489;
  assign n491 = pi04 ? n350 : n490;
  assign n492 = pi13 ? n406 : ~n130;
  assign n493 = pi12 ? n26 : n492;
  assign n494 = pi14 ? n73 : ~n26;
  assign n495 = pi13 ? n494 : ~n57;
  assign n496 = pi12 ? n26 : n495;
  assign n497 = pi11 ? n493 : n496;
  assign n498 = pi10 ? n405 : n497;
  assign n499 = pi09 ? n26 : n498;
  assign n500 = pi08 ? n26 : n499;
  assign n501 = pi14 ? n131 : ~n26;
  assign n502 = pi13 ? n501 : ~n72;
  assign n503 = pi12 ? n26 : n502;
  assign n504 = pi13 ? n126 : ~n38;
  assign n505 = pi12 ? n26 : n504;
  assign n506 = pi11 ? n503 : n505;
  assign n507 = pi14 ? n168 : ~n26;
  assign n508 = pi13 ? n507 : ~n126;
  assign n509 = pi12 ? n26 : n508;
  assign n510 = pi11 ? n505 : n509;
  assign n511 = pi10 ? n506 : n510;
  assign n512 = pi11 ? n26 : n178;
  assign n513 = pi10 ? n26 : n512;
  assign n514 = pi09 ? n511 : n513;
  assign n515 = pi13 ? n57 : ~n130;
  assign n516 = pi12 ? n26 : n515;
  assign n517 = pi15 ? n26 : n291;
  assign n518 = pi14 ? n517 : ~n26;
  assign n519 = pi13 ? n518 : ~n130;
  assign n520 = pi12 ? n26 : n519;
  assign n521 = pi11 ? n516 : n520;
  assign n522 = pi13 ? n79 : ~n72;
  assign n523 = pi12 ? n26 : n522;
  assign n524 = pi11 ? n523 : n368;
  assign n525 = pi10 ? n521 : n524;
  assign n526 = pi09 ? n516 : n525;
  assign n527 = pi08 ? n514 : n526;
  assign n528 = pi07 ? n500 : n527;
  assign n529 = pi09 ? n513 : n516;
  assign n530 = pi09 ? n525 : n513;
  assign n531 = pi08 ? n529 : n530;
  assign n532 = pi13 ? n57 : ~n169;
  assign n533 = pi12 ? n26 : n532;
  assign n534 = pi11 ? n533 : n238;
  assign n535 = pi11 ? n238 : n311;
  assign n536 = pi10 ? n534 : n535;
  assign n537 = pi11 ? n410 : n300;
  assign n538 = pi11 ? n395 : n424;
  assign n539 = pi10 ? n537 : n538;
  assign n540 = pi09 ? n536 : n539;
  assign n541 = pi08 ? n516 : n540;
  assign n542 = pi07 ? n531 : n541;
  assign n543 = pi06 ? n528 : n542;
  assign n544 = pi14 ? n233 : ~n26;
  assign n545 = pi13 ? n544 : ~n79;
  assign n546 = pi12 ? n26 : n545;
  assign n547 = pi11 ? n516 : n546;
  assign n548 = pi10 ? n405 : n547;
  assign n549 = pi09 ? n26 : n548;
  assign n550 = pi08 ? n26 : n549;
  assign n551 = pi13 ? n544 : ~n72;
  assign n552 = pi12 ? n26 : n551;
  assign n553 = pi14 ? n152 : ~n26;
  assign n554 = pi13 ? n553 : ~n38;
  assign n555 = pi12 ? n26 : n554;
  assign n556 = pi11 ? n552 : n555;
  assign n557 = pi13 ? n507 : ~n38;
  assign n558 = pi12 ? n26 : n557;
  assign n559 = pi13 ? n26 : n126;
  assign n560 = pi12 ? n26 : ~n559;
  assign n561 = pi11 ? n558 : n560;
  assign n562 = pi10 ? n556 : n561;
  assign n563 = pi09 ? n562 : n26;
  assign n564 = pi08 ? n563 : n26;
  assign n565 = pi07 ? n550 : n564;
  assign n566 = pi06 ? n565 : n26;
  assign n567 = pi05 ? n543 : n566;
  assign n568 = pi11 ? n238 : n410;
  assign n569 = pi10 ? n405 : n568;
  assign n570 = pi09 ? n26 : n569;
  assign n571 = pi08 ? n26 : n570;
  assign n572 = pi14 ? n163 : ~n26;
  assign n573 = pi13 ? n572 : ~n38;
  assign n574 = pi12 ? n26 : n573;
  assign n575 = pi11 ? n300 : n574;
  assign n576 = pi12 ? n26 : ~n39;
  assign n577 = pi12 ? n124 : ~n559;
  assign n578 = pi11 ? n576 : n577;
  assign n579 = pi10 ? n575 : n578;
  assign n580 = pi09 ? n579 : n26;
  assign n581 = pi08 ? n580 : n26;
  assign n582 = pi07 ? n571 : n581;
  assign n583 = pi06 ? n582 : n26;
  assign n584 = pi14 ? n61 : ~n26;
  assign n585 = pi13 ? n584 : ~n72;
  assign n586 = pi12 ? n26 : n585;
  assign n587 = pi11 ? n516 : n586;
  assign n588 = pi10 ? n405 : n587;
  assign n589 = pi09 ? n26 : n588;
  assign n590 = pi08 ? n26 : n589;
  assign n591 = pi14 ? n147 : n26;
  assign n592 = pi13 ? n591 : n38;
  assign n593 = pi12 ? n26 : ~n592;
  assign n594 = pi11 ? n586 : n593;
  assign n595 = pi13 ? n478 : n38;
  assign n596 = pi12 ? n124 : ~n595;
  assign n597 = pi12 ? n69 : ~n559;
  assign n598 = pi11 ? n596 : n597;
  assign n599 = pi10 ? n594 : n598;
  assign n600 = pi12 ? n78 : ~n95;
  assign n601 = pi11 ? n600 : n136;
  assign n602 = pi10 ? n601 : n136;
  assign n603 = pi09 ? n599 : n602;
  assign n604 = pi08 ? n603 : n136;
  assign n605 = pi07 ? n590 : n604;
  assign n606 = pi06 ? n605 : n136;
  assign n607 = pi05 ? n583 : n606;
  assign n608 = pi04 ? n567 : n607;
  assign n609 = pi03 ? n491 : n608;
  assign n610 = pi14 ? n152 : n26;
  assign n611 = pi13 ? n610 : n38;
  assign n612 = pi12 ? n26 : ~n611;
  assign n613 = pi11 ? n586 : n612;
  assign n614 = pi12 ? n124 : ~n592;
  assign n615 = pi11 ? n614 : n597;
  assign n616 = pi10 ? n613 : n615;
  assign n617 = pi12 ? n78 : ~n373;
  assign n618 = pi11 ? n617 : n275;
  assign n619 = pi10 ? n618 : n275;
  assign n620 = pi09 ? n616 : n619;
  assign n621 = pi12 ? n78 : ~n273;
  assign n622 = pi08 ? n620 : n621;
  assign n623 = pi07 ? n590 : n622;
  assign n624 = pi11 ? n621 : n275;
  assign n625 = pi10 ? n621 : n624;
  assign n626 = pi09 ? n621 : n625;
  assign n627 = pi08 ? n621 : n626;
  assign n628 = pi07 ? n621 : n627;
  assign n629 = pi06 ? n623 : n628;
  assign n630 = pi14 ? n168 : n26;
  assign n631 = pi13 ? n630 : n72;
  assign n632 = pi12 ? n26 : ~n631;
  assign n633 = pi11 ? n516 : n632;
  assign n634 = pi10 ? n405 : n633;
  assign n635 = pi09 ? n26 : n634;
  assign n636 = pi08 ? n26 : n635;
  assign n637 = pi12 ? n124 : n365;
  assign n638 = pi11 ? n300 : n637;
  assign n639 = pi14 ? n320 : n26;
  assign n640 = pi13 ? n639 : n38;
  assign n641 = pi12 ? n26 : ~n640;
  assign n642 = pi11 ? n641 : n597;
  assign n643 = pi10 ? n638 : n642;
  assign n644 = pi11 ? n509 : n560;
  assign n645 = pi13 ? n507 : n26;
  assign n646 = pi12 ? n26 : n645;
  assign n647 = pi12 ? n26 : ~n89;
  assign n648 = pi11 ? n646 : n647;
  assign n649 = pi10 ? n644 : n648;
  assign n650 = pi09 ? n643 : n649;
  assign n651 = pi08 ? n650 : n647;
  assign n652 = pi07 ? n636 : n651;
  assign n653 = pi14 ? n26 : n327;
  assign n654 = pi13 ? n26 : n653;
  assign n655 = pi12 ? n654 : ~n89;
  assign n656 = pi12 ? n654 : ~n212;
  assign n657 = pi10 ? n655 : n656;
  assign n658 = pi09 ? n647 : n657;
  assign n659 = pi08 ? n647 : n658;
  assign n660 = pi07 ? n647 : n659;
  assign n661 = pi06 ? n652 : n660;
  assign n662 = pi05 ? n629 : n661;
  assign n663 = pi11 ? n516 : n300;
  assign n664 = pi10 ? n512 : n663;
  assign n665 = pi09 ? n26 : n664;
  assign n666 = pi08 ? n26 : n665;
  assign n667 = pi11 ? n300 : n523;
  assign n668 = pi11 ? n523 : n395;
  assign n669 = pi10 ? n667 : n668;
  assign n670 = pi13 ? n30 : ~n72;
  assign n671 = pi12 ? n26 : n670;
  assign n672 = pi10 ? n395 : n671;
  assign n673 = pi09 ? n669 : n672;
  assign n674 = pi08 ? n673 : n671;
  assign n675 = pi07 ? n666 : n674;
  assign n676 = pi12 ? n654 : n508;
  assign n677 = pi11 ? n671 : n676;
  assign n678 = pi10 ? n677 : n646;
  assign n679 = pi09 ? n671 : n678;
  assign n680 = pi08 ? n671 : n679;
  assign n681 = pi07 ? n671 : n680;
  assign n682 = pi06 ? n675 : n681;
  assign n683 = pi13 ? n240 : ~n169;
  assign n684 = pi12 ? n26 : n683;
  assign n685 = pi11 ? n26 : n684;
  assign n686 = pi10 ? n26 : n685;
  assign n687 = pi13 ? n38 : ~n415;
  assign n688 = pi12 ? n26 : n687;
  assign n689 = pi11 ? n392 : n688;
  assign n690 = pi13 ? n38 : n26;
  assign n691 = pi12 ? n26 : n690;
  assign n692 = pi11 ? n691 : n646;
  assign n693 = pi10 ? n689 : n692;
  assign n694 = pi09 ? n686 : n693;
  assign n695 = pi08 ? n26 : n694;
  assign n696 = pi07 ? n26 : n695;
  assign n697 = pi06 ? n26 : n696;
  assign n698 = pi05 ? n682 : n697;
  assign n699 = pi04 ? n662 : n698;
  assign n700 = pi13 ? n176 : ~n176;
  assign n701 = pi12 ? n26 : n700;
  assign n702 = pi11 ? n26 : n701;
  assign n703 = pi10 ? n26 : n702;
  assign n704 = pi14 ? n37 : n125;
  assign n705 = pi13 ? n79 : ~n704;
  assign n706 = pi12 ? n26 : n705;
  assign n707 = pi11 ? n516 : n706;
  assign n708 = pi13 ? n79 : ~n126;
  assign n709 = pi12 ? n26 : n708;
  assign n710 = pi11 ? n709 : n509;
  assign n711 = pi10 ? n707 : n710;
  assign n712 = pi09 ? n703 : n711;
  assign n713 = pi08 ? n26 : n712;
  assign n714 = pi07 ? n26 : n713;
  assign n715 = pi06 ? n26 : n714;
  assign n716 = pi07 ? n36 : n32;
  assign n717 = pi14 ? n29 : ~n63;
  assign n718 = pi13 ? n26 : n717;
  assign n719 = pi12 ? n26 : n718;
  assign n720 = pi11 ? n32 : n719;
  assign n721 = pi10 ? n32 : n720;
  assign n722 = pi09 ? n32 : n721;
  assign n723 = pi14 ? n29 : ~n45;
  assign n724 = pi13 ? n26 : n723;
  assign n725 = pi12 ? n26 : n724;
  assign n726 = pi14 ? n29 : ~n71;
  assign n727 = pi13 ? n26 : n726;
  assign n728 = pi12 ? n26 : n727;
  assign n729 = pi11 ? n725 : n728;
  assign n730 = pi13 ? n97 : ~n143;
  assign n731 = pi12 ? n26 : n730;
  assign n732 = pi11 ? n731 : n376;
  assign n733 = pi10 ? n729 : n732;
  assign n734 = pi13 ? n57 : ~n176;
  assign n735 = pi12 ? n26 : n734;
  assign n736 = pi14 ? n320 : ~n292;
  assign n737 = pi13 ? n57 : ~n736;
  assign n738 = pi12 ? n26 : n737;
  assign n739 = pi11 ? n735 : n738;
  assign n740 = pi13 ? n478 : n126;
  assign n741 = pi12 ? n26 : ~n740;
  assign n742 = pi11 ? n741 : n509;
  assign n743 = pi10 ? n739 : n742;
  assign n744 = pi09 ? n733 : n743;
  assign n745 = pi08 ? n722 : n744;
  assign n746 = pi07 ? n32 : n745;
  assign n747 = pi06 ? n716 : n746;
  assign n748 = pi05 ? n715 : n747;
  assign n749 = pi07 ? n94 : n90;
  assign n750 = pi13 ? n26 : ~n97;
  assign n751 = pi12 ? n26 : n750;
  assign n752 = pi11 ? n90 : n751;
  assign n753 = pi10 ? n90 : n752;
  assign n754 = pi09 ? n90 : n753;
  assign n755 = pi13 ? n26 : ~n77;
  assign n756 = pi12 ? n26 : n755;
  assign n757 = pi11 ? n263 : n756;
  assign n758 = pi11 ? n326 : n376;
  assign n759 = pi10 ? n757 : n758;
  assign n760 = pi11 ? n419 : n560;
  assign n761 = pi10 ? n238 : n760;
  assign n762 = pi09 ? n759 : n761;
  assign n763 = pi08 ? n754 : n762;
  assign n764 = pi07 ? n90 : n763;
  assign n765 = pi06 ? n749 : n764;
  assign n766 = pi10 ? n405 : n457;
  assign n767 = pi09 ? n26 : n766;
  assign n768 = pi08 ? n26 : n767;
  assign n769 = pi11 ? n457 : n435;
  assign n770 = pi10 ? n457 : n769;
  assign n771 = pi13 ? n68 : ~n77;
  assign n772 = pi12 ? n26 : n771;
  assign n773 = pi14 ? n26 : n517;
  assign n774 = pi13 ? n773 : ~n77;
  assign n775 = pi12 ? n26 : n774;
  assign n776 = pi11 ? n772 : n775;
  assign n777 = pi13 ? n68 : ~n321;
  assign n778 = pi12 ? n26 : n777;
  assign n779 = pi13 ? n433 : ~n321;
  assign n780 = pi12 ? n26 : n779;
  assign n781 = pi11 ? n778 : n780;
  assign n782 = pi10 ? n776 : n781;
  assign n783 = pi09 ? n770 : n782;
  assign n784 = pi08 ? n457 : n783;
  assign n785 = pi07 ? n768 : n784;
  assign n786 = pi15 ? n26 : ~n60;
  assign n787 = pi14 ? n26 : n786;
  assign n788 = pi13 ? n433 : ~n787;
  assign n789 = pi12 ? n26 : n788;
  assign n790 = pi11 ? n457 : n789;
  assign n791 = pi11 ? n376 : n428;
  assign n792 = pi10 ? n790 : n791;
  assign n793 = pi14 ? n327 : ~n26;
  assign n794 = pi13 ? n494 : ~n793;
  assign n795 = pi12 ? n26 : n794;
  assign n796 = pi11 ? n238 : n795;
  assign n797 = pi11 ? n480 : n509;
  assign n798 = pi10 ? n796 : n797;
  assign n799 = pi09 ? n792 : n798;
  assign n800 = pi08 ? n457 : n799;
  assign n801 = pi07 ? n457 : n800;
  assign n802 = pi06 ? n785 : n801;
  assign n803 = pi05 ? n765 : n802;
  assign n804 = pi04 ? n748 : n803;
  assign n805 = pi03 ? n699 : n804;
  assign n806 = pi02 ? n609 : n805;
  assign n807 = pi01 ? n223 : n806;
  assign n808 = pi10 ? n512 : n516;
  assign n809 = pi09 ? n26 : n808;
  assign n810 = pi08 ? n26 : n809;
  assign n811 = pi14 ? n327 : ~n233;
  assign n812 = pi13 ? n811 : ~n143;
  assign n813 = pi12 ? n26 : n812;
  assign n814 = pi11 ? n813 : n516;
  assign n815 = pi10 ? n145 : n814;
  assign n816 = pi09 ? n516 : n815;
  assign n817 = pi08 ? n516 : n816;
  assign n818 = pi07 ? n810 : n817;
  assign n819 = pi11 ? n516 : n311;
  assign n820 = pi10 ? n516 : n819;
  assign n821 = pi09 ? n820 : n539;
  assign n822 = pi08 ? n516 : n821;
  assign n823 = pi07 ? n516 : n822;
  assign n824 = pi06 ? n818 : n823;
  assign n825 = pi13 ? n351 : ~n57;
  assign n826 = pi12 ? n26 : n825;
  assign n827 = pi11 ? n26 : n826;
  assign n828 = pi13 ? n79 : ~n240;
  assign n829 = pi12 ? n26 : n828;
  assign n830 = pi11 ? n392 : n829;
  assign n831 = pi10 ? n827 : n830;
  assign n832 = pi09 ? n26 : n831;
  assign n833 = pi08 ? n26 : n832;
  assign n834 = pi07 ? n26 : n833;
  assign n835 = pi13 ? n38 : ~n79;
  assign n836 = pi12 ? n26 : n835;
  assign n837 = pi11 ? n836 : n26;
  assign n838 = pi10 ? n837 : n26;
  assign n839 = pi09 ? n838 : n26;
  assign n840 = pi08 ? n839 : n26;
  assign n841 = pi07 ? n840 : n26;
  assign n842 = pi06 ? n834 : n841;
  assign n843 = pi05 ? n824 : n842;
  assign n844 = pi14 ? n432 : ~n26;
  assign n845 = pi13 ? n844 : ~n72;
  assign n846 = pi12 ? n26 : n845;
  assign n847 = pi11 ? n392 : n846;
  assign n848 = pi10 ? n405 : n847;
  assign n849 = pi09 ? n26 : n848;
  assign n850 = pi08 ? n26 : n849;
  assign n851 = pi07 ? n26 : n850;
  assign n852 = pi11 ? n424 : n26;
  assign n853 = pi10 ? n852 : n26;
  assign n854 = pi09 ? n853 : n26;
  assign n855 = pi08 ? n854 : n26;
  assign n856 = pi07 ? n855 : n26;
  assign n857 = pi06 ? n851 : n856;
  assign n858 = pi14 ? n44 : ~n26;
  assign n859 = pi13 ? n858 : ~n38;
  assign n860 = pi12 ? n26 : n859;
  assign n861 = pi11 ? n238 : n860;
  assign n862 = pi10 ? n377 : n861;
  assign n863 = pi09 ? n32 : n862;
  assign n864 = pi08 ? n32 : n863;
  assign n865 = pi07 ? n36 : n864;
  assign n866 = pi13 ? n126 : ~n126;
  assign n867 = pi12 ? n26 : n866;
  assign n868 = pi11 ? n867 : n398;
  assign n869 = pi14 ? n168 : ~n125;
  assign n870 = pi13 ? n869 : n26;
  assign n871 = pi12 ? n26 : n870;
  assign n872 = pi12 ? n26 : ~n135;
  assign n873 = pi11 ? n871 : n872;
  assign n874 = pi10 ? n868 : n873;
  assign n875 = pi12 ? n124 : ~n135;
  assign n876 = pi12 ? n69 : ~n135;
  assign n877 = pi11 ? n875 : n876;
  assign n878 = pi10 ? n877 : n136;
  assign n879 = pi09 ? n874 : n878;
  assign n880 = pi08 ? n879 : n136;
  assign n881 = pi07 ? n880 : n136;
  assign n882 = pi06 ? n865 : n881;
  assign n883 = pi05 ? n857 : n882;
  assign n884 = pi04 ? n843 : n883;
  assign n885 = pi11 ? n96 : n376;
  assign n886 = pi13 ? n415 : ~n38;
  assign n887 = pi12 ? n26 : n886;
  assign n888 = pi11 ? n516 : n887;
  assign n889 = pi10 ? n885 : n888;
  assign n890 = pi09 ? n90 : n889;
  assign n891 = pi08 ? n90 : n890;
  assign n892 = pi07 ? n94 : n891;
  assign n893 = pi13 ? n481 : n26;
  assign n894 = pi12 ? n26 : n893;
  assign n895 = pi11 ? n867 : n894;
  assign n896 = pi14 ? n168 : ~n71;
  assign n897 = pi13 ? n896 : n26;
  assign n898 = pi12 ? n26 : n897;
  assign n899 = pi11 ? n898 : n274;
  assign n900 = pi10 ? n895 : n899;
  assign n901 = pi12 ? n124 : ~n273;
  assign n902 = pi12 ? n69 : ~n273;
  assign n903 = pi11 ? n901 : n902;
  assign n904 = pi10 ? n903 : n621;
  assign n905 = pi09 ? n900 : n904;
  assign n906 = pi08 ? n905 : n621;
  assign n907 = pi07 ? n906 : n627;
  assign n908 = pi06 ? n892 : n907;
  assign n909 = pi13 ? n584 : ~n38;
  assign n910 = pi12 ? n26 : n909;
  assign n911 = pi11 ? n410 : n910;
  assign n912 = pi10 ? n411 : n911;
  assign n913 = pi09 ? n457 : n912;
  assign n914 = pi08 ? n457 : n913;
  assign n915 = pi07 ? n768 : n914;
  assign n916 = pi15 ? n60 : ~n26;
  assign n917 = pi14 ? n916 : ~n26;
  assign n918 = pi13 ? n917 : ~n126;
  assign n919 = pi12 ? n26 : n918;
  assign n920 = pi11 ? n919 : n741;
  assign n921 = pi12 ? n124 : ~n89;
  assign n922 = pi11 ? n647 : n921;
  assign n923 = pi10 ? n920 : n922;
  assign n924 = pi09 ? n923 : n647;
  assign n925 = pi08 ? n924 : n647;
  assign n926 = pi07 ? n925 : n659;
  assign n927 = pi06 ? n915 : n926;
  assign n928 = pi05 ? n908 : n927;
  assign n929 = pi10 ? n238 : n667;
  assign n930 = pi09 ? n516 : n929;
  assign n931 = pi08 ? n516 : n930;
  assign n932 = pi07 ? n810 : n931;
  assign n933 = pi09 ? n672 : n671;
  assign n934 = pi08 ? n933 : n671;
  assign n935 = pi07 ? n934 : n680;
  assign n936 = pi06 ? n932 : n935;
  assign n937 = pi13 ? n72 : ~n415;
  assign n938 = pi12 ? n26 : n937;
  assign n939 = pi11 ? n392 : n938;
  assign n940 = pi10 ? n939 : n692;
  assign n941 = pi09 ? n686 : n940;
  assign n942 = pi08 ? n26 : n941;
  assign n943 = pi07 ? n26 : n942;
  assign n944 = pi06 ? n26 : n943;
  assign n945 = pi05 ? n936 : n944;
  assign n946 = pi04 ? n928 : n945;
  assign n947 = pi03 ? n884 : n946;
  assign n948 = pi13 ? n321 : ~n77;
  assign n949 = pi12 ? n26 : n948;
  assign n950 = pi11 ? n26 : n949;
  assign n951 = pi13 ? n773 : ~n653;
  assign n952 = pi12 ? n26 : n951;
  assign n953 = pi11 ? n952 : n778;
  assign n954 = pi10 ? n950 : n953;
  assign n955 = pi09 ? n26 : n954;
  assign n956 = pi08 ? n26 : n955;
  assign n957 = pi07 ? n956 : n457;
  assign n958 = pi06 ? n957 : n801;
  assign n959 = pi05 ? n765 : n958;
  assign n960 = pi04 ? n748 : n959;
  assign n961 = pi13 ? n351 : ~n143;
  assign n962 = pi12 ? n26 : n961;
  assign n963 = pi11 ? n962 : n813;
  assign n964 = pi10 ? n146 : n963;
  assign n965 = pi09 ? n26 : n964;
  assign n966 = pi08 ? n26 : n965;
  assign n967 = pi07 ? n966 : n516;
  assign n968 = pi06 ? n967 : n823;
  assign n969 = pi10 ? n146 : n238;
  assign n970 = pi09 ? n26 : n969;
  assign n971 = pi08 ? n26 : n970;
  assign n972 = pi13 ? n38 : ~n240;
  assign n973 = pi12 ? n26 : n972;
  assign n974 = pi11 ? n973 : n836;
  assign n975 = pi10 ? n974 : n26;
  assign n976 = pi09 ? n975 : n26;
  assign n977 = pi08 ? n976 : n26;
  assign n978 = pi07 ? n971 : n977;
  assign n979 = pi06 ? n978 : n26;
  assign n980 = pi05 ? n968 : n979;
  assign n981 = pi13 ? n494 : ~n79;
  assign n982 = pi12 ? n26 : n981;
  assign n983 = pi11 ? n311 : n982;
  assign n984 = pi10 ? n146 : n983;
  assign n985 = pi09 ? n26 : n984;
  assign n986 = pi08 ? n26 : n985;
  assign n987 = pi11 ? n671 : n867;
  assign n988 = pi10 ? n987 : n26;
  assign n989 = pi09 ? n988 : n26;
  assign n990 = pi08 ? n989 : n26;
  assign n991 = pi07 ? n986 : n990;
  assign n992 = pi06 ? n991 : n26;
  assign n993 = pi11 ? n238 : n552;
  assign n994 = pi10 ? n146 : n993;
  assign n995 = pi09 ? n26 : n994;
  assign n996 = pi08 ? n26 : n995;
  assign n997 = pi11 ? n398 : n872;
  assign n998 = pi10 ? n510 : n997;
  assign n999 = pi09 ? n998 : n878;
  assign n1000 = pi08 ? n999 : n136;
  assign n1001 = pi07 ? n996 : n1000;
  assign n1002 = pi06 ? n1001 : n136;
  assign n1003 = pi05 ? n992 : n1002;
  assign n1004 = pi04 ? n980 : n1003;
  assign n1005 = pi03 ? n960 : n1004;
  assign n1006 = pi02 ? n947 : n1005;
  assign n1007 = pi13 ? n544 : ~n38;
  assign n1008 = pi12 ? n26 : n1007;
  assign n1009 = pi11 ? n238 : n1008;
  assign n1010 = pi10 ? n405 : n1009;
  assign n1011 = pi09 ? n26 : n1010;
  assign n1012 = pi08 ? n26 : n1011;
  assign n1013 = pi11 ? n894 : n343;
  assign n1014 = pi10 ? n510 : n1013;
  assign n1015 = pi12 ? n124 : ~n212;
  assign n1016 = pi11 ? n1015 : n902;
  assign n1017 = pi10 ? n1016 : n621;
  assign n1018 = pi09 ? n1014 : n1017;
  assign n1019 = pi08 ? n1018 : n621;
  assign n1020 = pi07 ? n1012 : n1019;
  assign n1021 = pi06 ? n1020 : n628;
  assign n1022 = pi11 ? n516 : n910;
  assign n1023 = pi10 ? n405 : n1022;
  assign n1024 = pi09 ? n26 : n1023;
  assign n1025 = pi08 ? n26 : n1024;
  assign n1026 = pi11 ? n574 : n741;
  assign n1027 = pi11 ? n560 : n577;
  assign n1028 = pi10 ? n1026 : n1027;
  assign n1029 = pi09 ? n1028 : n647;
  assign n1030 = pi08 ? n1029 : n647;
  assign n1031 = pi07 ? n1025 : n1030;
  assign n1032 = pi11 ? n647 : n655;
  assign n1033 = pi10 ? n647 : n1032;
  assign n1034 = pi13 ? n653 : ~n26;
  assign n1035 = pi12 ? n654 : ~n1034;
  assign n1036 = pi11 ? n655 : n1035;
  assign n1037 = pi10 ? n1036 : n647;
  assign n1038 = pi09 ? n1033 : n1037;
  assign n1039 = pi08 ? n1038 : n647;
  assign n1040 = pi07 ? n1039 : n647;
  assign n1041 = pi06 ? n1031 : n1040;
  assign n1042 = pi05 ? n1021 : n1041;
  assign n1043 = pi13 ? n57 : ~n793;
  assign n1044 = pi12 ? n26 : n1043;
  assign n1045 = pi11 ? n238 : n1044;
  assign n1046 = pi10 ? n512 : n1045;
  assign n1047 = pi09 ? n26 : n1046;
  assign n1048 = pi08 ? n26 : n1047;
  assign n1049 = pi11 ? n395 : n671;
  assign n1050 = pi10 ? n523 : n1049;
  assign n1051 = pi09 ? n1050 : n671;
  assign n1052 = pi08 ? n1051 : n671;
  assign n1053 = pi07 ? n1048 : n1052;
  assign n1054 = pi12 ? n654 : n645;
  assign n1055 = pi11 ? n1054 : n646;
  assign n1056 = pi13 ? n507 : ~n507;
  assign n1057 = pi12 ? n26 : n1056;
  assign n1058 = pi11 ? n1057 : n671;
  assign n1059 = pi10 ? n1055 : n1058;
  assign n1060 = pi09 ? n671 : n1059;
  assign n1061 = pi08 ? n1060 : n671;
  assign n1062 = pi11 ? n671 : n424;
  assign n1063 = pi10 ? n671 : n1062;
  assign n1064 = pi09 ? n671 : n1063;
  assign n1065 = pi08 ? n671 : n1064;
  assign n1066 = pi07 ? n1061 : n1065;
  assign n1067 = pi06 ? n1053 : n1066;
  assign n1068 = pi11 ? n684 : n392;
  assign n1069 = pi10 ? n26 : n1068;
  assign n1070 = pi13 ? n72 : n26;
  assign n1071 = pi12 ? n26 : n1070;
  assign n1072 = pi10 ? n1071 : n26;
  assign n1073 = pi09 ? n1069 : n1072;
  assign n1074 = pi08 ? n1073 : n26;
  assign n1075 = pi07 ? n1074 : n26;
  assign n1076 = pi06 ? n26 : n1075;
  assign n1077 = pi05 ? n1067 : n1076;
  assign n1078 = pi04 ? n1042 : n1077;
  assign n1079 = pi11 ? n178 : n516;
  assign n1080 = pi10 ? n26 : n1079;
  assign n1081 = pi11 ? n419 : n509;
  assign n1082 = pi10 ? n1081 : n26;
  assign n1083 = pi09 ? n1080 : n1082;
  assign n1084 = pi08 ? n1083 : n26;
  assign n1085 = pi07 ? n1084 : n26;
  assign n1086 = pi06 ? n26 : n1085;
  assign n1087 = pi10 ? n720 : n729;
  assign n1088 = pi09 ? n32 : n1087;
  assign n1089 = pi08 ? n32 : n1088;
  assign n1090 = pi07 ? n36 : n1089;
  assign n1091 = pi14 ? n29 : ~n37;
  assign n1092 = pi13 ? n26 : n1091;
  assign n1093 = pi12 ? n26 : n1092;
  assign n1094 = pi11 ? n1093 : n731;
  assign n1095 = pi13 ? n130 : ~n176;
  assign n1096 = pi12 ? n26 : n1095;
  assign n1097 = pi11 ? n701 : n1096;
  assign n1098 = pi10 ? n1094 : n1097;
  assign n1099 = pi10 ? n760 : n601;
  assign n1100 = pi09 ? n1098 : n1099;
  assign n1101 = pi08 ? n1100 : n136;
  assign n1102 = pi07 ? n1101 : n136;
  assign n1103 = pi06 ? n1090 : n1102;
  assign n1104 = pi05 ? n1086 : n1103;
  assign n1105 = pi10 ? n752 : n757;
  assign n1106 = pi09 ? n90 : n1105;
  assign n1107 = pi08 ? n90 : n1106;
  assign n1108 = pi07 ? n94 : n1107;
  assign n1109 = pi13 ? n26 : ~n143;
  assign n1110 = pi12 ? n26 : n1109;
  assign n1111 = pi11 ? n1110 : n326;
  assign n1112 = pi11 ? n701 : n173;
  assign n1113 = pi10 ? n1111 : n1112;
  assign n1114 = pi11 ? n480 : n560;
  assign n1115 = pi10 ? n1114 : n618;
  assign n1116 = pi09 ? n1113 : n1115;
  assign n1117 = pi08 ? n1116 : n621;
  assign n1118 = pi07 ? n1117 : n627;
  assign n1119 = pi06 ? n1108 : n1118;
  assign n1120 = pi11 ? n26 : n756;
  assign n1121 = pi13 ? n68 : ~n653;
  assign n1122 = pi12 ? n26 : n1121;
  assign n1123 = pi11 ? n1122 : n778;
  assign n1124 = pi10 ? n1120 : n1123;
  assign n1125 = pi09 ? n26 : n1124;
  assign n1126 = pi08 ? n26 : n1125;
  assign n1127 = pi10 ? n457 : n790;
  assign n1128 = pi09 ? n457 : n1127;
  assign n1129 = pi08 ? n457 : n1128;
  assign n1130 = pi07 ? n1126 : n1129;
  assign n1131 = pi13 ? n130 : ~n57;
  assign n1132 = pi12 ? n26 : n1131;
  assign n1133 = pi11 ? n178 : n1132;
  assign n1134 = pi10 ? n791 : n1133;
  assign n1135 = pi14 ? n125 : n26;
  assign n1136 = pi13 ? n1135 : n72;
  assign n1137 = pi12 ? n26 : ~n1136;
  assign n1138 = pi15 ? n291 : ~n26;
  assign n1139 = pi14 ? n1138 : ~n26;
  assign n1140 = pi13 ? n591 : n1139;
  assign n1141 = pi12 ? n26 : ~n1140;
  assign n1142 = pi11 ? n1137 : n1141;
  assign n1143 = pi13 ? n591 : n126;
  assign n1144 = pi12 ? n26 : ~n1143;
  assign n1145 = pi11 ? n1144 : n741;
  assign n1146 = pi10 ? n1142 : n1145;
  assign n1147 = pi09 ? n1134 : n1146;
  assign n1148 = pi08 ? n1147 : n647;
  assign n1149 = pi07 ? n1148 : n647;
  assign n1150 = pi06 ? n1130 : n1149;
  assign n1151 = pi05 ? n1119 : n1150;
  assign n1152 = pi04 ? n1104 : n1151;
  assign n1153 = pi03 ? n1078 : n1152;
  assign n1154 = pi10 ? n516 : n238;
  assign n1155 = pi11 ? n417 : n395;
  assign n1156 = pi10 ? n1155 : n395;
  assign n1157 = pi09 ? n1154 : n1156;
  assign n1158 = pi08 ? n1157 : n671;
  assign n1159 = pi07 ? n1158 : n1065;
  assign n1160 = pi06 ? n967 : n1159;
  assign n1161 = pi11 ? n826 : n238;
  assign n1162 = pi10 ? n146 : n1161;
  assign n1163 = pi09 ? n26 : n1162;
  assign n1164 = pi08 ? n26 : n1163;
  assign n1165 = pi07 ? n1164 : n977;
  assign n1166 = pi06 ? n1165 : n26;
  assign n1167 = pi05 ? n1160 : n1166;
  assign n1168 = pi11 ? n408 : n982;
  assign n1169 = pi10 ? n146 : n1168;
  assign n1170 = pi09 ? n26 : n1169;
  assign n1171 = pi08 ? n26 : n1170;
  assign n1172 = pi07 ? n1171 : n990;
  assign n1173 = pi06 ? n1172 : n26;
  assign n1174 = pi11 ? n876 : n136;
  assign n1175 = pi10 ? n1174 : n136;
  assign n1176 = pi09 ? n998 : n1175;
  assign n1177 = pi08 ? n1176 : n136;
  assign n1178 = pi07 ? n996 : n1177;
  assign n1179 = pi06 ? n1178 : n136;
  assign n1180 = pi05 ? n1173 : n1179;
  assign n1181 = pi04 ? n1167 : n1180;
  assign n1182 = pi13 ? n57 : ~n38;
  assign n1183 = pi12 ? n26 : n1182;
  assign n1184 = pi11 ? n238 : n1183;
  assign n1185 = pi10 ? n405 : n1184;
  assign n1186 = pi09 ? n26 : n1185;
  assign n1187 = pi08 ? n26 : n1186;
  assign n1188 = pi12 ? n26 : ~n373;
  assign n1189 = pi11 ? n1188 : n1015;
  assign n1190 = pi10 ? n510 : n1189;
  assign n1191 = pi09 ? n1190 : n621;
  assign n1192 = pi08 ? n1191 : n621;
  assign n1193 = pi07 ? n1187 : n1192;
  assign n1194 = pi06 ? n1193 : n628;
  assign n1195 = pi13 ? n26 : n507;
  assign n1196 = pi12 ? n124 : ~n1195;
  assign n1197 = pi12 ? n69 : ~n95;
  assign n1198 = pi11 ? n1196 : n1197;
  assign n1199 = pi10 ? n561 : n1198;
  assign n1200 = pi16 ? n27 : ~n27;
  assign n1201 = pi15 ? n26 : n1200;
  assign n1202 = pi14 ? n26 : n1201;
  assign n1203 = pi13 ? n26 : n1202;
  assign n1204 = pi12 ? n1203 : ~n212;
  assign n1205 = pi11 ? n1204 : n275;
  assign n1206 = pi12 ? n654 : ~n273;
  assign n1207 = pi11 ? n656 : n1206;
  assign n1208 = pi10 ? n1205 : n1207;
  assign n1209 = pi09 ? n1199 : n1208;
  assign n1210 = pi08 ? n1209 : n1206;
  assign n1211 = pi07 ? n1025 : n1210;
  assign n1212 = pi11 ? n1206 : n656;
  assign n1213 = pi10 ? n1206 : n1212;
  assign n1214 = pi09 ? n1206 : n1213;
  assign n1215 = pi08 ? n1206 : n1214;
  assign n1216 = pi07 ? n1206 : n1215;
  assign n1217 = pi06 ? n1211 : n1216;
  assign n1218 = pi05 ? n1194 : n1217;
  assign n1219 = pi13 ? n584 : ~n415;
  assign n1220 = pi12 ? n26 : n1219;
  assign n1221 = pi11 ? n238 : n1220;
  assign n1222 = pi10 ? n405 : n1221;
  assign n1223 = pi09 ? n26 : n1222;
  assign n1224 = pi08 ? n26 : n1223;
  assign n1225 = pi11 ? n574 : n1144;
  assign n1226 = pi12 ? n69 : n482;
  assign n1227 = pi11 ? n577 : n1226;
  assign n1228 = pi10 ? n1225 : n1227;
  assign n1229 = pi11 ? n560 : n509;
  assign n1230 = pi10 ? n1229 : n560;
  assign n1231 = pi09 ? n1228 : n1230;
  assign n1232 = pi08 ? n1231 : n560;
  assign n1233 = pi07 ? n1224 : n1232;
  assign n1234 = pi06 ? n1233 : n560;
  assign n1235 = pi10 ? n523 : n395;
  assign n1236 = pi10 ? n1049 : n671;
  assign n1237 = pi09 ? n1235 : n1236;
  assign n1238 = pi08 ? n1237 : n671;
  assign n1239 = pi07 ? n666 : n1238;
  assign n1240 = pi07 ? n671 : n1065;
  assign n1241 = pi06 ? n1239 : n1240;
  assign n1242 = pi05 ? n1234 : n1241;
  assign n1243 = pi04 ? n1218 : n1242;
  assign n1244 = pi03 ? n1181 : n1243;
  assign n1245 = pi02 ? n1153 : n1244;
  assign n1246 = pi01 ? n1006 : n1245;
  assign n1247 = pi00 ? n807 : n1246;
  assign n1248 = pi11 ? n26 : n725;
  assign n1249 = pi10 ? n1248 : n725;
  assign n1250 = pi09 ? n26 : n1249;
  assign n1251 = pi08 ? n26 : n1250;
  assign n1252 = pi14 ? n37 : ~n45;
  assign n1253 = pi13 ? n26 : n1252;
  assign n1254 = pi12 ? n26 : n1253;
  assign n1255 = pi11 ? n59 : n307;
  assign n1256 = pi10 ? n1254 : n1255;
  assign n1257 = pi09 ? n725 : n1256;
  assign n1258 = pi09 ? n50 : n1249;
  assign n1259 = pi08 ? n1257 : n1258;
  assign n1260 = pi07 ? n1251 : n1259;
  assign n1261 = pi09 ? n1256 : n50;
  assign n1262 = pi09 ? n1249 : n1256;
  assign n1263 = pi08 ? n1261 : n1262;
  assign n1264 = pi10 ? n33 : n41;
  assign n1265 = pi09 ? n50 : n1264;
  assign n1266 = pi11 ? n307 : n123;
  assign n1267 = pi10 ? n40 : n1266;
  assign n1268 = pi13 ? n72 : ~n26;
  assign n1269 = pi12 ? n78 : ~n1268;
  assign n1270 = pi11 ? n76 : n1269;
  assign n1271 = pi10 ? n67 : n1270;
  assign n1272 = pi09 ? n1267 : n1271;
  assign n1273 = pi08 ? n1265 : n1272;
  assign n1274 = pi07 ? n1263 : n1273;
  assign n1275 = pi06 ? n1260 : n1274;
  assign n1276 = pi05 ? n26 : n1275;
  assign n1277 = pi09 ? n26 : n265;
  assign n1278 = pi08 ? n26 : n1277;
  assign n1279 = pi10 ? n263 : n756;
  assign n1280 = pi14 ? n45 : n26;
  assign n1281 = pi13 ? n26 : ~n1280;
  assign n1282 = pi12 ? n26 : n1281;
  assign n1283 = pi11 ? n263 : n1282;
  assign n1284 = pi10 ? n756 : n1283;
  assign n1285 = pi09 ? n1279 : n1284;
  assign n1286 = pi13 ? n26 : n64;
  assign n1287 = pi12 ? n26 : n1286;
  assign n1288 = pi11 ? n1287 : n109;
  assign n1289 = pi10 ? n1288 : n26;
  assign n1290 = pi10 ? n264 : n756;
  assign n1291 = pi09 ? n1289 : n1290;
  assign n1292 = pi08 ? n1285 : n1291;
  assign n1293 = pi07 ? n1278 : n1292;
  assign n1294 = pi09 ? n1284 : n1289;
  assign n1295 = pi09 ? n1290 : n1284;
  assign n1296 = pi08 ? n1294 : n1295;
  assign n1297 = pi10 ? n264 : n32;
  assign n1298 = pi09 ? n1289 : n1297;
  assign n1299 = pi10 ? n40 : n308;
  assign n1300 = pi11 ? n59 : n128;
  assign n1301 = pi13 ? n79 : ~n132;
  assign n1302 = pi12 ? n78 : ~n1301;
  assign n1303 = pi12 ? n69 : ~n1268;
  assign n1304 = pi11 ? n1302 : n1303;
  assign n1305 = pi10 ? n1300 : n1304;
  assign n1306 = pi09 ? n1299 : n1305;
  assign n1307 = pi08 ? n1298 : n1306;
  assign n1308 = pi07 ? n1296 : n1307;
  assign n1309 = pi06 ? n1293 : n1308;
  assign n1310 = pi11 ? n26 : n731;
  assign n1311 = pi13 ? n97 : ~n130;
  assign n1312 = pi12 ? n26 : n1311;
  assign n1313 = pi10 ? n1310 : n1312;
  assign n1314 = pi09 ? n26 : n1313;
  assign n1315 = pi08 ? n26 : n1314;
  assign n1316 = pi13 ? n160 : ~n130;
  assign n1317 = pi12 ? n26 : n1316;
  assign n1318 = pi13 ? n68 : ~n130;
  assign n1319 = pi12 ? n26 : n1318;
  assign n1320 = pi11 ? n1317 : n1319;
  assign n1321 = pi13 ? n336 : ~n130;
  assign n1322 = pi12 ? n26 : n1321;
  assign n1323 = pi10 ? n1320 : n1322;
  assign n1324 = pi13 ? n433 : ~n130;
  assign n1325 = pi12 ? n26 : n1324;
  assign n1326 = pi10 ? n1325 : n1283;
  assign n1327 = pi09 ? n1323 : n1326;
  assign n1328 = pi11 ? n59 : n186;
  assign n1329 = pi10 ? n1328 : n26;
  assign n1330 = pi15 ? n70 : n44;
  assign n1331 = pi14 ? n26 : n1330;
  assign n1332 = pi13 ? n1331 : ~n130;
  assign n1333 = pi12 ? n26 : n1332;
  assign n1334 = pi11 ? n1333 : n1322;
  assign n1335 = pi10 ? n1310 : n1334;
  assign n1336 = pi09 ? n1329 : n1335;
  assign n1337 = pi08 ? n1327 : n1336;
  assign n1338 = pi07 ? n1315 : n1337;
  assign n1339 = pi09 ? n1326 : n1329;
  assign n1340 = pi09 ? n1335 : n1326;
  assign n1341 = pi08 ? n1339 : n1340;
  assign n1342 = pi10 ? n264 : n41;
  assign n1343 = pi09 ? n1329 : n1342;
  assign n1344 = pi14 ? n45 : ~n45;
  assign n1345 = pi13 ? n26 : n1344;
  assign n1346 = pi12 ? n26 : n1345;
  assign n1347 = pi14 ? n63 : ~n45;
  assign n1348 = pi13 ? n26 : n1347;
  assign n1349 = pi12 ? n26 : n1348;
  assign n1350 = pi11 ? n1346 : n1349;
  assign n1351 = pi10 ? n40 : n1350;
  assign n1352 = pi11 ? n1346 : n208;
  assign n1353 = pi13 ? n79 : ~n64;
  assign n1354 = pi12 ? n78 : ~n1353;
  assign n1355 = pi15 ? n44 : ~n70;
  assign n1356 = pi14 ? n45 : ~n1355;
  assign n1357 = pi13 ? n1356 : ~n26;
  assign n1358 = pi12 ? n124 : ~n1357;
  assign n1359 = pi11 ? n1354 : n1358;
  assign n1360 = pi10 ? n1352 : n1359;
  assign n1361 = pi09 ? n1351 : n1360;
  assign n1362 = pi08 ? n1343 : n1361;
  assign n1363 = pi07 ? n1341 : n1362;
  assign n1364 = pi06 ? n1338 : n1363;
  assign n1365 = pi05 ? n1309 : n1364;
  assign n1366 = pi04 ? n1276 : n1365;
  assign n1367 = pi03 ? n26 : n1366;
  assign n1368 = pi02 ? n26 : n1367;
  assign n1369 = pi11 ? n26 : n1110;
  assign n1370 = pi13 ? n26 : ~n169;
  assign n1371 = pi12 ? n26 : n1370;
  assign n1372 = pi13 ? n26 : ~n57;
  assign n1373 = pi12 ? n26 : n1372;
  assign n1374 = pi11 ? n1371 : n1373;
  assign n1375 = pi10 ? n1369 : n1374;
  assign n1376 = pi09 ? n26 : n1375;
  assign n1377 = pi08 ? n26 : n1376;
  assign n1378 = pi14 ? n26 : ~n61;
  assign n1379 = pi13 ? n1378 : ~n57;
  assign n1380 = pi12 ? n26 : n1379;
  assign n1381 = pi11 ? n826 : n1380;
  assign n1382 = pi13 ? n169 : ~n79;
  assign n1383 = pi12 ? n26 : n1382;
  assign n1384 = pi11 ? n1383 : n244;
  assign n1385 = pi10 ? n1381 : n1384;
  assign n1386 = pi13 ? n26 : ~n591;
  assign n1387 = pi12 ? n26 : n1386;
  assign n1388 = pi11 ? n26 : n1387;
  assign n1389 = pi10 ? n26 : n1388;
  assign n1390 = pi09 ? n1385 : n1389;
  assign n1391 = pi11 ? n59 : n252;
  assign n1392 = pi10 ? n1391 : n26;
  assign n1393 = pi10 ? n1369 : n244;
  assign n1394 = pi09 ? n1392 : n1393;
  assign n1395 = pi08 ? n1390 : n1394;
  assign n1396 = pi07 ? n1377 : n1395;
  assign n1397 = pi09 ? n1389 : n1392;
  assign n1398 = pi09 ? n1393 : n1389;
  assign n1399 = pi08 ? n1397 : n1398;
  assign n1400 = pi15 ? n291 : n44;
  assign n1401 = pi14 ? n26 : n1400;
  assign n1402 = pi13 ? n26 : ~n1401;
  assign n1403 = pi12 ? n26 : n1402;
  assign n1404 = pi11 ? n26 : n1403;
  assign n1405 = pi10 ? n1404 : n1403;
  assign n1406 = pi09 ? n1392 : n1405;
  assign n1407 = pi11 ? n274 : n1015;
  assign n1408 = pi10 ? n272 : n1407;
  assign n1409 = pi09 ? n1403 : n1408;
  assign n1410 = pi08 ? n1406 : n1409;
  assign n1411 = pi07 ? n1399 : n1410;
  assign n1412 = pi06 ? n1396 : n1411;
  assign n1413 = pi11 ? n26 : n326;
  assign n1414 = pi13 ? n68 : ~n57;
  assign n1415 = pi12 ? n26 : n1414;
  assign n1416 = pi10 ? n1413 : n1415;
  assign n1417 = pi09 ? n26 : n1416;
  assign n1418 = pi08 ? n26 : n1417;
  assign n1419 = pi13 ? n351 : ~n79;
  assign n1420 = pi12 ? n26 : n1419;
  assign n1421 = pi11 ? n1420 : n410;
  assign n1422 = pi13 ? n176 : ~n126;
  assign n1423 = pi12 ? n26 : n1422;
  assign n1424 = pi11 ? n300 : n1423;
  assign n1425 = pi10 ? n1421 : n1424;
  assign n1426 = pi11 ? n26 : n271;
  assign n1427 = pi10 ? n26 : n1426;
  assign n1428 = pi09 ? n1425 : n1427;
  assign n1429 = pi14 ? n63 : ~n327;
  assign n1430 = pi13 ? n26 : n1429;
  assign n1431 = pi12 ? n26 : n1430;
  assign n1432 = pi11 ? n1431 : n307;
  assign n1433 = pi10 ? n1432 : n26;
  assign n1434 = pi13 ? n68 : ~n284;
  assign n1435 = pi12 ? n26 : n1434;
  assign n1436 = pi11 ? n26 : n1435;
  assign n1437 = pi15 ? n27 : ~n26;
  assign n1438 = pi14 ? n26 : n1437;
  assign n1439 = pi13 ? n1438 : ~n126;
  assign n1440 = pi12 ? n26 : n1439;
  assign n1441 = pi11 ? n300 : n1440;
  assign n1442 = pi10 ? n1436 : n1441;
  assign n1443 = pi09 ? n1433 : n1442;
  assign n1444 = pi08 ? n1428 : n1443;
  assign n1445 = pi07 ? n1418 : n1444;
  assign n1446 = pi09 ? n1427 : n1433;
  assign n1447 = pi09 ? n1442 : n1427;
  assign n1448 = pi08 ? n1446 : n1447;
  assign n1449 = pi10 ? n1369 : n731;
  assign n1450 = pi09 ? n1433 : n1449;
  assign n1451 = pi13 ? n97 : ~n68;
  assign n1452 = pi12 ? n26 : n1451;
  assign n1453 = pi11 ? n1452 : n338;
  assign n1454 = pi10 ? n1453 : n344;
  assign n1455 = pi09 ? n731 : n1454;
  assign n1456 = pi08 ? n1450 : n1455;
  assign n1457 = pi07 ? n1448 : n1456;
  assign n1458 = pi06 ? n1445 : n1457;
  assign n1459 = pi05 ? n1412 : n1458;
  assign n1460 = pi11 ? n353 : n410;
  assign n1461 = pi10 ? n1413 : n1460;
  assign n1462 = pi09 ? n26 : n1461;
  assign n1463 = pi08 ? n26 : n1462;
  assign n1464 = pi14 ? n1201 : ~n26;
  assign n1465 = pi13 ? n1464 : ~n72;
  assign n1466 = pi12 ? n26 : n1465;
  assign n1467 = pi11 ? n410 : n1466;
  assign n1468 = pi13 ? n518 : ~n38;
  assign n1469 = pi12 ? n26 : n1468;
  assign n1470 = pi11 ? n1469 : n368;
  assign n1471 = pi10 ? n1467 : n1470;
  assign n1472 = pi09 ? n1471 : n371;
  assign n1473 = pi14 ? n327 : n37;
  assign n1474 = pi13 ? n176 : ~n1473;
  assign n1475 = pi12 ? n26 : n1474;
  assign n1476 = pi11 ? n731 : n1475;
  assign n1477 = pi10 ? n1476 : n1424;
  assign n1478 = pi09 ? n725 : n1477;
  assign n1479 = pi08 ? n1472 : n1478;
  assign n1480 = pi07 ? n1463 : n1479;
  assign n1481 = pi09 ? n371 : n725;
  assign n1482 = pi09 ? n1477 : n371;
  assign n1483 = pi08 ? n1481 : n1482;
  assign n1484 = pi11 ? n1452 : n1110;
  assign n1485 = pi10 ? n1484 : n388;
  assign n1486 = pi09 ? n725 : n1485;
  assign n1487 = pi13 ? n143 : ~n79;
  assign n1488 = pi12 ? n26 : n1487;
  assign n1489 = pi11 ? n1488 : n410;
  assign n1490 = pi14 ? n1330 : ~n45;
  assign n1491 = pi13 ? n1490 : n26;
  assign n1492 = pi12 ? n26 : n1491;
  assign n1493 = pi11 ? n523 : n1492;
  assign n1494 = pi10 ? n1489 : n1493;
  assign n1495 = pi09 ? n283 : n1494;
  assign n1496 = pi08 ? n1486 : n1495;
  assign n1497 = pi07 ? n1483 : n1496;
  assign n1498 = pi06 ? n1480 : n1497;
  assign n1499 = pi13 ? n406 : ~n79;
  assign n1500 = pi12 ? n26 : n1499;
  assign n1501 = pi11 ? n1500 : n410;
  assign n1502 = pi10 ? n405 : n1501;
  assign n1503 = pi09 ? n26 : n1502;
  assign n1504 = pi08 ? n26 : n1503;
  assign n1505 = pi11 ? n300 : n1183;
  assign n1506 = pi13 ? n501 : ~n38;
  assign n1507 = pi12 ? n26 : n1506;
  assign n1508 = pi14 ? n249 : ~n26;
  assign n1509 = pi13 ? n1508 : ~n126;
  assign n1510 = pi12 ? n26 : n1509;
  assign n1511 = pi11 ? n1507 : n1510;
  assign n1512 = pi10 ? n1505 : n1511;
  assign n1513 = pi14 ? n26 : n28;
  assign n1514 = pi13 ? n1513 : ~n77;
  assign n1515 = pi12 ? n26 : n1514;
  assign n1516 = pi11 ? n26 : n1515;
  assign n1517 = pi10 ? n26 : n1516;
  assign n1518 = pi09 ? n1512 : n1517;
  assign n1519 = pi13 ? n74 : ~n77;
  assign n1520 = pi12 ? n26 : n1519;
  assign n1521 = pi11 ? n1520 : n756;
  assign n1522 = pi10 ? n1521 : n756;
  assign n1523 = pi14 ? n327 : n71;
  assign n1524 = pi13 ? n97 : ~n1523;
  assign n1525 = pi12 ? n26 : n1524;
  assign n1526 = pi11 ? n1525 : n1475;
  assign n1527 = pi11 ? n300 : n447;
  assign n1528 = pi10 ? n1526 : n1527;
  assign n1529 = pi09 ? n1522 : n1528;
  assign n1530 = pi08 ? n1518 : n1529;
  assign n1531 = pi07 ? n1504 : n1530;
  assign n1532 = pi09 ? n1517 : n1522;
  assign n1533 = pi09 ? n1528 : n1517;
  assign n1534 = pi08 ? n1532 : n1533;
  assign n1535 = pi13 ? n97 : ~n77;
  assign n1536 = pi12 ? n26 : n1535;
  assign n1537 = pi13 ? n1513 : ~n143;
  assign n1538 = pi12 ? n26 : n1537;
  assign n1539 = pi11 ? n1536 : n1538;
  assign n1540 = pi10 ? n1539 : n462;
  assign n1541 = pi09 ? n1522 : n1540;
  assign n1542 = pi11 ? n461 : n472;
  assign n1543 = pi10 ? n1542 : n472;
  assign n1544 = pi14 ? n1400 : ~n26;
  assign n1545 = pi13 ? n57 : ~n1544;
  assign n1546 = pi12 ? n26 : n1545;
  assign n1547 = pi11 ? n1500 : n1546;
  assign n1548 = pi15 ? n44 : ~n28;
  assign n1549 = pi14 ? n1548 : n292;
  assign n1550 = pi13 ? n1549 : n72;
  assign n1551 = pi12 ? n26 : ~n1550;
  assign n1552 = pi15 ? n70 : n28;
  assign n1553 = pi14 ? n1552 : ~n45;
  assign n1554 = pi13 ? n1553 : ~n126;
  assign n1555 = pi12 ? n26 : n1554;
  assign n1556 = pi11 ? n1551 : n1555;
  assign n1557 = pi10 ? n1547 : n1556;
  assign n1558 = pi09 ? n1543 : n1557;
  assign n1559 = pi08 ? n1541 : n1558;
  assign n1560 = pi07 ? n1534 : n1559;
  assign n1561 = pi06 ? n1531 : n1560;
  assign n1562 = pi05 ? n1498 : n1561;
  assign n1563 = pi04 ? n1459 : n1562;
  assign n1564 = pi13 ? n176 : ~n284;
  assign n1565 = pi12 ? n26 : n1564;
  assign n1566 = pi11 ? n26 : n1565;
  assign n1567 = pi14 ? n45 : n125;
  assign n1568 = pi13 ? n406 : ~n1567;
  assign n1569 = pi12 ? n26 : n1568;
  assign n1570 = pi11 ? n1569 : n300;
  assign n1571 = pi10 ? n1566 : n1570;
  assign n1572 = pi09 ? n26 : n1571;
  assign n1573 = pi08 ? n26 : n1572;
  assign n1574 = pi13 ? n494 : ~n38;
  assign n1575 = pi12 ? n26 : n1574;
  assign n1576 = pi11 ? n300 : n1575;
  assign n1577 = pi10 ? n1576 : n1511;
  assign n1578 = pi13 ? n74 : ~n130;
  assign n1579 = pi12 ? n26 : n1578;
  assign n1580 = pi11 ? n26 : n1579;
  assign n1581 = pi10 ? n26 : n1580;
  assign n1582 = pi09 ? n1577 : n1581;
  assign n1583 = pi14 ? n26 : ~n37;
  assign n1584 = pi13 ? n1583 : ~n130;
  assign n1585 = pi12 ? n26 : n1584;
  assign n1586 = pi14 ? n26 : ~n320;
  assign n1587 = pi13 ? n1586 : ~n130;
  assign n1588 = pi12 ? n26 : n1587;
  assign n1589 = pi11 ? n1585 : n1588;
  assign n1590 = pi10 ? n1585 : n1589;
  assign n1591 = pi14 ? n44 : n125;
  assign n1592 = pi13 ? n57 : ~n1591;
  assign n1593 = pi12 ? n26 : n1592;
  assign n1594 = pi13 ? n57 : ~n1567;
  assign n1595 = pi12 ? n26 : n1594;
  assign n1596 = pi11 ? n1593 : n1595;
  assign n1597 = pi13 ? n240 : ~n72;
  assign n1598 = pi12 ? n26 : n1597;
  assign n1599 = pi11 ? n1598 : n447;
  assign n1600 = pi10 ? n1596 : n1599;
  assign n1601 = pi09 ? n1590 : n1600;
  assign n1602 = pi08 ? n1582 : n1601;
  assign n1603 = pi07 ? n1573 : n1602;
  assign n1604 = pi09 ? n1581 : n1590;
  assign n1605 = pi09 ? n1600 : n1581;
  assign n1606 = pi08 ? n1604 : n1605;
  assign n1607 = pi10 ? n516 : n1588;
  assign n1608 = pi09 ? n1590 : n1607;
  assign n1609 = pi13 ? n1586 : ~n57;
  assign n1610 = pi12 ? n26 : n1609;
  assign n1611 = pi13 ? n1586 : ~n79;
  assign n1612 = pi12 ? n26 : n1611;
  assign n1613 = pi11 ? n1610 : n1612;
  assign n1614 = pi10 ? n1610 : n1613;
  assign n1615 = pi15 ? n291 : n70;
  assign n1616 = pi14 ? n1615 : ~n26;
  assign n1617 = pi13 ? n57 : ~n1616;
  assign n1618 = pi12 ? n26 : n1617;
  assign n1619 = pi11 ? n410 : n1618;
  assign n1620 = pi14 ? n63 : ~n292;
  assign n1621 = pi13 ? n1620 : ~n72;
  assign n1622 = pi12 ? n26 : n1621;
  assign n1623 = pi13 ? n494 : ~n126;
  assign n1624 = pi12 ? n26 : n1623;
  assign n1625 = pi11 ? n1622 : n1624;
  assign n1626 = pi10 ? n1619 : n1625;
  assign n1627 = pi09 ? n1614 : n1626;
  assign n1628 = pi08 ? n1608 : n1627;
  assign n1629 = pi07 ? n1606 : n1628;
  assign n1630 = pi06 ? n1603 : n1629;
  assign n1631 = pi13 ? n494 : ~n72;
  assign n1632 = pi12 ? n26 : n1631;
  assign n1633 = pi11 ? n1595 : n1632;
  assign n1634 = pi10 ? n1566 : n1633;
  assign n1635 = pi09 ? n26 : n1634;
  assign n1636 = pi08 ? n26 : n1635;
  assign n1637 = pi11 ? n1632 : n1008;
  assign n1638 = pi15 ? n26 : ~n291;
  assign n1639 = pi14 ? n1638 : ~n26;
  assign n1640 = pi13 ? n1639 : ~n126;
  assign n1641 = pi12 ? n26 : n1640;
  assign n1642 = pi11 ? n419 : n1641;
  assign n1643 = pi10 ? n1637 : n1642;
  assign n1644 = pi09 ? n1643 : n26;
  assign n1645 = pi08 ? n1644 : n26;
  assign n1646 = pi07 ? n1636 : n1645;
  assign n1647 = pi06 ? n1646 : n26;
  assign n1648 = pi05 ? n1630 : n1647;
  assign n1649 = pi10 ? n1566 : n410;
  assign n1650 = pi09 ? n26 : n1649;
  assign n1651 = pi08 ? n26 : n1650;
  assign n1652 = pi13 ? n62 : n38;
  assign n1653 = pi12 ? n26 : ~n1652;
  assign n1654 = pi11 ? n1653 : n560;
  assign n1655 = pi10 ? n1505 : n1654;
  assign n1656 = pi09 ? n1655 : n26;
  assign n1657 = pi08 ? n1656 : n26;
  assign n1658 = pi07 ? n1651 : n1657;
  assign n1659 = pi06 ? n1658 : n26;
  assign n1660 = pi11 ? n1595 : n300;
  assign n1661 = pi10 ? n1566 : n1660;
  assign n1662 = pi09 ? n26 : n1661;
  assign n1663 = pi08 ? n26 : n1662;
  assign n1664 = pi12 ? n26 : ~n595;
  assign n1665 = pi11 ? n1664 : n560;
  assign n1666 = pi10 ? n1505 : n1665;
  assign n1667 = pi12 ? n26 : ~n95;
  assign n1668 = pi11 ? n1667 : n872;
  assign n1669 = pi10 ? n1668 : n872;
  assign n1670 = pi09 ? n1666 : n1669;
  assign n1671 = pi08 ? n1670 : n872;
  assign n1672 = pi07 ? n1663 : n1671;
  assign n1673 = pi10 ? n872 : n876;
  assign n1674 = pi09 ? n872 : n1673;
  assign n1675 = pi08 ? n872 : n1674;
  assign n1676 = pi07 ? n872 : n1675;
  assign n1677 = pi06 ? n1672 : n1676;
  assign n1678 = pi05 ? n1659 : n1677;
  assign n1679 = pi04 ? n1648 : n1678;
  assign n1680 = pi03 ? n1563 : n1679;
  assign n1681 = pi13 ? n630 : n38;
  assign n1682 = pi12 ? n26 : ~n1681;
  assign n1683 = pi11 ? n586 : n1682;
  assign n1684 = pi14 ? n1548 : n26;
  assign n1685 = pi13 ? n1684 : n38;
  assign n1686 = pi12 ? n26 : ~n1685;
  assign n1687 = pi11 ? n1686 : n741;
  assign n1688 = pi10 ? n1683 : n1687;
  assign n1689 = pi11 ? n1667 : n343;
  assign n1690 = pi10 ? n1689 : n343;
  assign n1691 = pi09 ? n1688 : n1690;
  assign n1692 = pi08 ? n1691 : n274;
  assign n1693 = pi07 ? n1663 : n1692;
  assign n1694 = pi11 ? n274 : n343;
  assign n1695 = pi10 ? n274 : n1694;
  assign n1696 = pi09 ? n274 : n1695;
  assign n1697 = pi08 ? n274 : n1696;
  assign n1698 = pi07 ? n274 : n1697;
  assign n1699 = pi06 ? n1693 : n1698;
  assign n1700 = pi11 ? n1595 : n632;
  assign n1701 = pi10 ? n1566 : n1700;
  assign n1702 = pi09 ? n26 : n1701;
  assign n1703 = pi08 ? n26 : n1702;
  assign n1704 = pi15 ? n26 : ~n28;
  assign n1705 = pi14 ? n1704 : n26;
  assign n1706 = pi13 ? n1705 : n38;
  assign n1707 = pi12 ? n26 : ~n1706;
  assign n1708 = pi11 ? n1707 : n560;
  assign n1709 = pi10 ? n1505 : n1708;
  assign n1710 = pi13 ? n68 : n126;
  assign n1711 = pi12 ? n26 : ~n1710;
  assign n1712 = pi11 ? n509 : n1711;
  assign n1713 = pi11 ? n898 : n343;
  assign n1714 = pi10 ? n1712 : n1713;
  assign n1715 = pi09 ? n1709 : n1714;
  assign n1716 = pi09 ? n1690 : n343;
  assign n1717 = pi08 ? n1715 : n1716;
  assign n1718 = pi07 ? n1703 : n1717;
  assign n1719 = pi06 ? n1718 : n343;
  assign n1720 = pi05 ? n1699 : n1719;
  assign n1721 = pi13 ? n176 : ~n1567;
  assign n1722 = pi12 ? n26 : n1721;
  assign n1723 = pi11 ? n26 : n1722;
  assign n1724 = pi10 ? n1723 : n1660;
  assign n1725 = pi09 ? n26 : n1724;
  assign n1726 = pi08 ? n26 : n1725;
  assign n1727 = pi11 ? n1598 : n395;
  assign n1728 = pi10 ? n300 : n1727;
  assign n1729 = pi13 ? n1252 : ~n38;
  assign n1730 = pi12 ? n26 : n1729;
  assign n1731 = pi11 ? n395 : n1730;
  assign n1732 = pi13 ? n723 : ~n72;
  assign n1733 = pi12 ? n26 : n1732;
  assign n1734 = pi13 ? n723 : ~n38;
  assign n1735 = pi12 ? n26 : n1734;
  assign n1736 = pi11 ? n1733 : n1735;
  assign n1737 = pi10 ? n1731 : n1736;
  assign n1738 = pi09 ? n1728 : n1737;
  assign n1739 = pi08 ? n1738 : n1735;
  assign n1740 = pi07 ? n1726 : n1739;
  assign n1741 = pi11 ? n671 : n509;
  assign n1742 = pi10 ? n1741 : n398;
  assign n1743 = pi09 ? n1735 : n1742;
  assign n1744 = pi08 ? n1735 : n1743;
  assign n1745 = pi07 ? n1735 : n1744;
  assign n1746 = pi06 ? n1740 : n1745;
  assign n1747 = pi11 ? n26 : n297;
  assign n1748 = pi10 ? n26 : n1747;
  assign n1749 = pi13 ? n240 : ~n38;
  assign n1750 = pi12 ? n26 : n1749;
  assign n1751 = pi14 ? n37 : ~n320;
  assign n1752 = pi13 ? n1751 : ~n38;
  assign n1753 = pi12 ? n26 : n1752;
  assign n1754 = pi11 ? n1750 : n1753;
  assign n1755 = pi13 ? n1252 : n26;
  assign n1756 = pi12 ? n26 : n1755;
  assign n1757 = pi11 ? n1756 : n398;
  assign n1758 = pi10 ? n1754 : n1757;
  assign n1759 = pi09 ? n1748 : n1758;
  assign n1760 = pi08 ? n26 : n1759;
  assign n1761 = pi07 ? n26 : n1760;
  assign n1762 = pi06 ? n26 : n1761;
  assign n1763 = pi05 ? n1746 : n1762;
  assign n1764 = pi04 ? n1720 : n1763;
  assign n1765 = pi13 ? n176 : ~n1591;
  assign n1766 = pi12 ? n26 : n1765;
  assign n1767 = pi11 ? n26 : n1766;
  assign n1768 = pi10 ? n26 : n1767;
  assign n1769 = pi13 ? n240 : ~n704;
  assign n1770 = pi12 ? n26 : n1769;
  assign n1771 = pi11 ? n1595 : n1770;
  assign n1772 = pi11 ? n368 : n509;
  assign n1773 = pi10 ? n1771 : n1772;
  assign n1774 = pi09 ? n1768 : n1773;
  assign n1775 = pi08 ? n26 : n1774;
  assign n1776 = pi07 ? n26 : n1775;
  assign n1777 = pi06 ? n26 : n1776;
  assign n1778 = pi07 ? n1251 : n725;
  assign n1779 = pi11 ? n728 : n1093;
  assign n1780 = pi14 ? n327 : n125;
  assign n1781 = pi13 ? n176 : ~n1780;
  assign n1782 = pi12 ? n26 : n1781;
  assign n1783 = pi11 ? n1312 : n1782;
  assign n1784 = pi10 ? n1779 : n1783;
  assign n1785 = pi11 ? n1595 : n1183;
  assign n1786 = pi13 ? n1684 : n126;
  assign n1787 = pi12 ? n26 : ~n1786;
  assign n1788 = pi14 ? n1552 : ~n26;
  assign n1789 = pi13 ? n1788 : ~n126;
  assign n1790 = pi12 ? n26 : n1789;
  assign n1791 = pi11 ? n1787 : n1790;
  assign n1792 = pi10 ? n1785 : n1791;
  assign n1793 = pi09 ? n1784 : n1792;
  assign n1794 = pi08 ? n725 : n1793;
  assign n1795 = pi07 ? n725 : n1794;
  assign n1796 = pi06 ? n1778 : n1795;
  assign n1797 = pi05 ? n1777 : n1796;
  assign n1798 = pi07 ? n1278 : n263;
  assign n1799 = pi11 ? n756 : n1110;
  assign n1800 = pi13 ? n97 : ~n57;
  assign n1801 = pi12 ? n26 : n1800;
  assign n1802 = pi13 ? n176 : ~n415;
  assign n1803 = pi12 ? n26 : n1802;
  assign n1804 = pi11 ? n1801 : n1803;
  assign n1805 = pi10 ? n1799 : n1804;
  assign n1806 = pi13 ? n639 : n126;
  assign n1807 = pi12 ? n26 : ~n1806;
  assign n1808 = pi11 ? n1750 : n1807;
  assign n1809 = pi10 ? n1183 : n1808;
  assign n1810 = pi09 ? n1805 : n1809;
  assign n1811 = pi08 ? n263 : n1810;
  assign n1812 = pi07 ? n263 : n1811;
  assign n1813 = pi06 ? n1798 : n1812;
  assign n1814 = pi13 ? n74 : ~n143;
  assign n1815 = pi12 ? n26 : n1814;
  assign n1816 = pi11 ? n26 : n1815;
  assign n1817 = pi10 ? n1816 : n1815;
  assign n1818 = pi09 ? n26 : n1817;
  assign n1819 = pi08 ? n26 : n1818;
  assign n1820 = pi11 ? n1815 : n1520;
  assign n1821 = pi10 ? n1815 : n1820;
  assign n1822 = pi11 ? n1110 : n1815;
  assign n1823 = pi10 ? n756 : n1822;
  assign n1824 = pi09 ? n1821 : n1823;
  assign n1825 = pi08 ? n1815 : n1824;
  assign n1826 = pi07 ? n1819 : n1825;
  assign n1827 = pi11 ? n1815 : n1538;
  assign n1828 = pi10 ? n1827 : n472;
  assign n1829 = pi11 ? n1183 : n1632;
  assign n1830 = pi13 ? n1684 : n72;
  assign n1831 = pi12 ? n26 : ~n1830;
  assign n1832 = pi15 ? n70 : n26;
  assign n1833 = pi14 ? n1832 : ~n26;
  assign n1834 = pi13 ? n1833 : ~n126;
  assign n1835 = pi12 ? n26 : n1834;
  assign n1836 = pi11 ? n1831 : n1835;
  assign n1837 = pi10 ? n1829 : n1836;
  assign n1838 = pi09 ? n1828 : n1837;
  assign n1839 = pi08 ? n1815 : n1838;
  assign n1840 = pi07 ? n1815 : n1839;
  assign n1841 = pi06 ? n1826 : n1840;
  assign n1842 = pi05 ? n1813 : n1841;
  assign n1843 = pi04 ? n1797 : n1842;
  assign n1844 = pi03 ? n1764 : n1843;
  assign n1845 = pi02 ? n1680 : n1844;
  assign n1846 = pi01 ? n1368 : n1845;
  assign n1847 = pi10 ? n1580 : n1585;
  assign n1848 = pi09 ? n26 : n1847;
  assign n1849 = pi08 ? n26 : n1848;
  assign n1850 = pi14 ? n26 : ~n125;
  assign n1851 = pi13 ? n1850 : ~n143;
  assign n1852 = pi12 ? n26 : n1851;
  assign n1853 = pi11 ? n1852 : n1585;
  assign n1854 = pi10 ? n1110 : n1853;
  assign n1855 = pi09 ? n1585 : n1854;
  assign n1856 = pi08 ? n1585 : n1855;
  assign n1857 = pi07 ? n1849 : n1856;
  assign n1858 = pi10 ? n1585 : n1588;
  assign n1859 = pi09 ? n1585 : n1858;
  assign n1860 = pi14 ? n26 : ~n1704;
  assign n1861 = pi13 ? n1860 : ~n130;
  assign n1862 = pi12 ? n26 : n1861;
  assign n1863 = pi11 ? n1588 : n1862;
  assign n1864 = pi11 ? n516 : n410;
  assign n1865 = pi10 ? n1863 : n1864;
  assign n1866 = pi11 ? n300 : n1624;
  assign n1867 = pi10 ? n537 : n1866;
  assign n1868 = pi09 ? n1865 : n1867;
  assign n1869 = pi08 ? n1859 : n1868;
  assign n1870 = pi07 ? n1585 : n1869;
  assign n1871 = pi06 ? n1857 : n1870;
  assign n1872 = pi15 ? n44 : ~n291;
  assign n1873 = pi14 ? n26 : ~n1872;
  assign n1874 = pi13 ? n1873 : ~n57;
  assign n1875 = pi12 ? n26 : n1874;
  assign n1876 = pi11 ? n26 : n1875;
  assign n1877 = pi10 ? n1876 : n1613;
  assign n1878 = pi09 ? n26 : n1877;
  assign n1879 = pi08 ? n26 : n1878;
  assign n1880 = pi07 ? n26 : n1879;
  assign n1881 = pi13 ? n79 : ~n79;
  assign n1882 = pi12 ? n26 : n1881;
  assign n1883 = pi11 ? n1882 : n26;
  assign n1884 = pi10 ? n1883 : n26;
  assign n1885 = pi09 ? n1884 : n26;
  assign n1886 = pi08 ? n1885 : n26;
  assign n1887 = pi07 ? n1886 : n26;
  assign n1888 = pi06 ? n1880 : n1887;
  assign n1889 = pi05 ? n1871 : n1888;
  assign n1890 = pi10 ? n1566 : n537;
  assign n1891 = pi09 ? n26 : n1890;
  assign n1892 = pi08 ? n26 : n1891;
  assign n1893 = pi07 ? n26 : n1892;
  assign n1894 = pi13 ? n406 : ~n126;
  assign n1895 = pi12 ? n26 : n1894;
  assign n1896 = pi11 ? n1895 : n26;
  assign n1897 = pi10 ? n1896 : n26;
  assign n1898 = pi09 ? n1897 : n26;
  assign n1899 = pi08 ? n1898 : n26;
  assign n1900 = pi07 ? n1899 : n26;
  assign n1901 = pi06 ? n1893 : n1900;
  assign n1902 = pi14 ? n29 : ~n44;
  assign n1903 = pi13 ? n26 : n1902;
  assign n1904 = pi12 ? n26 : n1903;
  assign n1905 = pi11 ? n725 : n1904;
  assign n1906 = pi10 ? n725 : n1905;
  assign n1907 = pi11 ? n1452 : n376;
  assign n1908 = pi10 ? n1907 : n1576;
  assign n1909 = pi09 ? n1906 : n1908;
  assign n1910 = pi08 ? n725 : n1909;
  assign n1911 = pi07 ? n1251 : n1910;
  assign n1912 = pi13 ? n501 : ~n126;
  assign n1913 = pi12 ? n26 : n1912;
  assign n1914 = pi14 ? n125 : ~n45;
  assign n1915 = pi13 ? n1914 : n26;
  assign n1916 = pi12 ? n26 : n1915;
  assign n1917 = pi11 ? n1913 : n1916;
  assign n1918 = pi10 ? n1917 : n873;
  assign n1919 = pi09 ? n1918 : n872;
  assign n1920 = pi08 ? n1919 : n872;
  assign n1921 = pi07 ? n1920 : n1675;
  assign n1922 = pi06 ? n1911 : n1921;
  assign n1923 = pi05 ? n1901 : n1922;
  assign n1924 = pi04 ? n1889 : n1923;
  assign n1925 = pi14 ? n71 : n125;
  assign n1926 = pi13 ? n57 : ~n1925;
  assign n1927 = pi12 ? n26 : n1926;
  assign n1928 = pi11 ? n1927 : n1183;
  assign n1929 = pi10 ? n732 : n1928;
  assign n1930 = pi09 ? n263 : n1929;
  assign n1931 = pi08 ? n263 : n1930;
  assign n1932 = pi07 ? n1278 : n1931;
  assign n1933 = pi13 ? n544 : ~n126;
  assign n1934 = pi12 ? n26 : n1933;
  assign n1935 = pi14 ? n1832 : ~n45;
  assign n1936 = pi13 ? n1935 : n26;
  assign n1937 = pi12 ? n26 : n1936;
  assign n1938 = pi11 ? n1934 : n1937;
  assign n1939 = pi14 ? n125 : ~n71;
  assign n1940 = pi13 ? n1939 : n26;
  assign n1941 = pi12 ? n26 : n1940;
  assign n1942 = pi14 ? n125 : ~n37;
  assign n1943 = pi13 ? n1942 : n26;
  assign n1944 = pi12 ? n26 : n1943;
  assign n1945 = pi11 ? n1941 : n1944;
  assign n1946 = pi10 ? n1938 : n1945;
  assign n1947 = pi09 ? n1946 : n274;
  assign n1948 = pi08 ? n1947 : n274;
  assign n1949 = pi07 ? n1948 : n1697;
  assign n1950 = pi06 ? n1932 : n1949;
  assign n1951 = pi10 ? n1815 : n1827;
  assign n1952 = pi11 ? n410 : n1183;
  assign n1953 = pi10 ? n1501 : n1952;
  assign n1954 = pi09 ? n1951 : n1953;
  assign n1955 = pi08 ? n1815 : n1954;
  assign n1956 = pi07 ? n1819 : n1955;
  assign n1957 = pi13 ? n584 : ~n126;
  assign n1958 = pi12 ? n26 : n1957;
  assign n1959 = pi11 ? n1958 : n368;
  assign n1960 = pi10 ? n1959 : n1689;
  assign n1961 = pi11 ? n343 : n1667;
  assign n1962 = pi10 ? n1961 : n343;
  assign n1963 = pi09 ? n1960 : n1962;
  assign n1964 = pi08 ? n1963 : n343;
  assign n1965 = pi07 ? n1964 : n343;
  assign n1966 = pi06 ? n1956 : n1965;
  assign n1967 = pi05 ? n1950 : n1966;
  assign n1968 = pi11 ? n26 : n1325;
  assign n1969 = pi10 ? n1968 : n1588;
  assign n1970 = pi09 ? n26 : n1969;
  assign n1971 = pi08 ? n26 : n1970;
  assign n1972 = pi10 ? n1588 : n1863;
  assign n1973 = pi10 ? n410 : n300;
  assign n1974 = pi09 ? n1972 : n1973;
  assign n1975 = pi08 ? n1588 : n1974;
  assign n1976 = pi07 ? n1971 : n1975;
  assign n1977 = pi10 ? n523 : n1733;
  assign n1978 = pi09 ? n1977 : n1735;
  assign n1979 = pi08 ? n1978 : n1735;
  assign n1980 = pi07 ? n1979 : n1744;
  assign n1981 = pi06 ? n1976 : n1980;
  assign n1982 = pi14 ? n45 : ~n320;
  assign n1983 = pi13 ? n1982 : ~n38;
  assign n1984 = pi12 ? n26 : n1983;
  assign n1985 = pi11 ? n1750 : n1984;
  assign n1986 = pi10 ? n1985 : n1757;
  assign n1987 = pi09 ? n1748 : n1986;
  assign n1988 = pi08 ? n26 : n1987;
  assign n1989 = pi07 ? n26 : n1988;
  assign n1990 = pi06 ? n26 : n1989;
  assign n1991 = pi05 ? n1981 : n1990;
  assign n1992 = pi04 ? n1967 : n1991;
  assign n1993 = pi03 ? n1924 : n1992;
  assign n1994 = pi10 ? n1120 : n1799;
  assign n1995 = pi09 ? n26 : n1994;
  assign n1996 = pi08 ? n26 : n1995;
  assign n1997 = pi07 ? n1996 : n1815;
  assign n1998 = pi06 ? n1997 : n1840;
  assign n1999 = pi05 ? n1813 : n1998;
  assign n2000 = pi04 ? n1797 : n1999;
  assign n2001 = pi10 ? n1369 : n1852;
  assign n2002 = pi09 ? n26 : n2001;
  assign n2003 = pi08 ? n26 : n2002;
  assign n2004 = pi13 ? n46 : ~n130;
  assign n2005 = pi12 ? n26 : n2004;
  assign n2006 = pi10 ? n2005 : n1585;
  assign n2007 = pi09 ? n2006 : n1585;
  assign n2008 = pi08 ? n2007 : n1585;
  assign n2009 = pi07 ? n2003 : n2008;
  assign n2010 = pi06 ? n2009 : n1870;
  assign n2011 = pi14 ? n26 : ~n1638;
  assign n2012 = pi13 ? n2011 : ~n57;
  assign n2013 = pi12 ? n26 : n2012;
  assign n2014 = pi11 ? n2013 : n1610;
  assign n2015 = pi10 ? n1413 : n2014;
  assign n2016 = pi09 ? n26 : n2015;
  assign n2017 = pi08 ? n26 : n2016;
  assign n2018 = pi10 ? n1882 : n26;
  assign n2019 = pi09 ? n2018 : n26;
  assign n2020 = pi08 ? n2019 : n26;
  assign n2021 = pi07 ? n2017 : n2020;
  assign n2022 = pi06 ? n2021 : n26;
  assign n2023 = pi05 ? n2010 : n2022;
  assign n2024 = pi10 ? n1413 : n410;
  assign n2025 = pi09 ? n26 : n2024;
  assign n2026 = pi08 ? n26 : n2025;
  assign n2027 = pi11 ? n300 : n1895;
  assign n2028 = pi10 ? n2027 : n26;
  assign n2029 = pi09 ? n2028 : n26;
  assign n2030 = pi08 ? n2029 : n26;
  assign n2031 = pi07 ? n2026 : n2030;
  assign n2032 = pi06 ? n2031 : n26;
  assign n2033 = pi13 ? n143 : ~n284;
  assign n2034 = pi12 ? n26 : n2033;
  assign n2035 = pi11 ? n26 : n2034;
  assign n2036 = pi10 ? n2035 : n537;
  assign n2037 = pi09 ? n26 : n2036;
  assign n2038 = pi08 ? n26 : n2037;
  assign n2039 = pi11 ? n1183 : n447;
  assign n2040 = pi11 ? n1916 : n872;
  assign n2041 = pi10 ? n2039 : n2040;
  assign n2042 = pi09 ? n2041 : n872;
  assign n2043 = pi08 ? n2042 : n872;
  assign n2044 = pi07 ? n2038 : n2043;
  assign n2045 = pi10 ? n876 : n872;
  assign n2046 = pi09 ? n2045 : n872;
  assign n2047 = pi08 ? n1674 : n2046;
  assign n2048 = pi07 ? n2047 : n872;
  assign n2049 = pi06 ? n2044 : n2048;
  assign n2050 = pi05 ? n2032 : n2049;
  assign n2051 = pi04 ? n2023 : n2050;
  assign n2052 = pi03 ? n2000 : n2051;
  assign n2053 = pi02 ? n1993 : n2052;
  assign n2054 = pi10 ? n1566 : n1952;
  assign n2055 = pi09 ? n26 : n2054;
  assign n2056 = pi08 ? n26 : n2055;
  assign n2057 = pi11 ? n1008 : n1934;
  assign n2058 = pi15 ? n70 : ~n28;
  assign n2059 = pi14 ? n2058 : ~n45;
  assign n2060 = pi13 ? n2059 : n26;
  assign n2061 = pi12 ? n26 : n2060;
  assign n2062 = pi11 ? n2061 : n1941;
  assign n2063 = pi10 ? n2057 : n2062;
  assign n2064 = pi11 ? n343 : n274;
  assign n2065 = pi10 ? n2064 : n274;
  assign n2066 = pi09 ? n2063 : n2065;
  assign n2067 = pi08 ? n2066 : n274;
  assign n2068 = pi07 ? n2056 : n2067;
  assign n2069 = pi06 ? n2068 : n1698;
  assign n2070 = pi14 ? n71 : n37;
  assign n2071 = pi13 ? n176 : ~n2070;
  assign n2072 = pi12 ? n26 : n2071;
  assign n2073 = pi11 ? n26 : n2072;
  assign n2074 = pi10 ? n2073 : n1785;
  assign n2075 = pi09 ? n26 : n2074;
  assign n2076 = pi08 ? n26 : n2075;
  assign n2077 = pi11 ? n366 : n1144;
  assign n2078 = pi13 ? n1914 : ~n126;
  assign n2079 = pi12 ? n26 : n2078;
  assign n2080 = pi11 ? n867 : n2079;
  assign n2081 = pi10 ? n2077 : n2080;
  assign n2082 = pi10 ? n343 : n1689;
  assign n2083 = pi09 ? n2081 : n2082;
  assign n2084 = pi08 ? n2083 : n343;
  assign n2085 = pi07 ? n2076 : n2084;
  assign n2086 = pi06 ? n2085 : n343;
  assign n2087 = pi05 ? n2069 : n2086;
  assign n2088 = pi13 ? n176 : ~n1925;
  assign n2089 = pi12 ? n26 : n2088;
  assign n2090 = pi11 ? n26 : n2089;
  assign n2091 = pi10 ? n2090 : n537;
  assign n2092 = pi09 ? n26 : n2091;
  assign n2093 = pi08 ? n26 : n2092;
  assign n2094 = pi11 ? n523 : n1598;
  assign n2095 = pi11 ? n395 : n1733;
  assign n2096 = pi10 ? n2094 : n2095;
  assign n2097 = pi10 ? n1736 : n1735;
  assign n2098 = pi09 ? n2096 : n2097;
  assign n2099 = pi08 ? n2098 : n1735;
  assign n2100 = pi07 ? n2093 : n2099;
  assign n2101 = pi11 ? n422 : n671;
  assign n2102 = pi10 ? n1735 : n2101;
  assign n2103 = pi11 ? n398 : n1735;
  assign n2104 = pi10 ? n646 : n2103;
  assign n2105 = pi09 ? n2102 : n2104;
  assign n2106 = pi08 ? n2105 : n1735;
  assign n2107 = pi13 ? n723 : ~n126;
  assign n2108 = pi12 ? n26 : n2107;
  assign n2109 = pi11 ? n1733 : n2108;
  assign n2110 = pi10 ? n1735 : n2109;
  assign n2111 = pi09 ? n1735 : n2110;
  assign n2112 = pi08 ? n1735 : n2111;
  assign n2113 = pi07 ? n2106 : n2112;
  assign n2114 = pi06 ? n2100 : n2113;
  assign n2115 = pi10 ? n26 : n297;
  assign n2116 = pi13 ? n79 : n26;
  assign n2117 = pi12 ? n26 : n2116;
  assign n2118 = pi11 ? n2117 : n1071;
  assign n2119 = pi10 ? n2118 : n26;
  assign n2120 = pi09 ? n2115 : n2119;
  assign n2121 = pi08 ? n2120 : n26;
  assign n2122 = pi07 ? n2121 : n26;
  assign n2123 = pi06 ? n26 : n2122;
  assign n2124 = pi05 ? n2114 : n2123;
  assign n2125 = pi04 ? n2087 : n2124;
  assign n2126 = pi11 ? n1766 : n1595;
  assign n2127 = pi10 ? n26 : n2126;
  assign n2128 = pi11 ? n1750 : n1790;
  assign n2129 = pi10 ? n2128 : n26;
  assign n2130 = pi09 ? n2127 : n2129;
  assign n2131 = pi08 ? n2130 : n26;
  assign n2132 = pi07 ? n2131 : n26;
  assign n2133 = pi06 ? n26 : n2132;
  assign n2134 = pi10 ? n725 : n1779;
  assign n2135 = pi09 ? n725 : n2134;
  assign n2136 = pi08 ? n725 : n2135;
  assign n2137 = pi07 ? n1251 : n2136;
  assign n2138 = pi11 ? n1093 : n1312;
  assign n2139 = pi13 ? n130 : ~n1591;
  assign n2140 = pi12 ? n26 : n2139;
  assign n2141 = pi11 ? n2089 : n2140;
  assign n2142 = pi10 ? n2138 : n2141;
  assign n2143 = pi11 ? n447 : n1807;
  assign n2144 = pi14 ? n292 : n125;
  assign n2145 = pi13 ? n2144 : ~n26;
  assign n2146 = pi12 ? n69 : ~n2145;
  assign n2147 = pi11 ? n1197 : n2146;
  assign n2148 = pi10 ? n2143 : n2147;
  assign n2149 = pi09 ? n2142 : n2148;
  assign n2150 = pi08 ? n2149 : n872;
  assign n2151 = pi07 ? n2150 : n872;
  assign n2152 = pi06 ? n2137 : n2151;
  assign n2153 = pi05 ? n2133 : n2152;
  assign n2154 = pi10 ? n263 : n1799;
  assign n2155 = pi09 ? n263 : n2154;
  assign n2156 = pi08 ? n263 : n2155;
  assign n2157 = pi07 ? n1278 : n2156;
  assign n2158 = pi11 ? n1110 : n731;
  assign n2159 = pi14 ? n233 : n125;
  assign n2160 = pi13 ? n130 : ~n2159;
  assign n2161 = pi12 ? n26 : n2160;
  assign n2162 = pi11 ? n178 : n2161;
  assign n2163 = pi10 ? n2158 : n2162;
  assign n2164 = pi11 ? n1137 : n1807;
  assign n2165 = pi14 ? n63 : n45;
  assign n2166 = pi13 ? n2165 : ~n26;
  assign n2167 = pi12 ? n26 : ~n2166;
  assign n2168 = pi11 ? n2167 : n343;
  assign n2169 = pi10 ? n2164 : n2168;
  assign n2170 = pi09 ? n2163 : n2169;
  assign n2171 = pi08 ? n2170 : n274;
  assign n2172 = pi07 ? n2171 : n1697;
  assign n2173 = pi06 ? n2157 : n2172;
  assign n2174 = pi15 ? n28 : ~n291;
  assign n2175 = pi14 ? n26 : n2174;
  assign n2176 = pi13 ? n2175 : ~n143;
  assign n2177 = pi12 ? n26 : n2176;
  assign n2178 = pi11 ? n2177 : n1475;
  assign n2179 = pi10 ? n2178 : n1133;
  assign n2180 = pi13 ? n1135 : n38;
  assign n2181 = pi12 ? n26 : ~n2180;
  assign n2182 = pi11 ? n2181 : n1141;
  assign n2183 = pi13 ? n269 : n126;
  assign n2184 = pi12 ? n26 : ~n2183;
  assign n2185 = pi11 ? n1787 : n2184;
  assign n2186 = pi10 ? n2182 : n2185;
  assign n2187 = pi09 ? n2179 : n2186;
  assign n2188 = pi09 ? n2082 : n343;
  assign n2189 = pi08 ? n2187 : n2188;
  assign n2190 = pi07 ? n2189 : n343;
  assign n2191 = pi06 ? n1997 : n2190;
  assign n2192 = pi05 ? n2173 : n2191;
  assign n2193 = pi04 ? n2153 : n2192;
  assign n2194 = pi03 ? n2125 : n2193;
  assign n2195 = pi10 ? n1310 : n962;
  assign n2196 = pi09 ? n26 : n2195;
  assign n2197 = pi08 ? n26 : n2196;
  assign n2198 = pi09 ? n1607 : n1588;
  assign n2199 = pi08 ? n2198 : n1588;
  assign n2200 = pi07 ? n2197 : n2199;
  assign n2201 = pi14 ? n26 : ~n517;
  assign n2202 = pi13 ? n2201 : ~n130;
  assign n2203 = pi12 ? n26 : n2202;
  assign n2204 = pi11 ? n2203 : n516;
  assign n2205 = pi10 ? n2204 : n537;
  assign n2206 = pi14 ? n45 : ~n163;
  assign n2207 = pi13 ? n2206 : ~n72;
  assign n2208 = pi12 ? n26 : n2207;
  assign n2209 = pi11 ? n523 : n2208;
  assign n2210 = pi10 ? n300 : n2209;
  assign n2211 = pi09 ? n2205 : n2210;
  assign n2212 = pi09 ? n2097 : n1735;
  assign n2213 = pi08 ? n2211 : n2212;
  assign n2214 = pi07 ? n2213 : n2112;
  assign n2215 = pi06 ? n2200 : n2214;
  assign n2216 = pi10 ? n1369 : n1161;
  assign n2217 = pi09 ? n26 : n2216;
  assign n2218 = pi08 ? n26 : n2217;
  assign n2219 = pi07 ? n2218 : n2020;
  assign n2220 = pi06 ? n2219 : n26;
  assign n2221 = pi05 ? n2215 : n2220;
  assign n2222 = pi10 ? n1413 : n1421;
  assign n2223 = pi09 ? n26 : n2222;
  assign n2224 = pi08 ? n26 : n2223;
  assign n2225 = pi14 ? n28 : ~n26;
  assign n2226 = pi13 ? n2225 : ~n72;
  assign n2227 = pi12 ? n26 : n2226;
  assign n2228 = pi14 ? n73 : ~n292;
  assign n2229 = pi13 ? n2228 : ~n126;
  assign n2230 = pi12 ? n26 : n2229;
  assign n2231 = pi11 ? n2227 : n2230;
  assign n2232 = pi10 ? n2231 : n26;
  assign n2233 = pi09 ? n2232 : n26;
  assign n2234 = pi08 ? n2233 : n26;
  assign n2235 = pi07 ? n2224 : n2234;
  assign n2236 = pi06 ? n2235 : n26;
  assign n2237 = pi11 ? n410 : n1632;
  assign n2238 = pi10 ? n2035 : n2237;
  assign n2239 = pi09 ? n26 : n2238;
  assign n2240 = pi08 ? n26 : n2239;
  assign n2241 = pi11 ? n1575 : n447;
  assign n2242 = pi10 ? n2241 : n2040;
  assign n2243 = pi13 ? n26 : n773;
  assign n2244 = pi12 ? n2243 : ~n135;
  assign n2245 = pi11 ? n2244 : n136;
  assign n2246 = pi10 ? n2245 : n875;
  assign n2247 = pi09 ? n2242 : n2246;
  assign n2248 = pi08 ? n2247 : n875;
  assign n2249 = pi07 ? n2240 : n2248;
  assign n2250 = pi06 ? n2249 : n875;
  assign n2251 = pi05 ? n2236 : n2250;
  assign n2252 = pi04 ? n2221 : n2251;
  assign n2253 = pi15 ? n60 : n28;
  assign n2254 = pi14 ? n2253 : n45;
  assign n2255 = pi13 ? n2254 : ~n26;
  assign n2256 = pi12 ? n26 : ~n2255;
  assign n2257 = pi11 ? n2256 : n1941;
  assign n2258 = pi10 ? n2039 : n2257;
  assign n2259 = pi11 ? n1206 : n274;
  assign n2260 = pi10 ? n2259 : n274;
  assign n2261 = pi09 ? n2258 : n2260;
  assign n2262 = pi08 ? n2261 : n274;
  assign n2263 = pi07 ? n2056 : n2262;
  assign n2264 = pi06 ? n2263 : n1698;
  assign n2265 = pi12 ? n26 : ~n1195;
  assign n2266 = pi11 ? n2265 : n1667;
  assign n2267 = pi10 ? n2039 : n2266;
  assign n2268 = pi10 ? n343 : n2064;
  assign n2269 = pi09 ? n2267 : n2268;
  assign n2270 = pi08 ? n2269 : n274;
  assign n2271 = pi07 ? n2076 : n2270;
  assign n2272 = pi06 ? n2271 : n1698;
  assign n2273 = pi05 ? n2264 : n2272;
  assign n2274 = pi10 ? n2073 : n1952;
  assign n2275 = pi09 ? n26 : n2274;
  assign n2276 = pi08 ? n26 : n2275;
  assign n2277 = pi13 ? n396 : ~n126;
  assign n2278 = pi12 ? n26 : n2277;
  assign n2279 = pi11 ? n560 : n2278;
  assign n2280 = pi10 ? n369 : n2279;
  assign n2281 = pi11 ? n1711 : n2278;
  assign n2282 = pi10 ? n2281 : n1711;
  assign n2283 = pi09 ? n2280 : n2282;
  assign n2284 = pi08 ? n2283 : n560;
  assign n2285 = pi07 ? n2276 : n2284;
  assign n2286 = pi06 ? n2285 : n560;
  assign n2287 = pi11 ? n395 : n419;
  assign n2288 = pi10 ? n2094 : n2287;
  assign n2289 = pi13 ? n1252 : ~n72;
  assign n2290 = pi12 ? n26 : n2289;
  assign n2291 = pi11 ? n2290 : n1733;
  assign n2292 = pi10 ? n2291 : n1735;
  assign n2293 = pi09 ? n2288 : n2292;
  assign n2294 = pi08 ? n2293 : n422;
  assign n2295 = pi07 ? n1726 : n2294;
  assign n2296 = pi10 ? n422 : n1062;
  assign n2297 = pi09 ? n422 : n2296;
  assign n2298 = pi08 ? n422 : n2297;
  assign n2299 = pi07 ? n422 : n2298;
  assign n2300 = pi06 ? n2295 : n2299;
  assign n2301 = pi05 ? n2286 : n2300;
  assign n2302 = pi04 ? n2273 : n2301;
  assign n2303 = pi03 ? n2252 : n2302;
  assign n2304 = pi02 ? n2194 : n2303;
  assign n2305 = pi01 ? n2053 : n2304;
  assign n2306 = pi00 ? n1846 : n2305;
  assign n2307 = pi12 ? n26 : n69;
  assign n2308 = pi11 ? n26 : n2307;
  assign n2309 = pi10 ? n2308 : n2307;
  assign n2310 = pi09 ? n26 : n2309;
  assign n2311 = pi08 ? n26 : n2310;
  assign n2312 = pi14 ? n73 : n45;
  assign n2313 = pi13 ? n26 : n2312;
  assign n2314 = pi12 ? n26 : n2313;
  assign n2315 = pi14 ? n233 : n45;
  assign n2316 = pi13 ? n26 : n2315;
  assign n2317 = pi12 ? n26 : n2316;
  assign n2318 = pi11 ? n2314 : n2317;
  assign n2319 = pi14 ? n37 : n26;
  assign n2320 = pi13 ? n321 : n2319;
  assign n2321 = pi12 ? n26 : n2320;
  assign n2322 = pi13 ? n653 : n1705;
  assign n2323 = pi12 ? n26 : n2322;
  assign n2324 = pi11 ? n2321 : n2323;
  assign n2325 = pi10 ? n2318 : n2324;
  assign n2326 = pi09 ? n2307 : n2325;
  assign n2327 = pi08 ? n2326 : n2310;
  assign n2328 = pi07 ? n2311 : n2327;
  assign n2329 = pi09 ? n2325 : n26;
  assign n2330 = pi09 ? n2309 : n2325;
  assign n2331 = pi08 ? n2329 : n2330;
  assign n2332 = pi14 ? n73 : n26;
  assign n2333 = pi13 ? n26 : n2332;
  assign n2334 = pi12 ? n26 : n2333;
  assign n2335 = pi11 ? n26 : n2334;
  assign n2336 = pi10 ? n26 : n2335;
  assign n2337 = pi09 ? n26 : n2336;
  assign n2338 = pi13 ? n26 : n1705;
  assign n2339 = pi12 ? n26 : n2338;
  assign n2340 = pi13 ? n26 : n639;
  assign n2341 = pi12 ? n26 : n2340;
  assign n2342 = pi11 ? n2339 : n2341;
  assign n2343 = pi10 ? n26 : n2342;
  assign n2344 = pi13 ? n653 : n26;
  assign n2345 = pi12 ? n26 : n2344;
  assign n2346 = pi11 ? n26 : n2345;
  assign n2347 = pi14 ? n327 : n26;
  assign n2348 = pi13 ? n2347 : n26;
  assign n2349 = pi12 ? n26 : n2348;
  assign n2350 = pi11 ? n26 : n2349;
  assign n2351 = pi10 ? n2346 : n2350;
  assign n2352 = pi09 ? n2343 : n2351;
  assign n2353 = pi08 ? n2337 : n2352;
  assign n2354 = pi07 ? n2331 : n2353;
  assign n2355 = pi06 ? n2328 : n2354;
  assign n2356 = pi05 ? n26 : n2355;
  assign n2357 = pi13 ? n143 : n68;
  assign n2358 = pi12 ? n26 : n2357;
  assign n2359 = pi13 ? n176 : n77;
  assign n2360 = pi12 ? n26 : n2359;
  assign n2361 = pi10 ? n2358 : n2360;
  assign n2362 = pi13 ? n143 : n77;
  assign n2363 = pi12 ? n26 : n2362;
  assign n2364 = pi11 ? n2360 : n2363;
  assign n2365 = pi13 ? n26 : n1280;
  assign n2366 = pi12 ? n26 : n2365;
  assign n2367 = pi11 ? n2358 : n2366;
  assign n2368 = pi10 ? n2364 : n2367;
  assign n2369 = pi09 ? n2361 : n2368;
  assign n2370 = pi14 ? n29 : n26;
  assign n2371 = pi13 ? n26 : n2370;
  assign n2372 = pi12 ? n26 : n2371;
  assign n2373 = pi11 ? n2372 : n2341;
  assign n2374 = pi10 ? n2373 : n26;
  assign n2375 = pi10 ? n2308 : n2360;
  assign n2376 = pi09 ? n2374 : n2375;
  assign n2377 = pi08 ? n2369 : n2376;
  assign n2378 = pi07 ? n2311 : n2377;
  assign n2379 = pi09 ? n2368 : n2374;
  assign n2380 = pi09 ? n2375 : n2368;
  assign n2381 = pi08 ? n2379 : n2380;
  assign n2382 = pi10 ? n2308 : n26;
  assign n2383 = pi09 ? n2374 : n2382;
  assign n2384 = pi11 ? n2341 : n2339;
  assign n2385 = pi10 ? n2334 : n2384;
  assign n2386 = pi15 ? n26 : ~n70;
  assign n2387 = pi14 ? n26 : n2386;
  assign n2388 = pi13 ? n2387 : n1280;
  assign n2389 = pi12 ? n26 : n2388;
  assign n2390 = pi11 ? n2389 : n26;
  assign n2391 = pi14 ? n45 : ~n125;
  assign n2392 = pi13 ? n2391 : n26;
  assign n2393 = pi12 ? n26 : n2392;
  assign n2394 = pi14 ? n71 : ~n125;
  assign n2395 = pi13 ? n2394 : n26;
  assign n2396 = pi12 ? n654 : n2395;
  assign n2397 = pi11 ? n2393 : n2396;
  assign n2398 = pi10 ? n2390 : n2397;
  assign n2399 = pi09 ? n2385 : n2398;
  assign n2400 = pi08 ? n2383 : n2399;
  assign n2401 = pi07 ? n2381 : n2400;
  assign n2402 = pi06 ? n2378 : n2401;
  assign n2403 = pi14 ? n26 : n1704;
  assign n2404 = pi13 ? n2403 : n2387;
  assign n2405 = pi12 ? n26 : n2404;
  assign n2406 = pi11 ? n26 : n2405;
  assign n2407 = pi14 ? n63 : ~n1872;
  assign n2408 = pi13 ? n2407 : n787;
  assign n2409 = pi12 ? n26 : n2408;
  assign n2410 = pi15 ? n70 : ~n291;
  assign n2411 = pi14 ? n26 : ~n2410;
  assign n2412 = pi13 ? n2411 : n787;
  assign n2413 = pi12 ? n26 : n2412;
  assign n2414 = pi11 ? n2409 : n2413;
  assign n2415 = pi10 ? n2406 : n2414;
  assign n2416 = pi09 ? n26 : n2415;
  assign n2417 = pi08 ? n26 : n2416;
  assign n2418 = pi13 ? n321 : n787;
  assign n2419 = pi12 ? n26 : n2418;
  assign n2420 = pi15 ? n60 : ~n44;
  assign n2421 = pi14 ? n26 : n2420;
  assign n2422 = pi13 ? n2421 : n787;
  assign n2423 = pi12 ? n26 : n2422;
  assign n2424 = pi11 ? n2419 : n2423;
  assign n2425 = pi13 ? n2421 : n2387;
  assign n2426 = pi12 ? n26 : n2425;
  assign n2427 = pi13 ? n321 : n2387;
  assign n2428 = pi12 ? n26 : n2427;
  assign n2429 = pi11 ? n2426 : n2428;
  assign n2430 = pi10 ? n2424 : n2429;
  assign n2431 = pi15 ? n291 : ~n44;
  assign n2432 = pi14 ? n26 : n2431;
  assign n2433 = pi13 ? n2432 : n2387;
  assign n2434 = pi12 ? n26 : n2433;
  assign n2435 = pi11 ? n2434 : n2428;
  assign n2436 = pi10 ? n2435 : n2367;
  assign n2437 = pi09 ? n2430 : n2436;
  assign n2438 = pi10 ? n2406 : n2428;
  assign n2439 = pi09 ? n2374 : n2438;
  assign n2440 = pi08 ? n2437 : n2439;
  assign n2441 = pi07 ? n2417 : n2440;
  assign n2442 = pi09 ? n2436 : n2374;
  assign n2443 = pi09 ? n2438 : n2436;
  assign n2444 = pi08 ? n2442 : n2443;
  assign n2445 = pi13 ? n198 : n26;
  assign n2446 = pi12 ? n26 : n2445;
  assign n2447 = pi11 ? n2446 : n26;
  assign n2448 = pi14 ? n320 : n45;
  assign n2449 = pi13 ? n26 : n2448;
  assign n2450 = pi12 ? n26 : n2449;
  assign n2451 = pi14 ? n1704 : n45;
  assign n2452 = pi13 ? n26 : n2451;
  assign n2453 = pi12 ? n26 : n2452;
  assign n2454 = pi11 ? n2450 : n2453;
  assign n2455 = pi10 ? n2447 : n2454;
  assign n2456 = pi11 ? n2307 : n26;
  assign n2457 = pi12 ? n1203 : n2392;
  assign n2458 = pi11 ? n2393 : n2457;
  assign n2459 = pi10 ? n2456 : n2458;
  assign n2460 = pi09 ? n2455 : n2459;
  assign n2461 = pi08 ? n2383 : n2460;
  assign n2462 = pi07 ? n2444 : n2461;
  assign n2463 = pi06 ? n2441 : n2462;
  assign n2464 = pi05 ? n2402 : n2463;
  assign n2465 = pi04 ? n2356 : n2464;
  assign n2466 = pi03 ? n26 : n2465;
  assign n2467 = pi02 ? n26 : n2466;
  assign n2468 = pi13 ? n143 : n2387;
  assign n2469 = pi12 ? n26 : n2468;
  assign n2470 = pi11 ? n26 : n2469;
  assign n2471 = pi13 ? n224 : n26;
  assign n2472 = pi12 ? n26 : n2471;
  assign n2473 = pi10 ? n2470 : n2472;
  assign n2474 = pi09 ? n26 : n2473;
  assign n2475 = pi08 ? n26 : n2474;
  assign n2476 = pi14 ? n26 : n61;
  assign n2477 = pi13 ? n2476 : n26;
  assign n2478 = pi12 ? n26 : n2477;
  assign n2479 = pi11 ? n2446 : n2478;
  assign n2480 = pi11 ? n2366 : n26;
  assign n2481 = pi10 ? n2479 : n2480;
  assign n2482 = pi13 ? n26 : n591;
  assign n2483 = pi12 ? n26 : n2482;
  assign n2484 = pi11 ? n26 : n2483;
  assign n2485 = pi10 ? n26 : n2484;
  assign n2486 = pi09 ? n2481 : n2485;
  assign n2487 = pi14 ? n45 : ~n168;
  assign n2488 = pi13 ? n2476 : n2487;
  assign n2489 = pi12 ? n26 : n2488;
  assign n2490 = pi11 ? n2489 : n26;
  assign n2491 = pi10 ? n2470 : n2490;
  assign n2492 = pi09 ? n2374 : n2491;
  assign n2493 = pi08 ? n2486 : n2492;
  assign n2494 = pi07 ? n2475 : n2493;
  assign n2495 = pi09 ? n2485 : n2374;
  assign n2496 = pi09 ? n2491 : n2485;
  assign n2497 = pi08 ? n2495 : n2496;
  assign n2498 = pi14 ? n26 : n292;
  assign n2499 = pi13 ? n26 : n2498;
  assign n2500 = pi12 ? n26 : n2499;
  assign n2501 = pi11 ? n26 : n2500;
  assign n2502 = pi10 ? n2501 : n2500;
  assign n2503 = pi09 ? n2374 : n2502;
  assign n2504 = pi13 ? n2347 : n2498;
  assign n2505 = pi12 ? n26 : n2504;
  assign n2506 = pi11 ? n2500 : n2505;
  assign n2507 = pi13 ? n26 : n1401;
  assign n2508 = pi12 ? n26 : n2507;
  assign n2509 = pi11 ? n2508 : n2500;
  assign n2510 = pi10 ? n2506 : n2509;
  assign n2511 = pi12 ? n1203 : n26;
  assign n2512 = pi11 ? n26 : n2511;
  assign n2513 = pi10 ? n2307 : n2512;
  assign n2514 = pi09 ? n2510 : n2513;
  assign n2515 = pi08 ? n2503 : n2514;
  assign n2516 = pi07 ? n2497 : n2515;
  assign n2517 = pi06 ? n2494 : n2516;
  assign n2518 = pi11 ? n26 : n2428;
  assign n2519 = pi14 ? n26 : ~n168;
  assign n2520 = pi13 ? n321 : n2519;
  assign n2521 = pi12 ? n26 : n2520;
  assign n2522 = pi14 ? n45 : n320;
  assign n2523 = pi13 ? n2522 : n2387;
  assign n2524 = pi12 ? n26 : n2523;
  assign n2525 = pi11 ? n2521 : n2524;
  assign n2526 = pi10 ? n2518 : n2525;
  assign n2527 = pi09 ? n26 : n2526;
  assign n2528 = pi08 ? n26 : n2527;
  assign n2529 = pi14 ? n45 : n73;
  assign n2530 = pi14 ? n45 : n2386;
  assign n2531 = pi13 ? n2529 : n2530;
  assign n2532 = pi12 ? n26 : n2531;
  assign n2533 = pi13 ? n198 : n2387;
  assign n2534 = pi12 ? n26 : n2533;
  assign n2535 = pi11 ? n2532 : n2534;
  assign n2536 = pi13 ? n26 : n2387;
  assign n2537 = pi12 ? n26 : n2536;
  assign n2538 = pi15 ? n1200 : n26;
  assign n2539 = pi14 ? n26 : n2538;
  assign n2540 = pi13 ? n2539 : n26;
  assign n2541 = pi12 ? n26 : n2540;
  assign n2542 = pi11 ? n2537 : n2541;
  assign n2543 = pi10 ? n2535 : n2542;
  assign n2544 = pi13 ? n26 : n269;
  assign n2545 = pi12 ? n26 : n2544;
  assign n2546 = pi11 ? n26 : n2545;
  assign n2547 = pi10 ? n26 : n2546;
  assign n2548 = pi09 ? n2543 : n2547;
  assign n2549 = pi14 ? n249 : n327;
  assign n2550 = pi13 ? n321 : n2549;
  assign n2551 = pi12 ? n26 : n2550;
  assign n2552 = pi11 ? n2551 : n2341;
  assign n2553 = pi10 ? n2552 : n26;
  assign n2554 = pi13 ? n149 : n2530;
  assign n2555 = pi12 ? n26 : n2554;
  assign n2556 = pi11 ? n26 : n2555;
  assign n2557 = pi14 ? n71 : ~n168;
  assign n2558 = pi13 ? n26 : n2557;
  assign n2559 = pi12 ? n26 : n2558;
  assign n2560 = pi13 ? n2498 : n26;
  assign n2561 = pi12 ? n26 : n2560;
  assign n2562 = pi11 ? n2559 : n2561;
  assign n2563 = pi10 ? n2556 : n2562;
  assign n2564 = pi09 ? n2553 : n2563;
  assign n2565 = pi08 ? n2548 : n2564;
  assign n2566 = pi07 ? n2528 : n2565;
  assign n2567 = pi09 ? n2547 : n2553;
  assign n2568 = pi09 ? n2563 : n2547;
  assign n2569 = pi08 ? n2567 : n2568;
  assign n2570 = pi14 ? n327 : n320;
  assign n2571 = pi13 ? n2570 : n2387;
  assign n2572 = pi12 ? n26 : n2571;
  assign n2573 = pi11 ? n26 : n2572;
  assign n2574 = pi14 ? n327 : n517;
  assign n2575 = pi13 ? n2574 : n2387;
  assign n2576 = pi12 ? n26 : n2575;
  assign n2577 = pi10 ? n2573 : n2576;
  assign n2578 = pi09 ? n2553 : n2577;
  assign n2579 = pi14 ? n2386 : n517;
  assign n2580 = pi13 ? n2579 : n2387;
  assign n2581 = pi12 ? n26 : n2580;
  assign n2582 = pi11 ? n2576 : n2581;
  assign n2583 = pi13 ? n773 : n2387;
  assign n2584 = pi12 ? n26 : n2583;
  assign n2585 = pi13 ? n773 : n321;
  assign n2586 = pi12 ? n26 : n2585;
  assign n2587 = pi11 ? n2584 : n2586;
  assign n2588 = pi10 ? n2582 : n2587;
  assign n2589 = pi13 ? n773 : n26;
  assign n2590 = pi12 ? n26 : n2589;
  assign n2591 = pi11 ? n2590 : n26;
  assign n2592 = pi10 ? n2591 : n26;
  assign n2593 = pi09 ? n2588 : n2592;
  assign n2594 = pi08 ? n2578 : n2593;
  assign n2595 = pi07 ? n2569 : n2594;
  assign n2596 = pi06 ? n2566 : n2595;
  assign n2597 = pi05 ? n2517 : n2596;
  assign n2598 = pi14 ? n71 : n26;
  assign n2599 = pi13 ? n2598 : n2530;
  assign n2600 = pi12 ? n26 : n2599;
  assign n2601 = pi11 ? n2349 : n2600;
  assign n2602 = pi10 ? n2573 : n2601;
  assign n2603 = pi09 ? n26 : n2602;
  assign n2604 = pi08 ? n26 : n2603;
  assign n2605 = pi13 ? n2598 : n26;
  assign n2606 = pi12 ? n26 : n2605;
  assign n2607 = pi11 ? n2606 : n2446;
  assign n2608 = pi10 ? n2607 : n2447;
  assign n2609 = pi10 ? n26 : n2308;
  assign n2610 = pi09 ? n2608 : n2609;
  assign n2611 = pi13 ? n321 : n68;
  assign n2612 = pi12 ? n26 : n2611;
  assign n2613 = pi13 ? n2387 : n143;
  assign n2614 = pi12 ? n26 : n2613;
  assign n2615 = pi14 ? n327 : n2386;
  assign n2616 = pi13 ? n26 : n2615;
  assign n2617 = pi12 ? n26 : n2616;
  assign n2618 = pi11 ? n2614 : n2617;
  assign n2619 = pi11 ? n2559 : n2541;
  assign n2620 = pi10 ? n2618 : n2619;
  assign n2621 = pi09 ? n2612 : n2620;
  assign n2622 = pi08 ? n2610 : n2621;
  assign n2623 = pi07 ? n2604 : n2622;
  assign n2624 = pi09 ? n2609 : n2612;
  assign n2625 = pi09 ? n2620 : n2609;
  assign n2626 = pi08 ? n2624 : n2625;
  assign n2627 = pi14 ? n2386 : n786;
  assign n2628 = pi13 ? n2627 : n2387;
  assign n2629 = pi12 ? n26 : n2628;
  assign n2630 = pi11 ? n2307 : n2629;
  assign n2631 = pi14 ? n2386 : n26;
  assign n2632 = pi13 ? n2631 : n26;
  assign n2633 = pi12 ? n26 : n2632;
  assign n2634 = pi10 ? n2630 : n2633;
  assign n2635 = pi09 ? n2612 : n2634;
  assign n2636 = pi11 ? n2633 : n26;
  assign n2637 = pi10 ? n2636 : n26;
  assign n2638 = pi12 ? n26 : n1280;
  assign n2639 = pi11 ? n2366 : n2638;
  assign n2640 = pi13 ? n639 : n26;
  assign n2641 = pi12 ? n26 : n2640;
  assign n2642 = pi14 ? n1330 : ~n26;
  assign n2643 = pi13 ? n2642 : n507;
  assign n2644 = pi12 ? n26 : ~n2643;
  assign n2645 = pi11 ? n2641 : n2644;
  assign n2646 = pi10 ? n2639 : n2645;
  assign n2647 = pi09 ? n2637 : n2646;
  assign n2648 = pi08 ? n2635 : n2647;
  assign n2649 = pi07 ? n2626 : n2648;
  assign n2650 = pi06 ? n2623 : n2649;
  assign n2651 = pi13 ? n2631 : n2387;
  assign n2652 = pi12 ? n26 : n2651;
  assign n2653 = pi11 ? n26 : n2652;
  assign n2654 = pi13 ? n639 : n2487;
  assign n2655 = pi12 ? n26 : n2654;
  assign n2656 = pi11 ? n2655 : n2641;
  assign n2657 = pi10 ? n2653 : n2656;
  assign n2658 = pi09 ? n26 : n2657;
  assign n2659 = pi08 ? n26 : n2658;
  assign n2660 = pi13 ? n2319 : n97;
  assign n2661 = pi12 ? n26 : n2660;
  assign n2662 = pi11 ? n2641 : n2661;
  assign n2663 = pi13 ? n1280 : n26;
  assign n2664 = pi12 ? n26 : n2663;
  assign n2665 = pi11 ? n2664 : n2446;
  assign n2666 = pi10 ? n2662 : n2665;
  assign n2667 = pi13 ? n2403 : n26;
  assign n2668 = pi12 ? n26 : n2667;
  assign n2669 = pi11 ? n26 : n2668;
  assign n2670 = pi10 ? n26 : n2669;
  assign n2671 = pi09 ? n2666 : n2670;
  assign n2672 = pi11 ? n2358 : n2360;
  assign n2673 = pi10 ? n2672 : n2360;
  assign n2674 = pi13 ? n250 : n1523;
  assign n2675 = pi12 ? n26 : n2674;
  assign n2676 = pi14 ? n327 : n1638;
  assign n2677 = pi13 ? n198 : n2676;
  assign n2678 = pi12 ? n26 : n2677;
  assign n2679 = pi11 ? n2675 : n2678;
  assign n2680 = pi13 ? n198 : n2391;
  assign n2681 = pi12 ? n26 : n2680;
  assign n2682 = pi13 ? n26 : n1850;
  assign n2683 = pi12 ? n26 : n2682;
  assign n2684 = pi11 ? n2681 : n2683;
  assign n2685 = pi10 ? n2679 : n2684;
  assign n2686 = pi09 ? n2673 : n2685;
  assign n2687 = pi08 ? n2671 : n2686;
  assign n2688 = pi07 ? n2659 : n2687;
  assign n2689 = pi09 ? n2670 : n2673;
  assign n2690 = pi09 ? n2685 : n2670;
  assign n2691 = pi08 ? n2689 : n2690;
  assign n2692 = pi13 ? n250 : n77;
  assign n2693 = pi12 ? n26 : n2692;
  assign n2694 = pi11 ? n2693 : n2405;
  assign n2695 = pi11 ? n26 : n2537;
  assign n2696 = pi10 ? n2694 : n2695;
  assign n2697 = pi09 ? n2673 : n2696;
  assign n2698 = pi14 ? n292 : n26;
  assign n2699 = pi14 ? n26 : ~n70;
  assign n2700 = pi13 ? n2698 : n2699;
  assign n2701 = pi12 ? n26 : n2700;
  assign n2702 = pi11 ? n2537 : n2701;
  assign n2703 = pi13 ? n2698 : n2387;
  assign n2704 = pi12 ? n26 : n2703;
  assign n2705 = pi11 ? n2704 : n2537;
  assign n2706 = pi10 ? n2702 : n2705;
  assign n2707 = pi13 ? n26 : n2530;
  assign n2708 = pi12 ? n26 : n2707;
  assign n2709 = pi14 ? n1400 : n2386;
  assign n2710 = pi13 ? n26 : n2709;
  assign n2711 = pi12 ? n26 : n2710;
  assign n2712 = pi11 ? n2708 : n2711;
  assign n2713 = pi14 ? n1704 : n292;
  assign n2714 = pi13 ? n2713 : n26;
  assign n2715 = pi12 ? n26 : n2714;
  assign n2716 = pi13 ? n1553 : ~n26;
  assign n2717 = pi12 ? n26 : ~n2716;
  assign n2718 = pi11 ? n2715 : n2717;
  assign n2719 = pi10 ? n2712 : n2718;
  assign n2720 = pi09 ? n2706 : n2719;
  assign n2721 = pi08 ? n2697 : n2720;
  assign n2722 = pi07 ? n2691 : n2721;
  assign n2723 = pi06 ? n2688 : n2722;
  assign n2724 = pi05 ? n2650 : n2723;
  assign n2725 = pi04 ? n2597 : n2724;
  assign n2726 = pi11 ? n26 : n2708;
  assign n2727 = pi14 ? n71 : n2386;
  assign n2728 = pi13 ? n2332 : n2727;
  assign n2729 = pi12 ? n26 : n2728;
  assign n2730 = pi11 ? n2366 : n2729;
  assign n2731 = pi10 ? n2726 : n2730;
  assign n2732 = pi09 ? n26 : n2731;
  assign n2733 = pi08 ? n26 : n2732;
  assign n2734 = pi14 ? n131 : n26;
  assign n2735 = pi13 ? n2734 : n26;
  assign n2736 = pi12 ? n26 : n2735;
  assign n2737 = pi14 ? n1138 : n26;
  assign n2738 = pi13 ? n2737 : n26;
  assign n2739 = pi12 ? n26 : n2738;
  assign n2740 = pi11 ? n2736 : n2739;
  assign n2741 = pi14 ? n1400 : n26;
  assign n2742 = pi13 ? n2741 : n26;
  assign n2743 = pi12 ? n26 : n2742;
  assign n2744 = pi15 ? n1200 : n28;
  assign n2745 = pi14 ? n2744 : n26;
  assign n2746 = pi13 ? n2745 : n26;
  assign n2747 = pi12 ? n26 : n2746;
  assign n2748 = pi11 ? n2743 : n2747;
  assign n2749 = pi10 ? n2740 : n2748;
  assign n2750 = pi13 ? n143 : n26;
  assign n2751 = pi12 ? n26 : n2750;
  assign n2752 = pi11 ? n26 : n2751;
  assign n2753 = pi10 ? n26 : n2752;
  assign n2754 = pi09 ? n2749 : n2753;
  assign n2755 = pi13 ? n321 : n26;
  assign n2756 = pi12 ? n26 : n2755;
  assign n2757 = pi11 ? n2751 : n2756;
  assign n2758 = pi10 ? n2751 : n2757;
  assign n2759 = pi14 ? n44 : n26;
  assign n2760 = pi13 ? n26 : n2759;
  assign n2761 = pi12 ? n26 : n2760;
  assign n2762 = pi14 ? n517 : n26;
  assign n2763 = pi13 ? n2762 : n1280;
  assign n2764 = pi12 ? n26 : n2763;
  assign n2765 = pi11 ? n2761 : n2764;
  assign n2766 = pi13 ? n2762 : n26;
  assign n2767 = pi12 ? n26 : n2766;
  assign n2768 = pi11 ? n2767 : n2446;
  assign n2769 = pi10 ? n2765 : n2768;
  assign n2770 = pi09 ? n2758 : n2769;
  assign n2771 = pi08 ? n2754 : n2770;
  assign n2772 = pi07 ? n2733 : n2771;
  assign n2773 = pi09 ? n2753 : n2758;
  assign n2774 = pi09 ? n2769 : n2753;
  assign n2775 = pi08 ? n2773 : n2774;
  assign n2776 = pi13 ? n1473 : n26;
  assign n2777 = pi12 ? n26 : n2776;
  assign n2778 = pi11 ? n2751 : n2777;
  assign n2779 = pi10 ? n2778 : n2757;
  assign n2780 = pi10 ? n26 : n2756;
  assign n2781 = pi09 ? n2779 : n2780;
  assign n2782 = pi11 ? n2521 : n2756;
  assign n2783 = pi13 ? n321 : n1280;
  assign n2784 = pi12 ? n26 : n2783;
  assign n2785 = pi11 ? n2756 : n2784;
  assign n2786 = pi10 ? n2782 : n2785;
  assign n2787 = pi12 ? n26 : n124;
  assign n2788 = pi13 ? n507 : ~n2698;
  assign n2789 = pi12 ? n26 : ~n2788;
  assign n2790 = pi11 ? n2787 : n2789;
  assign n2791 = pi13 ? n2319 : n26;
  assign n2792 = pi12 ? n654 : n2791;
  assign n2793 = pi11 ? n2715 : n2792;
  assign n2794 = pi10 ? n2790 : n2793;
  assign n2795 = pi09 ? n2786 : n2794;
  assign n2796 = pi08 ? n2781 : n2795;
  assign n2797 = pi07 ? n2775 : n2796;
  assign n2798 = pi06 ? n2772 : n2797;
  assign n2799 = pi13 ? n2698 : n2347;
  assign n2800 = pi12 ? n26 : n2799;
  assign n2801 = pi11 ? n2366 : n2800;
  assign n2802 = pi10 ? n2726 : n2801;
  assign n2803 = pi09 ? n26 : n2802;
  assign n2804 = pi08 ? n26 : n2803;
  assign n2805 = pi13 ? n2698 : n97;
  assign n2806 = pi12 ? n26 : n2805;
  assign n2807 = pi14 ? n2420 : n26;
  assign n2808 = pi13 ? n2807 : n2387;
  assign n2809 = pi12 ? n26 : n2808;
  assign n2810 = pi11 ? n2806 : n2809;
  assign n2811 = pi14 ? n1832 : n26;
  assign n2812 = pi13 ? n2811 : n26;
  assign n2813 = pi12 ? n26 : n2812;
  assign n2814 = pi13 ? n1639 : ~n26;
  assign n2815 = pi12 ? n26 : ~n2814;
  assign n2816 = pi11 ? n2813 : n2815;
  assign n2817 = pi10 ? n2810 : n2816;
  assign n2818 = pi09 ? n2817 : n26;
  assign n2819 = pi08 ? n2818 : n26;
  assign n2820 = pi07 ? n2804 : n2819;
  assign n2821 = pi06 ? n2820 : n26;
  assign n2822 = pi05 ? n2798 : n2821;
  assign n2823 = pi13 ? n26 : n2487;
  assign n2824 = pi12 ? n26 : n2823;
  assign n2825 = pi11 ? n2824 : n26;
  assign n2826 = pi10 ? n2726 : n2825;
  assign n2827 = pi09 ? n26 : n2826;
  assign n2828 = pi08 ? n26 : n2827;
  assign n2829 = pi14 ? n163 : n26;
  assign n2830 = pi13 ? n2829 : n26;
  assign n2831 = pi12 ? n26 : n2830;
  assign n2832 = pi11 ? n2787 : n2831;
  assign n2833 = pi13 ? n62 : n26;
  assign n2834 = pi12 ? n26 : n2833;
  assign n2835 = pi12 ? n124 : n26;
  assign n2836 = pi11 ? n2834 : n2835;
  assign n2837 = pi10 ? n2832 : n2836;
  assign n2838 = pi09 ? n2837 : n26;
  assign n2839 = pi08 ? n2838 : n26;
  assign n2840 = pi07 ? n2828 : n2839;
  assign n2841 = pi06 ? n2840 : n26;
  assign n2842 = pi13 ? n62 : n2387;
  assign n2843 = pi12 ? n26 : n2842;
  assign n2844 = pi11 ? n2366 : n2843;
  assign n2845 = pi10 ? n2726 : n2844;
  assign n2846 = pi09 ? n26 : n2845;
  assign n2847 = pi08 ? n26 : n2846;
  assign n2848 = pi13 ? n62 : n97;
  assign n2849 = pi12 ? n26 : n2848;
  assign n2850 = pi14 ? n147 : ~n26;
  assign n2851 = pi13 ? n2850 : ~n26;
  assign n2852 = pi12 ? n26 : ~n2851;
  assign n2853 = pi11 ? n2849 : n2852;
  assign n2854 = pi12 ? n69 : n26;
  assign n2855 = pi11 ? n2835 : n2854;
  assign n2856 = pi10 ? n2853 : n2855;
  assign n2857 = pi13 ? n26 : ~n507;
  assign n2858 = pi12 ? n78 : n2857;
  assign n2859 = pi12 ? n78 : n26;
  assign n2860 = pi11 ? n2858 : n2859;
  assign n2861 = pi13 ? n26 : n2631;
  assign n2862 = pi12 ? n78 : n2861;
  assign n2863 = pi11 ? n2862 : n2859;
  assign n2864 = pi10 ? n2860 : n2863;
  assign n2865 = pi09 ? n2856 : n2864;
  assign n2866 = pi08 ? n2865 : n2859;
  assign n2867 = pi07 ? n2847 : n2866;
  assign n2868 = pi12 ? n654 : n26;
  assign n2869 = pi10 ? n2859 : n2868;
  assign n2870 = pi09 ? n2859 : n2869;
  assign n2871 = pi08 ? n2859 : n2870;
  assign n2872 = pi07 ? n2859 : n2871;
  assign n2873 = pi06 ? n2867 : n2872;
  assign n2874 = pi05 ? n2841 : n2873;
  assign n2875 = pi04 ? n2822 : n2874;
  assign n2876 = pi03 ? n2725 : n2875;
  assign n2877 = pi11 ? n2366 : n2834;
  assign n2878 = pi10 ? n2726 : n2877;
  assign n2879 = pi09 ? n26 : n2878;
  assign n2880 = pi08 ? n26 : n2879;
  assign n2881 = pi11 ? n2787 : n2664;
  assign n2882 = pi13 ? n1705 : n26;
  assign n2883 = pi12 ? n124 : n2882;
  assign n2884 = pi13 ? n478 : n26;
  assign n2885 = pi12 ? n69 : n2884;
  assign n2886 = pi11 ? n2883 : n2885;
  assign n2887 = pi10 ? n2881 : n2886;
  assign n2888 = pi13 ? n68 : n26;
  assign n2889 = pi12 ? n78 : n2888;
  assign n2890 = pi11 ? n2889 : n2859;
  assign n2891 = pi13 ? n26 : n2347;
  assign n2892 = pi12 ? n78 : n2891;
  assign n2893 = pi11 ? n2892 : n2859;
  assign n2894 = pi10 ? n2890 : n2893;
  assign n2895 = pi09 ? n2887 : n2894;
  assign n2896 = pi08 ? n2895 : n2859;
  assign n2897 = pi07 ? n2880 : n2896;
  assign n2898 = pi06 ? n2897 : n2859;
  assign n2899 = pi10 ? n2726 : n2480;
  assign n2900 = pi09 ? n26 : n2899;
  assign n2901 = pi08 ? n26 : n2900;
  assign n2902 = pi12 ? n124 : n2663;
  assign n2903 = pi11 ? n2787 : n2902;
  assign n2904 = pi14 ? n1201 : n26;
  assign n2905 = pi13 ? n2904 : n26;
  assign n2906 = pi12 ? n26 : n2905;
  assign n2907 = pi11 ? n2906 : n2854;
  assign n2908 = pi10 ? n2903 : n2907;
  assign n2909 = pi13 ? n507 : ~n26;
  assign n2910 = pi12 ? n654 : ~n2909;
  assign n2911 = pi12 ? n26 : n2888;
  assign n2912 = pi11 ? n2910 : n2911;
  assign n2913 = pi13 ? n896 : n126;
  assign n2914 = pi12 ? n26 : ~n2913;
  assign n2915 = pi13 ? n77 : ~n126;
  assign n2916 = pi12 ? n26 : n2915;
  assign n2917 = pi11 ? n2914 : n2916;
  assign n2918 = pi10 ? n2912 : n2917;
  assign n2919 = pi09 ? n2908 : n2918;
  assign n2920 = pi14 ? n1548 : ~n26;
  assign n2921 = pi13 ? n68 : ~n2920;
  assign n2922 = pi12 ? n26 : n2921;
  assign n2923 = pi11 ? n2922 : n2916;
  assign n2924 = pi10 ? n2923 : n2916;
  assign n2925 = pi09 ? n2924 : n2916;
  assign n2926 = pi08 ? n2919 : n2925;
  assign n2927 = pi07 ? n2901 : n2926;
  assign n2928 = pi12 ? n654 : n2915;
  assign n2929 = pi13 ? n77 : n26;
  assign n2930 = pi12 ? n654 : n2929;
  assign n2931 = pi11 ? n2928 : n2930;
  assign n2932 = pi10 ? n2931 : n2868;
  assign n2933 = pi09 ? n2916 : n2932;
  assign n2934 = pi08 ? n2916 : n2933;
  assign n2935 = pi07 ? n2916 : n2934;
  assign n2936 = pi06 ? n2927 : n2935;
  assign n2937 = pi05 ? n2898 : n2936;
  assign n2938 = pi11 ? n26 : n2366;
  assign n2939 = pi10 ? n2938 : n2480;
  assign n2940 = pi09 ? n26 : n2939;
  assign n2941 = pi08 ? n26 : n2940;
  assign n2942 = pi11 ? n2906 : n26;
  assign n2943 = pi10 ? n2881 : n2942;
  assign n2944 = pi13 ? n68 : n2631;
  assign n2945 = pi12 ? n26 : n2944;
  assign n2946 = pi11 ? n2868 : n2945;
  assign n2947 = pi11 ? n2911 : n2945;
  assign n2948 = pi10 ? n2946 : n2947;
  assign n2949 = pi09 ? n2943 : n2948;
  assign n2950 = pi14 ? n2386 : ~n168;
  assign n2951 = pi13 ? n68 : n2950;
  assign n2952 = pi12 ? n26 : n2951;
  assign n2953 = pi11 ? n2952 : n2945;
  assign n2954 = pi15 ? n26 : ~n1200;
  assign n2955 = pi14 ? n2954 : n26;
  assign n2956 = pi13 ? n68 : n2955;
  assign n2957 = pi12 ? n26 : n2956;
  assign n2958 = pi10 ? n2953 : n2957;
  assign n2959 = pi09 ? n2958 : n2957;
  assign n2960 = pi08 ? n2949 : n2959;
  assign n2961 = pi07 ? n2941 : n2960;
  assign n2962 = pi13 ? n26 : n198;
  assign n2963 = pi12 ? n26 : n2962;
  assign n2964 = pi13 ? n507 : ~n1280;
  assign n2965 = pi12 ? n654 : ~n2964;
  assign n2966 = pi11 ? n2963 : n2965;
  assign n2967 = pi13 ? n396 : ~n1280;
  assign n2968 = pi12 ? n26 : ~n2967;
  assign n2969 = pi13 ? n396 : ~n198;
  assign n2970 = pi12 ? n26 : ~n2969;
  assign n2971 = pi11 ? n2968 : n2970;
  assign n2972 = pi10 ? n2966 : n2971;
  assign n2973 = pi09 ? n2957 : n2972;
  assign n2974 = pi08 ? n2957 : n2973;
  assign n2975 = pi07 ? n2957 : n2974;
  assign n2976 = pi06 ? n2961 : n2975;
  assign n2977 = pi11 ? n26 : n2824;
  assign n2978 = pi10 ? n26 : n2977;
  assign n2979 = pi14 ? n37 : ~n168;
  assign n2980 = pi13 ? n2904 : n2979;
  assign n2981 = pi12 ? n26 : n2980;
  assign n2982 = pi13 ? n321 : n2487;
  assign n2983 = pi12 ? n26 : n2982;
  assign n2984 = pi11 ? n2981 : n2983;
  assign n2985 = pi13 ? n68 : n2519;
  assign n2986 = pi12 ? n26 : n2985;
  assign n2987 = pi13 ? n396 : ~n2519;
  assign n2988 = pi12 ? n26 : ~n2987;
  assign n2989 = pi11 ? n2986 : n2988;
  assign n2990 = pi10 ? n2984 : n2989;
  assign n2991 = pi09 ? n2978 : n2990;
  assign n2992 = pi08 ? n26 : n2991;
  assign n2993 = pi07 ? n26 : n2992;
  assign n2994 = pi06 ? n26 : n2993;
  assign n2995 = pi05 ? n2976 : n2994;
  assign n2996 = pi04 ? n2937 : n2995;
  assign n2997 = pi14 ? n44 : n292;
  assign n2998 = pi13 ? n26 : n2997;
  assign n2999 = pi12 ? n26 : n2998;
  assign n3000 = pi11 ? n26 : n2999;
  assign n3001 = pi10 ? n26 : n3000;
  assign n3002 = pi12 ? n26 : ~n2964;
  assign n3003 = pi14 ? n2410 : ~n26;
  assign n3004 = pi13 ? n3003 : ~n26;
  assign n3005 = pi12 ? n26 : ~n3004;
  assign n3006 = pi11 ? n3002 : n3005;
  assign n3007 = pi12 ? n26 : n2882;
  assign n3008 = pi12 ? n26 : ~n2909;
  assign n3009 = pi11 ? n3007 : n3008;
  assign n3010 = pi10 ? n3006 : n3009;
  assign n3011 = pi09 ? n3001 : n3010;
  assign n3012 = pi08 ? n26 : n3011;
  assign n3013 = pi07 ? n26 : n3012;
  assign n3014 = pi06 ? n26 : n3013;
  assign n3015 = pi07 ? n2311 : n2307;
  assign n3016 = pi12 ? n26 : n2243;
  assign n3017 = pi11 ? n2307 : n3016;
  assign n3018 = pi10 ? n2307 : n3017;
  assign n3019 = pi09 ? n2307 : n3018;
  assign n3020 = pi13 ? n2519 : n653;
  assign n3021 = pi12 ? n26 : n3020;
  assign n3022 = pi11 ? n3021 : n2537;
  assign n3023 = pi14 ? n26 : n233;
  assign n3024 = pi13 ? n2387 : n3023;
  assign n3025 = pi12 ? n26 : n3024;
  assign n3026 = pi14 ? n327 : n233;
  assign n3027 = pi13 ? n26 : n3026;
  assign n3028 = pi12 ? n26 : n3027;
  assign n3029 = pi11 ? n3025 : n3028;
  assign n3030 = pi10 ? n3022 : n3029;
  assign n3031 = pi14 ? n45 : n292;
  assign n3032 = pi13 ? n26 : n3031;
  assign n3033 = pi12 ? n26 : n3032;
  assign n3034 = pi13 ? n507 : ~n3031;
  assign n3035 = pi12 ? n26 : ~n3034;
  assign n3036 = pi11 ? n3033 : n3035;
  assign n3037 = pi13 ? n1788 : ~n26;
  assign n3038 = pi12 ? n26 : ~n3037;
  assign n3039 = pi11 ? n3007 : n3038;
  assign n3040 = pi10 ? n3036 : n3039;
  assign n3041 = pi09 ? n3030 : n3040;
  assign n3042 = pi08 ? n3019 : n3041;
  assign n3043 = pi07 ? n2307 : n3042;
  assign n3044 = pi06 ? n3015 : n3043;
  assign n3045 = pi05 ? n3014 : n3044;
  assign n3046 = pi10 ? n2308 : n2612;
  assign n3047 = pi09 ? n26 : n3046;
  assign n3048 = pi08 ? n26 : n3047;
  assign n3049 = pi07 ? n3048 : n2612;
  assign n3050 = pi13 ? n321 : n773;
  assign n3051 = pi12 ? n26 : n3050;
  assign n3052 = pi11 ? n2612 : n3051;
  assign n3053 = pi10 ? n2612 : n3052;
  assign n3054 = pi09 ? n2612 : n3053;
  assign n3055 = pi14 ? n63 : n320;
  assign n3056 = pi13 ? n3055 : n653;
  assign n3057 = pi12 ? n26 : n3056;
  assign n3058 = pi11 ? n3057 : n2428;
  assign n3059 = pi13 ? n2403 : n1583;
  assign n3060 = pi12 ? n26 : n3059;
  assign n3061 = pi14 ? n320 : ~n37;
  assign n3062 = pi13 ? n26 : n3061;
  assign n3063 = pi12 ? n26 : n3062;
  assign n3064 = pi11 ? n3060 : n3063;
  assign n3065 = pi10 ? n3058 : n3064;
  assign n3066 = pi14 ? n37 : ~n125;
  assign n3067 = pi13 ? n26 : n3066;
  assign n3068 = pi12 ? n26 : n3067;
  assign n3069 = pi13 ? n507 : ~n3066;
  assign n3070 = pi12 ? n654 : ~n3069;
  assign n3071 = pi11 ? n3068 : n3070;
  assign n3072 = pi11 ? n3007 : n2641;
  assign n3073 = pi10 ? n3071 : n3072;
  assign n3074 = pi09 ? n3065 : n3073;
  assign n3075 = pi08 ? n3054 : n3074;
  assign n3076 = pi07 ? n2612 : n3075;
  assign n3077 = pi06 ? n3049 : n3076;
  assign n3078 = pi10 ? n2470 : n2469;
  assign n3079 = pi09 ? n26 : n3078;
  assign n3080 = pi08 ? n26 : n3079;
  assign n3081 = pi11 ? n2469 : n2751;
  assign n3082 = pi10 ? n2469 : n3081;
  assign n3083 = pi11 ? n2751 : n2668;
  assign n3084 = pi13 ? n143 : n787;
  assign n3085 = pi12 ? n26 : n3084;
  assign n3086 = pi10 ? n3083 : n3085;
  assign n3087 = pi09 ? n3082 : n3086;
  assign n3088 = pi08 ? n2469 : n3087;
  assign n3089 = pi07 ? n3080 : n3088;
  assign n3090 = pi13 ? n1473 : n787;
  assign n3091 = pi12 ? n26 : n3090;
  assign n3092 = pi11 ? n3091 : n2469;
  assign n3093 = pi10 ? n2469 : n3092;
  assign n3094 = pi09 ? n2469 : n3093;
  assign n3095 = pi13 ? n2403 : n321;
  assign n3096 = pi12 ? n26 : n3095;
  assign n3097 = pi11 ? n2469 : n3096;
  assign n3098 = pi13 ? n26 : n1583;
  assign n3099 = pi12 ? n26 : n3098;
  assign n3100 = pi14 ? n26 : ~n71;
  assign n3101 = pi13 ? n26 : n3100;
  assign n3102 = pi12 ? n26 : n3101;
  assign n3103 = pi11 ? n3099 : n3102;
  assign n3104 = pi10 ? n3097 : n3103;
  assign n3105 = pi13 ? n507 : ~n2391;
  assign n3106 = pi12 ? n26 : ~n3105;
  assign n3107 = pi11 ? n3068 : n3106;
  assign n3108 = pi13 ? n1833 : ~n26;
  assign n3109 = pi12 ? n26 : ~n3108;
  assign n3110 = pi11 ? n3007 : n3109;
  assign n3111 = pi10 ? n3107 : n3110;
  assign n3112 = pi09 ? n3104 : n3111;
  assign n3113 = pi08 ? n3094 : n3112;
  assign n3114 = pi07 ? n2469 : n3113;
  assign n3115 = pi06 ? n3089 : n3114;
  assign n3116 = pi05 ? n3077 : n3115;
  assign n3117 = pi04 ? n3045 : n3116;
  assign n3118 = pi03 ? n2996 : n3117;
  assign n3119 = pi02 ? n2876 : n3118;
  assign n3120 = pi01 ? n2467 : n3119;
  assign n3121 = pi11 ? n26 : n2777;
  assign n3122 = pi10 ? n3121 : n2777;
  assign n3123 = pi09 ? n26 : n3122;
  assign n3124 = pi08 ? n26 : n3123;
  assign n3125 = pi13 ? n1473 : n2387;
  assign n3126 = pi12 ? n26 : n3125;
  assign n3127 = pi13 ? n1473 : n321;
  assign n3128 = pi12 ? n26 : n3127;
  assign n3129 = pi11 ? n3128 : n2777;
  assign n3130 = pi10 ? n3126 : n3129;
  assign n3131 = pi09 ? n2777 : n3130;
  assign n3132 = pi08 ? n2777 : n3131;
  assign n3133 = pi07 ? n3124 : n3132;
  assign n3134 = pi11 ? n2777 : n2751;
  assign n3135 = pi14 ? n2386 : n320;
  assign n3136 = pi13 ? n3135 : n68;
  assign n3137 = pi12 ? n26 : n3136;
  assign n3138 = pi11 ? n3137 : n2756;
  assign n3139 = pi10 ? n3134 : n3138;
  assign n3140 = pi09 ? n2777 : n3139;
  assign n3141 = pi11 ? n2756 : n2668;
  assign n3142 = pi10 ? n3141 : n2938;
  assign n3143 = pi12 ? n26 : n2791;
  assign n3144 = pi11 ? n2792 : n3143;
  assign n3145 = pi10 ? n26 : n3144;
  assign n3146 = pi09 ? n3142 : n3145;
  assign n3147 = pi08 ? n3140 : n3146;
  assign n3148 = pi07 ? n2777 : n3147;
  assign n3149 = pi06 ? n3133 : n3148;
  assign n3150 = pi14 ? n320 : n1872;
  assign n3151 = pi13 ? n3150 : n26;
  assign n3152 = pi12 ? n26 : n3151;
  assign n3153 = pi11 ? n26 : n3152;
  assign n3154 = pi14 ? n37 : n320;
  assign n3155 = pi13 ? n3154 : n26;
  assign n3156 = pi12 ? n26 : n3155;
  assign n3157 = pi13 ? n3154 : n1280;
  assign n3158 = pi12 ? n26 : n3157;
  assign n3159 = pi11 ? n3156 : n3158;
  assign n3160 = pi10 ? n3153 : n3159;
  assign n3161 = pi09 ? n26 : n3160;
  assign n3162 = pi08 ? n26 : n3161;
  assign n3163 = pi07 ? n26 : n3162;
  assign n3164 = pi11 ? n2641 : n26;
  assign n3165 = pi10 ? n3164 : n26;
  assign n3166 = pi09 ? n3165 : n26;
  assign n3167 = pi08 ? n3166 : n26;
  assign n3168 = pi07 ? n3167 : n26;
  assign n3169 = pi06 ? n3163 : n3168;
  assign n3170 = pi05 ? n3149 : n3169;
  assign n3171 = pi14 ? n45 : ~n70;
  assign n3172 = pi13 ? n2319 : n3171;
  assign n3173 = pi12 ? n26 : n3172;
  assign n3174 = pi13 ? n2370 : n2387;
  assign n3175 = pi12 ? n26 : n3174;
  assign n3176 = pi11 ? n3173 : n3175;
  assign n3177 = pi10 ? n2726 : n3176;
  assign n3178 = pi09 ? n26 : n3177;
  assign n3179 = pi08 ? n26 : n3178;
  assign n3180 = pi07 ? n26 : n3179;
  assign n3181 = pi14 ? n29 : n292;
  assign n3182 = pi13 ? n3181 : n26;
  assign n3183 = pi12 ? n26 : n3182;
  assign n3184 = pi11 ? n3183 : n26;
  assign n3185 = pi10 ? n3184 : n26;
  assign n3186 = pi09 ? n3185 : n26;
  assign n3187 = pi08 ? n3186 : n26;
  assign n3188 = pi07 ? n3187 : n26;
  assign n3189 = pi06 ? n3180 : n3188;
  assign n3190 = pi13 ? n26 : n336;
  assign n3191 = pi12 ? n26 : n3190;
  assign n3192 = pi11 ? n2307 : n3191;
  assign n3193 = pi10 ? n2307 : n3192;
  assign n3194 = pi13 ? n2387 : n68;
  assign n3195 = pi12 ? n26 : n3194;
  assign n3196 = pi11 ? n3195 : n2537;
  assign n3197 = pi13 ? n639 : n2557;
  assign n3198 = pi12 ? n26 : n3197;
  assign n3199 = pi11 ? n3198 : n2739;
  assign n3200 = pi10 ? n3196 : n3199;
  assign n3201 = pi09 ? n3193 : n3200;
  assign n3202 = pi08 ? n2307 : n3201;
  assign n3203 = pi07 ? n2311 : n3202;
  assign n3204 = pi13 ? n62 : ~n507;
  assign n3205 = pi12 ? n26 : n3204;
  assign n3206 = pi11 ? n2743 : n3205;
  assign n3207 = pi12 ? n26 : n2861;
  assign n3208 = pi11 ? n26 : n3207;
  assign n3209 = pi10 ? n3206 : n3208;
  assign n3210 = pi10 ? n2855 : n2859;
  assign n3211 = pi09 ? n3209 : n3210;
  assign n3212 = pi08 ? n3211 : n2859;
  assign n3213 = pi07 ? n3212 : n2871;
  assign n3214 = pi06 ? n3203 : n3213;
  assign n3215 = pi05 ? n3189 : n3214;
  assign n3216 = pi04 ? n3170 : n3215;
  assign n3217 = pi14 ? n320 : n1704;
  assign n3218 = pi13 ? n3217 : n143;
  assign n3219 = pi12 ? n26 : n3218;
  assign n3220 = pi11 ? n3219 : n2537;
  assign n3221 = pi14 ? n71 : n63;
  assign n3222 = pi13 ? n26 : n3221;
  assign n3223 = pi12 ? n26 : n3222;
  assign n3224 = pi13 ? n639 : n2387;
  assign n3225 = pi12 ? n26 : n3224;
  assign n3226 = pi11 ? n3223 : n3225;
  assign n3227 = pi10 ? n3220 : n3226;
  assign n3228 = pi09 ? n2612 : n3227;
  assign n3229 = pi08 ? n2612 : n3228;
  assign n3230 = pi07 ? n3048 : n3229;
  assign n3231 = pi14 ? n37 : n45;
  assign n3232 = pi13 ? n3231 : n2519;
  assign n3233 = pi12 ? n26 : n3232;
  assign n3234 = pi11 ? n3143 : n3233;
  assign n3235 = pi13 ? n126 : ~n2347;
  assign n3236 = pi12 ? n26 : ~n3235;
  assign n3237 = pi11 ? n2834 : n3236;
  assign n3238 = pi10 ? n3234 : n3237;
  assign n3239 = pi09 ? n3238 : n3210;
  assign n3240 = pi08 ? n3239 : n2859;
  assign n3241 = pi07 ? n3240 : n2859;
  assign n3242 = pi06 ? n3230 : n3241;
  assign n3243 = pi11 ? n2469 : n3128;
  assign n3244 = pi10 ? n3243 : n3083;
  assign n3245 = pi11 ? n26 : n2834;
  assign n3246 = pi10 ? n2825 : n3245;
  assign n3247 = pi09 ? n3244 : n3246;
  assign n3248 = pi08 ? n2469 : n3247;
  assign n3249 = pi07 ? n3080 : n3248;
  assign n3250 = pi15 ? n44 : n28;
  assign n3251 = pi14 ? n3250 : ~n26;
  assign n3252 = pi13 ? n3251 : ~n26;
  assign n3253 = pi12 ? n26 : ~n3252;
  assign n3254 = pi11 ? n3143 : n3253;
  assign n3255 = pi13 ? n68 : ~n126;
  assign n3256 = pi12 ? n26 : n3255;
  assign n3257 = pi12 ? n124 : n2915;
  assign n3258 = pi11 ? n3256 : n3257;
  assign n3259 = pi10 ? n3254 : n3258;
  assign n3260 = pi11 ? n2916 : n2922;
  assign n3261 = pi11 ? n2928 : n2916;
  assign n3262 = pi10 ? n3260 : n3261;
  assign n3263 = pi09 ? n3259 : n3262;
  assign n3264 = pi08 ? n3263 : n2916;
  assign n3265 = pi07 ? n3264 : n2934;
  assign n3266 = pi06 ? n3249 : n3265;
  assign n3267 = pi05 ? n3242 : n3266;
  assign n3268 = pi13 ? n2570 : n26;
  assign n3269 = pi12 ? n26 : n3268;
  assign n3270 = pi11 ? n26 : n3269;
  assign n3271 = pi10 ? n3270 : n3269;
  assign n3272 = pi09 ? n26 : n3271;
  assign n3273 = pi08 ? n26 : n3272;
  assign n3274 = pi10 ? n2756 : n3141;
  assign n3275 = pi13 ? n26 : n45;
  assign n3276 = pi12 ? n26 : n3275;
  assign n3277 = pi13 ? n26 : n321;
  assign n3278 = pi12 ? n26 : n3277;
  assign n3279 = pi11 ? n3278 : n2664;
  assign n3280 = pi10 ? n3276 : n3279;
  assign n3281 = pi09 ? n3274 : n3280;
  assign n3282 = pi08 ? n3269 : n3281;
  assign n3283 = pi07 ? n3273 : n3282;
  assign n3284 = pi10 ? n2641 : n2911;
  assign n3285 = pi11 ? n2945 : n2952;
  assign n3286 = pi12 ? n654 : n2944;
  assign n3287 = pi11 ? n3286 : n2957;
  assign n3288 = pi10 ? n3285 : n3287;
  assign n3289 = pi09 ? n3284 : n3288;
  assign n3290 = pi08 ? n3289 : n2957;
  assign n3291 = pi07 ? n3290 : n2974;
  assign n3292 = pi06 ? n3283 : n3291;
  assign n3293 = pi13 ? n2570 : n2487;
  assign n3294 = pi12 ? n26 : n3293;
  assign n3295 = pi11 ? n2981 : n3294;
  assign n3296 = pi10 ? n3295 : n2989;
  assign n3297 = pi09 ? n2978 : n3296;
  assign n3298 = pi08 ? n26 : n3297;
  assign n3299 = pi07 ? n26 : n3298;
  assign n3300 = pi06 ? n26 : n3299;
  assign n3301 = pi05 ? n3292 : n3300;
  assign n3302 = pi04 ? n3267 : n3301;
  assign n3303 = pi03 ? n3216 : n3302;
  assign n3304 = pi07 ? n2311 : n2612;
  assign n3305 = pi06 ? n3304 : n3076;
  assign n3306 = pi11 ? n26 : n2756;
  assign n3307 = pi13 ? n773 : n68;
  assign n3308 = pi12 ? n26 : n3307;
  assign n3309 = pi13 ? n68 : n787;
  assign n3310 = pi12 ? n26 : n3309;
  assign n3311 = pi11 ? n3308 : n3310;
  assign n3312 = pi10 ? n3306 : n3311;
  assign n3313 = pi09 ? n26 : n3312;
  assign n3314 = pi08 ? n26 : n3313;
  assign n3315 = pi07 ? n3314 : n2469;
  assign n3316 = pi06 ? n3315 : n3114;
  assign n3317 = pi05 ? n3305 : n3316;
  assign n3318 = pi04 ? n3045 : n3317;
  assign n3319 = pi11 ? n26 : n3126;
  assign n3320 = pi11 ? n3126 : n3128;
  assign n3321 = pi10 ? n3319 : n3320;
  assign n3322 = pi09 ? n26 : n3321;
  assign n3323 = pi08 ? n26 : n3322;
  assign n3324 = pi13 ? n328 : n26;
  assign n3325 = pi12 ? n26 : n3324;
  assign n3326 = pi10 ? n3325 : n2777;
  assign n3327 = pi09 ? n3326 : n2777;
  assign n3328 = pi08 ? n3327 : n2777;
  assign n3329 = pi07 ? n3323 : n3328;
  assign n3330 = pi06 ? n3329 : n3148;
  assign n3331 = pi13 ? n320 : n2387;
  assign n3332 = pi12 ? n26 : n3331;
  assign n3333 = pi11 ? n26 : n3332;
  assign n3334 = pi14 ? n320 : n1638;
  assign n3335 = pi13 ? n3334 : n2519;
  assign n3336 = pi12 ? n26 : n3335;
  assign n3337 = pi13 ? n320 : n26;
  assign n3338 = pi12 ? n26 : n3337;
  assign n3339 = pi11 ? n3336 : n3338;
  assign n3340 = pi10 ? n3333 : n3339;
  assign n3341 = pi09 ? n26 : n3340;
  assign n3342 = pi08 ? n26 : n3341;
  assign n3343 = pi13 ? n639 : n1280;
  assign n3344 = pi12 ? n26 : n3343;
  assign n3345 = pi11 ? n3344 : n2641;
  assign n3346 = pi10 ? n3345 : n26;
  assign n3347 = pi09 ? n3346 : n26;
  assign n3348 = pi08 ? n3347 : n26;
  assign n3349 = pi07 ? n3342 : n3348;
  assign n3350 = pi06 ? n3349 : n26;
  assign n3351 = pi05 ? n3330 : n3350;
  assign n3352 = pi13 ? n2332 : n2387;
  assign n3353 = pi12 ? n26 : n3352;
  assign n3354 = pi11 ? n2824 : n3353;
  assign n3355 = pi10 ? n2518 : n3354;
  assign n3356 = pi09 ? n26 : n3355;
  assign n3357 = pi08 ? n26 : n3356;
  assign n3358 = pi14 ? n125 : n292;
  assign n3359 = pi13 ? n3358 : n26;
  assign n3360 = pi12 ? n26 : n3359;
  assign n3361 = pi11 ? n3175 : n3360;
  assign n3362 = pi10 ? n3361 : n26;
  assign n3363 = pi09 ? n3362 : n26;
  assign n3364 = pi08 ? n3363 : n26;
  assign n3365 = pi07 ? n3357 : n3364;
  assign n3366 = pi06 ? n3365 : n26;
  assign n3367 = pi13 ? n3023 : n2530;
  assign n3368 = pi12 ? n26 : n3367;
  assign n3369 = pi11 ? n26 : n3368;
  assign n3370 = pi13 ? n478 : n2387;
  assign n3371 = pi12 ? n26 : n3370;
  assign n3372 = pi11 ? n2824 : n3371;
  assign n3373 = pi10 ? n3369 : n3372;
  assign n3374 = pi09 ? n26 : n3373;
  assign n3375 = pi08 ? n26 : n3374;
  assign n3376 = pi13 ? n1135 : n26;
  assign n3377 = pi12 ? n26 : n3376;
  assign n3378 = pi13 ? n630 : n26;
  assign n3379 = pi12 ? n26 : n3378;
  assign n3380 = pi11 ? n3377 : n3379;
  assign n3381 = pi11 ? n3205 : n26;
  assign n3382 = pi10 ? n3380 : n3381;
  assign n3383 = pi12 ? n124 : n2861;
  assign n3384 = pi11 ? n3383 : n2854;
  assign n3385 = pi10 ? n3384 : n2859;
  assign n3386 = pi09 ? n3382 : n3385;
  assign n3387 = pi08 ? n3386 : n2859;
  assign n3388 = pi07 ? n3375 : n3387;
  assign n3389 = pi10 ? n2868 : n2859;
  assign n3390 = pi09 ? n3389 : n2859;
  assign n3391 = pi08 ? n2870 : n3390;
  assign n3392 = pi07 ? n3391 : n2859;
  assign n3393 = pi06 ? n3388 : n3392;
  assign n3394 = pi05 ? n3366 : n3393;
  assign n3395 = pi04 ? n3351 : n3394;
  assign n3396 = pi03 ? n3318 : n3395;
  assign n3397 = pi02 ? n3303 : n3396;
  assign n3398 = pi14 ? n26 : n2954;
  assign n3399 = pi13 ? n478 : n3398;
  assign n3400 = pi12 ? n26 : n3399;
  assign n3401 = pi11 ? n2824 : n3400;
  assign n3402 = pi10 ? n2726 : n3401;
  assign n3403 = pi09 ? n26 : n3402;
  assign n3404 = pi08 ? n26 : n3403;
  assign n3405 = pi14 ? n916 : n26;
  assign n3406 = pi13 ? n3405 : n26;
  assign n3407 = pi12 ? n26 : n3406;
  assign n3408 = pi11 ? n3143 : n3407;
  assign n3409 = pi13 ? n2165 : n26;
  assign n3410 = pi12 ? n26 : n3409;
  assign n3411 = pi13 ? n126 : ~n26;
  assign n3412 = pi12 ? n26 : ~n3411;
  assign n3413 = pi11 ? n3410 : n3412;
  assign n3414 = pi10 ? n3408 : n3413;
  assign n3415 = pi12 ? n124 : n2891;
  assign n3416 = pi11 ? n3415 : n2854;
  assign n3417 = pi10 ? n3416 : n2859;
  assign n3418 = pi09 ? n3414 : n3417;
  assign n3419 = pi08 ? n3418 : n2859;
  assign n3420 = pi07 ? n3404 : n3419;
  assign n3421 = pi06 ? n3420 : n2859;
  assign n3422 = pi13 ? n26 : n2727;
  assign n3423 = pi12 ? n26 : n3422;
  assign n3424 = pi11 ? n26 : n3423;
  assign n3425 = pi10 ? n3424 : n2844;
  assign n3426 = pi09 ? n26 : n3425;
  assign n3427 = pi08 ? n26 : n3426;
  assign n3428 = pi11 ? n2834 : n2641;
  assign n3429 = pi13 ? n1914 : ~n26;
  assign n3430 = pi12 ? n124 : ~n3429;
  assign n3431 = pi11 ? n3412 : n3430;
  assign n3432 = pi10 ? n3428 : n3431;
  assign n3433 = pi12 ? n654 : n2921;
  assign n3434 = pi11 ? n3433 : n2916;
  assign n3435 = pi10 ? n2916 : n3434;
  assign n3436 = pi09 ? n3432 : n3435;
  assign n3437 = pi08 ? n3436 : n2916;
  assign n3438 = pi07 ? n3427 : n3437;
  assign n3439 = pi11 ? n2916 : n2928;
  assign n3440 = pi10 ? n2916 : n3439;
  assign n3441 = pi12 ? n654 : n2888;
  assign n3442 = pi11 ? n2930 : n3441;
  assign n3443 = pi13 ? n77 : ~n507;
  assign n3444 = pi12 ? n26 : n3443;
  assign n3445 = pi11 ? n3444 : n2916;
  assign n3446 = pi10 ? n3442 : n3445;
  assign n3447 = pi09 ? n3440 : n3446;
  assign n3448 = pi08 ? n3447 : n2916;
  assign n3449 = pi07 ? n3448 : n2916;
  assign n3450 = pi06 ? n3438 : n3449;
  assign n3451 = pi05 ? n3421 : n3450;
  assign n3452 = pi13 ? n26 : n2598;
  assign n3453 = pi12 ? n26 : n3452;
  assign n3454 = pi11 ? n26 : n3453;
  assign n3455 = pi14 ? n45 : ~n2058;
  assign n3456 = pi13 ? n26 : n3455;
  assign n3457 = pi12 ? n26 : n3456;
  assign n3458 = pi11 ? n3457 : n2366;
  assign n3459 = pi10 ? n3454 : n3458;
  assign n3460 = pi09 ? n26 : n3459;
  assign n3461 = pi08 ? n26 : n3460;
  assign n3462 = pi11 ? n26 : n2906;
  assign n3463 = pi11 ? n26 : n2911;
  assign n3464 = pi10 ? n3462 : n3463;
  assign n3465 = pi12 ? n654 : n2951;
  assign n3466 = pi11 ? n3465 : n2945;
  assign n3467 = pi10 ? n2947 : n3466;
  assign n3468 = pi09 ? n3464 : n3467;
  assign n3469 = pi08 ? n3468 : n2957;
  assign n3470 = pi07 ? n3461 : n3469;
  assign n3471 = pi13 ? n26 : n2955;
  assign n3472 = pi12 ? n26 : n3471;
  assign n3473 = pi11 ? n3472 : n2963;
  assign n3474 = pi10 ? n2957 : n3473;
  assign n3475 = pi13 ? n507 : n2850;
  assign n3476 = pi12 ? n654 : ~n3475;
  assign n3477 = pi11 ? n3476 : n3002;
  assign n3478 = pi14 ? n2058 : ~n26;
  assign n3479 = pi13 ? n396 : n3478;
  assign n3480 = pi12 ? n26 : ~n3479;
  assign n3481 = pi11 ? n3480 : n2957;
  assign n3482 = pi10 ? n3477 : n3481;
  assign n3483 = pi09 ? n3474 : n3482;
  assign n3484 = pi08 ? n3483 : n2957;
  assign n3485 = pi13 ? n68 : n198;
  assign n3486 = pi12 ? n26 : n3485;
  assign n3487 = pi10 ? n2957 : n3486;
  assign n3488 = pi09 ? n2957 : n3487;
  assign n3489 = pi08 ? n2957 : n3488;
  assign n3490 = pi07 ? n3484 : n3489;
  assign n3491 = pi06 ? n3470 : n3490;
  assign n3492 = pi13 ? n2904 : n2487;
  assign n3493 = pi12 ? n26 : n3492;
  assign n3494 = pi11 ? n2824 : n3493;
  assign n3495 = pi10 ? n26 : n3494;
  assign n3496 = pi14 ? n147 : n168;
  assign n3497 = pi13 ? n2347 : ~n3496;
  assign n3498 = pi12 ? n26 : n3497;
  assign n3499 = pi13 ? n26 : ~n3496;
  assign n3500 = pi12 ? n26 : n3499;
  assign n3501 = pi11 ? n3498 : n3500;
  assign n3502 = pi10 ? n3501 : n26;
  assign n3503 = pi09 ? n3495 : n3502;
  assign n3504 = pi08 ? n3503 : n26;
  assign n3505 = pi07 ? n3504 : n26;
  assign n3506 = pi06 ? n26 : n3505;
  assign n3507 = pi05 ? n3491 : n3506;
  assign n3508 = pi04 ? n3451 : n3507;
  assign n3509 = pi11 ? n2761 : n3002;
  assign n3510 = pi10 ? n26 : n3509;
  assign n3511 = pi10 ? n3038 : n26;
  assign n3512 = pi09 ? n3510 : n3511;
  assign n3513 = pi08 ? n3512 : n26;
  assign n3514 = pi07 ? n3513 : n26;
  assign n3515 = pi06 ? n26 : n3514;
  assign n3516 = pi12 ? n26 : n654;
  assign n3517 = pi13 ? n2519 : n2387;
  assign n3518 = pi12 ? n26 : n3517;
  assign n3519 = pi11 ? n3516 : n3518;
  assign n3520 = pi10 ? n3017 : n3519;
  assign n3521 = pi09 ? n2307 : n3520;
  assign n3522 = pi08 ? n2307 : n3521;
  assign n3523 = pi07 ? n2311 : n3522;
  assign n3524 = pi11 ? n26 : n3025;
  assign n3525 = pi14 ? n71 : n292;
  assign n3526 = pi13 ? n26 : n3525;
  assign n3527 = pi12 ? n26 : n3526;
  assign n3528 = pi11 ? n3527 : n2999;
  assign n3529 = pi10 ? n3524 : n3528;
  assign n3530 = pi13 ? n2319 : n478;
  assign n3531 = pi12 ? n26 : n3530;
  assign n3532 = pi11 ? n3531 : n2641;
  assign n3533 = pi12 ? n654 : n2857;
  assign n3534 = pi13 ? n2698 : n26;
  assign n3535 = pi12 ? n654 : n3534;
  assign n3536 = pi11 ? n3533 : n3535;
  assign n3537 = pi10 ? n3532 : n3536;
  assign n3538 = pi09 ? n3529 : n3537;
  assign n3539 = pi08 ? n3538 : n2859;
  assign n3540 = pi07 ? n3539 : n2859;
  assign n3541 = pi06 ? n3523 : n3540;
  assign n3542 = pi05 ? n3515 : n3541;
  assign n3543 = pi13 ? n321 : n653;
  assign n3544 = pi12 ? n26 : n3543;
  assign n3545 = pi13 ? n3055 : n2387;
  assign n3546 = pi12 ? n26 : n3545;
  assign n3547 = pi11 ? n3544 : n3546;
  assign n3548 = pi10 ? n3052 : n3547;
  assign n3549 = pi09 ? n2612 : n3548;
  assign n3550 = pi08 ? n2612 : n3549;
  assign n3551 = pi07 ? n2311 : n3550;
  assign n3552 = pi13 ? n507 : ~n478;
  assign n3553 = pi12 ? n26 : ~n3552;
  assign n3554 = pi11 ? n2500 : n3553;
  assign n3555 = pi10 ? n3141 : n3554;
  assign n3556 = pi11 ? n2792 : n2641;
  assign n3557 = pi13 ? n2165 : n2519;
  assign n3558 = pi12 ? n78 : n3557;
  assign n3559 = pi11 ? n3558 : n2859;
  assign n3560 = pi10 ? n3556 : n3559;
  assign n3561 = pi09 ? n3555 : n3560;
  assign n3562 = pi08 ? n3561 : n2859;
  assign n3563 = pi07 ? n3562 : n2859;
  assign n3564 = pi06 ? n3551 : n3563;
  assign n3565 = pi12 ? n26 : n68;
  assign n3566 = pi11 ? n3565 : n3310;
  assign n3567 = pi10 ? n26 : n3566;
  assign n3568 = pi09 ? n26 : n3567;
  assign n3569 = pi08 ? n26 : n3568;
  assign n3570 = pi11 ? n3085 : n3126;
  assign n3571 = pi13 ? n143 : n321;
  assign n3572 = pi12 ? n26 : n3571;
  assign n3573 = pi11 ? n2469 : n3572;
  assign n3574 = pi10 ? n3570 : n3573;
  assign n3575 = pi09 ? n2469 : n3574;
  assign n3576 = pi08 ? n2469 : n3575;
  assign n3577 = pi07 ? n3569 : n3576;
  assign n3578 = pi11 ? n2590 : n2617;
  assign n3579 = pi10 ? n3578 : n26;
  assign n3580 = pi11 ? n3207 : n26;
  assign n3581 = pi13 ? n2448 : n2519;
  assign n3582 = pi12 ? n26 : n3581;
  assign n3583 = pi11 ? n3007 : n3582;
  assign n3584 = pi10 ? n3580 : n3583;
  assign n3585 = pi09 ? n3579 : n3584;
  assign n3586 = pi13 ? n77 : ~n2920;
  assign n3587 = pi12 ? n26 : n3586;
  assign n3588 = pi11 ? n2916 : n3587;
  assign n3589 = pi11 ? n3256 : n2916;
  assign n3590 = pi10 ? n3588 : n3589;
  assign n3591 = pi09 ? n3590 : n2916;
  assign n3592 = pi08 ? n3585 : n3591;
  assign n3593 = pi07 ? n3592 : n2916;
  assign n3594 = pi06 ? n3577 : n3593;
  assign n3595 = pi05 ? n3564 : n3594;
  assign n3596 = pi04 ? n3542 : n3595;
  assign n3597 = pi03 ? n3508 : n3596;
  assign n3598 = pi14 ? n327 : n1704;
  assign n3599 = pi13 ? n3598 : n2387;
  assign n3600 = pi12 ? n26 : n3599;
  assign n3601 = pi11 ? n26 : n3600;
  assign n3602 = pi13 ? n2347 : n2387;
  assign n3603 = pi12 ? n26 : n3602;
  assign n3604 = pi13 ? n2347 : n321;
  assign n3605 = pi12 ? n26 : n3604;
  assign n3606 = pi11 ? n3603 : n3605;
  assign n3607 = pi10 ? n3601 : n3606;
  assign n3608 = pi09 ? n26 : n3607;
  assign n3609 = pi08 ? n26 : n3608;
  assign n3610 = pi10 ? n2349 : n3269;
  assign n3611 = pi09 ? n3610 : n3269;
  assign n3612 = pi13 ? n3135 : n26;
  assign n3613 = pi12 ? n26 : n3612;
  assign n3614 = pi11 ? n2612 : n3613;
  assign n3615 = pi10 ? n3614 : n2756;
  assign n3616 = pi09 ? n3269 : n3615;
  assign n3617 = pi08 ? n3611 : n3616;
  assign n3618 = pi07 ? n3609 : n3617;
  assign n3619 = pi11 ? n2366 : n3453;
  assign n3620 = pi10 ? n2591 : n3619;
  assign n3621 = pi13 ? n2642 : ~n26;
  assign n3622 = pi12 ? n26 : ~n3621;
  assign n3623 = pi11 ? n3622 : n2792;
  assign n3624 = pi14 ? n320 : n163;
  assign n3625 = pi13 ? n3624 : n26;
  assign n3626 = pi12 ? n26 : n3625;
  assign n3627 = pi11 ? n2641 : n3626;
  assign n3628 = pi10 ? n3623 : n3627;
  assign n3629 = pi09 ? n3620 : n3628;
  assign n3630 = pi11 ? n2945 : n2957;
  assign n3631 = pi10 ? n2947 : n3630;
  assign n3632 = pi09 ? n3631 : n2957;
  assign n3633 = pi08 ? n3629 : n3632;
  assign n3634 = pi07 ? n3633 : n3489;
  assign n3635 = pi06 ? n3618 : n3634;
  assign n3636 = pi14 ? n320 : n37;
  assign n3637 = pi13 ? n3636 : n2387;
  assign n3638 = pi12 ? n26 : n3637;
  assign n3639 = pi11 ? n26 : n3638;
  assign n3640 = pi13 ? n639 : n2519;
  assign n3641 = pi12 ? n26 : n3640;
  assign n3642 = pi11 ? n3641 : n2641;
  assign n3643 = pi10 ? n3639 : n3642;
  assign n3644 = pi09 ? n26 : n3643;
  assign n3645 = pi08 ? n26 : n3644;
  assign n3646 = pi07 ? n3645 : n3348;
  assign n3647 = pi06 ? n3646 : n26;
  assign n3648 = pi05 ? n3635 : n3647;
  assign n3649 = pi13 ? n74 : n2487;
  assign n3650 = pi12 ? n26 : n3649;
  assign n3651 = pi11 ? n3650 : n3353;
  assign n3652 = pi10 ? n2518 : n3651;
  assign n3653 = pi09 ? n26 : n3652;
  assign n3654 = pi08 ? n26 : n3653;
  assign n3655 = pi13 ? n1705 : n2387;
  assign n3656 = pi12 ? n26 : n3655;
  assign n3657 = pi14 ? n1138 : n292;
  assign n3658 = pi13 ? n3657 : n26;
  assign n3659 = pi12 ? n26 : n3658;
  assign n3660 = pi11 ? n3656 : n3659;
  assign n3661 = pi10 ? n3660 : n26;
  assign n3662 = pi09 ? n3661 : n26;
  assign n3663 = pi08 ? n3662 : n26;
  assign n3664 = pi07 ? n3654 : n3663;
  assign n3665 = pi06 ? n3664 : n26;
  assign n3666 = pi11 ? n2824 : n2704;
  assign n3667 = pi10 ? n3369 : n3666;
  assign n3668 = pi09 ? n26 : n3667;
  assign n3669 = pi08 ? n26 : n3668;
  assign n3670 = pi11 ? n2739 : n3379;
  assign n3671 = pi10 ? n3670 : n3381;
  assign n3672 = pi11 ? n2835 : n26;
  assign n3673 = pi10 ? n3672 : n2511;
  assign n3674 = pi09 ? n3671 : n3673;
  assign n3675 = pi08 ? n3674 : n2511;
  assign n3676 = pi07 ? n3669 : n3675;
  assign n3677 = pi06 ? n3676 : n2511;
  assign n3678 = pi05 ? n3665 : n3677;
  assign n3679 = pi04 ? n3648 : n3678;
  assign n3680 = pi13 ? n26 : n3398;
  assign n3681 = pi12 ? n26 : n3680;
  assign n3682 = pi11 ? n2824 : n3681;
  assign n3683 = pi10 ? n2726 : n3682;
  assign n3684 = pi09 ? n26 : n3683;
  assign n3685 = pi08 ? n26 : n3684;
  assign n3686 = pi13 ? n2254 : n26;
  assign n3687 = pi12 ? n26 : n3686;
  assign n3688 = pi12 ? n124 : ~n3411;
  assign n3689 = pi11 ? n3687 : n3688;
  assign n3690 = pi10 ? n3380 : n3689;
  assign n3691 = pi11 ? n2854 : n2859;
  assign n3692 = pi10 ? n3691 : n2859;
  assign n3693 = pi09 ? n3690 : n3692;
  assign n3694 = pi08 ? n3693 : n2859;
  assign n3695 = pi07 ? n3685 : n3694;
  assign n3696 = pi06 ? n3695 : n2859;
  assign n3697 = pi13 ? n57 : ~n26;
  assign n3698 = pi12 ? n26 : ~n3697;
  assign n3699 = pi11 ? n3379 : n3698;
  assign n3700 = pi12 ? n69 : n2857;
  assign n3701 = pi11 ? n2835 : n3700;
  assign n3702 = pi10 ? n3699 : n3701;
  assign n3703 = pi12 ? n1203 : n2891;
  assign n3704 = pi11 ? n3703 : n2892;
  assign n3705 = pi12 ? n654 : n2962;
  assign n3706 = pi11 ? n3705 : n2868;
  assign n3707 = pi10 ? n3704 : n3706;
  assign n3708 = pi09 ? n3702 : n3707;
  assign n3709 = pi08 ? n3708 : n2868;
  assign n3710 = pi07 ? n3427 : n3709;
  assign n3711 = pi06 ? n3710 : n2868;
  assign n3712 = pi05 ? n3696 : n3711;
  assign n3713 = pi13 ? n62 : n1280;
  assign n3714 = pi12 ? n26 : n3713;
  assign n3715 = pi11 ? n3457 : n3714;
  assign n3716 = pi10 ? n3424 : n3715;
  assign n3717 = pi09 ? n26 : n3716;
  assign n3718 = pi08 ? n26 : n3717;
  assign n3719 = pi15 ? n44 : ~n1200;
  assign n3720 = pi14 ? n3719 : ~n26;
  assign n3721 = pi13 ? n3720 : ~n26;
  assign n3722 = pi12 ? n26 : ~n3721;
  assign n3723 = pi11 ? n2834 : n3722;
  assign n3724 = pi13 ? n396 : ~n26;
  assign n3725 = pi12 ? n69 : ~n3724;
  assign n3726 = pi11 ? n2835 : n3725;
  assign n3727 = pi10 ? n3723 : n3726;
  assign n3728 = pi12 ? n654 : ~n3724;
  assign n3729 = pi11 ? n3441 : n3728;
  assign n3730 = pi11 ? n2986 : n2911;
  assign n3731 = pi10 ? n3729 : n3730;
  assign n3732 = pi09 ? n3727 : n3731;
  assign n3733 = pi08 ? n3732 : n2963;
  assign n3734 = pi07 ? n3718 : n3733;
  assign n3735 = pi06 ? n3734 : n2963;
  assign n3736 = pi14 ? n45 : n63;
  assign n3737 = pi13 ? n26 : n3736;
  assign n3738 = pi12 ? n26 : n3737;
  assign n3739 = pi11 ? n3738 : n2537;
  assign n3740 = pi10 ? n2938 : n3739;
  assign n3741 = pi09 ? n26 : n3740;
  assign n3742 = pi08 ? n26 : n3741;
  assign n3743 = pi10 ? n3462 : n3208;
  assign n3744 = pi11 ? n3441 : n2911;
  assign n3745 = pi10 ? n3744 : n2945;
  assign n3746 = pi09 ? n3743 : n3745;
  assign n3747 = pi13 ? n26 : n2950;
  assign n3748 = pi12 ? n26 : n3747;
  assign n3749 = pi08 ? n3746 : n3748;
  assign n3750 = pi07 ? n3742 : n3749;
  assign n3751 = pi13 ? n26 : n2519;
  assign n3752 = pi12 ? n26 : n3751;
  assign n3753 = pi10 ? n3748 : n3752;
  assign n3754 = pi09 ? n3748 : n3753;
  assign n3755 = pi08 ? n3748 : n3754;
  assign n3756 = pi07 ? n3748 : n3755;
  assign n3757 = pi06 ? n3750 : n3756;
  assign n3758 = pi05 ? n3735 : n3757;
  assign n3759 = pi04 ? n3712 : n3758;
  assign n3760 = pi03 ? n3679 : n3759;
  assign n3761 = pi02 ? n3597 : n3760;
  assign n3762 = pi01 ? n3397 : n3761;
  assign n3763 = pi00 ? n3120 : n3762;
  assign n3764 = pi13 ? n169 : n57;
  assign n3765 = pi12 ? n26 : n3764;
  assign n3766 = pi11 ? n26 : n3765;
  assign n3767 = pi13 ? n169 : ~n2370;
  assign n3768 = pi12 ? n26 : n3767;
  assign n3769 = pi10 ? n3766 : n3768;
  assign n3770 = pi09 ? n26 : n3769;
  assign n3771 = pi08 ? n26 : n3770;
  assign n3772 = pi13 ? n130 : ~n2370;
  assign n3773 = pi12 ? n26 : n3772;
  assign n3774 = pi11 ? n3768 : n3773;
  assign n3775 = pi13 ? n176 : ~n2370;
  assign n3776 = pi12 ? n26 : n3775;
  assign n3777 = pi11 ? n3773 : n3776;
  assign n3778 = pi10 ? n3774 : n3777;
  assign n3779 = pi13 ? n143 : ~n2319;
  assign n3780 = pi12 ? n26 : n3779;
  assign n3781 = pi11 ? n3776 : n3780;
  assign n3782 = pi14 ? n37 : ~n37;
  assign n3783 = pi13 ? n143 : ~n3782;
  assign n3784 = pi12 ? n26 : n3783;
  assign n3785 = pi13 ? n77 : ~n3782;
  assign n3786 = pi12 ? n26 : n3785;
  assign n3787 = pi11 ? n3784 : n3786;
  assign n3788 = pi10 ? n3781 : n3787;
  assign n3789 = pi09 ? n3778 : n3788;
  assign n3790 = pi13 ? n26 : n630;
  assign n3791 = pi12 ? n26 : n3790;
  assign n3792 = pi11 ? n1415 : n3791;
  assign n3793 = pi10 ? n3792 : n26;
  assign n3794 = pi13 ? n130 : n57;
  assign n3795 = pi12 ? n26 : n3794;
  assign n3796 = pi11 ? n26 : n3795;
  assign n3797 = pi10 ? n3796 : n3777;
  assign n3798 = pi09 ? n3793 : n3797;
  assign n3799 = pi08 ? n3789 : n3798;
  assign n3800 = pi07 ? n3771 : n3799;
  assign n3801 = pi09 ? n3788 : n3793;
  assign n3802 = pi09 ? n3797 : n3788;
  assign n3803 = pi08 ? n3801 : n3802;
  assign n3804 = pi14 ? n26 : n916;
  assign n3805 = pi13 ? n3804 : n143;
  assign n3806 = pi12 ? n26 : n3805;
  assign n3807 = pi11 ? n26 : n3806;
  assign n3808 = pi13 ? n3804 : ~n1091;
  assign n3809 = pi12 ? n26 : n3808;
  assign n3810 = pi15 ? n60 : ~n28;
  assign n3811 = pi14 ? n26 : n3810;
  assign n3812 = pi13 ? n3811 : ~n1091;
  assign n3813 = pi12 ? n26 : n3812;
  assign n3814 = pi11 ? n3809 : n3813;
  assign n3815 = pi10 ? n3807 : n3814;
  assign n3816 = pi09 ? n3793 : n3815;
  assign n3817 = pi13 ? n3804 : ~n3782;
  assign n3818 = pi12 ? n26 : n3817;
  assign n3819 = pi11 ? n3818 : n3784;
  assign n3820 = pi10 ? n3818 : n3819;
  assign n3821 = pi13 ? n77 : ~n1583;
  assign n3822 = pi12 ? n26 : n3821;
  assign n3823 = pi14 ? n61 : n71;
  assign n3824 = pi14 ? n292 : ~n320;
  assign n3825 = pi13 ? n3823 : ~n3824;
  assign n3826 = pi12 ? n26 : n3825;
  assign n3827 = pi11 ? n3822 : n3826;
  assign n3828 = pi14 ? n71 : ~n517;
  assign n3829 = pi14 ? n292 : ~n26;
  assign n3830 = pi13 ? n3828 : n3829;
  assign n3831 = pi12 ? n2243 : ~n3830;
  assign n3832 = pi13 ? n79 : n2225;
  assign n3833 = pi12 ? n26 : ~n3832;
  assign n3834 = pi11 ? n3831 : n3833;
  assign n3835 = pi10 ? n3827 : n3834;
  assign n3836 = pi09 ? n3820 : n3835;
  assign n3837 = pi08 ? n3816 : n3836;
  assign n3838 = pi07 ? n3803 : n3837;
  assign n3839 = pi06 ? n3800 : n3838;
  assign n3840 = pi05 ? n26 : n3839;
  assign n3841 = pi12 ? n26 : n57;
  assign n3842 = pi11 ? n26 : n3841;
  assign n3843 = pi13 ? n57 : n79;
  assign n3844 = pi12 ? n26 : n3843;
  assign n3845 = pi13 ? n169 : n79;
  assign n3846 = pi12 ? n26 : n3845;
  assign n3847 = pi11 ? n3844 : n3846;
  assign n3848 = pi10 ? n3842 : n3847;
  assign n3849 = pi09 ? n26 : n3848;
  assign n3850 = pi08 ? n26 : n3849;
  assign n3851 = pi14 ? n26 : n152;
  assign n3852 = pi13 ? n3851 : n79;
  assign n3853 = pi12 ? n26 : n3852;
  assign n3854 = pi13 ? n149 : n79;
  assign n3855 = pi12 ? n26 : n3854;
  assign n3856 = pi11 ? n3853 : n3855;
  assign n3857 = pi13 ? n149 : n57;
  assign n3858 = pi12 ? n26 : n3857;
  assign n3859 = pi13 ? n132 : n64;
  assign n3860 = pi12 ? n26 : n3859;
  assign n3861 = pi11 ? n3858 : n3860;
  assign n3862 = pi10 ? n3856 : n3861;
  assign n3863 = pi13 ? n321 : n64;
  assign n3864 = pi12 ? n26 : n3863;
  assign n3865 = pi11 ? n3860 : n3864;
  assign n3866 = pi13 ? n77 : n143;
  assign n3867 = pi12 ? n26 : n3866;
  assign n3868 = pi11 ? n3864 : n3867;
  assign n3869 = pi10 ? n3865 : n3868;
  assign n3870 = pi09 ? n3862 : n3869;
  assign n3871 = pi13 ? n68 : ~n79;
  assign n3872 = pi12 ? n26 : n3871;
  assign n3873 = pi14 ? n168 : ~n29;
  assign n3874 = pi13 ? n26 : n3873;
  assign n3875 = pi12 ? n26 : n3874;
  assign n3876 = pi11 ? n3872 : n3875;
  assign n3877 = pi10 ? n3876 : n26;
  assign n3878 = pi10 ? n3796 : n3861;
  assign n3879 = pi09 ? n3877 : n3878;
  assign n3880 = pi08 ? n3870 : n3879;
  assign n3881 = pi07 ? n3850 : n3880;
  assign n3882 = pi09 ? n3869 : n3877;
  assign n3883 = pi09 ? n3878 : n3869;
  assign n3884 = pi08 ? n3882 : n3883;
  assign n3885 = pi13 ? n57 : n143;
  assign n3886 = pi12 ? n26 : n3885;
  assign n3887 = pi11 ? n26 : n3886;
  assign n3888 = pi14 ? n29 : ~n125;
  assign n3889 = pi13 ? n57 : ~n3888;
  assign n3890 = pi12 ? n26 : n3889;
  assign n3891 = pi10 ? n3887 : n3890;
  assign n3892 = pi09 ? n3877 : n3891;
  assign n3893 = pi13 ? n169 : ~n3782;
  assign n3894 = pi12 ? n26 : n3893;
  assign n3895 = pi13 ? n143 : ~n1091;
  assign n3896 = pi12 ? n26 : n3895;
  assign n3897 = pi11 ? n3894 : n3896;
  assign n3898 = pi10 ? n3890 : n3897;
  assign n3899 = pi14 ? n432 : ~n71;
  assign n3900 = pi13 ? n143 : ~n3899;
  assign n3901 = pi12 ? n26 : n3900;
  assign n3902 = pi14 ? n73 : ~n45;
  assign n3903 = pi13 ? n1942 : n3902;
  assign n3904 = pi12 ? n124 : ~n3903;
  assign n3905 = pi11 ? n3901 : n3904;
  assign n3906 = pi15 ? n1200 : ~n26;
  assign n3907 = pi14 ? n3906 : ~n29;
  assign n3908 = pi13 ? n130 : ~n3907;
  assign n3909 = pi12 ? n26 : ~n3908;
  assign n3910 = pi13 ? n130 : n3251;
  assign n3911 = pi12 ? n26 : ~n3910;
  assign n3912 = pi11 ? n3909 : n3911;
  assign n3913 = pi10 ? n3905 : n3912;
  assign n3914 = pi09 ? n3898 : n3913;
  assign n3915 = pi08 ? n3892 : n3914;
  assign n3916 = pi07 ? n3884 : n3915;
  assign n3917 = pi06 ? n3881 : n3916;
  assign n3918 = pi14 ? n45 : ~n37;
  assign n3919 = pi13 ? n1583 : n3918;
  assign n3920 = pi12 ? n26 : n3919;
  assign n3921 = pi11 ? n26 : n3920;
  assign n3922 = pi14 ? n45 : ~n147;
  assign n3923 = pi13 ? n149 : n3922;
  assign n3924 = pi12 ? n26 : n3923;
  assign n3925 = pi13 ? n3851 : n3922;
  assign n3926 = pi12 ? n26 : n3925;
  assign n3927 = pi11 ? n3924 : n3926;
  assign n3928 = pi10 ? n3921 : n3927;
  assign n3929 = pi09 ? n26 : n3928;
  assign n3930 = pi08 ? n26 : n3929;
  assign n3931 = pi13 ? n26 : n2391;
  assign n3932 = pi12 ? n26 : n3931;
  assign n3933 = pi10 ? n3924 : n3932;
  assign n3934 = pi12 ? n26 : n143;
  assign n3935 = pi11 ? n48 : n3934;
  assign n3936 = pi10 ? n3932 : n3935;
  assign n3937 = pi09 ? n3933 : n3936;
  assign n3938 = pi13 ? n77 : ~n105;
  assign n3939 = pi12 ? n26 : n3938;
  assign n3940 = pi11 ? n3939 : n3875;
  assign n3941 = pi10 ? n3940 : n26;
  assign n3942 = pi14 ? n26 : n1832;
  assign n3943 = pi13 ? n3942 : n3918;
  assign n3944 = pi12 ? n26 : n3943;
  assign n3945 = pi11 ? n26 : n3944;
  assign n3946 = pi10 ? n3945 : n3932;
  assign n3947 = pi09 ? n3941 : n3946;
  assign n3948 = pi08 ? n3937 : n3947;
  assign n3949 = pi07 ? n3930 : n3948;
  assign n3950 = pi09 ? n3936 : n3941;
  assign n3951 = pi09 ? n3946 : n3936;
  assign n3952 = pi08 ? n3950 : n3951;
  assign n3953 = pi13 ? n240 : n130;
  assign n3954 = pi12 ? n26 : n3953;
  assign n3955 = pi11 ? n26 : n3954;
  assign n3956 = pi13 ? n240 : ~n3888;
  assign n3957 = pi12 ? n26 : n3956;
  assign n3958 = pi13 ? n240 : ~n3066;
  assign n3959 = pi12 ? n26 : n3958;
  assign n3960 = pi11 ? n3957 : n3959;
  assign n3961 = pi10 ? n3955 : n3960;
  assign n3962 = pi09 ? n3941 : n3961;
  assign n3963 = pi13 ? n57 : ~n3066;
  assign n3964 = pi12 ? n26 : n3963;
  assign n3965 = pi14 ? n517 : n125;
  assign n3966 = pi13 ? n3965 : ~n3066;
  assign n3967 = pi12 ? n26 : n3966;
  assign n3968 = pi11 ? n3964 : n3967;
  assign n3969 = pi14 ? n37 : ~n249;
  assign n3970 = pi13 ? n3804 : ~n3969;
  assign n3971 = pi12 ? n26 : n3970;
  assign n3972 = pi11 ? n3964 : n3971;
  assign n3973 = pi10 ? n3968 : n3972;
  assign n3974 = pi14 ? n45 : ~n249;
  assign n3975 = pi13 ? n143 : ~n3974;
  assign n3976 = pi12 ? n26 : n3975;
  assign n3977 = pi13 ? n1252 : n46;
  assign n3978 = pi12 ? n69 : ~n3977;
  assign n3979 = pi11 ? n3976 : n3978;
  assign n3980 = pi14 ? n125 : ~n125;
  assign n3981 = pi13 ? n3980 : ~n57;
  assign n3982 = pi12 ? n26 : n3981;
  assign n3983 = pi14 ? n916 : ~n29;
  assign n3984 = pi13 ? n1939 : n3983;
  assign n3985 = pi12 ? n654 : n3984;
  assign n3986 = pi11 ? n3982 : n3985;
  assign n3987 = pi10 ? n3979 : n3986;
  assign n3988 = pi09 ? n3973 : n3987;
  assign n3989 = pi08 ? n3962 : n3988;
  assign n3990 = pi07 ? n3952 : n3989;
  assign n3991 = pi06 ? n3949 : n3990;
  assign n3992 = pi05 ? n3917 : n3991;
  assign n3993 = pi04 ? n3840 : n3992;
  assign n3994 = pi03 ? n26 : n3993;
  assign n3995 = pi02 ? n26 : n3994;
  assign n3996 = pi14 ? n63 : ~n37;
  assign n3997 = pi13 ? n3996 : n3782;
  assign n3998 = pi12 ? n26 : n3997;
  assign n3999 = pi11 ? n26 : n3998;
  assign n4000 = pi13 ? n1583 : n2979;
  assign n4001 = pi12 ? n26 : n4000;
  assign n4002 = pi13 ? n1583 : n2319;
  assign n4003 = pi12 ? n26 : n4002;
  assign n4004 = pi11 ? n4001 : n4003;
  assign n4005 = pi10 ? n3999 : n4004;
  assign n4006 = pi09 ? n26 : n4005;
  assign n4007 = pi08 ? n26 : n4006;
  assign n4008 = pi13 ? n3023 : n1135;
  assign n4009 = pi12 ? n26 : n4008;
  assign n4010 = pi13 ? n26 : n1135;
  assign n4011 = pi12 ? n26 : n4010;
  assign n4012 = pi11 ? n4009 : n4011;
  assign n4013 = pi13 ? n26 : ~n240;
  assign n4014 = pi12 ? n26 : n4013;
  assign n4015 = pi13 ? n26 : ~n79;
  assign n4016 = pi12 ? n26 : n4015;
  assign n4017 = pi11 ? n4014 : n4016;
  assign n4018 = pi10 ? n4012 : n4017;
  assign n4019 = pi11 ? n26 : n3934;
  assign n4020 = pi10 ? n26 : n4019;
  assign n4021 = pi09 ? n4018 : n4020;
  assign n4022 = pi13 ? n143 : ~n3918;
  assign n4023 = pi12 ? n26 : n4022;
  assign n4024 = pi11 ? n4023 : n3875;
  assign n4025 = pi10 ? n4024 : n26;
  assign n4026 = pi13 ? n3942 : n3782;
  assign n4027 = pi12 ? n26 : n4026;
  assign n4028 = pi11 ? n26 : n4027;
  assign n4029 = pi10 ? n4028 : n4017;
  assign n4030 = pi09 ? n4025 : n4029;
  assign n4031 = pi08 ? n4021 : n4030;
  assign n4032 = pi07 ? n4007 : n4031;
  assign n4033 = pi09 ? n4020 : n4025;
  assign n4034 = pi09 ? n4029 : n4020;
  assign n4035 = pi08 ? n4033 : n4034;
  assign n4036 = pi13 ? n79 : n46;
  assign n4037 = pi12 ? n26 : n4036;
  assign n4038 = pi11 ? n26 : n4037;
  assign n4039 = pi10 ? n4038 : n4037;
  assign n4040 = pi09 ? n4025 : n4039;
  assign n4041 = pi13 ? n1464 : n46;
  assign n4042 = pi12 ? n26 : n4041;
  assign n4043 = pi11 ? n4037 : n4042;
  assign n4044 = pi13 ? n169 : n46;
  assign n4045 = pi12 ? n26 : n4044;
  assign n4046 = pi11 ? n3841 : n4045;
  assign n4047 = pi10 ? n4043 : n4046;
  assign n4048 = pi13 ? n130 : n46;
  assign n4049 = pi12 ? n26 : n4048;
  assign n4050 = pi12 ? n26 : n3918;
  assign n4051 = pi14 ? n45 : ~n71;
  assign n4052 = pi13 ? n4051 : n3918;
  assign n4053 = pi12 ? n26 : n4052;
  assign n4054 = pi11 ? n4050 : n4053;
  assign n4055 = pi10 ? n4049 : n4054;
  assign n4056 = pi09 ? n4047 : n4055;
  assign n4057 = pi08 ? n4040 : n4056;
  assign n4058 = pi07 ? n4035 : n4057;
  assign n4059 = pi06 ? n4032 : n4058;
  assign n4060 = pi11 ? n26 : n4050;
  assign n4061 = pi13 ? n3918 : n2319;
  assign n4062 = pi12 ? n26 : n4061;
  assign n4063 = pi11 ? n4062 : n4003;
  assign n4064 = pi10 ? n4060 : n4063;
  assign n4065 = pi09 ? n26 : n4064;
  assign n4066 = pi08 ? n26 : n4065;
  assign n4067 = pi13 ? n2498 : ~n240;
  assign n4068 = pi12 ? n26 : n4067;
  assign n4069 = pi11 ? n4068 : n4016;
  assign n4070 = pi14 ? n71 : ~n61;
  assign n4071 = pi13 ? n26 : ~n4070;
  assign n4072 = pi12 ? n26 : n4071;
  assign n4073 = pi15 ? n60 : n291;
  assign n4074 = pi14 ? n125 : ~n4073;
  assign n4075 = pi13 ? n68 : ~n4074;
  assign n4076 = pi12 ? n26 : n4075;
  assign n4077 = pi11 ? n4072 : n4076;
  assign n4078 = pi10 ? n4069 : n4077;
  assign n4079 = pi13 ? n169 : n406;
  assign n4080 = pi12 ? n26 : n4079;
  assign n4081 = pi11 ? n26 : n4080;
  assign n4082 = pi10 ? n26 : n4081;
  assign n4083 = pi09 ? n4078 : n4082;
  assign n4084 = pi13 ? n143 : ~n3996;
  assign n4085 = pi12 ? n26 : n4084;
  assign n4086 = pi11 ? n4023 : n4085;
  assign n4087 = pi10 ? n4086 : n26;
  assign n4088 = pi13 ? n3942 : ~n143;
  assign n4089 = pi12 ? n26 : n4088;
  assign n4090 = pi11 ? n26 : n4089;
  assign n4091 = pi14 ? n125 : ~n517;
  assign n4092 = pi13 ? n68 : ~n4091;
  assign n4093 = pi12 ? n26 : n4092;
  assign n4094 = pi11 ? n4014 : n4093;
  assign n4095 = pi10 ? n4090 : n4094;
  assign n4096 = pi09 ? n4087 : n4095;
  assign n4097 = pi08 ? n4083 : n4096;
  assign n4098 = pi07 ? n4066 : n4097;
  assign n4099 = pi09 ? n4082 : n4087;
  assign n4100 = pi09 ? n4095 : n4082;
  assign n4101 = pi08 ? n4099 : n4100;
  assign n4102 = pi14 ? n71 : ~n320;
  assign n4103 = pi13 ? n4102 : n3918;
  assign n4104 = pi12 ? n26 : n4103;
  assign n4105 = pi11 ? n26 : n4104;
  assign n4106 = pi14 ? n71 : ~n45;
  assign n4107 = pi13 ? n4106 : n3918;
  assign n4108 = pi12 ? n26 : n4107;
  assign n4109 = pi13 ? n1344 : n3918;
  assign n4110 = pi12 ? n26 : n4109;
  assign n4111 = pi11 ? n4108 : n4110;
  assign n4112 = pi10 ? n4105 : n4111;
  assign n4113 = pi09 ? n4087 : n4112;
  assign n4114 = pi13 ? n1252 : n3918;
  assign n4115 = pi12 ? n26 : n4114;
  assign n4116 = pi11 ? n4108 : n4115;
  assign n4117 = pi10 ? n4116 : n4115;
  assign n4118 = pi12 ? n26 : n1344;
  assign n4119 = pi14 ? n45 : ~n44;
  assign n4120 = pi13 ? n1344 : n4119;
  assign n4121 = pi12 ? n26 : n4120;
  assign n4122 = pi11 ? n4118 : n4121;
  assign n4123 = pi13 ? n3023 : n1583;
  assign n4124 = pi12 ? n69 : n4123;
  assign n4125 = pi14 ? n26 : n1355;
  assign n4126 = pi13 ? n4125 : n1583;
  assign n4127 = pi12 ? n78 : n4126;
  assign n4128 = pi11 ? n4124 : n4127;
  assign n4129 = pi10 ? n4122 : n4128;
  assign n4130 = pi09 ? n4117 : n4129;
  assign n4131 = pi08 ? n4113 : n4130;
  assign n4132 = pi07 ? n4101 : n4131;
  assign n4133 = pi06 ? n4098 : n4132;
  assign n4134 = pi05 ? n4059 : n4133;
  assign n4135 = pi14 ? n71 : ~n37;
  assign n4136 = pi13 ? n4135 : n3918;
  assign n4137 = pi12 ? n26 : n4136;
  assign n4138 = pi11 ? n26 : n4137;
  assign n4139 = pi14 ? n71 : n233;
  assign n4140 = pi15 ? n44 : ~n60;
  assign n4141 = pi14 ? n26 : n4140;
  assign n4142 = pi13 ? n4139 : ~n4141;
  assign n4143 = pi12 ? n26 : n4142;
  assign n4144 = pi11 ? n4143 : n4014;
  assign n4145 = pi10 ? n4138 : n4144;
  assign n4146 = pi09 ? n26 : n4145;
  assign n4147 = pi08 ? n26 : n4146;
  assign n4148 = pi13 ? n26 : ~n72;
  assign n4149 = pi12 ? n26 : n4148;
  assign n4150 = pi11 ? n4016 : n4149;
  assign n4151 = pi13 ? n2762 : ~n38;
  assign n4152 = pi12 ? n26 : n4151;
  assign n4153 = pi14 ? n125 : ~n61;
  assign n4154 = pi13 ? n2165 : ~n4153;
  assign n4155 = pi12 ? n26 : n4154;
  assign n4156 = pi11 ? n4152 : n4155;
  assign n4157 = pi10 ? n4150 : n4156;
  assign n4158 = pi13 ? n57 : n46;
  assign n4159 = pi12 ? n26 : n4158;
  assign n4160 = pi11 ? n26 : n4159;
  assign n4161 = pi10 ? n26 : n4160;
  assign n4162 = pi09 ? n4157 : n4161;
  assign n4163 = pi13 ? n57 : ~n2370;
  assign n4164 = pi12 ? n26 : n4163;
  assign n4165 = pi13 ? n64 : n38;
  assign n4166 = pi12 ? n26 : n4165;
  assign n4167 = pi14 ? n26 : ~n29;
  assign n4168 = pi13 ? n4167 : ~n143;
  assign n4169 = pi12 ? n26 : n4168;
  assign n4170 = pi11 ? n4166 : n4169;
  assign n4171 = pi13 ? n26 : ~n1429;
  assign n4172 = pi12 ? n26 : n4171;
  assign n4173 = pi14 ? n125 : ~n320;
  assign n4174 = pi13 ? n68 : ~n4173;
  assign n4175 = pi12 ? n26 : n4174;
  assign n4176 = pi11 ? n4172 : n4175;
  assign n4177 = pi10 ? n4170 : n4176;
  assign n4178 = pi09 ? n4164 : n4177;
  assign n4179 = pi08 ? n4162 : n4178;
  assign n4180 = pi07 ? n4147 : n4179;
  assign n4181 = pi09 ? n4161 : n4164;
  assign n4182 = pi09 ? n4177 : n4161;
  assign n4183 = pi08 ? n4181 : n4182;
  assign n4184 = pi11 ? n4164 : n3768;
  assign n4185 = pi10 ? n4184 : n3768;
  assign n4186 = pi14 ? n327 : ~n63;
  assign n4187 = pi13 ? n4186 : n79;
  assign n4188 = pi12 ? n26 : n4187;
  assign n4189 = pi14 ? n320 : ~n45;
  assign n4190 = pi13 ? n4189 : n4135;
  assign n4191 = pi12 ? n26 : n4190;
  assign n4192 = pi11 ? n4188 : n4191;
  assign n4193 = pi13 ? n3782 : n2979;
  assign n4194 = pi12 ? n26 : n4193;
  assign n4195 = pi13 ? n3782 : n2319;
  assign n4196 = pi12 ? n26 : n4195;
  assign n4197 = pi11 ? n4194 : n4196;
  assign n4198 = pi10 ? n4192 : n4197;
  assign n4199 = pi09 ? n4185 : n4198;
  assign n4200 = pi13 ? n3061 : n2319;
  assign n4201 = pi12 ? n26 : n4200;
  assign n4202 = pi13 ? n4135 : n2319;
  assign n4203 = pi12 ? n26 : n4202;
  assign n4204 = pi10 ? n4201 : n4203;
  assign n4205 = pi14 ? n916 : ~n37;
  assign n4206 = pi13 ? n4205 : n1135;
  assign n4207 = pi12 ? n26 : n4206;
  assign n4208 = pi13 ? n591 : ~n57;
  assign n4209 = pi12 ? n26 : n4208;
  assign n4210 = pi11 ? n4207 : n4209;
  assign n4211 = pi13 ? n1252 : n3828;
  assign n4212 = pi12 ? n78 : ~n4211;
  assign n4213 = pi14 ? n168 : ~n147;
  assign n4214 = pi13 ? n4213 : ~n2539;
  assign n4215 = pi12 ? n78 : ~n4214;
  assign n4216 = pi11 ? n4212 : n4215;
  assign n4217 = pi10 ? n4210 : n4216;
  assign n4218 = pi09 ? n4204 : n4217;
  assign n4219 = pi08 ? n4199 : n4218;
  assign n4220 = pi07 ? n4183 : n4219;
  assign n4221 = pi06 ? n4180 : n4220;
  assign n4222 = pi14 ? n37 : ~n29;
  assign n4223 = pi13 ? n4222 : ~n340;
  assign n4224 = pi12 ? n26 : n4223;
  assign n4225 = pi11 ? n26 : n4224;
  assign n4226 = pi14 ? n37 : n292;
  assign n4227 = pi13 ? n4226 : ~n1429;
  assign n4228 = pi12 ? n26 : n4227;
  assign n4229 = pi14 ? n45 : ~n327;
  assign n4230 = pi13 ? n2319 : ~n4229;
  assign n4231 = pi12 ? n26 : n4230;
  assign n4232 = pi11 ? n4228 : n4231;
  assign n4233 = pi10 ? n4225 : n4232;
  assign n4234 = pi09 ? n26 : n4233;
  assign n4235 = pi08 ? n26 : n4234;
  assign n4236 = pi13 ? n1280 : ~n72;
  assign n4237 = pi12 ? n26 : n4236;
  assign n4238 = pi13 ? n26 : ~n38;
  assign n4239 = pi12 ? n26 : n4238;
  assign n4240 = pi11 ? n4237 : n4239;
  assign n4241 = pi13 ? n2312 : ~n38;
  assign n4242 = pi12 ? n26 : n4241;
  assign n4243 = pi15 ? n28 : n291;
  assign n4244 = pi14 ? n4243 : n45;
  assign n4245 = pi13 ? n4244 : ~n126;
  assign n4246 = pi12 ? n26 : n4245;
  assign n4247 = pi11 ? n4242 : n4246;
  assign n4248 = pi10 ? n4240 : n4247;
  assign n4249 = pi14 ? n63 : ~n29;
  assign n4250 = pi13 ? n4249 : n3100;
  assign n4251 = pi12 ? n26 : n4250;
  assign n4252 = pi11 ? n26 : n4251;
  assign n4253 = pi10 ? n26 : n4252;
  assign n4254 = pi09 ? n4248 : n4253;
  assign n4255 = pi14 ? n63 : ~n432;
  assign n4256 = pi13 ? n4255 : n3100;
  assign n4257 = pi12 ? n26 : n4256;
  assign n4258 = pi13 ? n1347 : n64;
  assign n4259 = pi12 ? n26 : n4258;
  assign n4260 = pi11 ? n4257 : n4259;
  assign n4261 = pi14 ? n1638 : ~n63;
  assign n4262 = pi13 ? n1347 : n4261;
  assign n4263 = pi12 ? n26 : n4262;
  assign n4264 = pi13 ? n1347 : n202;
  assign n4265 = pi12 ? n26 : n4264;
  assign n4266 = pi11 ? n4263 : n4265;
  assign n4267 = pi10 ? n4260 : n4266;
  assign n4268 = pi11 ? n4265 : n4169;
  assign n4269 = pi13 ? n68 : ~n443;
  assign n4270 = pi12 ? n26 : n4269;
  assign n4271 = pi11 ? n4270 : n3256;
  assign n4272 = pi10 ? n4268 : n4271;
  assign n4273 = pi09 ? n4267 : n4272;
  assign n4274 = pi08 ? n4254 : n4273;
  assign n4275 = pi07 ? n4235 : n4274;
  assign n4276 = pi09 ? n4253 : n4267;
  assign n4277 = pi13 ? n4249 : n4051;
  assign n4278 = pi12 ? n26 : n4277;
  assign n4279 = pi11 ? n26 : n4278;
  assign n4280 = pi10 ? n26 : n4279;
  assign n4281 = pi09 ? n4272 : n4280;
  assign n4282 = pi08 ? n4276 : n4281;
  assign n4283 = pi13 ? n4255 : n4051;
  assign n4284 = pi12 ? n26 : n4283;
  assign n4285 = pi13 ? n1344 : n105;
  assign n4286 = pi12 ? n26 : n4285;
  assign n4287 = pi11 ? n4284 : n4286;
  assign n4288 = pi13 ? n4106 : n105;
  assign n4289 = pi12 ? n26 : n4288;
  assign n4290 = pi11 ? n4286 : n4289;
  assign n4291 = pi10 ? n4287 : n4290;
  assign n4292 = pi13 ? n1252 : n105;
  assign n4293 = pi12 ? n26 : n4292;
  assign n4294 = pi14 ? n37 : ~n432;
  assign n4295 = pi13 ? n4294 : n3918;
  assign n4296 = pi12 ? n26 : n4295;
  assign n4297 = pi11 ? n4293 : n4296;
  assign n4298 = pi13 ? n4222 : n3066;
  assign n4299 = pi12 ? n26 : n4298;
  assign n4300 = pi10 ? n4297 : n4299;
  assign n4301 = pi09 ? n4291 : n4300;
  assign n4302 = pi14 ? n786 : ~n29;
  assign n4303 = pi13 ? n4302 : n3066;
  assign n4304 = pi12 ? n26 : n4303;
  assign n4305 = pi14 ? n432 : ~n29;
  assign n4306 = pi13 ? n4305 : n2979;
  assign n4307 = pi12 ? n26 : n4306;
  assign n4308 = pi11 ? n4304 : n4307;
  assign n4309 = pi13 ? n4302 : n2319;
  assign n4310 = pi12 ? n26 : n4309;
  assign n4311 = pi13 ? n3983 : n2319;
  assign n4312 = pi12 ? n26 : n4311;
  assign n4313 = pi11 ? n4310 : n4312;
  assign n4314 = pi10 ? n4308 : n4313;
  assign n4315 = pi14 ? n168 : n292;
  assign n4316 = pi14 ? n125 : n61;
  assign n4317 = pi13 ? n4315 : n4316;
  assign n4318 = pi12 ? n26 : n4317;
  assign n4319 = pi13 ? n630 : ~n1378;
  assign n4320 = pi12 ? n26 : n4319;
  assign n4321 = pi11 ? n4318 : n4320;
  assign n4322 = pi14 ? n71 : ~n2420;
  assign n4323 = pi13 ? n2315 : ~n4322;
  assign n4324 = pi12 ? n69 : n4323;
  assign n4325 = pi14 ? n168 : ~n1704;
  assign n4326 = pi13 ? n4325 : n4153;
  assign n4327 = pi12 ? n78 : ~n4326;
  assign n4328 = pi11 ? n4324 : n4327;
  assign n4329 = pi10 ? n4321 : n4328;
  assign n4330 = pi09 ? n4314 : n4329;
  assign n4331 = pi08 ? n4301 : n4330;
  assign n4332 = pi07 ? n4282 : n4331;
  assign n4333 = pi06 ? n4275 : n4332;
  assign n4334 = pi05 ? n4221 : n4333;
  assign n4335 = pi04 ? n4134 : n4334;
  assign n4336 = pi13 ? n4222 : ~n143;
  assign n4337 = pi12 ? n26 : n4336;
  assign n4338 = pi11 ? n26 : n4337;
  assign n4339 = pi13 ? n4226 : ~n130;
  assign n4340 = pi12 ? n26 : n4339;
  assign n4341 = pi14 ? n26 : ~n327;
  assign n4342 = pi13 ? n2319 : ~n4341;
  assign n4343 = pi12 ? n26 : n4342;
  assign n4344 = pi11 ? n4340 : n4343;
  assign n4345 = pi10 ? n4338 : n4344;
  assign n4346 = pi09 ? n26 : n4345;
  assign n4347 = pi08 ? n26 : n4346;
  assign n4348 = pi14 ? n71 : ~n327;
  assign n4349 = pi13 ? n45 : ~n4348;
  assign n4350 = pi12 ? n26 : n4349;
  assign n4351 = pi13 ? n68 : ~n1751;
  assign n4352 = pi12 ? n26 : n4351;
  assign n4353 = pi11 ? n4350 : n4352;
  assign n4354 = pi13 ? n68 : ~n4153;
  assign n4355 = pi12 ? n26 : n4354;
  assign n4356 = pi11 ? n4352 : n4355;
  assign n4357 = pi10 ? n4353 : n4356;
  assign n4358 = pi13 ? n1280 : n3066;
  assign n4359 = pi12 ? n26 : n4358;
  assign n4360 = pi11 ? n26 : n4359;
  assign n4361 = pi10 ? n26 : n4360;
  assign n4362 = pi09 ? n4357 : n4361;
  assign n4363 = pi13 ? n1280 : ~n130;
  assign n4364 = pi12 ? n26 : n4363;
  assign n4365 = pi13 ? n198 : ~n130;
  assign n4366 = pi12 ? n26 : n4365;
  assign n4367 = pi11 ? n4364 : n4366;
  assign n4368 = pi13 ? n68 : ~n72;
  assign n4369 = pi12 ? n26 : n4368;
  assign n4370 = pi11 ? n4369 : n3256;
  assign n4371 = pi10 ? n4367 : n4370;
  assign n4372 = pi09 ? n4359 : n4371;
  assign n4373 = pi08 ? n4362 : n4372;
  assign n4374 = pi07 ? n4347 : n4373;
  assign n4375 = pi09 ? n4361 : n4359;
  assign n4376 = pi13 ? n1280 : n2391;
  assign n4377 = pi12 ? n26 : n4376;
  assign n4378 = pi11 ? n26 : n4377;
  assign n4379 = pi10 ? n26 : n4378;
  assign n4380 = pi09 ? n4371 : n4379;
  assign n4381 = pi08 ? n4375 : n4380;
  assign n4382 = pi13 ? n2598 : n2391;
  assign n4383 = pi12 ? n26 : n4382;
  assign n4384 = pi11 ? n4377 : n4383;
  assign n4385 = pi14 ? n786 : n26;
  assign n4386 = pi13 ? n4385 : n2391;
  assign n4387 = pi12 ? n26 : n4386;
  assign n4388 = pi11 ? n4383 : n4387;
  assign n4389 = pi10 ? n4384 : n4388;
  assign n4390 = pi13 ? n2370 : n2391;
  assign n4391 = pi12 ? n26 : n4390;
  assign n4392 = pi11 ? n4387 : n4391;
  assign n4393 = pi14 ? n45 : ~n4140;
  assign n4394 = pi13 ? n2370 : n4393;
  assign n4395 = pi12 ? n26 : n4394;
  assign n4396 = pi11 ? n4395 : n4391;
  assign n4397 = pi10 ? n4392 : n4396;
  assign n4398 = pi09 ? n4389 : n4397;
  assign n4399 = pi13 ? n2370 : n2487;
  assign n4400 = pi12 ? n26 : n4399;
  assign n4401 = pi14 ? n432 : n26;
  assign n4402 = pi13 ? n4401 : n1280;
  assign n4403 = pi12 ? n26 : n4402;
  assign n4404 = pi11 ? n4400 : n4403;
  assign n4405 = pi13 ? n2759 : n2319;
  assign n4406 = pi12 ? n26 : n4405;
  assign n4407 = pi13 ? n630 : n1705;
  assign n4408 = pi12 ? n26 : n4407;
  assign n4409 = pi11 ? n4406 : n4408;
  assign n4410 = pi10 ? n4404 : n4409;
  assign n4411 = pi13 ? n630 : ~n79;
  assign n4412 = pi12 ? n26 : n4411;
  assign n4413 = pi13 ? n57 : n72;
  assign n4414 = pi12 ? n26 : ~n4413;
  assign n4415 = pi11 ? n4412 : n4414;
  assign n4416 = pi13 ? n1252 : n72;
  assign n4417 = pi12 ? n69 : ~n4416;
  assign n4418 = pi12 ? n78 : n2915;
  assign n4419 = pi11 ? n4417 : n4418;
  assign n4420 = pi10 ? n4415 : n4419;
  assign n4421 = pi09 ? n4410 : n4420;
  assign n4422 = pi08 ? n4398 : n4421;
  assign n4423 = pi07 ? n4381 : n4422;
  assign n4424 = pi06 ? n4374 : n4423;
  assign n4425 = pi14 ? n29 : ~n29;
  assign n4426 = pi13 ? n4425 : ~n143;
  assign n4427 = pi12 ? n26 : n4426;
  assign n4428 = pi11 ? n26 : n4427;
  assign n4429 = pi13 ? n2370 : ~n4141;
  assign n4430 = pi12 ? n26 : n4429;
  assign n4431 = pi13 ? n2319 : ~n79;
  assign n4432 = pi12 ? n26 : n4431;
  assign n4433 = pi11 ? n4430 : n4432;
  assign n4434 = pi10 ? n4428 : n4433;
  assign n4435 = pi09 ? n26 : n4434;
  assign n4436 = pi08 ? n26 : n4435;
  assign n4437 = pi13 ? n3231 : ~n4348;
  assign n4438 = pi12 ? n26 : n4437;
  assign n4439 = pi13 ? n45 : ~n1751;
  assign n4440 = pi12 ? n26 : n4439;
  assign n4441 = pi11 ? n4438 : n4440;
  assign n4442 = pi14 ? n37 : ~n2386;
  assign n4443 = pi13 ? n68 : ~n4442;
  assign n4444 = pi12 ? n26 : n4443;
  assign n4445 = pi11 ? n4444 : n3256;
  assign n4446 = pi10 ? n4441 : n4445;
  assign n4447 = pi09 ? n4446 : n26;
  assign n4448 = pi08 ? n4447 : n26;
  assign n4449 = pi07 ? n4436 : n4448;
  assign n4450 = pi06 ? n4449 : n26;
  assign n4451 = pi05 ? n4424 : n4450;
  assign n4452 = pi13 ? n2370 : ~n57;
  assign n4453 = pi12 ? n26 : n4452;
  assign n4454 = pi13 ? n1135 : ~n4229;
  assign n4455 = pi12 ? n26 : n4454;
  assign n4456 = pi11 ? n4453 : n4455;
  assign n4457 = pi10 ? n4428 : n4456;
  assign n4458 = pi09 ? n26 : n4457;
  assign n4459 = pi08 ? n26 : n4458;
  assign n4460 = pi14 ? n125 : n45;
  assign n4461 = pi13 ? n4460 : ~n4348;
  assign n4462 = pi12 ? n26 : n4461;
  assign n4463 = pi13 ? n269 : ~n1751;
  assign n4464 = pi12 ? n26 : n4463;
  assign n4465 = pi11 ? n4462 : n4464;
  assign n4466 = pi10 ? n4465 : n4445;
  assign n4467 = pi09 ? n4466 : n26;
  assign n4468 = pi08 ? n4467 : n26;
  assign n4469 = pi07 ? n4459 : n4468;
  assign n4470 = pi06 ? n4469 : n26;
  assign n4471 = pi14 ? n125 : ~n29;
  assign n4472 = pi13 ? n4471 : ~n143;
  assign n4473 = pi12 ? n26 : n4472;
  assign n4474 = pi11 ? n26 : n4473;
  assign n4475 = pi13 ? n1135 : ~n130;
  assign n4476 = pi12 ? n26 : n4475;
  assign n4477 = pi13 ? n1135 : ~n72;
  assign n4478 = pi12 ? n26 : n4477;
  assign n4479 = pi11 ? n4476 : n4478;
  assign n4480 = pi10 ? n4474 : n4479;
  assign n4481 = pi09 ? n26 : n4480;
  assign n4482 = pi08 ? n26 : n4481;
  assign n4483 = pi14 ? n37 : ~n327;
  assign n4484 = pi13 ? n269 : ~n4483;
  assign n4485 = pi12 ? n26 : n4484;
  assign n4486 = pi11 ? n4462 : n4485;
  assign n4487 = pi13 ? n2315 : ~n4442;
  assign n4488 = pi12 ? n26 : n4487;
  assign n4489 = pi11 ? n4488 : n3256;
  assign n4490 = pi10 ? n4486 : n4489;
  assign n4491 = pi13 ? n149 : n2539;
  assign n4492 = pi12 ? n26 : n4491;
  assign n4493 = pi13 ? n2391 : n1280;
  assign n4494 = pi12 ? n26 : n4493;
  assign n4495 = pi11 ? n4492 : n4494;
  assign n4496 = pi13 ? n2391 : n1705;
  assign n4497 = pi12 ? n26 : n4496;
  assign n4498 = pi13 ? n2391 : n639;
  assign n4499 = pi12 ? n26 : n4498;
  assign n4500 = pi11 ? n4497 : n4499;
  assign n4501 = pi10 ? n4495 : n4500;
  assign n4502 = pi09 ? n4490 : n4501;
  assign n4503 = pi08 ? n4502 : n2393;
  assign n4504 = pi07 ? n4482 : n4503;
  assign n4505 = pi06 ? n4504 : n2393;
  assign n4506 = pi05 ? n4470 : n4505;
  assign n4507 = pi04 ? n4451 : n4506;
  assign n4508 = pi03 ? n4335 : n4507;
  assign n4509 = pi13 ? n4460 : ~n72;
  assign n4510 = pi12 ? n26 : n4509;
  assign n4511 = pi14 ? n152 : n45;
  assign n4512 = pi13 ? n4511 : ~n38;
  assign n4513 = pi12 ? n26 : n4512;
  assign n4514 = pi11 ? n4510 : n4513;
  assign n4515 = pi13 ? n269 : ~n38;
  assign n4516 = pi12 ? n26 : n4515;
  assign n4517 = pi11 ? n4516 : n3256;
  assign n4518 = pi10 ? n4514 : n4517;
  assign n4519 = pi14 ? n26 : n1548;
  assign n4520 = pi13 ? n4519 : n4167;
  assign n4521 = pi12 ? n26 : n4520;
  assign n4522 = pi13 ? n4125 : n1850;
  assign n4523 = pi12 ? n26 : n4522;
  assign n4524 = pi11 ? n4521 : n4523;
  assign n4525 = pi13 ? n3100 : n2347;
  assign n4526 = pi12 ? n26 : n4525;
  assign n4527 = pi13 ? n4051 : n2762;
  assign n4528 = pi12 ? n26 : n4527;
  assign n4529 = pi11 ? n4526 : n4528;
  assign n4530 = pi10 ? n4524 : n4529;
  assign n4531 = pi09 ? n4518 : n4530;
  assign n4532 = pi13 ? n3918 : n26;
  assign n4533 = pi12 ? n26 : n4532;
  assign n4534 = pi13 ? n1583 : n26;
  assign n4535 = pi12 ? n26 : n4534;
  assign n4536 = pi10 ? n4533 : n4535;
  assign n4537 = pi09 ? n4536 : n4535;
  assign n4538 = pi08 ? n4531 : n4537;
  assign n4539 = pi07 ? n4482 : n4538;
  assign n4540 = pi13 ? n3100 : n26;
  assign n4541 = pi12 ? n26 : n4540;
  assign n4542 = pi11 ? n4535 : n4541;
  assign n4543 = pi10 ? n4535 : n4542;
  assign n4544 = pi09 ? n4535 : n4543;
  assign n4545 = pi08 ? n4535 : n4544;
  assign n4546 = pi07 ? n4535 : n4545;
  assign n4547 = pi06 ? n4539 : n4546;
  assign n4548 = pi13 ? n3873 : ~n143;
  assign n4549 = pi12 ? n26 : n4548;
  assign n4550 = pi11 ? n26 : n4549;
  assign n4551 = pi13 ? n630 : ~n130;
  assign n4552 = pi12 ? n26 : n4551;
  assign n4553 = pi13 ? n630 : ~n72;
  assign n4554 = pi12 ? n26 : n4553;
  assign n4555 = pi11 ? n4552 : n4554;
  assign n4556 = pi10 ? n4550 : n4555;
  assign n4557 = pi09 ? n26 : n4556;
  assign n4558 = pi08 ? n26 : n4557;
  assign n4559 = pi13 ? n46 : n72;
  assign n4560 = pi12 ? n26 : ~n4559;
  assign n4561 = pi13 ? n1344 : n38;
  assign n4562 = pi12 ? n26 : ~n4561;
  assign n4563 = pi11 ? n4560 : n4562;
  assign n4564 = pi13 ? n2448 : ~n38;
  assign n4565 = pi12 ? n124 : n4564;
  assign n4566 = pi11 ? n4565 : n3256;
  assign n4567 = pi10 ? n4563 : n4566;
  assign n4568 = pi13 ? n869 : n125;
  assign n4569 = pi12 ? n78 : ~n4568;
  assign n4570 = pi13 ? n130 : ~n125;
  assign n4571 = pi12 ? n78 : n4570;
  assign n4572 = pi11 ? n4569 : n4571;
  assign n4573 = pi13 ? n630 : ~n2762;
  assign n4574 = pi12 ? n78 : ~n4573;
  assign n4575 = pi13 ? n57 : n2762;
  assign n4576 = pi12 ? n78 : n4575;
  assign n4577 = pi11 ? n4574 : n4576;
  assign n4578 = pi10 ? n4572 : n4577;
  assign n4579 = pi09 ? n4567 : n4578;
  assign n4580 = pi13 ? n57 : n26;
  assign n4581 = pi12 ? n78 : n4580;
  assign n4582 = pi08 ? n4579 : n4581;
  assign n4583 = pi07 ? n4558 : n4582;
  assign n4584 = pi12 ? n69 : n4580;
  assign n4585 = pi12 ? n69 : n4540;
  assign n4586 = pi10 ? n4584 : n4585;
  assign n4587 = pi09 ? n4581 : n4586;
  assign n4588 = pi08 ? n4581 : n4587;
  assign n4589 = pi07 ? n4581 : n4588;
  assign n4590 = pi06 ? n4583 : n4589;
  assign n4591 = pi05 ? n4547 : n4590;
  assign n4592 = pi11 ? n26 : n4552;
  assign n4593 = pi10 ? n4592 : n4555;
  assign n4594 = pi09 ? n26 : n4593;
  assign n4595 = pi08 ? n26 : n4594;
  assign n4596 = pi13 ? n1344 : n72;
  assign n4597 = pi12 ? n26 : ~n4596;
  assign n4598 = pi11 ? n4560 : n4597;
  assign n4599 = pi12 ? n124 : ~n4596;
  assign n4600 = pi11 ? n4599 : n4417;
  assign n4601 = pi10 ? n4598 : n4600;
  assign n4602 = pi13 ? n3782 : n72;
  assign n4603 = pi12 ? n78 : ~n4602;
  assign n4604 = pi13 ? n3888 : n1464;
  assign n4605 = pi12 ? n78 : ~n4604;
  assign n4606 = pi10 ? n4603 : n4605;
  assign n4607 = pi09 ? n4601 : n4606;
  assign n4608 = pi13 ? n3888 : n72;
  assign n4609 = pi12 ? n78 : ~n4608;
  assign n4610 = pi08 ? n4607 : n4609;
  assign n4611 = pi07 ? n4595 : n4610;
  assign n4612 = pi13 ? n869 : n126;
  assign n4613 = pi12 ? n69 : ~n4612;
  assign n4614 = pi11 ? n4609 : n4613;
  assign n4615 = pi13 ? n869 : ~n26;
  assign n4616 = pi12 ? n78 : ~n4615;
  assign n4617 = pi10 ? n4614 : n4616;
  assign n4618 = pi09 ? n4609 : n4617;
  assign n4619 = pi08 ? n4609 : n4618;
  assign n4620 = pi07 ? n4609 : n4619;
  assign n4621 = pi06 ? n4611 : n4620;
  assign n4622 = pi14 ? n63 : ~n71;
  assign n4623 = pi13 ? n4622 : n169;
  assign n4624 = pi12 ? n78 : ~n4623;
  assign n4625 = pi11 ? n26 : n4624;
  assign n4626 = pi10 ? n26 : n4625;
  assign n4627 = pi13 ? n4051 : n57;
  assign n4628 = pi12 ? n78 : ~n4627;
  assign n4629 = pi13 ? n4222 : n415;
  assign n4630 = pi12 ? n78 : ~n4629;
  assign n4631 = pi11 ? n4628 : n4630;
  assign n4632 = pi13 ? n4222 : ~n26;
  assign n4633 = pi12 ? n78 : ~n4632;
  assign n4634 = pi11 ? n4633 : n4616;
  assign n4635 = pi10 ? n4631 : n4634;
  assign n4636 = pi09 ? n4626 : n4635;
  assign n4637 = pi08 ? n26 : n4636;
  assign n4638 = pi07 ? n26 : n4637;
  assign n4639 = pi06 ? n26 : n4638;
  assign n4640 = pi05 ? n4621 : n4639;
  assign n4641 = pi04 ? n4591 : n4640;
  assign n4642 = pi12 ? n26 : ~n176;
  assign n4643 = pi11 ? n26 : n4642;
  assign n4644 = pi10 ? n26 : n4643;
  assign n4645 = pi13 ? n46 : n130;
  assign n4646 = pi12 ? n78 : ~n4645;
  assign n4647 = pi13 ? n1344 : n704;
  assign n4648 = pi12 ? n78 : ~n4647;
  assign n4649 = pi11 ? n4646 : n4648;
  assign n4650 = pi13 ? n4051 : n126;
  assign n4651 = pi12 ? n78 : ~n4650;
  assign n4652 = pi12 ? n78 : ~n2913;
  assign n4653 = pi11 ? n4651 : n4652;
  assign n4654 = pi10 ? n4649 : n4653;
  assign n4655 = pi09 ? n4644 : n4654;
  assign n4656 = pi08 ? n26 : n4655;
  assign n4657 = pi07 ? n26 : n4656;
  assign n4658 = pi06 ? n26 : n4657;
  assign n4659 = pi10 ? n3842 : n4164;
  assign n4660 = pi09 ? n26 : n4659;
  assign n4661 = pi08 ? n26 : n4660;
  assign n4662 = pi07 ? n4661 : n4164;
  assign n4663 = pi14 ? n29 : n63;
  assign n4664 = pi13 ? n57 : ~n4663;
  assign n4665 = pi12 ? n26 : n4664;
  assign n4666 = pi11 ? n4164 : n4665;
  assign n4667 = pi10 ? n4164 : n4666;
  assign n4668 = pi09 ? n4164 : n4667;
  assign n4669 = pi14 ? n29 : n45;
  assign n4670 = pi13 ? n169 : ~n4669;
  assign n4671 = pi12 ? n26 : n4670;
  assign n4672 = pi14 ? n29 : n71;
  assign n4673 = pi13 ? n169 : ~n4672;
  assign n4674 = pi12 ? n26 : n4673;
  assign n4675 = pi11 ? n4671 : n4674;
  assign n4676 = pi13 ? n105 : n3782;
  assign n4677 = pi12 ? n26 : n4676;
  assign n4678 = pi13 ? n176 : n143;
  assign n4679 = pi12 ? n26 : ~n4678;
  assign n4680 = pi11 ? n4677 : n4679;
  assign n4681 = pi10 ? n4675 : n4680;
  assign n4682 = pi14 ? n26 : ~n442;
  assign n4683 = pi13 ? n4682 : n176;
  assign n4684 = pi12 ? n69 : ~n4683;
  assign n4685 = pi13 ? n46 : n736;
  assign n4686 = pi12 ? n78 : ~n4685;
  assign n4687 = pi11 ? n4684 : n4686;
  assign n4688 = pi13 ? n2315 : ~n126;
  assign n4689 = pi12 ? n1203 : n4688;
  assign n4690 = pi13 ? n396 : n126;
  assign n4691 = pi12 ? n78 : ~n4690;
  assign n4692 = pi11 ? n4689 : n4691;
  assign n4693 = pi10 ? n4687 : n4692;
  assign n4694 = pi09 ? n4681 : n4693;
  assign n4695 = pi08 ? n4668 : n4694;
  assign n4696 = pi07 ? n4164 : n4695;
  assign n4697 = pi06 ? n4662 : n4696;
  assign n4698 = pi05 ? n4658 : n4697;
  assign n4699 = pi13 ? n240 : n57;
  assign n4700 = pi12 ? n26 : n4699;
  assign n4701 = pi11 ? n26 : n4700;
  assign n4702 = pi10 ? n4701 : n4700;
  assign n4703 = pi09 ? n26 : n4702;
  assign n4704 = pi08 ? n26 : n4703;
  assign n4705 = pi07 ? n4704 : n4700;
  assign n4706 = pi11 ? n4700 : n3841;
  assign n4707 = pi13 ? n79 : n57;
  assign n4708 = pi12 ? n26 : n4707;
  assign n4709 = pi13 ? n57 : n64;
  assign n4710 = pi12 ? n26 : n4709;
  assign n4711 = pi11 ? n4708 : n4710;
  assign n4712 = pi10 ? n4706 : n4711;
  assign n4713 = pi09 ? n4700 : n4712;
  assign n4714 = pi13 ? n1464 : n4189;
  assign n4715 = pi12 ? n26 : n4714;
  assign n4716 = pi14 ? n37 : ~n71;
  assign n4717 = pi13 ? n79 : n4716;
  assign n4718 = pi12 ? n26 : n4717;
  assign n4719 = pi11 ? n4715 : n4718;
  assign n4720 = pi13 ? n1344 : n3782;
  assign n4721 = pi12 ? n26 : n4720;
  assign n4722 = pi11 ? n4721 : n4679;
  assign n4723 = pi10 ? n4719 : n4722;
  assign n4724 = pi12 ? n69 : ~n57;
  assign n4725 = pi13 ? n46 : n57;
  assign n4726 = pi12 ? n1203 : ~n4725;
  assign n4727 = pi11 ? n4724 : n4726;
  assign n4728 = pi13 ? n1252 : n38;
  assign n4729 = pi12 ? n1203 : ~n4728;
  assign n4730 = pi12 ? n78 : n3255;
  assign n4731 = pi11 ? n4729 : n4730;
  assign n4732 = pi10 ? n4727 : n4731;
  assign n4733 = pi09 ? n4723 : n4732;
  assign n4734 = pi08 ? n4713 : n4733;
  assign n4735 = pi07 ? n4700 : n4734;
  assign n4736 = pi06 ? n4705 : n4735;
  assign n4737 = pi14 ? n45 : ~n29;
  assign n4738 = pi13 ? n4737 : n1583;
  assign n4739 = pi12 ? n26 : n4738;
  assign n4740 = pi11 ? n26 : n4739;
  assign n4741 = pi14 ? n45 : ~n432;
  assign n4742 = pi13 ? n4741 : n1583;
  assign n4743 = pi12 ? n26 : n4742;
  assign n4744 = pi10 ? n4740 : n4743;
  assign n4745 = pi09 ? n26 : n4744;
  assign n4746 = pi08 ? n26 : n4745;
  assign n4747 = pi13 ? n4741 : n3100;
  assign n4748 = pi12 ? n26 : n4747;
  assign n4749 = pi11 ? n4743 : n4748;
  assign n4750 = pi10 ? n4743 : n4749;
  assign n4751 = pi13 ? n1344 : n3100;
  assign n4752 = pi12 ? n26 : n4751;
  assign n4753 = pi14 ? n45 : ~n517;
  assign n4754 = pi13 ? n4753 : n3100;
  assign n4755 = pi12 ? n26 : n4754;
  assign n4756 = pi11 ? n4752 : n4755;
  assign n4757 = pi13 ? n1344 : n1586;
  assign n4758 = pi12 ? n26 : n4757;
  assign n4759 = pi13 ? n4741 : n1586;
  assign n4760 = pi12 ? n26 : n4759;
  assign n4761 = pi11 ? n4758 : n4760;
  assign n4762 = pi10 ? n4756 : n4761;
  assign n4763 = pi09 ? n4750 : n4762;
  assign n4764 = pi08 ? n4743 : n4763;
  assign n4765 = pi07 ? n4746 : n4764;
  assign n4766 = pi14 ? n71 : ~n432;
  assign n4767 = pi13 ? n4766 : n1583;
  assign n4768 = pi12 ? n26 : n4767;
  assign n4769 = pi14 ? n442 : ~n432;
  assign n4770 = pi13 ? n4769 : n3996;
  assign n4771 = pi12 ? n26 : n4770;
  assign n4772 = pi11 ? n4768 : n4771;
  assign n4773 = pi10 ? n4743 : n4772;
  assign n4774 = pi09 ? n4743 : n4773;
  assign n4775 = pi13 ? n4255 : n3782;
  assign n4776 = pi12 ? n26 : n4775;
  assign n4777 = pi14 ? n37 : ~n786;
  assign n4778 = pi13 ? n4255 : n4777;
  assign n4779 = pi12 ? n26 : n4778;
  assign n4780 = pi11 ? n4776 : n4779;
  assign n4781 = pi15 ? n1200 : ~n28;
  assign n4782 = pi14 ? n4781 : ~n29;
  assign n4783 = pi13 ? n4782 : ~n340;
  assign n4784 = pi12 ? n26 : n4783;
  assign n4785 = pi12 ? n26 : ~n2359;
  assign n4786 = pi11 ? n4784 : n4785;
  assign n4787 = pi10 ? n4780 : n4786;
  assign n4788 = pi12 ? n26 : ~n57;
  assign n4789 = pi13 ? n494 : n793;
  assign n4790 = pi12 ? n2243 : ~n4789;
  assign n4791 = pi11 ? n4788 : n4790;
  assign n4792 = pi13 ? n2315 : ~n72;
  assign n4793 = pi12 ? n1203 : n4792;
  assign n4794 = pi11 ? n4793 : n4691;
  assign n4795 = pi10 ? n4791 : n4794;
  assign n4796 = pi09 ? n4787 : n4795;
  assign n4797 = pi08 ? n4774 : n4796;
  assign n4798 = pi07 ? n4743 : n4797;
  assign n4799 = pi06 ? n4765 : n4798;
  assign n4800 = pi05 ? n4736 : n4799;
  assign n4801 = pi04 ? n4698 : n4800;
  assign n4802 = pi03 ? n4641 : n4801;
  assign n4803 = pi02 ? n4508 : n4802;
  assign n4804 = pi01 ? n3995 : n4803;
  assign n4805 = pi11 ? n26 : n4383;
  assign n4806 = pi10 ? n4805 : n4383;
  assign n4807 = pi09 ? n26 : n4806;
  assign n4808 = pi08 ? n26 : n4807;
  assign n4809 = pi14 ? n45 : n233;
  assign n4810 = pi13 ? n4809 : n3918;
  assign n4811 = pi12 ? n26 : n4810;
  assign n4812 = pi11 ? n4811 : n4383;
  assign n4813 = pi10 ? n4137 : n4812;
  assign n4814 = pi09 ? n4383 : n4813;
  assign n4815 = pi08 ? n4383 : n4814;
  assign n4816 = pi07 ? n4808 : n4815;
  assign n4817 = pi13 ? n2598 : n3066;
  assign n4818 = pi12 ? n26 : n4817;
  assign n4819 = pi13 ? n2319 : n2391;
  assign n4820 = pi12 ? n26 : n4819;
  assign n4821 = pi11 ? n4820 : n4387;
  assign n4822 = pi10 ? n4818 : n4821;
  assign n4823 = pi09 ? n4383 : n4822;
  assign n4824 = pi13 ? n57 : n240;
  assign n4825 = pi12 ? n26 : ~n4824;
  assign n4826 = pi11 ? n4552 : n4825;
  assign n4827 = pi10 ? n4377 : n4826;
  assign n4828 = pi12 ? n124 : ~n3843;
  assign n4829 = pi12 ? n69 : ~n4413;
  assign n4830 = pi11 ? n4828 : n4829;
  assign n4831 = pi12 ? n1203 : ~n4416;
  assign n4832 = pi11 ? n4831 : n4730;
  assign n4833 = pi10 ? n4830 : n4832;
  assign n4834 = pi09 ? n4827 : n4833;
  assign n4835 = pi08 ? n4823 : n4834;
  assign n4836 = pi07 ? n4383 : n4835;
  assign n4837 = pi06 ? n4816 : n4836;
  assign n4838 = pi14 ? n37 : n233;
  assign n4839 = pi13 ? n4838 : n1280;
  assign n4840 = pi12 ? n26 : n4839;
  assign n4841 = pi11 ? n26 : n4840;
  assign n4842 = pi13 ? n639 : n1135;
  assign n4843 = pi12 ? n26 : n4842;
  assign n4844 = pi13 ? n639 : ~n240;
  assign n4845 = pi12 ? n26 : n4844;
  assign n4846 = pi11 ? n4843 : n4845;
  assign n4847 = pi10 ? n4841 : n4846;
  assign n4848 = pi09 ? n26 : n4847;
  assign n4849 = pi08 ? n26 : n4848;
  assign n4850 = pi07 ? n26 : n4849;
  assign n4851 = pi11 ? n4016 : n26;
  assign n4852 = pi10 ? n4851 : n26;
  assign n4853 = pi09 ? n4852 : n26;
  assign n4854 = pi08 ? n4853 : n26;
  assign n4855 = pi07 ? n4854 : n26;
  assign n4856 = pi06 ? n4850 : n4855;
  assign n4857 = pi05 ? n4837 : n4856;
  assign n4858 = pi13 ? n4222 : n3782;
  assign n4859 = pi12 ? n26 : n4858;
  assign n4860 = pi11 ? n26 : n4859;
  assign n4861 = pi13 ? n639 : ~n57;
  assign n4862 = pi12 ? n26 : n4861;
  assign n4863 = pi13 ? n639 : ~n72;
  assign n4864 = pi12 ? n26 : n4863;
  assign n4865 = pi11 ? n4862 : n4864;
  assign n4866 = pi10 ? n4860 : n4865;
  assign n4867 = pi09 ? n26 : n4866;
  assign n4868 = pi08 ? n26 : n4867;
  assign n4869 = pi07 ? n26 : n4868;
  assign n4870 = pi11 ? n4093 : n26;
  assign n4871 = pi10 ? n4870 : n26;
  assign n4872 = pi09 ? n4871 : n26;
  assign n4873 = pi08 ? n4872 : n26;
  assign n4874 = pi07 ? n4873 : n26;
  assign n4875 = pi06 ? n4869 : n4874;
  assign n4876 = pi13 ? n202 : n38;
  assign n4877 = pi12 ? n26 : n4876;
  assign n4878 = pi11 ? n4877 : n4427;
  assign n4879 = pi13 ? n639 : ~n38;
  assign n4880 = pi12 ? n26 : n4879;
  assign n4881 = pi11 ? n4453 : n4880;
  assign n4882 = pi10 ? n4878 : n4881;
  assign n4883 = pi09 ? n4164 : n4882;
  assign n4884 = pi08 ? n4164 : n4883;
  assign n4885 = pi07 ? n4661 : n4884;
  assign n4886 = pi13 ? n149 : n1583;
  assign n4887 = pi12 ? n26 : n4886;
  assign n4888 = pi11 ? n3256 : n4887;
  assign n4889 = pi11 ? n4494 : n4497;
  assign n4890 = pi10 ? n4888 : n4889;
  assign n4891 = pi11 ? n4499 : n2393;
  assign n4892 = pi10 ? n4891 : n2393;
  assign n4893 = pi09 ? n4890 : n4892;
  assign n4894 = pi08 ? n4893 : n2393;
  assign n4895 = pi07 ? n4894 : n2393;
  assign n4896 = pi06 ? n4885 : n4895;
  assign n4897 = pi05 ? n4875 : n4896;
  assign n4898 = pi04 ? n4857 : n4897;
  assign n4899 = pi11 ? n3841 : n4708;
  assign n4900 = pi13 ? n57 : n38;
  assign n4901 = pi12 ? n26 : n4900;
  assign n4902 = pi12 ? n26 : n38;
  assign n4903 = pi11 ? n4901 : n4902;
  assign n4904 = pi10 ? n4899 : n4903;
  assign n4905 = pi12 ? n26 : n4728;
  assign n4906 = pi11 ? n4905 : n4427;
  assign n4907 = pi13 ? n4669 : ~n4141;
  assign n4908 = pi12 ? n26 : n4907;
  assign n4909 = pi14 ? n44 : n45;
  assign n4910 = pi13 ? n4909 : ~n4442;
  assign n4911 = pi12 ? n26 : n4910;
  assign n4912 = pi11 ? n4908 : n4911;
  assign n4913 = pi10 ? n4906 : n4912;
  assign n4914 = pi09 ? n4904 : n4913;
  assign n4915 = pi08 ? n4700 : n4914;
  assign n4916 = pi07 ? n4704 : n4915;
  assign n4917 = pi13 ? n4519 : n2539;
  assign n4918 = pi12 ? n26 : n4917;
  assign n4919 = pi11 ? n3256 : n4918;
  assign n4920 = pi13 ? n1583 : n2347;
  assign n4921 = pi12 ? n26 : n4920;
  assign n4922 = pi11 ? n4523 : n4921;
  assign n4923 = pi10 ? n4919 : n4922;
  assign n4924 = pi13 ? n3918 : n2762;
  assign n4925 = pi12 ? n26 : n4924;
  assign n4926 = pi11 ? n4925 : n4533;
  assign n4927 = pi10 ? n4926 : n4533;
  assign n4928 = pi09 ? n4923 : n4927;
  assign n4929 = pi08 ? n4928 : n4533;
  assign n4930 = pi13 ? n4051 : n26;
  assign n4931 = pi12 ? n26 : n4930;
  assign n4932 = pi11 ? n4533 : n4931;
  assign n4933 = pi10 ? n4533 : n4932;
  assign n4934 = pi09 ? n4533 : n4933;
  assign n4935 = pi08 ? n4533 : n4934;
  assign n4936 = pi07 ? n4929 : n4935;
  assign n4937 = pi06 ? n4916 : n4936;
  assign n4938 = pi13 ? n4741 : n3061;
  assign n4939 = pi12 ? n26 : n4938;
  assign n4940 = pi13 ? n4769 : n3782;
  assign n4941 = pi12 ? n26 : n4940;
  assign n4942 = pi11 ? n4939 : n4941;
  assign n4943 = pi14 ? n1638 : ~n432;
  assign n4944 = pi13 ? n4943 : n3782;
  assign n4945 = pi12 ? n26 : n4944;
  assign n4946 = pi13 ? n4294 : n3782;
  assign n4947 = pi12 ? n26 : n4946;
  assign n4948 = pi11 ? n4945 : n4947;
  assign n4949 = pi10 ? n4942 : n4948;
  assign n4950 = pi15 ? n291 : n28;
  assign n4951 = pi14 ? n4950 : ~n26;
  assign n4952 = pi13 ? n3181 : ~n4951;
  assign n4953 = pi12 ? n26 : n4952;
  assign n4954 = pi13 ? n1135 : ~n79;
  assign n4955 = pi12 ? n26 : n4954;
  assign n4956 = pi11 ? n4953 : n4955;
  assign n4957 = pi13 ? n4460 : ~n4229;
  assign n4958 = pi12 ? n26 : n4957;
  assign n4959 = pi13 ? n4460 : ~n4483;
  assign n4960 = pi12 ? n26 : n4959;
  assign n4961 = pi11 ? n4958 : n4960;
  assign n4962 = pi10 ? n4956 : n4961;
  assign n4963 = pi09 ? n4949 : n4962;
  assign n4964 = pi08 ? n4743 : n4963;
  assign n4965 = pi07 ? n4746 : n4964;
  assign n4966 = pi12 ? n26 : n4688;
  assign n4967 = pi13 ? n340 : ~n126;
  assign n4968 = pi12 ? n26 : n4967;
  assign n4969 = pi11 ? n4966 : n4968;
  assign n4970 = pi13 ? n130 : n1850;
  assign n4971 = pi12 ? n26 : n4970;
  assign n4972 = pi13 ? n130 : n2762;
  assign n4973 = pi12 ? n26 : n4972;
  assign n4974 = pi11 ? n4971 : n4973;
  assign n4975 = pi10 ? n4969 : n4974;
  assign n4976 = pi13 ? n79 : n2762;
  assign n4977 = pi12 ? n124 : n4976;
  assign n4978 = pi12 ? n69 : n2116;
  assign n4979 = pi11 ? n4977 : n4978;
  assign n4980 = pi12 ? n78 : n2116;
  assign n4981 = pi10 ? n4979 : n4980;
  assign n4982 = pi09 ? n4975 : n4981;
  assign n4983 = pi08 ? n4982 : n4980;
  assign n4984 = pi12 ? n69 : n4930;
  assign n4985 = pi10 ? n4978 : n4984;
  assign n4986 = pi09 ? n4980 : n4985;
  assign n4987 = pi08 ? n4980 : n4986;
  assign n4988 = pi07 ? n4983 : n4987;
  assign n4989 = pi06 ? n4965 : n4988;
  assign n4990 = pi05 ? n4937 : n4989;
  assign n4991 = pi13 ? n4385 : n3066;
  assign n4992 = pi12 ? n26 : n4991;
  assign n4993 = pi11 ? n4818 : n4992;
  assign n4994 = pi13 ? n2370 : n3066;
  assign n4995 = pi12 ? n26 : n4994;
  assign n4996 = pi11 ? n4992 : n4995;
  assign n4997 = pi10 ? n4993 : n4996;
  assign n4998 = pi13 ? n1135 : ~n57;
  assign n4999 = pi12 ? n26 : n4998;
  assign n5000 = pi11 ? n4453 : n4999;
  assign n5001 = pi13 ? n4511 : ~n72;
  assign n5002 = pi12 ? n26 : n5001;
  assign n5003 = pi11 ? n4510 : n5002;
  assign n5004 = pi10 ? n5000 : n5003;
  assign n5005 = pi09 ? n4997 : n5004;
  assign n5006 = pi08 ? n4383 : n5005;
  assign n5007 = pi07 ? n4808 : n5006;
  assign n5008 = pi14 ? n1832 : n45;
  assign n5009 = pi13 ? n5008 : ~n72;
  assign n5010 = pi12 ? n26 : n5009;
  assign n5011 = pi14 ? n1832 : n37;
  assign n5012 = pi13 ? n5011 : ~n72;
  assign n5013 = pi12 ? n26 : n5012;
  assign n5014 = pi11 ? n5010 : n5013;
  assign n5015 = pi12 ? n26 : ~n4608;
  assign n5016 = pi12 ? n26 : ~n4604;
  assign n5017 = pi11 ? n5015 : n5016;
  assign n5018 = pi10 ? n5014 : n5017;
  assign n5019 = pi12 ? n124 : ~n4604;
  assign n5020 = pi12 ? n69 : ~n4608;
  assign n5021 = pi11 ? n5019 : n5020;
  assign n5022 = pi13 ? n2370 : n72;
  assign n5023 = pi12 ? n78 : ~n5022;
  assign n5024 = pi10 ? n5021 : n5023;
  assign n5025 = pi09 ? n5018 : n5024;
  assign n5026 = pi08 ? n5025 : n5023;
  assign n5027 = pi13 ? n630 : n126;
  assign n5028 = pi12 ? n69 : ~n5027;
  assign n5029 = pi11 ? n5023 : n5028;
  assign n5030 = pi13 ? n630 : ~n26;
  assign n5031 = pi12 ? n78 : ~n5030;
  assign n5032 = pi10 ? n5029 : n5031;
  assign n5033 = pi09 ? n5023 : n5032;
  assign n5034 = pi08 ? n5023 : n5033;
  assign n5035 = pi07 ? n5026 : n5034;
  assign n5036 = pi06 ? n5007 : n5035;
  assign n5037 = pi14 ? n71 : ~n29;
  assign n5038 = pi13 ? n5037 : n415;
  assign n5039 = pi12 ? n78 : ~n5038;
  assign n5040 = pi11 ? n4628 : n5039;
  assign n5041 = pi13 ? n4226 : ~n26;
  assign n5042 = pi12 ? n78 : ~n5041;
  assign n5043 = pi11 ? n5042 : n5031;
  assign n5044 = pi10 ? n5040 : n5043;
  assign n5045 = pi09 ? n4626 : n5044;
  assign n5046 = pi08 ? n26 : n5045;
  assign n5047 = pi07 ? n26 : n5046;
  assign n5048 = pi06 ? n26 : n5047;
  assign n5049 = pi05 ? n5036 : n5048;
  assign n5050 = pi04 ? n4990 : n5049;
  assign n5051 = pi03 ? n4898 : n5050;
  assign n5052 = pi13 ? n1982 : n3100;
  assign n5053 = pi12 ? n26 : n5052;
  assign n5054 = pi11 ? n26 : n5053;
  assign n5055 = pi13 ? n4753 : n4341;
  assign n5056 = pi12 ? n26 : n5055;
  assign n5057 = pi11 ? n5056 : n4758;
  assign n5058 = pi10 ? n5054 : n5057;
  assign n5059 = pi09 ? n26 : n5058;
  assign n5060 = pi08 ? n26 : n5059;
  assign n5061 = pi07 ? n5060 : n4743;
  assign n5062 = pi06 ? n5061 : n4798;
  assign n5063 = pi05 ? n4736 : n5062;
  assign n5064 = pi04 ? n4698 : n5063;
  assign n5065 = pi13 ? n4139 : n3782;
  assign n5066 = pi12 ? n26 : n5065;
  assign n5067 = pi13 ? n4809 : n3782;
  assign n5068 = pi12 ? n26 : n5067;
  assign n5069 = pi11 ? n5066 : n5068;
  assign n5070 = pi10 ? n4138 : n5069;
  assign n5071 = pi09 ? n26 : n5070;
  assign n5072 = pi08 ? n26 : n5071;
  assign n5073 = pi07 ? n5072 : n4383;
  assign n5074 = pi06 ? n5073 : n4836;
  assign n5075 = pi13 ? n3782 : n3918;
  assign n5076 = pi12 ? n26 : n5075;
  assign n5077 = pi11 ? n26 : n5076;
  assign n5078 = pi12 ? n26 : n2319;
  assign n5079 = pi10 ? n5077 : n5078;
  assign n5080 = pi09 ? n26 : n5079;
  assign n5081 = pi08 ? n26 : n5080;
  assign n5082 = pi10 ? n4017 : n26;
  assign n5083 = pi09 ? n5082 : n26;
  assign n5084 = pi08 ? n5083 : n26;
  assign n5085 = pi07 ? n5081 : n5084;
  assign n5086 = pi06 ? n5085 : n26;
  assign n5087 = pi05 ? n5074 : n5086;
  assign n5088 = pi12 ? n26 : n3782;
  assign n5089 = pi11 ? n26 : n5088;
  assign n5090 = pi13 ? n2319 : ~n240;
  assign n5091 = pi12 ? n26 : n5090;
  assign n5092 = pi11 ? n5091 : n4432;
  assign n5093 = pi10 ? n5089 : n5092;
  assign n5094 = pi09 ? n26 : n5093;
  assign n5095 = pi08 ? n26 : n5094;
  assign n5096 = pi11 ? n4149 : n4093;
  assign n5097 = pi10 ? n5096 : n26;
  assign n5098 = pi09 ? n5097 : n26;
  assign n5099 = pi08 ? n5098 : n26;
  assign n5100 = pi07 ? n5095 : n5099;
  assign n5101 = pi06 ? n5100 : n26;
  assign n5102 = pi13 ? n1091 : ~n143;
  assign n5103 = pi12 ? n26 : n5102;
  assign n5104 = pi11 ? n26 : n5103;
  assign n5105 = pi13 ? n2319 : ~n72;
  assign n5106 = pi12 ? n26 : n5105;
  assign n5107 = pi11 ? n4453 : n5106;
  assign n5108 = pi10 ? n5104 : n5107;
  assign n5109 = pi09 ? n26 : n5108;
  assign n5110 = pi08 ? n26 : n5109;
  assign n5111 = pi11 ? n4239 : n3256;
  assign n5112 = pi11 ? n4887 : n4494;
  assign n5113 = pi10 ? n5111 : n5112;
  assign n5114 = pi10 ? n4500 : n2393;
  assign n5115 = pi09 ? n5113 : n5114;
  assign n5116 = pi08 ? n5115 : n2393;
  assign n5117 = pi07 ? n5110 : n5116;
  assign n5118 = pi06 ? n5117 : n2393;
  assign n5119 = pi05 ? n5101 : n5118;
  assign n5120 = pi04 ? n5087 : n5119;
  assign n5121 = pi03 ? n5064 : n5120;
  assign n5122 = pi02 ? n5051 : n5121;
  assign n5123 = pi13 ? n2370 : ~n4341;
  assign n5124 = pi12 ? n26 : n5123;
  assign n5125 = pi13 ? n2319 : ~n38;
  assign n5126 = pi12 ? n26 : n5125;
  assign n5127 = pi11 ? n5124 : n5126;
  assign n5128 = pi10 ? n4428 : n5127;
  assign n5129 = pi09 ? n26 : n5128;
  assign n5130 = pi08 ? n26 : n5129;
  assign n5131 = pi13 ? n68 : ~n38;
  assign n5132 = pi12 ? n26 : n5131;
  assign n5133 = pi11 ? n5132 : n3256;
  assign n5134 = pi10 ? n5133 : n4524;
  assign n5135 = pi13 ? n4051 : n2347;
  assign n5136 = pi12 ? n26 : n5135;
  assign n5137 = pi11 ? n5136 : n4925;
  assign n5138 = pi10 ? n5137 : n4533;
  assign n5139 = pi09 ? n5134 : n5138;
  assign n5140 = pi08 ? n5139 : n4533;
  assign n5141 = pi07 ? n5130 : n5140;
  assign n5142 = pi07 ? n4533 : n4935;
  assign n5143 = pi06 ? n5141 : n5142;
  assign n5144 = pi13 ? n1135 : ~n4483;
  assign n5145 = pi12 ? n26 : n5144;
  assign n5146 = pi11 ? n4476 : n5145;
  assign n5147 = pi10 ? n4474 : n5146;
  assign n5148 = pi09 ? n26 : n5147;
  assign n5149 = pi08 ? n26 : n5148;
  assign n5150 = pi11 ? n4516 : n4966;
  assign n5151 = pi13 ? n130 : ~n4153;
  assign n5152 = pi12 ? n26 : n5151;
  assign n5153 = pi12 ? n26 : n4570;
  assign n5154 = pi11 ? n5152 : n5153;
  assign n5155 = pi10 ? n5150 : n5154;
  assign n5156 = pi13 ? n130 : n1280;
  assign n5157 = pi12 ? n124 : n5156;
  assign n5158 = pi12 ? n69 : n4972;
  assign n5159 = pi11 ? n5157 : n5158;
  assign n5160 = pi10 ? n5159 : n4980;
  assign n5161 = pi09 ? n5155 : n5160;
  assign n5162 = pi08 ? n5161 : n4980;
  assign n5163 = pi07 ? n5149 : n5162;
  assign n5164 = pi11 ? n4980 : n4978;
  assign n5165 = pi10 ? n4980 : n5164;
  assign n5166 = pi13 ? n4229 : n26;
  assign n5167 = pi12 ? n69 : n5166;
  assign n5168 = pi11 ? n4978 : n5167;
  assign n5169 = pi10 ? n5168 : n4980;
  assign n5170 = pi09 ? n5165 : n5169;
  assign n5171 = pi08 ? n5170 : n4980;
  assign n5172 = pi07 ? n5171 : n4980;
  assign n5173 = pi06 ? n5163 : n5172;
  assign n5174 = pi05 ? n5143 : n5173;
  assign n5175 = pi11 ? n26 : n4476;
  assign n5176 = pi13 ? n4460 : ~n4341;
  assign n5177 = pi12 ? n26 : n5176;
  assign n5178 = pi14 ? n168 : n45;
  assign n5179 = pi13 ? n5178 : ~n793;
  assign n5180 = pi12 ? n26 : n5179;
  assign n5181 = pi11 ? n5177 : n5180;
  assign n5182 = pi10 ? n5175 : n5181;
  assign n5183 = pi09 ? n26 : n5182;
  assign n5184 = pi08 ? n26 : n5183;
  assign n5185 = pi12 ? n26 : ~n4602;
  assign n5186 = pi14 ? n71 : ~n2538;
  assign n5187 = pi13 ? n1091 : n5186;
  assign n5188 = pi12 ? n26 : ~n5187;
  assign n5189 = pi11 ? n5185 : n5188;
  assign n5190 = pi10 ? n5002 : n5189;
  assign n5191 = pi12 ? n69 : ~n4604;
  assign n5192 = pi11 ? n5019 : n5191;
  assign n5193 = pi10 ? n5192 : n4609;
  assign n5194 = pi09 ? n5190 : n5193;
  assign n5195 = pi08 ? n5194 : n5023;
  assign n5196 = pi07 ? n5184 : n5195;
  assign n5197 = pi12 ? n69 : ~n5030;
  assign n5198 = pi11 ? n5197 : n5031;
  assign n5199 = pi13 ? n630 : n507;
  assign n5200 = pi12 ? n78 : ~n5199;
  assign n5201 = pi11 ? n5200 : n5023;
  assign n5202 = pi10 ? n5198 : n5201;
  assign n5203 = pi09 ? n5023 : n5202;
  assign n5204 = pi08 ? n5203 : n5023;
  assign n5205 = pi12 ? n78 : n446;
  assign n5206 = pi11 ? n5023 : n5205;
  assign n5207 = pi10 ? n5023 : n5206;
  assign n5208 = pi09 ? n5023 : n5207;
  assign n5209 = pi08 ? n5023 : n5208;
  assign n5210 = pi07 ? n5204 : n5209;
  assign n5211 = pi06 ? n5196 : n5210;
  assign n5212 = pi11 ? n4624 : n4628;
  assign n5213 = pi10 ? n26 : n5212;
  assign n5214 = pi13 ? n3525 : ~n26;
  assign n5215 = pi12 ? n78 : ~n5214;
  assign n5216 = pi10 ? n5215 : n26;
  assign n5217 = pi09 ? n5213 : n5216;
  assign n5218 = pi08 ? n5217 : n26;
  assign n5219 = pi07 ? n5218 : n26;
  assign n5220 = pi06 ? n26 : n5219;
  assign n5221 = pi05 ? n5211 : n5220;
  assign n5222 = pi04 ? n5174 : n5221;
  assign n5223 = pi13 ? n176 : n130;
  assign n5224 = pi12 ? n26 : ~n5223;
  assign n5225 = pi11 ? n5224 : n4646;
  assign n5226 = pi10 ? n26 : n5225;
  assign n5227 = pi12 ? n78 : ~n4728;
  assign n5228 = pi11 ? n5227 : n4652;
  assign n5229 = pi10 ? n5228 : n26;
  assign n5230 = pi09 ? n5226 : n5229;
  assign n5231 = pi08 ? n5230 : n26;
  assign n5232 = pi07 ? n5231 : n26;
  assign n5233 = pi06 ? n26 : n5232;
  assign n5234 = pi13 ? n57 : ~n4669;
  assign n5235 = pi12 ? n26 : n5234;
  assign n5236 = pi11 ? n5235 : n4674;
  assign n5237 = pi10 ? n4666 : n5236;
  assign n5238 = pi09 ? n4164 : n5237;
  assign n5239 = pi08 ? n4164 : n5238;
  assign n5240 = pi07 ? n4661 : n5239;
  assign n5241 = pi14 ? n29 : n37;
  assign n5242 = pi13 ? n169 : ~n5241;
  assign n5243 = pi12 ? n26 : n5242;
  assign n5244 = pi14 ? n71 : ~n63;
  assign n5245 = pi13 ? n5244 : n3782;
  assign n5246 = pi12 ? n26 : n5245;
  assign n5247 = pi11 ? n5243 : n5246;
  assign n5248 = pi15 ? n44 : ~n27;
  assign n5249 = pi14 ? n26 : n5248;
  assign n5250 = pi13 ? n5249 : n176;
  assign n5251 = pi12 ? n69 : ~n5250;
  assign n5252 = pi11 ? n4642 : n5251;
  assign n5253 = pi10 ? n5247 : n5252;
  assign n5254 = pi11 ? n5227 : n4730;
  assign n5255 = pi13 ? n3851 : n26;
  assign n5256 = pi12 ? n26 : n5255;
  assign n5257 = pi13 ? n2391 : n2762;
  assign n5258 = pi12 ? n26 : n5257;
  assign n5259 = pi11 ? n5256 : n5258;
  assign n5260 = pi10 ? n5254 : n5259;
  assign n5261 = pi09 ? n5253 : n5260;
  assign n5262 = pi09 ? n4892 : n2393;
  assign n5263 = pi08 ? n5261 : n5262;
  assign n5264 = pi07 ? n5263 : n2393;
  assign n5265 = pi06 ? n5240 : n5264;
  assign n5266 = pi05 ? n5233 : n5265;
  assign n5267 = pi13 ? n79 : n64;
  assign n5268 = pi12 ? n26 : n5267;
  assign n5269 = pi11 ? n3841 : n5268;
  assign n5270 = pi13 ? n57 : n4189;
  assign n5271 = pi12 ? n26 : n5270;
  assign n5272 = pi14 ? n1638 : ~n71;
  assign n5273 = pi13 ? n1464 : n5272;
  assign n5274 = pi12 ? n26 : n5273;
  assign n5275 = pi11 ? n5271 : n5274;
  assign n5276 = pi10 ? n5269 : n5275;
  assign n5277 = pi09 ? n4700 : n5276;
  assign n5278 = pi08 ? n4700 : n5277;
  assign n5279 = pi07 ? n4704 : n5278;
  assign n5280 = pi13 ? n38 : n3782;
  assign n5281 = pi12 ? n26 : n5280;
  assign n5282 = pi13 ? n1252 : n3782;
  assign n5283 = pi12 ? n26 : n5282;
  assign n5284 = pi11 ? n5281 : n5283;
  assign n5285 = pi13 ? n869 : ~n130;
  assign n5286 = pi12 ? n69 : n5285;
  assign n5287 = pi11 ? n4642 : n5286;
  assign n5288 = pi10 ? n5284 : n5287;
  assign n5289 = pi11 ? n4793 : n4730;
  assign n5290 = pi13 ? n4519 : n26;
  assign n5291 = pi12 ? n26 : n5290;
  assign n5292 = pi13 ? n4125 : n26;
  assign n5293 = pi12 ? n26 : n5292;
  assign n5294 = pi11 ? n5291 : n5293;
  assign n5295 = pi10 ? n5289 : n5294;
  assign n5296 = pi09 ? n5288 : n5295;
  assign n5297 = pi11 ? n4535 : n4533;
  assign n5298 = pi10 ? n5297 : n4533;
  assign n5299 = pi09 ? n5298 : n4533;
  assign n5300 = pi08 ? n5296 : n5299;
  assign n5301 = pi07 ? n5300 : n4935;
  assign n5302 = pi06 ? n5279 : n5301;
  assign n5303 = pi13 ? n79 : n3100;
  assign n5304 = pi12 ? n26 : n5303;
  assign n5305 = pi11 ? n26 : n5304;
  assign n5306 = pi13 ? n1344 : n4341;
  assign n5307 = pi12 ? n26 : n5306;
  assign n5308 = pi11 ? n5307 : n4758;
  assign n5309 = pi10 ? n5305 : n5308;
  assign n5310 = pi09 ? n26 : n5309;
  assign n5311 = pi08 ? n26 : n5310;
  assign n5312 = pi11 ? n4743 : n4768;
  assign n5313 = pi13 ? n4769 : n3061;
  assign n5314 = pi12 ? n26 : n5313;
  assign n5315 = pi11 ? n5314 : n4779;
  assign n5316 = pi10 ? n5312 : n5315;
  assign n5317 = pi09 ? n4743 : n5316;
  assign n5318 = pi08 ? n4743 : n5317;
  assign n5319 = pi07 ? n5311 : n5318;
  assign n5320 = pi14 ? n1638 : ~n29;
  assign n5321 = pi13 ? n5320 : n3782;
  assign n5322 = pi12 ? n26 : n5321;
  assign n5323 = pi13 ? n3873 : n4716;
  assign n5324 = pi12 ? n26 : n5323;
  assign n5325 = pi11 ? n5322 : n5324;
  assign n5326 = pi12 ? n26 : ~n3794;
  assign n5327 = pi11 ? n5224 : n5326;
  assign n5328 = pi10 ? n5325 : n5327;
  assign n5329 = pi12 ? n2243 : n4477;
  assign n5330 = pi13 ? n269 : ~n1139;
  assign n5331 = pi12 ? n78 : n5330;
  assign n5332 = pi11 ? n5329 : n5331;
  assign n5333 = pi14 ? n147 : n125;
  assign n5334 = pi13 ? n5333 : ~n126;
  assign n5335 = pi12 ? n78 : n5334;
  assign n5336 = pi13 ? n2159 : ~n126;
  assign n5337 = pi12 ? n78 : n5336;
  assign n5338 = pi11 ? n5335 : n5337;
  assign n5339 = pi10 ? n5332 : n5338;
  assign n5340 = pi09 ? n5328 : n5339;
  assign n5341 = pi13 ? n130 : n26;
  assign n5342 = pi12 ? n78 : n5341;
  assign n5343 = pi12 ? n78 : n4972;
  assign n5344 = pi11 ? n5342 : n5343;
  assign n5345 = pi10 ? n5344 : n4980;
  assign n5346 = pi09 ? n5345 : n4980;
  assign n5347 = pi08 ? n5340 : n5346;
  assign n5348 = pi07 ? n5347 : n4980;
  assign n5349 = pi06 ? n5319 : n5348;
  assign n5350 = pi05 ? n5302 : n5349;
  assign n5351 = pi04 ? n5266 : n5350;
  assign n5352 = pi03 ? n5222 : n5351;
  assign n5353 = pi13 ? n4139 : n3918;
  assign n5354 = pi12 ? n26 : n5353;
  assign n5355 = pi11 ? n5354 : n4811;
  assign n5356 = pi10 ? n4138 : n5355;
  assign n5357 = pi09 ? n26 : n5356;
  assign n5358 = pi08 ? n26 : n5357;
  assign n5359 = pi13 ? n2319 : n3066;
  assign n5360 = pi12 ? n26 : n5359;
  assign n5361 = pi11 ? n4818 : n5360;
  assign n5362 = pi11 ? n4387 : n4377;
  assign n5363 = pi10 ? n5361 : n5362;
  assign n5364 = pi09 ? n4383 : n5363;
  assign n5365 = pi08 ? n4383 : n5364;
  assign n5366 = pi07 ? n5358 : n5365;
  assign n5367 = pi13 ? n1135 : n3066;
  assign n5368 = pi12 ? n26 : n5367;
  assign n5369 = pi13 ? n630 : n3066;
  assign n5370 = pi12 ? n26 : n5369;
  assign n5371 = pi11 ? n5368 : n5370;
  assign n5372 = pi12 ? n124 : ~n57;
  assign n5373 = pi11 ? n4788 : n5372;
  assign n5374 = pi10 ? n5371 : n5373;
  assign n5375 = pi13 ? n415 : n72;
  assign n5376 = pi12 ? n69 : ~n5375;
  assign n5377 = pi12 ? n78 : ~n4416;
  assign n5378 = pi11 ? n5376 : n5377;
  assign n5379 = pi13 ? n3066 : n72;
  assign n5380 = pi12 ? n78 : ~n5379;
  assign n5381 = pi11 ? n4603 : n5380;
  assign n5382 = pi10 ? n5378 : n5381;
  assign n5383 = pi09 ? n5374 : n5382;
  assign n5384 = pi10 ? n4605 : n4609;
  assign n5385 = pi09 ? n5384 : n5023;
  assign n5386 = pi08 ? n5383 : n5385;
  assign n5387 = pi07 ? n5386 : n5209;
  assign n5388 = pi06 ? n5366 : n5387;
  assign n5389 = pi13 ? n4838 : n2319;
  assign n5390 = pi12 ? n26 : n5389;
  assign n5391 = pi11 ? n5390 : n5078;
  assign n5392 = pi10 ? n5089 : n5391;
  assign n5393 = pi09 ? n26 : n5392;
  assign n5394 = pi08 ? n26 : n5393;
  assign n5395 = pi07 ? n5394 : n5084;
  assign n5396 = pi06 ? n5395 : n26;
  assign n5397 = pi05 ? n5388 : n5396;
  assign n5398 = pi13 ? n4226 : ~n240;
  assign n5399 = pi12 ? n26 : n5398;
  assign n5400 = pi11 ? n5399 : n4432;
  assign n5401 = pi10 ? n5089 : n5400;
  assign n5402 = pi09 ? n26 : n5401;
  assign n5403 = pi08 ? n26 : n5402;
  assign n5404 = pi07 ? n5403 : n5099;
  assign n5405 = pi06 ? n5404 : n26;
  assign n5406 = pi11 ? n5124 : n5106;
  assign n5407 = pi10 ? n5104 : n5406;
  assign n5408 = pi09 ? n26 : n5407;
  assign n5409 = pi08 ? n26 : n5408;
  assign n5410 = pi12 ? n2243 : n4496;
  assign n5411 = pi11 ? n5410 : n4499;
  assign n5412 = pi10 ? n5411 : n2393;
  assign n5413 = pi09 ? n5113 : n5412;
  assign n5414 = pi08 ? n5413 : n2393;
  assign n5415 = pi07 ? n5409 : n5414;
  assign n5416 = pi06 ? n5415 : n2393;
  assign n5417 = pi05 ? n5405 : n5416;
  assign n5418 = pi04 ? n5397 : n5417;
  assign n5419 = pi11 ? n5124 : n5145;
  assign n5420 = pi10 ? n4428 : n5419;
  assign n5421 = pi09 ? n26 : n5420;
  assign n5422 = pi08 ? n26 : n5421;
  assign n5423 = pi13 ? n3918 : n2347;
  assign n5424 = pi12 ? n26 : n5423;
  assign n5425 = pi11 ? n5424 : n4533;
  assign n5426 = pi10 ? n4533 : n5425;
  assign n5427 = pi09 ? n5134 : n5426;
  assign n5428 = pi08 ? n5427 : n4533;
  assign n5429 = pi07 ? n5422 : n5428;
  assign n5430 = pi06 ? n5429 : n5142;
  assign n5431 = pi14 ? n168 : ~n61;
  assign n5432 = pi13 ? n130 : ~n5431;
  assign n5433 = pi12 ? n26 : n5432;
  assign n5434 = pi13 ? n149 : n1850;
  assign n5435 = pi12 ? n26 : n5434;
  assign n5436 = pi11 ? n5433 : n5435;
  assign n5437 = pi10 ? n5133 : n5436;
  assign n5438 = pi14 ? n442 : n26;
  assign n5439 = pi13 ? n4125 : n5438;
  assign n5440 = pi12 ? n124 : n5439;
  assign n5441 = pi13 ? n4125 : n2904;
  assign n5442 = pi12 ? n26 : n5441;
  assign n5443 = pi11 ? n5440 : n5442;
  assign n5444 = pi12 ? n69 : n4527;
  assign n5445 = pi12 ? n69 : n4532;
  assign n5446 = pi11 ? n5444 : n5445;
  assign n5447 = pi10 ? n5443 : n5446;
  assign n5448 = pi09 ? n5437 : n5447;
  assign n5449 = pi08 ? n5448 : n5445;
  assign n5450 = pi07 ? n5149 : n5449;
  assign n5451 = pi11 ? n5445 : n4984;
  assign n5452 = pi10 ? n5445 : n5451;
  assign n5453 = pi09 ? n5445 : n5452;
  assign n5454 = pi08 ? n5445 : n5453;
  assign n5455 = pi07 ? n5445 : n5454;
  assign n5456 = pi06 ? n5450 : n5455;
  assign n5457 = pi05 ? n5430 : n5456;
  assign n5458 = pi13 ? n4460 : ~n415;
  assign n5459 = pi12 ? n26 : n5458;
  assign n5460 = pi11 ? n5177 : n5459;
  assign n5461 = pi10 ? n4474 : n5460;
  assign n5462 = pi09 ? n26 : n5461;
  assign n5463 = pi08 ? n26 : n5462;
  assign n5464 = pi13 ? n269 : ~n126;
  assign n5465 = pi12 ? n26 : n5464;
  assign n5466 = pi11 ? n4516 : n5465;
  assign n5467 = pi13 ? n143 : ~n126;
  assign n5468 = pi12 ? n26 : n5467;
  assign n5469 = pi14 ? n125 : ~n2538;
  assign n5470 = pi13 ? n4325 : n5469;
  assign n5471 = pi12 ? n26 : ~n5470;
  assign n5472 = pi11 ? n5468 : n5471;
  assign n5473 = pi10 ? n5466 : n5472;
  assign n5474 = pi13 ? n130 : ~n2850;
  assign n5475 = pi12 ? n78 : n5474;
  assign n5476 = pi13 ? n869 : n2850;
  assign n5477 = pi12 ? n78 : ~n5476;
  assign n5478 = pi11 ? n5475 : n5477;
  assign n5479 = pi14 ? n1872 : ~n26;
  assign n5480 = pi13 ? n130 : ~n5479;
  assign n5481 = pi12 ? n78 : n5480;
  assign n5482 = pi13 ? n130 : ~n126;
  assign n5483 = pi12 ? n78 : n5482;
  assign n5484 = pi11 ? n5481 : n5483;
  assign n5485 = pi10 ? n5478 : n5484;
  assign n5486 = pi09 ? n5473 : n5485;
  assign n5487 = pi10 ? n5205 : n5483;
  assign n5488 = pi09 ? n5487 : n5483;
  assign n5489 = pi08 ? n5486 : n5488;
  assign n5490 = pi07 ? n5463 : n5489;
  assign n5491 = pi06 ? n5490 : n5483;
  assign n5492 = pi13 ? n5178 : ~n130;
  assign n5493 = pi12 ? n26 : n5492;
  assign n5494 = pi13 ? n5178 : ~n72;
  assign n5495 = pi12 ? n26 : n5494;
  assign n5496 = pi11 ? n5493 : n5495;
  assign n5497 = pi10 ? n4592 : n5496;
  assign n5498 = pi09 ? n26 : n5497;
  assign n5499 = pi08 ? n26 : n5498;
  assign n5500 = pi12 ? n124 : ~n4602;
  assign n5501 = pi13 ? n3782 : n1925;
  assign n5502 = pi12 ? n69 : ~n5501;
  assign n5503 = pi11 ? n5500 : n5502;
  assign n5504 = pi10 ? n4597 : n5503;
  assign n5505 = pi14 ? n1201 : n125;
  assign n5506 = pi13 ? n3066 : n5505;
  assign n5507 = pi12 ? n78 : ~n5506;
  assign n5508 = pi11 ? n5507 : n4605;
  assign n5509 = pi11 ? n4605 : n4609;
  assign n5510 = pi10 ? n5508 : n5509;
  assign n5511 = pi09 ? n5504 : n5510;
  assign n5512 = pi10 ? n5023 : n4609;
  assign n5513 = pi09 ? n5512 : n4609;
  assign n5514 = pi08 ? n5511 : n5513;
  assign n5515 = pi07 ? n5499 : n5514;
  assign n5516 = pi11 ? n4609 : n5483;
  assign n5517 = pi10 ? n4609 : n5516;
  assign n5518 = pi09 ? n4609 : n5517;
  assign n5519 = pi08 ? n4609 : n5518;
  assign n5520 = pi07 ? n4609 : n5519;
  assign n5521 = pi06 ? n5515 : n5520;
  assign n5522 = pi05 ? n5491 : n5521;
  assign n5523 = pi04 ? n5457 : n5522;
  assign n5524 = pi03 ? n5418 : n5523;
  assign n5525 = pi02 ? n5352 : n5524;
  assign n5526 = pi01 ? n5122 : n5525;
  assign n5527 = pi00 ? n4804 : n5526;
  assign n5528 = pi14 ? n45 : n29;
  assign n5529 = pi13 ? n169 : n5528;
  assign n5530 = pi12 ? n26 : n5529;
  assign n5531 = pi11 ? n26 : n5530;
  assign n5532 = pi14 ? n131 : ~n29;
  assign n5533 = pi13 ? n169 : ~n5532;
  assign n5534 = pi12 ? n26 : n5533;
  assign n5535 = pi10 ? n5531 : n5534;
  assign n5536 = pi09 ? n26 : n5535;
  assign n5537 = pi08 ? n26 : n5536;
  assign n5538 = pi13 ? n130 : ~n5532;
  assign n5539 = pi12 ? n26 : n5538;
  assign n5540 = pi11 ? n5534 : n5539;
  assign n5541 = pi13 ? n176 : ~n5532;
  assign n5542 = pi12 ? n26 : n5541;
  assign n5543 = pi11 ? n5539 : n5542;
  assign n5544 = pi10 ? n5540 : n5543;
  assign n5545 = pi14 ? n131 : ~n37;
  assign n5546 = pi13 ? n176 : ~n5545;
  assign n5547 = pi12 ? n26 : n5546;
  assign n5548 = pi13 ? n143 : ~n3061;
  assign n5549 = pi12 ? n26 : n5548;
  assign n5550 = pi11 ? n5547 : n5549;
  assign n5551 = pi13 ? n143 : ~n1252;
  assign n5552 = pi12 ? n26 : n5551;
  assign n5553 = pi13 ? n77 : ~n202;
  assign n5554 = pi12 ? n26 : n5553;
  assign n5555 = pi11 ? n5552 : n5554;
  assign n5556 = pi10 ? n5550 : n5555;
  assign n5557 = pi09 ? n5544 : n5556;
  assign n5558 = pi13 ? n130 : n5528;
  assign n5559 = pi12 ? n26 : n5558;
  assign n5560 = pi11 ? n26 : n5559;
  assign n5561 = pi10 ? n5560 : n5543;
  assign n5562 = pi09 ? n3793 : n5561;
  assign n5563 = pi08 ? n5557 : n5562;
  assign n5564 = pi07 ? n5537 : n5563;
  assign n5565 = pi09 ? n5556 : n3793;
  assign n5566 = pi09 ? n5561 : n5556;
  assign n5567 = pi08 ? n5565 : n5566;
  assign n5568 = pi11 ? n26 : n3565;
  assign n5569 = pi13 ? n97 : ~n723;
  assign n5570 = pi12 ? n26 : n5569;
  assign n5571 = pi13 ? n26 : ~n723;
  assign n5572 = pi12 ? n26 : n5571;
  assign n5573 = pi11 ? n5570 : n5572;
  assign n5574 = pi10 ? n5568 : n5573;
  assign n5575 = pi09 ? n3793 : n5574;
  assign n5576 = pi13 ? n68 : ~n1252;
  assign n5577 = pi12 ? n26 : n5576;
  assign n5578 = pi14 ? n916 : ~n45;
  assign n5579 = pi13 ? n164 : ~n5578;
  assign n5580 = pi12 ? n26 : n5579;
  assign n5581 = pi11 ? n5577 : n5580;
  assign n5582 = pi13 ? n68 : ~n5578;
  assign n5583 = pi12 ? n26 : n5582;
  assign n5584 = pi11 ? n5580 : n5583;
  assign n5585 = pi10 ? n5581 : n5584;
  assign n5586 = pi14 ? n61 : ~n45;
  assign n5587 = pi13 ? n68 : ~n5586;
  assign n5588 = pi12 ? n26 : n5587;
  assign n5589 = pi14 ? n61 : n442;
  assign n5590 = pi14 ? n2538 : ~n26;
  assign n5591 = pi13 ? n5589 : ~n5590;
  assign n5592 = pi12 ? n26 : n5591;
  assign n5593 = pi11 ? n5588 : n5592;
  assign n5594 = pi14 ? n1355 : n517;
  assign n5595 = pi13 ? n5594 : n2370;
  assign n5596 = pi12 ? n26 : n5595;
  assign n5597 = pi12 ? n26 : n639;
  assign n5598 = pi11 ? n5596 : n5597;
  assign n5599 = pi10 ? n5593 : n5598;
  assign n5600 = pi09 ? n5585 : n5599;
  assign n5601 = pi08 ? n5575 : n5600;
  assign n5602 = pi07 ? n5567 : n5601;
  assign n5603 = pi06 ? n5564 : n5602;
  assign n5604 = pi05 ? n26 : n5603;
  assign n5605 = pi13 ? n57 : n1567;
  assign n5606 = pi12 ? n26 : n5605;
  assign n5607 = pi11 ? n26 : n5606;
  assign n5608 = pi11 ? n3841 : n3765;
  assign n5609 = pi10 ? n5607 : n5608;
  assign n5610 = pi09 ? n26 : n5609;
  assign n5611 = pi08 ? n26 : n5610;
  assign n5612 = pi13 ? n3851 : n57;
  assign n5613 = pi12 ? n26 : n5612;
  assign n5614 = pi11 ? n5613 : n3858;
  assign n5615 = pi14 ? n45 : n1548;
  assign n5616 = pi13 ? n132 : n5615;
  assign n5617 = pi12 ? n26 : n5616;
  assign n5618 = pi11 ? n3855 : n5617;
  assign n5619 = pi10 ? n5614 : n5618;
  assign n5620 = pi14 ? n45 : n1704;
  assign n5621 = pi13 ? n321 : n5620;
  assign n5622 = pi12 ? n26 : n5621;
  assign n5623 = pi11 ? n5617 : n5622;
  assign n5624 = pi11 ? n5622 : n2911;
  assign n5625 = pi10 ? n5623 : n5624;
  assign n5626 = pi09 ? n5619 : n5625;
  assign n5627 = pi13 ? n97 : ~n79;
  assign n5628 = pi12 ? n26 : n5627;
  assign n5629 = pi11 ? n5628 : n3875;
  assign n5630 = pi10 ? n5629 : n26;
  assign n5631 = pi13 ? n130 : n1567;
  assign n5632 = pi12 ? n26 : n5631;
  assign n5633 = pi11 ? n26 : n5632;
  assign n5634 = pi10 ? n5633 : n5618;
  assign n5635 = pi09 ? n5630 : n5634;
  assign n5636 = pi08 ? n5626 : n5635;
  assign n5637 = pi07 ? n5611 : n5636;
  assign n5638 = pi09 ? n5625 : n5630;
  assign n5639 = pi09 ? n5634 : n5625;
  assign n5640 = pi08 ? n5638 : n5639;
  assign n5641 = pi13 ? n130 : n143;
  assign n5642 = pi12 ? n26 : n5641;
  assign n5643 = pi11 ? n26 : n5642;
  assign n5644 = pi13 ? n57 : ~n1091;
  assign n5645 = pi12 ? n26 : n5644;
  assign n5646 = pi13 ? n57 : ~n1942;
  assign n5647 = pi12 ? n26 : n5646;
  assign n5648 = pi11 ? n5645 : n5647;
  assign n5649 = pi10 ? n5643 : n5648;
  assign n5650 = pi09 ? n5630 : n5649;
  assign n5651 = pi14 ? n1138 : ~n45;
  assign n5652 = pi13 ? n1438 : ~n5651;
  assign n5653 = pi12 ? n26 : n5652;
  assign n5654 = pi13 ? n143 : ~n1914;
  assign n5655 = pi12 ? n26 : n5654;
  assign n5656 = pi11 ? n5653 : n5655;
  assign n5657 = pi10 ? n5647 : n5656;
  assign n5658 = pi14 ? n44 : ~n37;
  assign n5659 = pi13 ? n143 : ~n5658;
  assign n5660 = pi12 ? n26 : n5659;
  assign n5661 = pi14 ? n125 : ~n63;
  assign n5662 = pi14 ? n233 : ~n1638;
  assign n5663 = pi13 ? n5661 : n5662;
  assign n5664 = pi12 ? n26 : ~n5663;
  assign n5665 = pi11 ? n5660 : n5664;
  assign n5666 = pi14 ? n916 : ~n125;
  assign n5667 = pi13 ? n3066 : n5666;
  assign n5668 = pi12 ? n26 : n5667;
  assign n5669 = pi13 ? n3066 : n639;
  assign n5670 = pi12 ? n26 : n5669;
  assign n5671 = pi11 ? n5668 : n5670;
  assign n5672 = pi10 ? n5665 : n5671;
  assign n5673 = pi09 ? n5657 : n5672;
  assign n5674 = pi08 ? n5650 : n5673;
  assign n5675 = pi07 ? n5640 : n5674;
  assign n5676 = pi06 ? n5637 : n5675;
  assign n5677 = pi14 ? n320 : ~n1138;
  assign n5678 = pi13 ? n1583 : n5677;
  assign n5679 = pi12 ? n26 : n5678;
  assign n5680 = pi11 ? n26 : n5679;
  assign n5681 = pi14 ? n320 : ~n147;
  assign n5682 = pi13 ? n149 : n5681;
  assign n5683 = pi12 ? n26 : n5682;
  assign n5684 = pi13 ? n3851 : n5681;
  assign n5685 = pi12 ? n26 : n5684;
  assign n5686 = pi11 ? n5683 : n5685;
  assign n5687 = pi10 ? n5680 : n5686;
  assign n5688 = pi09 ? n26 : n5687;
  assign n5689 = pi08 ? n26 : n5688;
  assign n5690 = pi14 ? n320 : ~n125;
  assign n5691 = pi13 ? n26 : n5690;
  assign n5692 = pi12 ? n26 : n5691;
  assign n5693 = pi10 ? n5683 : n5692;
  assign n5694 = pi13 ? n26 : n2522;
  assign n5695 = pi12 ? n26 : n5694;
  assign n5696 = pi13 ? n97 : n68;
  assign n5697 = pi12 ? n26 : n5696;
  assign n5698 = pi11 ? n5695 : n5697;
  assign n5699 = pi10 ? n5692 : n5698;
  assign n5700 = pi09 ? n5693 : n5699;
  assign n5701 = pi13 ? n97 : ~n105;
  assign n5702 = pi12 ? n26 : n5701;
  assign n5703 = pi13 ? n26 : n869;
  assign n5704 = pi12 ? n26 : n5703;
  assign n5705 = pi11 ? n5702 : n5704;
  assign n5706 = pi10 ? n5705 : n26;
  assign n5707 = pi13 ? n3942 : n5677;
  assign n5708 = pi12 ? n26 : n5707;
  assign n5709 = pi11 ? n26 : n5708;
  assign n5710 = pi10 ? n5709 : n5692;
  assign n5711 = pi09 ? n5706 : n5710;
  assign n5712 = pi08 ? n5700 : n5711;
  assign n5713 = pi07 ? n5689 : n5712;
  assign n5714 = pi09 ? n5699 : n5706;
  assign n5715 = pi09 ? n5710 : n5699;
  assign n5716 = pi08 ? n5714 : n5715;
  assign n5717 = pi13 ? n240 : n143;
  assign n5718 = pi12 ? n26 : n5717;
  assign n5719 = pi11 ? n26 : n5718;
  assign n5720 = pi13 ? n240 : ~n1091;
  assign n5721 = pi12 ? n26 : n5720;
  assign n5722 = pi13 ? n240 : ~n3782;
  assign n5723 = pi12 ? n26 : n5722;
  assign n5724 = pi11 ? n5721 : n5723;
  assign n5725 = pi10 ? n5719 : n5724;
  assign n5726 = pi09 ? n5706 : n5725;
  assign n5727 = pi13 ? n57 : ~n3782;
  assign n5728 = pi12 ? n26 : n5727;
  assign n5729 = pi13 ? n518 : ~n3782;
  assign n5730 = pi12 ? n26 : n5729;
  assign n5731 = pi11 ? n5728 : n5730;
  assign n5732 = pi13 ? n130 : ~n3782;
  assign n5733 = pi12 ? n26 : n5732;
  assign n5734 = pi13 ? n143 : ~n3969;
  assign n5735 = pi12 ? n26 : n5734;
  assign n5736 = pi11 ? n5733 : n5735;
  assign n5737 = pi10 ? n5731 : n5736;
  assign n5738 = pi14 ? n45 : ~n1704;
  assign n5739 = pi13 ? n143 : ~n5738;
  assign n5740 = pi12 ? n26 : n5739;
  assign n5741 = pi14 ? n1138 : ~n37;
  assign n5742 = pi13 ? n5741 : n1586;
  assign n5743 = pi12 ? n26 : ~n5742;
  assign n5744 = pi11 ? n5740 : n5743;
  assign n5745 = pi13 ? n2159 : ~n1135;
  assign n5746 = pi12 ? n26 : ~n5745;
  assign n5747 = pi13 ? n4716 : n4222;
  assign n5748 = pi12 ? n654 : n5747;
  assign n5749 = pi11 ? n5746 : n5748;
  assign n5750 = pi10 ? n5744 : n5749;
  assign n5751 = pi09 ? n5737 : n5750;
  assign n5752 = pi08 ? n5726 : n5751;
  assign n5753 = pi07 ? n5716 : n5752;
  assign n5754 = pi06 ? n5713 : n5753;
  assign n5755 = pi05 ? n5676 : n5754;
  assign n5756 = pi04 ? n5604 : n5755;
  assign n5757 = pi03 ? n26 : n5756;
  assign n5758 = pi02 ? n26 : n5757;
  assign n5759 = pi13 ? n3996 : n5677;
  assign n5760 = pi12 ? n26 : n5759;
  assign n5761 = pi11 ? n26 : n5760;
  assign n5762 = pi10 ? n5761 : n4004;
  assign n5763 = pi09 ? n26 : n5762;
  assign n5764 = pi08 ? n26 : n5763;
  assign n5765 = pi13 ? n3023 : n2319;
  assign n5766 = pi12 ? n26 : n5765;
  assign n5767 = pi13 ? n2519 : n2319;
  assign n5768 = pi12 ? n26 : n5767;
  assign n5769 = pi11 ? n5766 : n5768;
  assign n5770 = pi10 ? n5769 : n2342;
  assign n5771 = pi14 ? n26 : n1638;
  assign n5772 = pi13 ? n5771 : n68;
  assign n5773 = pi12 ? n26 : n5772;
  assign n5774 = pi11 ? n26 : n5773;
  assign n5775 = pi10 ? n26 : n5774;
  assign n5776 = pi09 ? n5770 : n5775;
  assign n5777 = pi14 ? n37 : ~n1138;
  assign n5778 = pi13 ? n3942 : n5777;
  assign n5779 = pi12 ? n26 : n5778;
  assign n5780 = pi11 ? n26 : n5779;
  assign n5781 = pi10 ? n5780 : n2342;
  assign n5782 = pi09 ? n5706 : n5781;
  assign n5783 = pi08 ? n5776 : n5782;
  assign n5784 = pi07 ? n5764 : n5783;
  assign n5785 = pi09 ? n5775 : n5706;
  assign n5786 = pi09 ? n5781 : n5775;
  assign n5787 = pi08 ? n5785 : n5786;
  assign n5788 = pi14 ? n45 : n2431;
  assign n5789 = pi13 ? n79 : n5788;
  assign n5790 = pi12 ? n26 : n5789;
  assign n5791 = pi11 ? n26 : n5790;
  assign n5792 = pi10 ? n5791 : n5790;
  assign n5793 = pi09 ? n5706 : n5792;
  assign n5794 = pi13 ? n1464 : n5788;
  assign n5795 = pi12 ? n26 : n5794;
  assign n5796 = pi11 ? n5790 : n5795;
  assign n5797 = pi14 ? n45 : n1138;
  assign n5798 = pi13 ? n130 : n5797;
  assign n5799 = pi12 ? n26 : n5798;
  assign n5800 = pi13 ? n1438 : n5788;
  assign n5801 = pi12 ? n26 : n5800;
  assign n5802 = pi11 ? n5799 : n5801;
  assign n5803 = pi10 ? n5796 : n5802;
  assign n5804 = pi13 ? n57 : n2522;
  assign n5805 = pi12 ? n26 : n5804;
  assign n5806 = pi13 ? n3061 : n3782;
  assign n5807 = pi12 ? n26 : n5806;
  assign n5808 = pi14 ? n320 : ~n71;
  assign n5809 = pi13 ? n5808 : n3782;
  assign n5810 = pi12 ? n26 : n5809;
  assign n5811 = pi11 ? n5807 : n5810;
  assign n5812 = pi10 ? n5805 : n5811;
  assign n5813 = pi09 ? n5803 : n5812;
  assign n5814 = pi08 ? n5793 : n5813;
  assign n5815 = pi07 ? n5787 : n5814;
  assign n5816 = pi06 ? n5784 : n5815;
  assign n5817 = pi13 ? n3918 : n3782;
  assign n5818 = pi12 ? n26 : n5817;
  assign n5819 = pi11 ? n26 : n5818;
  assign n5820 = pi10 ? n5819 : n4063;
  assign n5821 = pi09 ? n26 : n5820;
  assign n5822 = pi08 ? n26 : n5821;
  assign n5823 = pi13 ? n2498 : n1705;
  assign n5824 = pi12 ? n26 : n5823;
  assign n5825 = pi11 ? n5824 : n2341;
  assign n5826 = pi14 ? n2386 : n61;
  assign n5827 = pi13 ? n26 : n5826;
  assign n5828 = pi12 ? n26 : n5827;
  assign n5829 = pi14 ? n125 : ~n2420;
  assign n5830 = pi13 ? n321 : ~n5829;
  assign n5831 = pi12 ? n26 : n5830;
  assign n5832 = pi11 ? n5828 : n5831;
  assign n5833 = pi10 ? n5825 : n5832;
  assign n5834 = pi13 ? n169 : n176;
  assign n5835 = pi12 ? n26 : n5834;
  assign n5836 = pi11 ? n26 : n5835;
  assign n5837 = pi10 ? n26 : n5836;
  assign n5838 = pi09 ? n5833 : n5837;
  assign n5839 = pi13 ? n143 : ~n4051;
  assign n5840 = pi12 ? n26 : n5839;
  assign n5841 = pi13 ? n77 : ~n1347;
  assign n5842 = pi12 ? n26 : n5841;
  assign n5843 = pi11 ? n5840 : n5842;
  assign n5844 = pi10 ? n5843 : n26;
  assign n5845 = pi13 ? n321 : ~n4173;
  assign n5846 = pi12 ? n26 : n5845;
  assign n5847 = pi11 ? n2339 : n5846;
  assign n5848 = pi10 ? n4028 : n5847;
  assign n5849 = pi09 ? n5844 : n5848;
  assign n5850 = pi08 ? n5838 : n5849;
  assign n5851 = pi07 ? n5822 : n5850;
  assign n5852 = pi09 ? n5837 : n5844;
  assign n5853 = pi09 ? n5848 : n5837;
  assign n5854 = pi08 ? n5852 : n5853;
  assign n5855 = pi13 ? n4102 : n5677;
  assign n5856 = pi12 ? n26 : n5855;
  assign n5857 = pi11 ? n26 : n5856;
  assign n5858 = pi13 ? n4106 : n5677;
  assign n5859 = pi12 ? n26 : n5858;
  assign n5860 = pi13 ? n1344 : n5677;
  assign n5861 = pi12 ? n26 : n5860;
  assign n5862 = pi11 ? n5859 : n5861;
  assign n5863 = pi10 ? n5857 : n5862;
  assign n5864 = pi09 ? n5844 : n5863;
  assign n5865 = pi14 ? n2954 : ~n45;
  assign n5866 = pi13 ? n5865 : n5677;
  assign n5867 = pi12 ? n26 : n5866;
  assign n5868 = pi11 ? n5859 : n5867;
  assign n5869 = pi13 ? n1347 : n5677;
  assign n5870 = pi12 ? n26 : n5869;
  assign n5871 = pi14 ? n63 : ~n1400;
  assign n5872 = pi13 ? n5871 : n5677;
  assign n5873 = pi12 ? n26 : n5872;
  assign n5874 = pi11 ? n5870 : n5873;
  assign n5875 = pi10 ? n5868 : n5874;
  assign n5876 = pi14 ? n320 : ~n1400;
  assign n5877 = pi13 ? n1252 : n5876;
  assign n5878 = pi12 ? n26 : n5877;
  assign n5879 = pi14 ? n320 : ~n44;
  assign n5880 = pi13 ? n1252 : n5879;
  assign n5881 = pi12 ? n26 : n5880;
  assign n5882 = pi11 ? n5878 : n5881;
  assign n5883 = pi13 ? n1850 : n3023;
  assign n5884 = pi12 ? n69 : n5883;
  assign n5885 = pi15 ? n44 : n70;
  assign n5886 = pi14 ? n26 : ~n5885;
  assign n5887 = pi13 ? n5886 : n3023;
  assign n5888 = pi12 ? n78 : n5887;
  assign n5889 = pi11 ? n5884 : n5888;
  assign n5890 = pi10 ? n5882 : n5889;
  assign n5891 = pi09 ? n5875 : n5890;
  assign n5892 = pi08 ? n5864 : n5891;
  assign n5893 = pi07 ? n5854 : n5892;
  assign n5894 = pi06 ? n5851 : n5893;
  assign n5895 = pi05 ? n5816 : n5894;
  assign n5896 = pi13 ? n4135 : n5777;
  assign n5897 = pi12 ? n26 : n5896;
  assign n5898 = pi11 ? n26 : n5897;
  assign n5899 = pi14 ? n37 : ~n4140;
  assign n5900 = pi13 ? n4139 : n5899;
  assign n5901 = pi12 ? n26 : n5900;
  assign n5902 = pi11 ? n5901 : n2339;
  assign n5903 = pi10 ? n5898 : n5902;
  assign n5904 = pi09 ? n26 : n5903;
  assign n5905 = pi08 ? n26 : n5904;
  assign n5906 = pi11 ? n2341 : n3207;
  assign n5907 = pi13 ? n26 : n478;
  assign n5908 = pi12 ? n26 : n5907;
  assign n5909 = pi14 ? n26 : ~n1330;
  assign n5910 = pi14 ? n125 : ~n60;
  assign n5911 = pi13 ? n5909 : ~n5910;
  assign n5912 = pi12 ? n26 : n5911;
  assign n5913 = pi11 ? n5908 : n5912;
  assign n5914 = pi10 ? n5906 : n5913;
  assign n5915 = pi14 ? n45 : n131;
  assign n5916 = pi13 ? n169 : n5915;
  assign n5917 = pi12 ? n26 : n5916;
  assign n5918 = pi11 ? n26 : n5917;
  assign n5919 = pi10 ? n26 : n5918;
  assign n5920 = pi09 ? n5914 : n5919;
  assign n5921 = pi14 ? n147 : ~n29;
  assign n5922 = pi13 ? n169 : ~n5921;
  assign n5923 = pi12 ? n26 : n5922;
  assign n5924 = pi11 ? n5923 : n5534;
  assign n5925 = pi10 ? n5924 : n5923;
  assign n5926 = pi13 ? n46 : n79;
  assign n5927 = pi12 ? n26 : n5926;
  assign n5928 = pi13 ? n4167 : n3782;
  assign n5929 = pi12 ? n26 : n5928;
  assign n5930 = pi11 ? n5927 : n5929;
  assign n5931 = pi14 ? n1548 : n327;
  assign n5932 = pi13 ? n26 : n5931;
  assign n5933 = pi12 ? n26 : n5932;
  assign n5934 = pi13 ? n321 : ~n126;
  assign n5935 = pi12 ? n26 : n5934;
  assign n5936 = pi11 ? n5933 : n5935;
  assign n5937 = pi10 ? n5930 : n5936;
  assign n5938 = pi09 ? n5925 : n5937;
  assign n5939 = pi08 ? n5920 : n5938;
  assign n5940 = pi07 ? n5905 : n5939;
  assign n5941 = pi09 ? n5919 : n5925;
  assign n5942 = pi09 ? n5937 : n5919;
  assign n5943 = pi08 ? n5941 : n5942;
  assign n5944 = pi13 ? n64 : n415;
  assign n5945 = pi12 ? n26 : n5944;
  assign n5946 = pi14 ? n2386 : ~n45;
  assign n5947 = pi13 ? n5946 : n3061;
  assign n5948 = pi12 ? n26 : n5947;
  assign n5949 = pi11 ? n5945 : n5948;
  assign n5950 = pi14 ? n786 : ~n37;
  assign n5951 = pi13 ? n5950 : n2319;
  assign n5952 = pi12 ? n26 : n5951;
  assign n5953 = pi11 ? n4194 : n5952;
  assign n5954 = pi10 ? n5949 : n5953;
  assign n5955 = pi09 ? n5923 : n5954;
  assign n5956 = pi14 ? n2386 : ~n37;
  assign n5957 = pi13 ? n5956 : n2319;
  assign n5958 = pi12 ? n26 : n5957;
  assign n5959 = pi11 ? n5958 : n4003;
  assign n5960 = pi14 ? n327 : ~n37;
  assign n5961 = pi13 ? n5960 : n2319;
  assign n5962 = pi12 ? n26 : n5961;
  assign n5963 = pi11 ? n5962 : n4203;
  assign n5964 = pi10 ? n5959 : n5963;
  assign n5965 = pi13 ? n79 : ~n2319;
  assign n5966 = pi12 ? n26 : ~n5965;
  assign n5967 = pi11 ? n4196 : n5966;
  assign n5968 = pi14 ? n1615 : ~n320;
  assign n5969 = pi13 ? n1751 : n5968;
  assign n5970 = pi12 ? n69 : ~n5969;
  assign n5971 = pi14 ? n168 : n44;
  assign n5972 = pi13 ? n5971 : ~n26;
  assign n5973 = pi12 ? n78 : ~n5972;
  assign n5974 = pi11 ? n5970 : n5973;
  assign n5975 = pi10 ? n5967 : n5974;
  assign n5976 = pi09 ? n5964 : n5975;
  assign n5977 = pi08 ? n5955 : n5976;
  assign n5978 = pi07 ? n5943 : n5977;
  assign n5979 = pi06 ? n5940 : n5978;
  assign n5980 = pi13 ? n4222 : n3918;
  assign n5981 = pi12 ? n26 : n5980;
  assign n5982 = pi11 ? n26 : n5981;
  assign n5983 = pi14 ? n1704 : n327;
  assign n5984 = pi13 ? n4226 : n5983;
  assign n5985 = pi12 ? n26 : n5984;
  assign n5986 = pi14 ? n320 : n327;
  assign n5987 = pi13 ? n2319 : n5986;
  assign n5988 = pi12 ? n26 : n5987;
  assign n5989 = pi11 ? n5985 : n5988;
  assign n5990 = pi10 ? n5982 : n5989;
  assign n5991 = pi09 ? n26 : n5990;
  assign n5992 = pi08 ? n26 : n5991;
  assign n5993 = pi13 ? n1280 : n2631;
  assign n5994 = pi12 ? n26 : n5993;
  assign n5995 = pi11 ? n5994 : n5908;
  assign n5996 = pi13 ? n3135 : ~n126;
  assign n5997 = pi12 ? n26 : n5996;
  assign n5998 = pi11 ? n4239 : n5997;
  assign n5999 = pi10 ? n5995 : n5998;
  assign n6000 = pi14 ? n45 : n1355;
  assign n6001 = pi13 ? n4249 : n6000;
  assign n6002 = pi12 ? n26 : n6001;
  assign n6003 = pi11 ? n26 : n6002;
  assign n6004 = pi10 ? n26 : n6003;
  assign n6005 = pi09 ? n5999 : n6004;
  assign n6006 = pi13 ? n4255 : n6000;
  assign n6007 = pi12 ? n26 : n6006;
  assign n6008 = pi13 ? n1347 : n5615;
  assign n6009 = pi12 ? n26 : n6008;
  assign n6010 = pi11 ? n6007 : n6009;
  assign n6011 = pi14 ? n63 : ~n63;
  assign n6012 = pi13 ? n1347 : n6011;
  assign n6013 = pi12 ? n26 : n6012;
  assign n6014 = pi10 ? n6010 : n6013;
  assign n6015 = pi13 ? n1347 : n5244;
  assign n6016 = pi12 ? n26 : n6015;
  assign n6017 = pi13 ? n4167 : n1091;
  assign n6018 = pi12 ? n26 : n6017;
  assign n6019 = pi11 ? n6016 : n6018;
  assign n6020 = pi13 ? n26 : ~n443;
  assign n6021 = pi12 ? n26 : n6020;
  assign n6022 = pi11 ? n6021 : n5935;
  assign n6023 = pi10 ? n6019 : n6022;
  assign n6024 = pi09 ? n6014 : n6023;
  assign n6025 = pi08 ? n6005 : n6024;
  assign n6026 = pi07 ? n5992 : n6025;
  assign n6027 = pi09 ? n6004 : n6014;
  assign n6028 = pi13 ? n4249 : n5808;
  assign n6029 = pi12 ? n26 : n6028;
  assign n6030 = pi11 ? n26 : n6029;
  assign n6031 = pi10 ? n26 : n6030;
  assign n6032 = pi09 ? n6023 : n6031;
  assign n6033 = pi08 ? n6027 : n6032;
  assign n6034 = pi13 ? n4255 : n5808;
  assign n6035 = pi12 ? n26 : n6034;
  assign n6036 = pi14 ? n320 : ~n63;
  assign n6037 = pi13 ? n1344 : n6036;
  assign n6038 = pi12 ? n26 : n6037;
  assign n6039 = pi11 ? n6035 : n6038;
  assign n6040 = pi13 ? n1347 : n6036;
  assign n6041 = pi12 ? n26 : n6040;
  assign n6042 = pi11 ? n6041 : n6038;
  assign n6043 = pi10 ? n6039 : n6042;
  assign n6044 = pi11 ? n6041 : n4939;
  assign n6045 = pi13 ? n4737 : n3066;
  assign n6046 = pi12 ? n26 : n6045;
  assign n6047 = pi11 ? n4299 : n6046;
  assign n6048 = pi10 ? n6044 : n6047;
  assign n6049 = pi09 ? n6043 : n6048;
  assign n6050 = pi13 ? n5037 : n3066;
  assign n6051 = pi12 ? n26 : n6050;
  assign n6052 = pi13 ? n4425 : n2979;
  assign n6053 = pi12 ? n26 : n6052;
  assign n6054 = pi11 ? n6051 : n6053;
  assign n6055 = pi13 ? n4222 : n2319;
  assign n6056 = pi12 ? n26 : n6055;
  assign n6057 = pi15 ? n60 : ~n291;
  assign n6058 = pi14 ? n6057 : ~n29;
  assign n6059 = pi13 ? n6058 : n2319;
  assign n6060 = pi12 ? n26 : n6059;
  assign n6061 = pi11 ? n6056 : n6060;
  assign n6062 = pi10 ? n6054 : n6061;
  assign n6063 = pi14 ? n37 : n61;
  assign n6064 = pi13 ? n3358 : n6063;
  assign n6065 = pi12 ? n26 : n6064;
  assign n6066 = pi14 ? n1437 : n26;
  assign n6067 = pi14 ? n1138 : n61;
  assign n6068 = pi13 ? n6066 : n6067;
  assign n6069 = pi12 ? n26 : n6068;
  assign n6070 = pi11 ? n6065 : n6069;
  assign n6071 = pi14 ? n233 : n320;
  assign n6072 = pi14 ? n1615 : ~n61;
  assign n6073 = pi13 ? n6071 : ~n6072;
  assign n6074 = pi12 ? n124 : n6073;
  assign n6075 = pi14 ? n26 : n442;
  assign n6076 = pi13 ? n26 : n6075;
  assign n6077 = pi12 ? n6076 : ~n4326;
  assign n6078 = pi11 ? n6074 : n6077;
  assign n6079 = pi10 ? n6070 : n6078;
  assign n6080 = pi09 ? n6062 : n6079;
  assign n6081 = pi08 ? n6049 : n6080;
  assign n6082 = pi07 ? n6033 : n6081;
  assign n6083 = pi06 ? n6026 : n6082;
  assign n6084 = pi05 ? n5979 : n6083;
  assign n6085 = pi04 ? n5895 : n6084;
  assign n6086 = pi13 ? n4226 : n3066;
  assign n6087 = pi12 ? n26 : n6086;
  assign n6088 = pi14 ? n37 : n327;
  assign n6089 = pi13 ? n2319 : n6088;
  assign n6090 = pi12 ? n26 : n6089;
  assign n6091 = pi11 ? n6087 : n6090;
  assign n6092 = pi10 ? n4860 : n6091;
  assign n6093 = pi09 ? n26 : n6092;
  assign n6094 = pi08 ? n26 : n6093;
  assign n6095 = pi13 ? n1280 : ~n4348;
  assign n6096 = pi12 ? n26 : n6095;
  assign n6097 = pi13 ? n2387 : ~n4442;
  assign n6098 = pi12 ? n26 : n6097;
  assign n6099 = pi11 ? n6096 : n6098;
  assign n6100 = pi13 ? n321 : ~n4153;
  assign n6101 = pi12 ? n26 : n6100;
  assign n6102 = pi11 ? n4239 : n6101;
  assign n6103 = pi10 ? n6099 : n6102;
  assign n6104 = pi13 ? n1280 : n1850;
  assign n6105 = pi12 ? n26 : n6104;
  assign n6106 = pi11 ? n26 : n6105;
  assign n6107 = pi10 ? n26 : n6106;
  assign n6108 = pi09 ? n6103 : n6107;
  assign n6109 = pi14 ? n63 : ~n125;
  assign n6110 = pi13 ? n1280 : n6109;
  assign n6111 = pi12 ? n26 : n6110;
  assign n6112 = pi11 ? n6111 : n6105;
  assign n6113 = pi10 ? n6112 : n4377;
  assign n6114 = pi13 ? n1280 : n3980;
  assign n6115 = pi12 ? n26 : n6114;
  assign n6116 = pi13 ? n198 : n3888;
  assign n6117 = pi12 ? n26 : n6116;
  assign n6118 = pi11 ? n6115 : n6117;
  assign n6119 = pi11 ? n4149 : n5935;
  assign n6120 = pi10 ? n6118 : n6119;
  assign n6121 = pi09 ? n6113 : n6120;
  assign n6122 = pi08 ? n6108 : n6121;
  assign n6123 = pi07 ? n6094 : n6122;
  assign n6124 = pi09 ? n6107 : n6113;
  assign n6125 = pi13 ? n1280 : n5690;
  assign n6126 = pi12 ? n26 : n6125;
  assign n6127 = pi11 ? n26 : n6126;
  assign n6128 = pi10 ? n26 : n6127;
  assign n6129 = pi09 ? n6120 : n6128;
  assign n6130 = pi08 ? n6124 : n6129;
  assign n6131 = pi13 ? n2598 : n5690;
  assign n6132 = pi12 ? n26 : n6131;
  assign n6133 = pi11 ? n6126 : n6132;
  assign n6134 = pi13 ? n5438 : n5690;
  assign n6135 = pi12 ? n26 : n6134;
  assign n6136 = pi11 ? n6126 : n6135;
  assign n6137 = pi10 ? n6133 : n6136;
  assign n6138 = pi13 ? n2319 : n5690;
  assign n6139 = pi12 ? n26 : n6138;
  assign n6140 = pi14 ? n2174 : n26;
  assign n6141 = pi13 ? n6140 : n5690;
  assign n6142 = pi12 ? n26 : n6141;
  assign n6143 = pi11 ? n6139 : n6142;
  assign n6144 = pi14 ? n320 : ~n4140;
  assign n6145 = pi13 ? n2370 : n6144;
  assign n6146 = pi12 ? n26 : n6145;
  assign n6147 = pi13 ? n2370 : n5690;
  assign n6148 = pi12 ? n26 : n6147;
  assign n6149 = pi11 ? n6146 : n6148;
  assign n6150 = pi10 ? n6143 : n6149;
  assign n6151 = pi09 ? n6137 : n6150;
  assign n6152 = pi13 ? n2370 : n2979;
  assign n6153 = pi12 ? n26 : n6152;
  assign n6154 = pi13 ? n2370 : n2319;
  assign n6155 = pi12 ? n26 : n6154;
  assign n6156 = pi11 ? n6153 : n6155;
  assign n6157 = pi13 ? n1135 : n2319;
  assign n6158 = pi12 ? n26 : n6157;
  assign n6159 = pi11 ? n6158 : n4408;
  assign n6160 = pi10 ? n6156 : n6159;
  assign n6161 = pi13 ? n1135 : n639;
  assign n6162 = pi12 ? n26 : n6161;
  assign n6163 = pi15 ? n291 : ~n70;
  assign n6164 = pi14 ? n6163 : n26;
  assign n6165 = pi13 ? n57 : ~n6164;
  assign n6166 = pi12 ? n26 : ~n6165;
  assign n6167 = pi11 ? n6162 : n6166;
  assign n6168 = pi13 ? n1751 : n72;
  assign n6169 = pi12 ? n69 : ~n6168;
  assign n6170 = pi12 ? n6076 : n5467;
  assign n6171 = pi11 ? n6169 : n6170;
  assign n6172 = pi10 ? n6167 : n6171;
  assign n6173 = pi09 ? n6160 : n6172;
  assign n6174 = pi08 ? n6151 : n6173;
  assign n6175 = pi07 ? n6130 : n6174;
  assign n6176 = pi06 ? n6123 : n6175;
  assign n6177 = pi13 ? n3888 : n3782;
  assign n6178 = pi12 ? n26 : n6177;
  assign n6179 = pi11 ? n26 : n6178;
  assign n6180 = pi13 ? n2370 : n5899;
  assign n6181 = pi12 ? n26 : n6180;
  assign n6182 = pi13 ? n2319 : n639;
  assign n6183 = pi12 ? n26 : n6182;
  assign n6184 = pi11 ? n6181 : n6183;
  assign n6185 = pi10 ? n6179 : n6184;
  assign n6186 = pi09 ? n26 : n6185;
  assign n6187 = pi08 ? n26 : n6186;
  assign n6188 = pi13 ? n2319 : ~n4348;
  assign n6189 = pi12 ? n26 : n6188;
  assign n6190 = pi13 ? n2522 : ~n4442;
  assign n6191 = pi12 ? n26 : n6190;
  assign n6192 = pi11 ? n6189 : n6191;
  assign n6193 = pi11 ? n4239 : n5935;
  assign n6194 = pi10 ? n6192 : n6193;
  assign n6195 = pi09 ? n6194 : n26;
  assign n6196 = pi08 ? n6195 : n26;
  assign n6197 = pi07 ? n6187 : n6196;
  assign n6198 = pi06 ? n6197 : n26;
  assign n6199 = pi05 ? n6176 : n6198;
  assign n6200 = pi13 ? n1135 : n5986;
  assign n6201 = pi12 ? n26 : n6200;
  assign n6202 = pi11 ? n6155 : n6201;
  assign n6203 = pi10 ? n6179 : n6202;
  assign n6204 = pi09 ? n26 : n6203;
  assign n6205 = pi08 ? n26 : n6204;
  assign n6206 = pi13 ? n1135 : ~n4348;
  assign n6207 = pi12 ? n26 : n6206;
  assign n6208 = pi14 ? n147 : n320;
  assign n6209 = pi13 ? n6208 : ~n38;
  assign n6210 = pi12 ? n26 : n6209;
  assign n6211 = pi11 ? n6207 : n6210;
  assign n6212 = pi13 ? n507 : n38;
  assign n6213 = pi12 ? n26 : ~n6212;
  assign n6214 = pi11 ? n6213 : n5935;
  assign n6215 = pi10 ? n6211 : n6214;
  assign n6216 = pi09 ? n6215 : n26;
  assign n6217 = pi08 ? n6216 : n26;
  assign n6218 = pi07 ? n6205 : n6217;
  assign n6219 = pi06 ? n6218 : n26;
  assign n6220 = pi13 ? n3980 : n3782;
  assign n6221 = pi12 ? n26 : n6220;
  assign n6222 = pi11 ? n26 : n6221;
  assign n6223 = pi13 ? n1135 : n2631;
  assign n6224 = pi12 ? n26 : n6223;
  assign n6225 = pi11 ? n5368 : n6224;
  assign n6226 = pi10 ? n6222 : n6225;
  assign n6227 = pi09 ? n26 : n6226;
  assign n6228 = pi08 ? n26 : n6227;
  assign n6229 = pi13 ? n478 : ~n38;
  assign n6230 = pi12 ? n26 : n6229;
  assign n6231 = pi11 ? n6230 : n5935;
  assign n6232 = pi10 ? n6211 : n6231;
  assign n6233 = pi14 ? n26 : ~n44;
  assign n6234 = pi13 ? n6233 : n1850;
  assign n6235 = pi12 ? n26 : n6234;
  assign n6236 = pi13 ? n5690 : n2598;
  assign n6237 = pi12 ? n26 : n6236;
  assign n6238 = pi11 ? n6235 : n6237;
  assign n6239 = pi13 ? n5690 : n2631;
  assign n6240 = pi12 ? n26 : n6239;
  assign n6241 = pi13 ? n5690 : n26;
  assign n6242 = pi12 ? n26 : n6241;
  assign n6243 = pi11 ? n6240 : n6242;
  assign n6244 = pi10 ? n6238 : n6243;
  assign n6245 = pi09 ? n6232 : n6244;
  assign n6246 = pi08 ? n6245 : n6242;
  assign n6247 = pi07 ? n6228 : n6246;
  assign n6248 = pi06 ? n6247 : n6242;
  assign n6249 = pi05 ? n6219 : n6248;
  assign n6250 = pi04 ? n6199 : n6249;
  assign n6251 = pi03 ? n6085 : n6250;
  assign n6252 = pi15 ? n28 : ~n70;
  assign n6253 = pi14 ? n6252 : n26;
  assign n6254 = pi13 ? n1135 : n6253;
  assign n6255 = pi12 ? n26 : n6254;
  assign n6256 = pi11 ? n5368 : n6255;
  assign n6257 = pi10 ? n6222 : n6256;
  assign n6258 = pi09 ? n26 : n6257;
  assign n6259 = pi08 ? n26 : n6258;
  assign n6260 = pi14 ? n152 : n320;
  assign n6261 = pi13 ? n6260 : ~n38;
  assign n6262 = pi12 ? n26 : n6261;
  assign n6263 = pi11 ? n4478 : n6262;
  assign n6264 = pi13 ? n591 : ~n38;
  assign n6265 = pi12 ? n26 : n6264;
  assign n6266 = pi11 ? n6265 : n5935;
  assign n6267 = pi10 ? n6263 : n6266;
  assign n6268 = pi14 ? n26 : ~n3250;
  assign n6269 = pi13 ? n6268 : n2498;
  assign n6270 = pi12 ? n26 : n6269;
  assign n6271 = pi13 ? n5886 : n26;
  assign n6272 = pi12 ? n26 : n6271;
  assign n6273 = pi11 ? n6270 : n6272;
  assign n6274 = pi13 ? n4125 : n2347;
  assign n6275 = pi12 ? n26 : n6274;
  assign n6276 = pi11 ? n6275 : n5293;
  assign n6277 = pi10 ? n6273 : n6276;
  assign n6278 = pi09 ? n6267 : n6277;
  assign n6279 = pi08 ? n6278 : n4535;
  assign n6280 = pi07 ? n6259 : n6279;
  assign n6281 = pi06 ? n6280 : n4546;
  assign n6282 = pi13 ? n869 : n3782;
  assign n6283 = pi12 ? n26 : n6282;
  assign n6284 = pi11 ? n26 : n6283;
  assign n6285 = pi13 ? n630 : n6253;
  assign n6286 = pi12 ? n26 : n6285;
  assign n6287 = pi11 ? n5370 : n6286;
  assign n6288 = pi10 ? n6284 : n6287;
  assign n6289 = pi09 ? n26 : n6288;
  assign n6290 = pi08 ? n26 : n6289;
  assign n6291 = pi13 ? n1982 : n38;
  assign n6292 = pi12 ? n26 : ~n6291;
  assign n6293 = pi11 ? n4414 : n6292;
  assign n6294 = pi12 ? n124 : n4879;
  assign n6295 = pi11 ? n6294 : n5935;
  assign n6296 = pi10 ? n6293 : n6295;
  assign n6297 = pi14 ? n168 : n233;
  assign n6298 = pi13 ? n6297 : n126;
  assign n6299 = pi12 ? n78 : ~n6298;
  assign n6300 = pi13 ? n351 : ~n126;
  assign n6301 = pi12 ? n78 : n6300;
  assign n6302 = pi11 ? n6299 : n6301;
  assign n6303 = pi14 ? n168 : ~n37;
  assign n6304 = pi14 ? n517 : ~n168;
  assign n6305 = pi13 ? n6303 : ~n6304;
  assign n6306 = pi12 ? n78 : ~n6305;
  assign n6307 = pi13 ? n176 : n2762;
  assign n6308 = pi12 ? n78 : n6307;
  assign n6309 = pi11 ? n6306 : n6308;
  assign n6310 = pi10 ? n6302 : n6309;
  assign n6311 = pi09 ? n6296 : n6310;
  assign n6312 = pi13 ? n176 : n26;
  assign n6313 = pi12 ? n78 : n6312;
  assign n6314 = pi11 ? n6313 : n5342;
  assign n6315 = pi10 ? n6314 : n4581;
  assign n6316 = pi09 ? n6315 : n4581;
  assign n6317 = pi08 ? n6311 : n6316;
  assign n6318 = pi07 ? n6290 : n6317;
  assign n6319 = pi06 ? n6318 : n4589;
  assign n6320 = pi05 ? n6281 : n6319;
  assign n6321 = pi11 ? n26 : n5370;
  assign n6322 = pi11 ? n5370 : n6255;
  assign n6323 = pi10 ? n6321 : n6322;
  assign n6324 = pi09 ? n26 : n6323;
  assign n6325 = pi08 ? n26 : n6324;
  assign n6326 = pi13 ? n1982 : n72;
  assign n6327 = pi12 ? n26 : ~n6326;
  assign n6328 = pi11 ? n4414 : n6327;
  assign n6329 = pi13 ? n79 : n72;
  assign n6330 = pi12 ? n124 : ~n6329;
  assign n6331 = pi11 ? n6330 : n6169;
  assign n6332 = pi10 ? n6328 : n6331;
  assign n6333 = pi14 ? n29 : n233;
  assign n6334 = pi14 ? n71 : n168;
  assign n6335 = pi13 ? n6333 : n6334;
  assign n6336 = pi12 ? n78 : ~n6335;
  assign n6337 = pi10 ? n4603 : n6336;
  assign n6338 = pi09 ? n6332 : n6337;
  assign n6339 = pi13 ? n6333 : n72;
  assign n6340 = pi12 ? n78 : ~n6339;
  assign n6341 = pi08 ? n6338 : n6340;
  assign n6342 = pi07 ? n6325 : n6341;
  assign n6343 = pi12 ? n69 : ~n6298;
  assign n6344 = pi11 ? n6340 : n6343;
  assign n6345 = pi13 ? n6297 : ~n26;
  assign n6346 = pi12 ? n78 : ~n6345;
  assign n6347 = pi10 ? n6344 : n6346;
  assign n6348 = pi09 ? n6340 : n6347;
  assign n6349 = pi08 ? n6340 : n6348;
  assign n6350 = pi07 ? n6340 : n6349;
  assign n6351 = pi06 ? n6342 : n6350;
  assign n6352 = pi14 ? n45 : ~n786;
  assign n6353 = pi13 ? n6352 : n169;
  assign n6354 = pi12 ? n78 : ~n6353;
  assign n6355 = pi11 ? n26 : n6354;
  assign n6356 = pi10 ? n26 : n6355;
  assign n6357 = pi13 ? n6352 : n57;
  assign n6358 = pi12 ? n78 : ~n6357;
  assign n6359 = pi11 ? n6358 : n4630;
  assign n6360 = pi11 ? n5042 : n6346;
  assign n6361 = pi10 ? n6359 : n6360;
  assign n6362 = pi09 ? n6356 : n6361;
  assign n6363 = pi08 ? n26 : n6362;
  assign n6364 = pi07 ? n26 : n6363;
  assign n6365 = pi06 ? n26 : n6364;
  assign n6366 = pi05 ? n6351 : n6365;
  assign n6367 = pi04 ? n6320 : n6366;
  assign n6368 = pi14 ? n1437 : ~n125;
  assign n6369 = pi13 ? n6368 : n4471;
  assign n6370 = pi12 ? n26 : n6369;
  assign n6371 = pi11 ? n26 : n6370;
  assign n6372 = pi10 ? n26 : n6371;
  assign n6373 = pi14 ? n292 : ~n1638;
  assign n6374 = pi13 ? n6373 : n130;
  assign n6375 = pi12 ? n69 : ~n6374;
  assign n6376 = pi14 ? n1400 : ~n37;
  assign n6377 = pi13 ? n6376 : n704;
  assign n6378 = pi12 ? n78 : ~n6377;
  assign n6379 = pi11 ? n6375 : n6378;
  assign n6380 = pi13 ? n1344 : n126;
  assign n6381 = pi12 ? n78 : ~n6380;
  assign n6382 = pi14 ? n168 : ~n786;
  assign n6383 = pi13 ? n6382 : n126;
  assign n6384 = pi12 ? n6076 : ~n6383;
  assign n6385 = pi11 ? n6381 : n6384;
  assign n6386 = pi10 ? n6379 : n6385;
  assign n6387 = pi09 ? n6372 : n6386;
  assign n6388 = pi08 ? n26 : n6387;
  assign n6389 = pi07 ? n26 : n6388;
  assign n6390 = pi06 ? n26 : n6389;
  assign n6391 = pi13 ? n130 : n284;
  assign n6392 = pi12 ? n26 : n6391;
  assign n6393 = pi11 ? n26 : n6392;
  assign n6394 = pi13 ? n130 : ~n5545;
  assign n6395 = pi12 ? n26 : n6394;
  assign n6396 = pi10 ? n6393 : n6395;
  assign n6397 = pi09 ? n26 : n6396;
  assign n6398 = pi08 ? n26 : n6397;
  assign n6399 = pi13 ? n169 : ~n5545;
  assign n6400 = pi12 ? n26 : n6399;
  assign n6401 = pi11 ? n6395 : n6400;
  assign n6402 = pi10 ? n6395 : n6401;
  assign n6403 = pi11 ? n6400 : n6395;
  assign n6404 = pi10 ? n6403 : n6395;
  assign n6405 = pi09 ? n6402 : n6404;
  assign n6406 = pi08 ? n6395 : n6405;
  assign n6407 = pi07 ? n6398 : n6406;
  assign n6408 = pi14 ? n131 : ~n1704;
  assign n6409 = pi13 ? n176 : ~n6408;
  assign n6410 = pi12 ? n26 : n6409;
  assign n6411 = pi11 ? n6395 : n6410;
  assign n6412 = pi10 ? n6395 : n6411;
  assign n6413 = pi09 ? n6395 : n6412;
  assign n6414 = pi14 ? n131 : ~n320;
  assign n6415 = pi13 ? n176 : ~n6414;
  assign n6416 = pi12 ? n26 : n6415;
  assign n6417 = pi14 ? n147 : ~n6252;
  assign n6418 = pi13 ? n1438 : ~n6417;
  assign n6419 = pi12 ? n26 : n6418;
  assign n6420 = pi11 ? n6416 : n6419;
  assign n6421 = pi14 ? n1638 : ~n45;
  assign n6422 = pi13 ? n6421 : n3918;
  assign n6423 = pi12 ? n26 : n6422;
  assign n6424 = pi14 ? n1872 : ~n125;
  assign n6425 = pi13 ? n6424 : n1091;
  assign n6426 = pi12 ? n26 : n6425;
  assign n6427 = pi11 ? n6423 : n6426;
  assign n6428 = pi10 ? n6420 : n6427;
  assign n6429 = pi14 ? n61 : ~n2954;
  assign n6430 = pi13 ? n6429 : n176;
  assign n6431 = pi12 ? n69 : ~n6430;
  assign n6432 = pi13 ? n3829 : n736;
  assign n6433 = pi12 ? n69 : ~n6432;
  assign n6434 = pi11 ? n6431 : n6433;
  assign n6435 = pi13 ? n6303 : n126;
  assign n6436 = pi12 ? n124 : ~n6435;
  assign n6437 = pi11 ? n4968 : n6436;
  assign n6438 = pi10 ? n6434 : n6437;
  assign n6439 = pi09 ? n6428 : n6438;
  assign n6440 = pi08 ? n6413 : n6439;
  assign n6441 = pi07 ? n6395 : n6440;
  assign n6442 = pi06 ? n6407 : n6441;
  assign n6443 = pi05 ? n6390 : n6442;
  assign n6444 = pi13 ? n240 : n1567;
  assign n6445 = pi12 ? n26 : n6444;
  assign n6446 = pi11 ? n26 : n6445;
  assign n6447 = pi10 ? n6446 : n6445;
  assign n6448 = pi09 ? n26 : n6447;
  assign n6449 = pi08 ? n26 : n6448;
  assign n6450 = pi14 ? n63 : ~n61;
  assign n6451 = pi13 ? n6450 : n1567;
  assign n6452 = pi12 ? n26 : n6451;
  assign n6453 = pi11 ? n6452 : n6445;
  assign n6454 = pi10 ? n6445 : n6453;
  assign n6455 = pi09 ? n6454 : n6445;
  assign n6456 = pi08 ? n6445 : n6455;
  assign n6457 = pi07 ? n6449 : n6456;
  assign n6458 = pi11 ? n6445 : n5606;
  assign n6459 = pi13 ? n79 : n1567;
  assign n6460 = pi12 ? n26 : n6459;
  assign n6461 = pi13 ? n57 : n5615;
  assign n6462 = pi12 ? n26 : n6461;
  assign n6463 = pi11 ? n6460 : n6462;
  assign n6464 = pi10 ? n6458 : n6463;
  assign n6465 = pi09 ? n6445 : n6464;
  assign n6466 = pi14 ? n45 : n147;
  assign n6467 = pi13 ? n57 : n6466;
  assign n6468 = pi12 ? n26 : n6467;
  assign n6469 = pi13 ? n38 : n4622;
  assign n6470 = pi12 ? n26 : n6469;
  assign n6471 = pi11 ? n6468 : n6470;
  assign n6472 = pi13 ? n4471 : n1091;
  assign n6473 = pi12 ? n26 : n6472;
  assign n6474 = pi11 ? n4115 : n6473;
  assign n6475 = pi10 ? n6471 : n6474;
  assign n6476 = pi13 ? n584 : n57;
  assign n6477 = pi12 ? n69 : ~n6476;
  assign n6478 = pi12 ? n654 : ~n57;
  assign n6479 = pi11 ? n6477 : n6478;
  assign n6480 = pi13 ? n1751 : n38;
  assign n6481 = pi12 ? n26 : ~n6480;
  assign n6482 = pi12 ? n124 : n5934;
  assign n6483 = pi11 ? n6481 : n6482;
  assign n6484 = pi10 ? n6479 : n6483;
  assign n6485 = pi09 ? n6475 : n6484;
  assign n6486 = pi08 ? n6465 : n6485;
  assign n6487 = pi07 ? n6445 : n6486;
  assign n6488 = pi06 ? n6457 : n6487;
  assign n6489 = pi13 ? n4737 : n4809;
  assign n6490 = pi12 ? n26 : n6489;
  assign n6491 = pi11 ? n26 : n6490;
  assign n6492 = pi13 ? n4741 : n4809;
  assign n6493 = pi12 ? n26 : n6492;
  assign n6494 = pi10 ? n6491 : n6493;
  assign n6495 = pi09 ? n26 : n6494;
  assign n6496 = pi08 ? n26 : n6495;
  assign n6497 = pi13 ? n4119 : n6000;
  assign n6498 = pi12 ? n26 : n6497;
  assign n6499 = pi11 ? n6493 : n6498;
  assign n6500 = pi10 ? n6493 : n6499;
  assign n6501 = pi13 ? n1344 : n6000;
  assign n6502 = pi12 ? n26 : n6501;
  assign n6503 = pi13 ? n4753 : n6000;
  assign n6504 = pi12 ? n26 : n6503;
  assign n6505 = pi11 ? n6502 : n6504;
  assign n6506 = pi14 ? n45 : n44;
  assign n6507 = pi13 ? n1344 : n6506;
  assign n6508 = pi12 ? n26 : n6507;
  assign n6509 = pi13 ? n4741 : n6506;
  assign n6510 = pi12 ? n26 : n6509;
  assign n6511 = pi11 ? n6508 : n6510;
  assign n6512 = pi10 ? n6505 : n6511;
  assign n6513 = pi09 ? n6500 : n6512;
  assign n6514 = pi08 ? n6493 : n6513;
  assign n6515 = pi07 ? n6496 : n6514;
  assign n6516 = pi13 ? n4255 : n4809;
  assign n6517 = pi12 ? n26 : n6516;
  assign n6518 = pi11 ? n6493 : n6517;
  assign n6519 = pi13 ? n4769 : n3918;
  assign n6520 = pi12 ? n26 : n6519;
  assign n6521 = pi13 ? n4255 : n3996;
  assign n6522 = pi12 ? n26 : n6521;
  assign n6523 = pi11 ? n6520 : n6522;
  assign n6524 = pi10 ? n6518 : n6523;
  assign n6525 = pi09 ? n6493 : n6524;
  assign n6526 = pi13 ? n4943 : n3918;
  assign n6527 = pi12 ? n26 : n6526;
  assign n6528 = pi13 ? n4943 : n6352;
  assign n6529 = pi12 ? n26 : n6528;
  assign n6530 = pi11 ? n6527 : n6529;
  assign n6531 = pi14 ? n2420 : ~n29;
  assign n6532 = pi13 ? n6531 : n3918;
  assign n6533 = pi12 ? n26 : n6532;
  assign n6534 = pi13 ? n3980 : n4716;
  assign n6535 = pi12 ? n26 : n6534;
  assign n6536 = pi11 ? n6533 : n6535;
  assign n6537 = pi10 ? n6530 : n6536;
  assign n6538 = pi13 ? n57 : ~n1135;
  assign n6539 = pi12 ? n26 : ~n6538;
  assign n6540 = pi14 ? n4140 : n26;
  assign n6541 = pi13 ? n544 : ~n6540;
  assign n6542 = pi12 ? n26 : ~n6541;
  assign n6543 = pi11 ? n6539 : n6542;
  assign n6544 = pi13 ? n6071 : ~n72;
  assign n6545 = pi12 ? n26 : n6544;
  assign n6546 = pi14 ? n168 : ~n320;
  assign n6547 = pi13 ? n6546 : n126;
  assign n6548 = pi12 ? n124 : ~n6547;
  assign n6549 = pi11 ? n6545 : n6548;
  assign n6550 = pi10 ? n6543 : n6549;
  assign n6551 = pi09 ? n6537 : n6550;
  assign n6552 = pi08 ? n6525 : n6551;
  assign n6553 = pi07 ? n6493 : n6552;
  assign n6554 = pi06 ? n6515 : n6553;
  assign n6555 = pi05 ? n6488 : n6554;
  assign n6556 = pi04 ? n6443 : n6555;
  assign n6557 = pi03 ? n6367 : n6556;
  assign n6558 = pi02 ? n6251 : n6557;
  assign n6559 = pi01 ? n5758 : n6558;
  assign n6560 = pi11 ? n26 : n6132;
  assign n6561 = pi10 ? n6560 : n6132;
  assign n6562 = pi09 ? n26 : n6561;
  assign n6563 = pi08 ? n26 : n6562;
  assign n6564 = pi11 ? n6135 : n6132;
  assign n6565 = pi10 ? n6132 : n6564;
  assign n6566 = pi13 ? n4135 : n3061;
  assign n6567 = pi12 ? n26 : n6566;
  assign n6568 = pi13 ? n4809 : n3061;
  assign n6569 = pi12 ? n26 : n6568;
  assign n6570 = pi11 ? n6569 : n6132;
  assign n6571 = pi10 ? n6567 : n6570;
  assign n6572 = pi09 ? n6565 : n6571;
  assign n6573 = pi08 ? n6132 : n6572;
  assign n6574 = pi07 ? n6563 : n6573;
  assign n6575 = pi13 ? n2598 : n1850;
  assign n6576 = pi12 ? n26 : n6575;
  assign n6577 = pi11 ? n6576 : n6111;
  assign n6578 = pi13 ? n2955 : n5690;
  assign n6579 = pi12 ? n26 : n6578;
  assign n6580 = pi11 ? n6579 : n6135;
  assign n6581 = pi10 ? n6577 : n6580;
  assign n6582 = pi09 ? n6132 : n6581;
  assign n6583 = pi14 ? n1638 : n26;
  assign n6584 = pi13 ? n6583 : n3066;
  assign n6585 = pi12 ? n26 : n6584;
  assign n6586 = pi15 ? n27 : ~n291;
  assign n6587 = pi14 ? n6586 : n26;
  assign n6588 = pi13 ? n6587 : n3066;
  assign n6589 = pi12 ? n26 : n6588;
  assign n6590 = pi13 ? n1135 : n1705;
  assign n6591 = pi12 ? n26 : n6590;
  assign n6592 = pi11 ? n6589 : n6591;
  assign n6593 = pi10 ? n6585 : n6592;
  assign n6594 = pi13 ? n584 : ~n591;
  assign n6595 = pi12 ? n124 : ~n6594;
  assign n6596 = pi14 ? n1355 : n26;
  assign n6597 = pi13 ? n57 : ~n6596;
  assign n6598 = pi12 ? n69 : ~n6597;
  assign n6599 = pi11 ? n6595 : n6598;
  assign n6600 = pi12 ? n654 : ~n6168;
  assign n6601 = pi12 ? n69 : n5934;
  assign n6602 = pi11 ? n6600 : n6601;
  assign n6603 = pi10 ? n6599 : n6602;
  assign n6604 = pi09 ? n6593 : n6603;
  assign n6605 = pi08 ? n6582 : n6604;
  assign n6606 = pi07 ? n6132 : n6605;
  assign n6607 = pi06 ? n6574 : n6606;
  assign n6608 = pi11 ? n26 : n5390;
  assign n6609 = pi13 ? n639 : n2319;
  assign n6610 = pi12 ? n26 : n6609;
  assign n6611 = pi13 ? n639 : n1705;
  assign n6612 = pi12 ? n26 : n6611;
  assign n6613 = pi11 ? n6610 : n6612;
  assign n6614 = pi10 ? n6608 : n6613;
  assign n6615 = pi09 ? n26 : n6614;
  assign n6616 = pi08 ? n26 : n6615;
  assign n6617 = pi07 ? n26 : n6616;
  assign n6618 = pi11 ? n2341 : n26;
  assign n6619 = pi10 ? n6618 : n26;
  assign n6620 = pi09 ? n6619 : n26;
  assign n6621 = pi08 ? n6620 : n26;
  assign n6622 = pi07 ? n6621 : n26;
  assign n6623 = pi06 ? n6617 : n6622;
  assign n6624 = pi05 ? n6607 : n6623;
  assign n6625 = pi13 ? n4222 : n5777;
  assign n6626 = pi12 ? n26 : n6625;
  assign n6627 = pi11 ? n26 : n6626;
  assign n6628 = pi13 ? n639 : n2631;
  assign n6629 = pi12 ? n26 : n6628;
  assign n6630 = pi11 ? n6610 : n6629;
  assign n6631 = pi10 ? n6627 : n6630;
  assign n6632 = pi09 ? n26 : n6631;
  assign n6633 = pi08 ? n26 : n6632;
  assign n6634 = pi07 ? n26 : n6633;
  assign n6635 = pi14 ? n125 : ~n327;
  assign n6636 = pi13 ? n321 : ~n6635;
  assign n6637 = pi12 ? n26 : n6636;
  assign n6638 = pi11 ? n6637 : n26;
  assign n6639 = pi10 ? n6638 : n26;
  assign n6640 = pi09 ? n6639 : n26;
  assign n6641 = pi08 ? n6640 : n26;
  assign n6642 = pi07 ? n6641 : n26;
  assign n6643 = pi06 ? n6634 : n6642;
  assign n6644 = pi14 ? n147 : ~n37;
  assign n6645 = pi13 ? n130 : ~n6644;
  assign n6646 = pi12 ? n26 : n6645;
  assign n6647 = pi10 ? n6393 : n6646;
  assign n6648 = pi09 ? n26 : n6647;
  assign n6649 = pi08 ? n26 : n6648;
  assign n6650 = pi11 ? n6646 : n5542;
  assign n6651 = pi13 ? n176 : ~n5921;
  assign n6652 = pi12 ? n26 : n6651;
  assign n6653 = pi14 ? n147 : ~n125;
  assign n6654 = pi13 ? n1438 : ~n6653;
  assign n6655 = pi12 ? n26 : n6654;
  assign n6656 = pi11 ? n6652 : n6655;
  assign n6657 = pi10 ? n6650 : n6656;
  assign n6658 = pi13 ? n4106 : n79;
  assign n6659 = pi12 ? n26 : n6658;
  assign n6660 = pi13 ? n4425 : n3782;
  assign n6661 = pi12 ? n26 : n6660;
  assign n6662 = pi11 ? n6659 : n6661;
  assign n6663 = pi13 ? n639 : n478;
  assign n6664 = pi12 ? n26 : n6663;
  assign n6665 = pi11 ? n6155 : n6664;
  assign n6666 = pi10 ? n6662 : n6665;
  assign n6667 = pi09 ? n6657 : n6666;
  assign n6668 = pi08 ? n6646 : n6667;
  assign n6669 = pi07 ? n6649 : n6668;
  assign n6670 = pi13 ? n6233 : n3942;
  assign n6671 = pi12 ? n26 : n6670;
  assign n6672 = pi11 ? n6637 : n6671;
  assign n6673 = pi13 ? n5690 : n6583;
  assign n6674 = pi12 ? n26 : n6673;
  assign n6675 = pi11 ? n6674 : n6240;
  assign n6676 = pi10 ? n6672 : n6675;
  assign n6677 = pi09 ? n6676 : n6242;
  assign n6678 = pi08 ? n6677 : n6242;
  assign n6679 = pi07 ? n6678 : n6242;
  assign n6680 = pi06 ? n6669 : n6679;
  assign n6681 = pi05 ? n6643 : n6680;
  assign n6682 = pi04 ? n6624 : n6681;
  assign n6683 = pi12 ? n26 : n79;
  assign n6684 = pi11 ? n3844 : n6683;
  assign n6685 = pi12 ? n26 : n4824;
  assign n6686 = pi13 ? n79 : n240;
  assign n6687 = pi12 ? n26 : n6686;
  assign n6688 = pi11 ? n6685 : n6687;
  assign n6689 = pi10 ? n6684 : n6688;
  assign n6690 = pi13 ? n1252 : n79;
  assign n6691 = pi12 ? n26 : n6690;
  assign n6692 = pi11 ? n6691 : n6661;
  assign n6693 = pi13 ? n2759 : ~n4442;
  assign n6694 = pi12 ? n26 : n6693;
  assign n6695 = pi11 ? n4430 : n6694;
  assign n6696 = pi10 ? n6692 : n6695;
  assign n6697 = pi09 ? n6689 : n6696;
  assign n6698 = pi08 ? n6445 : n6697;
  assign n6699 = pi07 ? n6449 : n6698;
  assign n6700 = pi13 ? n6268 : n2476;
  assign n6701 = pi12 ? n26 : n6700;
  assign n6702 = pi11 ? n5935 : n6701;
  assign n6703 = pi11 ? n6272 : n4921;
  assign n6704 = pi10 ? n6702 : n6703;
  assign n6705 = pi09 ? n6704 : n4535;
  assign n6706 = pi08 ? n6705 : n4535;
  assign n6707 = pi07 ? n6706 : n4545;
  assign n6708 = pi06 ? n6699 : n6707;
  assign n6709 = pi13 ? n4769 : n1583;
  assign n6710 = pi12 ? n26 : n6709;
  assign n6711 = pi11 ? n6517 : n6710;
  assign n6712 = pi13 ? n4255 : n3918;
  assign n6713 = pi12 ? n26 : n6712;
  assign n6714 = pi11 ? n6713 : n6520;
  assign n6715 = pi10 ? n6711 : n6714;
  assign n6716 = pi14 ? n249 : n26;
  assign n6717 = pi13 ? n3181 : n6716;
  assign n6718 = pi12 ? n26 : n6717;
  assign n6719 = pi11 ? n6718 : n6162;
  assign n6720 = pi14 ? n125 : n2386;
  assign n6721 = pi13 ? n6720 : ~n4229;
  assign n6722 = pi12 ? n26 : n6721;
  assign n6723 = pi13 ? n1135 : ~n38;
  assign n6724 = pi12 ? n26 : n6723;
  assign n6725 = pi11 ? n6722 : n6724;
  assign n6726 = pi10 ? n6719 : n6725;
  assign n6727 = pi09 ? n6715 : n6726;
  assign n6728 = pi08 ? n6493 : n6727;
  assign n6729 = pi07 ? n6496 : n6728;
  assign n6730 = pi13 ? n351 : n26;
  assign n6731 = pi12 ? n26 : n6730;
  assign n6732 = pi13 ? n351 : n6304;
  assign n6733 = pi12 ? n26 : n6732;
  assign n6734 = pi11 ? n6731 : n6733;
  assign n6735 = pi10 ? n4968 : n6734;
  assign n6736 = pi12 ? n124 : n4575;
  assign n6737 = pi14 ? n2386 : ~n26;
  assign n6738 = pi13 ? n6737 : n26;
  assign n6739 = pi12 ? n69 : n6738;
  assign n6740 = pi11 ? n6736 : n6739;
  assign n6741 = pi13 ? n415 : n26;
  assign n6742 = pi12 ? n78 : n6741;
  assign n6743 = pi10 ? n6740 : n6742;
  assign n6744 = pi09 ? n6735 : n6743;
  assign n6745 = pi08 ? n6744 : n6742;
  assign n6746 = pi12 ? n69 : n6741;
  assign n6747 = pi13 ? n5808 : n26;
  assign n6748 = pi12 ? n69 : n6747;
  assign n6749 = pi10 ? n6746 : n6748;
  assign n6750 = pi09 ? n6742 : n6749;
  assign n6751 = pi08 ? n6742 : n6750;
  assign n6752 = pi07 ? n6745 : n6751;
  assign n6753 = pi06 ? n6729 : n6752;
  assign n6754 = pi05 ? n6708 : n6753;
  assign n6755 = pi13 ? n198 : n1850;
  assign n6756 = pi12 ? n26 : n6755;
  assign n6757 = pi13 ? n5438 : n1850;
  assign n6758 = pi12 ? n26 : n6757;
  assign n6759 = pi11 ? n6756 : n6758;
  assign n6760 = pi13 ? n5438 : n2391;
  assign n6761 = pi12 ? n26 : n6760;
  assign n6762 = pi15 ? n28 : ~n1200;
  assign n6763 = pi14 ? n6762 : n26;
  assign n6764 = pi13 ? n6763 : n2391;
  assign n6765 = pi12 ? n26 : n6764;
  assign n6766 = pi11 ? n6761 : n6765;
  assign n6767 = pi10 ? n6759 : n6766;
  assign n6768 = pi13 ? n6140 : n2370;
  assign n6769 = pi12 ? n26 : n6768;
  assign n6770 = pi11 ? n6769 : n6158;
  assign n6771 = pi14 ? n125 : n320;
  assign n6772 = pi13 ? n6771 : ~n72;
  assign n6773 = pi12 ? n26 : n6772;
  assign n6774 = pi13 ? n610 : ~n72;
  assign n6775 = pi12 ? n26 : n6774;
  assign n6776 = pi11 ? n6773 : n6775;
  assign n6777 = pi10 ? n6770 : n6776;
  assign n6778 = pi09 ? n6767 : n6777;
  assign n6779 = pi08 ? n6132 : n6778;
  assign n6780 = pi07 ? n6563 : n6779;
  assign n6781 = pi12 ? n26 : ~n6339;
  assign n6782 = pi12 ? n26 : ~n6335;
  assign n6783 = pi11 ? n6781 : n6782;
  assign n6784 = pi10 ? n5013 : n6783;
  assign n6785 = pi12 ? n124 : ~n6335;
  assign n6786 = pi12 ? n69 : ~n6339;
  assign n6787 = pi11 ? n6785 : n6786;
  assign n6788 = pi13 ? n1091 : n72;
  assign n6789 = pi12 ? n78 : ~n6788;
  assign n6790 = pi13 ? n4425 : n72;
  assign n6791 = pi12 ? n78 : ~n6790;
  assign n6792 = pi11 ? n6789 : n6791;
  assign n6793 = pi10 ? n6787 : n6792;
  assign n6794 = pi09 ? n6784 : n6793;
  assign n6795 = pi08 ? n6794 : n6789;
  assign n6796 = pi12 ? n69 : ~n6435;
  assign n6797 = pi11 ? n6789 : n6796;
  assign n6798 = pi13 ? n6303 : ~n26;
  assign n6799 = pi12 ? n78 : ~n6798;
  assign n6800 = pi10 ? n6797 : n6799;
  assign n6801 = pi09 ? n6789 : n6800;
  assign n6802 = pi08 ? n6789 : n6801;
  assign n6803 = pi07 ? n6795 : n6802;
  assign n6804 = pi06 ? n6780 : n6803;
  assign n6805 = pi11 ? n6358 : n5039;
  assign n6806 = pi11 ? n4633 : n6799;
  assign n6807 = pi10 ? n6805 : n6806;
  assign n6808 = pi09 ? n6356 : n6807;
  assign n6809 = pi08 ? n26 : n6808;
  assign n6810 = pi07 ? n26 : n6809;
  assign n6811 = pi06 ? n26 : n6810;
  assign n6812 = pi05 ? n6804 : n6811;
  assign n6813 = pi04 ? n6754 : n6812;
  assign n6814 = pi03 ? n6682 : n6813;
  assign n6815 = pi13 ? n869 : n4471;
  assign n6816 = pi12 ? n26 : n6815;
  assign n6817 = pi11 ? n26 : n6816;
  assign n6818 = pi10 ? n26 : n6817;
  assign n6819 = pi13 ? n2011 : n130;
  assign n6820 = pi12 ? n69 : ~n6819;
  assign n6821 = pi11 ? n6820 : n6378;
  assign n6822 = pi10 ? n6821 : n6385;
  assign n6823 = pi09 ? n6818 : n6822;
  assign n6824 = pi08 ? n26 : n6823;
  assign n6825 = pi07 ? n26 : n6824;
  assign n6826 = pi06 ? n26 : n6825;
  assign n6827 = pi13 ? n169 : n284;
  assign n6828 = pi12 ? n26 : n6827;
  assign n6829 = pi11 ? n26 : n6828;
  assign n6830 = pi10 ? n6829 : n6395;
  assign n6831 = pi09 ? n26 : n6830;
  assign n6832 = pi08 ? n26 : n6831;
  assign n6833 = pi07 ? n6832 : n6395;
  assign n6834 = pi06 ? n6833 : n6441;
  assign n6835 = pi05 ? n6826 : n6834;
  assign n6836 = pi07 ? n6449 : n6445;
  assign n6837 = pi06 ? n6836 : n6487;
  assign n6838 = pi13 ? n1982 : n6000;
  assign n6839 = pi12 ? n26 : n6838;
  assign n6840 = pi11 ? n26 : n6839;
  assign n6841 = pi14 ? n45 : n4140;
  assign n6842 = pi13 ? n4753 : n6841;
  assign n6843 = pi12 ? n26 : n6842;
  assign n6844 = pi11 ? n6843 : n6508;
  assign n6845 = pi10 ? n6840 : n6844;
  assign n6846 = pi09 ? n26 : n6845;
  assign n6847 = pi08 ? n26 : n6846;
  assign n6848 = pi07 ? n6847 : n6493;
  assign n6849 = pi06 ? n6848 : n6553;
  assign n6850 = pi05 ? n6837 : n6849;
  assign n6851 = pi04 ? n6835 : n6850;
  assign n6852 = pi11 ? n26 : n6567;
  assign n6853 = pi10 ? n6852 : n5355;
  assign n6854 = pi09 ? n26 : n6853;
  assign n6855 = pi08 ? n26 : n6854;
  assign n6856 = pi07 ? n6855 : n6132;
  assign n6857 = pi06 ? n6856 : n6606;
  assign n6858 = pi13 ? n3782 : n5777;
  assign n6859 = pi12 ? n26 : n6858;
  assign n6860 = pi11 ? n26 : n6859;
  assign n6861 = pi13 ? n2319 : n1280;
  assign n6862 = pi12 ? n26 : n6861;
  assign n6863 = pi10 ? n6860 : n6862;
  assign n6864 = pi09 ? n26 : n6863;
  assign n6865 = pi08 ? n26 : n6864;
  assign n6866 = pi10 ? n2342 : n26;
  assign n6867 = pi09 ? n6866 : n26;
  assign n6868 = pi08 ? n6867 : n26;
  assign n6869 = pi07 ? n6865 : n6868;
  assign n6870 = pi06 ? n6869 : n26;
  assign n6871 = pi05 ? n6857 : n6870;
  assign n6872 = pi13 ? n2319 : n1705;
  assign n6873 = pi12 ? n26 : n6872;
  assign n6874 = pi11 ? n6873 : n6183;
  assign n6875 = pi10 ? n5089 : n6874;
  assign n6876 = pi09 ? n26 : n6875;
  assign n6877 = pi08 ? n26 : n6876;
  assign n6878 = pi11 ? n3207 : n6637;
  assign n6879 = pi10 ? n6878 : n26;
  assign n6880 = pi09 ? n6879 : n26;
  assign n6881 = pi08 ? n6880 : n26;
  assign n6882 = pi07 ? n6877 : n6881;
  assign n6883 = pi06 ? n6882 : n26;
  assign n6884 = pi13 ? n1091 : n5777;
  assign n6885 = pi12 ? n26 : n6884;
  assign n6886 = pi11 ? n26 : n6885;
  assign n6887 = pi13 ? n2319 : n2631;
  assign n6888 = pi12 ? n26 : n6887;
  assign n6889 = pi11 ? n6155 : n6888;
  assign n6890 = pi10 ? n6886 : n6889;
  assign n6891 = pi09 ? n26 : n6890;
  assign n6892 = pi08 ? n26 : n6891;
  assign n6893 = pi11 ? n5908 : n6637;
  assign n6894 = pi13 ? n5690 : n2319;
  assign n6895 = pi12 ? n26 : n6894;
  assign n6896 = pi11 ? n6671 : n6895;
  assign n6897 = pi10 ? n6893 : n6896;
  assign n6898 = pi10 ? n6243 : n6242;
  assign n6899 = pi09 ? n6897 : n6898;
  assign n6900 = pi08 ? n6899 : n6242;
  assign n6901 = pi07 ? n6892 : n6900;
  assign n6902 = pi06 ? n6901 : n6242;
  assign n6903 = pi05 ? n6883 : n6902;
  assign n6904 = pi04 ? n6871 : n6903;
  assign n6905 = pi03 ? n6851 : n6904;
  assign n6906 = pi02 ? n6814 : n6905;
  assign n6907 = pi13 ? n2370 : n6088;
  assign n6908 = pi12 ? n26 : n6907;
  assign n6909 = pi11 ? n6908 : n3531;
  assign n6910 = pi10 ? n6179 : n6909;
  assign n6911 = pi09 ? n26 : n6910;
  assign n6912 = pi08 ? n26 : n6911;
  assign n6913 = pi10 ? n6193 : n6273;
  assign n6914 = pi11 ? n4526 : n4535;
  assign n6915 = pi10 ? n6914 : n4535;
  assign n6916 = pi09 ? n6913 : n6915;
  assign n6917 = pi08 ? n6916 : n4535;
  assign n6918 = pi07 ? n6912 : n6917;
  assign n6919 = pi06 ? n6918 : n4546;
  assign n6920 = pi13 ? n1135 : n3980;
  assign n6921 = pi12 ? n26 : n6920;
  assign n6922 = pi14 ? n233 : n327;
  assign n6923 = pi13 ? n6720 : n6922;
  assign n6924 = pi12 ? n26 : n6923;
  assign n6925 = pi11 ? n6921 : n6924;
  assign n6926 = pi10 ? n6222 : n6925;
  assign n6927 = pi09 ? n26 : n6926;
  assign n6928 = pi08 ? n26 : n6927;
  assign n6929 = pi13 ? n6071 : ~n126;
  assign n6930 = pi12 ? n26 : n6929;
  assign n6931 = pi11 ? n6265 : n6930;
  assign n6932 = pi13 ? n143 : ~n4153;
  assign n6933 = pi12 ? n26 : n6932;
  assign n6934 = pi12 ? n26 : n6300;
  assign n6935 = pi11 ? n6933 : n6934;
  assign n6936 = pi10 ? n6931 : n6935;
  assign n6937 = pi12 ? n124 : n6732;
  assign n6938 = pi13 ? n406 : n2762;
  assign n6939 = pi12 ? n69 : n6938;
  assign n6940 = pi11 ? n6937 : n6939;
  assign n6941 = pi12 ? n78 : n6738;
  assign n6942 = pi11 ? n6941 : n6742;
  assign n6943 = pi10 ? n6940 : n6942;
  assign n6944 = pi09 ? n6936 : n6943;
  assign n6945 = pi08 ? n6944 : n6742;
  assign n6946 = pi07 ? n6928 : n6945;
  assign n6947 = pi11 ? n6742 : n6746;
  assign n6948 = pi10 ? n6742 : n6947;
  assign n6949 = pi14 ? n320 : ~n327;
  assign n6950 = pi13 ? n6949 : n26;
  assign n6951 = pi12 ? n69 : n6950;
  assign n6952 = pi11 ? n6746 : n6951;
  assign n6953 = pi10 ? n6952 : n6742;
  assign n6954 = pi09 ? n6948 : n6953;
  assign n6955 = pi08 ? n6954 : n6742;
  assign n6956 = pi07 ? n6955 : n6742;
  assign n6957 = pi06 ? n6946 : n6956;
  assign n6958 = pi05 ? n6919 : n6957;
  assign n6959 = pi11 ? n26 : n5368;
  assign n6960 = pi14 ? n125 : n327;
  assign n6961 = pi13 ? n1135 : n6960;
  assign n6962 = pi12 ? n26 : n6961;
  assign n6963 = pi14 ? n168 : n320;
  assign n6964 = pi13 ? n6963 : n6540;
  assign n6965 = pi12 ? n26 : n6964;
  assign n6966 = pi11 ? n6962 : n6965;
  assign n6967 = pi10 ? n6959 : n6966;
  assign n6968 = pi09 ? n26 : n6967;
  assign n6969 = pi08 ? n26 : n6968;
  assign n6970 = pi13 ? n6260 : ~n72;
  assign n6971 = pi12 ? n26 : n6970;
  assign n6972 = pi11 ? n6775 : n6971;
  assign n6973 = pi13 ? n1091 : n1925;
  assign n6974 = pi12 ? n26 : ~n6973;
  assign n6975 = pi11 ? n5185 : n6974;
  assign n6976 = pi10 ? n6972 : n6975;
  assign n6977 = pi12 ? n69 : ~n6335;
  assign n6978 = pi11 ? n6785 : n6977;
  assign n6979 = pi10 ? n6978 : n6340;
  assign n6980 = pi09 ? n6976 : n6979;
  assign n6981 = pi11 ? n6791 : n6789;
  assign n6982 = pi10 ? n6981 : n6789;
  assign n6983 = pi09 ? n6982 : n6789;
  assign n6984 = pi08 ? n6980 : n6983;
  assign n6985 = pi07 ? n6969 : n6984;
  assign n6986 = pi12 ? n69 : ~n6798;
  assign n6987 = pi11 ? n6986 : n6799;
  assign n6988 = pi13 ? n6303 : n507;
  assign n6989 = pi12 ? n78 : ~n6988;
  assign n6990 = pi11 ? n6989 : n6789;
  assign n6991 = pi10 ? n6987 : n6990;
  assign n6992 = pi09 ? n6789 : n6991;
  assign n6993 = pi08 ? n6992 : n6789;
  assign n6994 = pi12 ? n78 : n5467;
  assign n6995 = pi11 ? n6789 : n6994;
  assign n6996 = pi10 ? n6789 : n6995;
  assign n6997 = pi09 ? n6789 : n6996;
  assign n6998 = pi08 ? n6789 : n6997;
  assign n6999 = pi07 ? n6993 : n6998;
  assign n7000 = pi06 ? n6985 : n6999;
  assign n7001 = pi11 ? n6354 : n6358;
  assign n7002 = pi10 ? n26 : n7001;
  assign n7003 = pi13 ? n5037 : ~n26;
  assign n7004 = pi12 ? n78 : ~n7003;
  assign n7005 = pi10 ? n7004 : n26;
  assign n7006 = pi09 ? n7002 : n7005;
  assign n7007 = pi08 ? n7006 : n26;
  assign n7008 = pi07 ? n7007 : n26;
  assign n7009 = pi06 ? n26 : n7008;
  assign n7010 = pi05 ? n7000 : n7009;
  assign n7011 = pi04 ? n6958 : n7010;
  assign n7012 = pi13 ? n869 : n3980;
  assign n7013 = pi12 ? n26 : n7012;
  assign n7014 = pi11 ? n7013 : n6820;
  assign n7015 = pi10 ? n26 : n7014;
  assign n7016 = pi13 ? n3782 : n38;
  assign n7017 = pi12 ? n78 : ~n7016;
  assign n7018 = pi12 ? n78 : ~n6383;
  assign n7019 = pi11 ? n7017 : n7018;
  assign n7020 = pi10 ? n7019 : n26;
  assign n7021 = pi09 ? n7015 : n7020;
  assign n7022 = pi08 ? n7021 : n26;
  assign n7023 = pi07 ? n7022 : n26;
  assign n7024 = pi06 ? n26 : n7023;
  assign n7025 = pi10 ? n6829 : n6646;
  assign n7026 = pi09 ? n26 : n7025;
  assign n7027 = pi08 ? n26 : n7026;
  assign n7028 = pi14 ? n147 : ~n1704;
  assign n7029 = pi13 ? n130 : ~n7028;
  assign n7030 = pi12 ? n26 : n7029;
  assign n7031 = pi11 ? n6646 : n7030;
  assign n7032 = pi13 ? n176 : ~n6417;
  assign n7033 = pi12 ? n26 : n7032;
  assign n7034 = pi11 ? n6416 : n7033;
  assign n7035 = pi10 ? n7031 : n7034;
  assign n7036 = pi09 ? n6646 : n7035;
  assign n7037 = pi08 ? n6646 : n7036;
  assign n7038 = pi07 ? n7027 : n7037;
  assign n7039 = pi14 ? n147 : ~n73;
  assign n7040 = pi13 ? n1438 : ~n7039;
  assign n7041 = pi12 ? n26 : n7040;
  assign n7042 = pi11 ? n7041 : n4108;
  assign n7043 = pi13 ? n3980 : n4425;
  assign n7044 = pi12 ? n26 : n7043;
  assign n7045 = pi15 ? n44 : n1200;
  assign n7046 = pi14 ? n292 : n7045;
  assign n7047 = pi13 ? n7046 : n176;
  assign n7048 = pi12 ? n69 : ~n7047;
  assign n7049 = pi11 ? n7044 : n7048;
  assign n7050 = pi10 ? n7042 : n7049;
  assign n7051 = pi12 ? n69 : ~n7016;
  assign n7052 = pi12 ? n124 : n5467;
  assign n7053 = pi11 ? n7051 : n7052;
  assign n7054 = pi15 ? n1200 : n44;
  assign n7055 = pi14 ? n26 : ~n7054;
  assign n7056 = pi13 ? n7055 : n2519;
  assign n7057 = pi12 ? n26 : n7056;
  assign n7058 = pi13 ? n5690 : n2347;
  assign n7059 = pi12 ? n26 : n7058;
  assign n7060 = pi11 ? n7057 : n7059;
  assign n7061 = pi10 ? n7053 : n7060;
  assign n7062 = pi09 ? n7050 : n7061;
  assign n7063 = pi08 ? n7062 : n6242;
  assign n7064 = pi07 ? n7063 : n6242;
  assign n7065 = pi06 ? n7038 : n7064;
  assign n7066 = pi05 ? n7024 : n7065;
  assign n7067 = pi13 ? n79 : n5615;
  assign n7068 = pi12 ? n26 : n7067;
  assign n7069 = pi11 ? n5606 : n7068;
  assign n7070 = pi13 ? n57 : n1344;
  assign n7071 = pi12 ? n26 : n7070;
  assign n7072 = pi13 ? n57 : n4622;
  assign n7073 = pi12 ? n26 : n7072;
  assign n7074 = pi11 ? n7071 : n7073;
  assign n7075 = pi10 ? n7069 : n7074;
  assign n7076 = pi09 ? n6445 : n7075;
  assign n7077 = pi08 ? n6445 : n7076;
  assign n7078 = pi07 ? n6449 : n7077;
  assign n7079 = pi13 ? n79 : n3996;
  assign n7080 = pi12 ? n26 : n7079;
  assign n7081 = pi11 ? n7080 : n4108;
  assign n7082 = pi13 ? n4471 : n4425;
  assign n7083 = pi12 ? n26 : n7082;
  assign n7084 = pi13 ? n6368 : n3980;
  assign n7085 = pi12 ? n69 : n7084;
  assign n7086 = pi11 ? n7083 : n7085;
  assign n7087 = pi10 ? n7081 : n7086;
  assign n7088 = pi12 ? n654 : n6544;
  assign n7089 = pi11 ? n7088 : n6482;
  assign n7090 = pi13 ? n6268 : n26;
  assign n7091 = pi12 ? n26 : n7090;
  assign n7092 = pi13 ? n5886 : n2519;
  assign n7093 = pi12 ? n26 : n7092;
  assign n7094 = pi11 ? n7091 : n7093;
  assign n7095 = pi10 ? n7089 : n7094;
  assign n7096 = pi09 ? n7087 : n7095;
  assign n7097 = pi08 ? n7096 : n4535;
  assign n7098 = pi07 ? n7097 : n4545;
  assign n7099 = pi06 ? n7078 : n7098;
  assign n7100 = pi13 ? n79 : n6000;
  assign n7101 = pi12 ? n26 : n7100;
  assign n7102 = pi11 ? n26 : n7101;
  assign n7103 = pi13 ? n1344 : n6841;
  assign n7104 = pi12 ? n26 : n7103;
  assign n7105 = pi11 ? n7104 : n6508;
  assign n7106 = pi10 ? n7102 : n7105;
  assign n7107 = pi09 ? n26 : n7106;
  assign n7108 = pi08 ? n26 : n7107;
  assign n7109 = pi13 ? n4769 : n4809;
  assign n7110 = pi12 ? n26 : n7109;
  assign n7111 = pi11 ? n6517 : n7110;
  assign n7112 = pi11 ? n6713 : n6529;
  assign n7113 = pi10 ? n7111 : n7112;
  assign n7114 = pi09 ? n6493 : n7113;
  assign n7115 = pi08 ? n6493 : n7114;
  assign n7116 = pi07 ? n7108 : n7115;
  assign n7117 = pi13 ? n5320 : n3918;
  assign n7118 = pi12 ? n26 : n7117;
  assign n7119 = pi14 ? n1437 : ~n29;
  assign n7120 = pi14 ? n71 : ~n71;
  assign n7121 = pi13 ? n7119 : n7120;
  assign n7122 = pi12 ? n26 : n7121;
  assign n7123 = pi11 ? n7118 : n7122;
  assign n7124 = pi13 ? n3980 : n3066;
  assign n7125 = pi12 ? n26 : n7124;
  assign n7126 = pi13 ? n130 : ~n1135;
  assign n7127 = pi12 ? n26 : ~n7126;
  assign n7128 = pi11 ? n7125 : n7127;
  assign n7129 = pi10 ? n7123 : n7128;
  assign n7130 = pi13 ? n6771 : n6596;
  assign n7131 = pi12 ? n26 : n7130;
  assign n7132 = pi13 ? n6208 : ~n1139;
  assign n7133 = pi12 ? n69 : n7132;
  assign n7134 = pi11 ? n7131 : n7133;
  assign n7135 = pi14 ? n147 : n37;
  assign n7136 = pi13 ? n7135 : ~n126;
  assign n7137 = pi12 ? n78 : n7136;
  assign n7138 = pi14 ? n233 : ~n233;
  assign n7139 = pi13 ? n7138 : ~n126;
  assign n7140 = pi12 ? n78 : n7139;
  assign n7141 = pi11 ? n7137 : n7140;
  assign n7142 = pi10 ? n7134 : n7141;
  assign n7143 = pi09 ? n7129 : n7142;
  assign n7144 = pi13 ? n351 : n2519;
  assign n7145 = pi12 ? n78 : n7144;
  assign n7146 = pi11 ? n7145 : n4576;
  assign n7147 = pi10 ? n7146 : n6942;
  assign n7148 = pi09 ? n7147 : n6742;
  assign n7149 = pi08 ? n7143 : n7148;
  assign n7150 = pi07 ? n7149 : n6742;
  assign n7151 = pi06 ? n7116 : n7150;
  assign n7152 = pi05 ? n7099 : n7151;
  assign n7153 = pi04 ? n7066 : n7152;
  assign n7154 = pi03 ? n7011 : n7153;
  assign n7155 = pi13 ? n4135 : n5677;
  assign n7156 = pi12 ? n26 : n7155;
  assign n7157 = pi11 ? n26 : n7156;
  assign n7158 = pi13 ? n4139 : n3061;
  assign n7159 = pi12 ? n26 : n7158;
  assign n7160 = pi11 ? n7159 : n6569;
  assign n7161 = pi10 ? n7157 : n7160;
  assign n7162 = pi09 ? n26 : n7161;
  assign n7163 = pi08 ? n26 : n7162;
  assign n7164 = pi13 ? n2955 : n6109;
  assign n7165 = pi12 ? n26 : n7164;
  assign n7166 = pi11 ? n6105 : n7165;
  assign n7167 = pi13 ? n5438 : n3066;
  assign n7168 = pi12 ? n26 : n7167;
  assign n7169 = pi11 ? n7168 : n6585;
  assign n7170 = pi10 ? n7166 : n7169;
  assign n7171 = pi09 ? n6132 : n7170;
  assign n7172 = pi08 ? n6132 : n7171;
  assign n7173 = pi07 ? n7163 : n7172;
  assign n7174 = pi14 ? n3250 : n26;
  assign n7175 = pi13 ? n7174 : n3066;
  assign n7176 = pi12 ? n26 : n7175;
  assign n7177 = pi14 ? n2410 : n26;
  assign n7178 = pi13 ? n7177 : n3066;
  assign n7179 = pi12 ? n26 : n7178;
  assign n7180 = pi11 ? n7176 : n7179;
  assign n7181 = pi13 ? n630 : n2319;
  assign n7182 = pi12 ? n26 : n7181;
  assign n7183 = pi12 ? n124 : ~n6538;
  assign n7184 = pi11 ? n7182 : n7183;
  assign n7185 = pi10 ? n7180 : n7184;
  assign n7186 = pi13 ? n415 : ~n6596;
  assign n7187 = pi12 ? n69 : ~n7186;
  assign n7188 = pi12 ? n78 : ~n6168;
  assign n7189 = pi11 ? n7187 : n7188;
  assign n7190 = pi14 ? n37 : n1832;
  assign n7191 = pi13 ? n7190 : n72;
  assign n7192 = pi12 ? n78 : ~n7191;
  assign n7193 = pi11 ? n4603 : n7192;
  assign n7194 = pi10 ? n7189 : n7193;
  assign n7195 = pi09 ? n7185 : n7194;
  assign n7196 = pi10 ? n6336 : n6340;
  assign n7197 = pi09 ? n7196 : n6982;
  assign n7198 = pi08 ? n7195 : n7197;
  assign n7199 = pi07 ? n7198 : n6998;
  assign n7200 = pi06 ? n7173 : n7199;
  assign n7201 = pi10 ? n6860 : n5391;
  assign n7202 = pi09 ? n26 : n7201;
  assign n7203 = pi08 ? n26 : n7202;
  assign n7204 = pi07 ? n7203 : n6868;
  assign n7205 = pi06 ? n7204 : n26;
  assign n7206 = pi05 ? n7200 : n7205;
  assign n7207 = pi13 ? n4226 : n1705;
  assign n7208 = pi12 ? n26 : n7207;
  assign n7209 = pi11 ? n7208 : n6183;
  assign n7210 = pi10 ? n5077 : n7209;
  assign n7211 = pi09 ? n26 : n7210;
  assign n7212 = pi08 ? n26 : n7211;
  assign n7213 = pi07 ? n7212 : n6881;
  assign n7214 = pi06 ? n7213 : n26;
  assign n7215 = pi11 ? n6908 : n6888;
  assign n7216 = pi10 ? n6886 : n7215;
  assign n7217 = pi09 ? n26 : n7216;
  assign n7218 = pi08 ? n26 : n7217;
  assign n7219 = pi09 ? n6897 : n6242;
  assign n7220 = pi08 ? n7219 : n6242;
  assign n7221 = pi07 ? n7218 : n7220;
  assign n7222 = pi06 ? n7221 : n6242;
  assign n7223 = pi05 ? n7214 : n7222;
  assign n7224 = pi04 ? n7206 : n7223;
  assign n7225 = pi13 ? n1135 : n6922;
  assign n7226 = pi12 ? n26 : n7225;
  assign n7227 = pi11 ? n6908 : n7226;
  assign n7228 = pi10 ? n6179 : n7227;
  assign n7229 = pi09 ? n26 : n7228;
  assign n7230 = pi08 ? n26 : n7229;
  assign n7231 = pi14 ? n168 : n3250;
  assign n7232 = pi13 ? n7231 : ~n2498;
  assign n7233 = pi12 ? n26 : ~n7232;
  assign n7234 = pi11 ? n7233 : n6272;
  assign n7235 = pi10 ? n6193 : n7234;
  assign n7236 = pi13 ? n5956 : n26;
  assign n7237 = pi12 ? n26 : n7236;
  assign n7238 = pi13 ? n3061 : n26;
  assign n7239 = pi12 ? n26 : n7238;
  assign n7240 = pi11 ? n7237 : n7239;
  assign n7241 = pi10 ? n7240 : n7239;
  assign n7242 = pi09 ? n7235 : n7241;
  assign n7243 = pi08 ? n7242 : n7239;
  assign n7244 = pi07 ? n7230 : n7243;
  assign n7245 = pi12 ? n26 : n6747;
  assign n7246 = pi11 ? n7239 : n7245;
  assign n7247 = pi10 ? n7239 : n7246;
  assign n7248 = pi09 ? n7239 : n7247;
  assign n7249 = pi08 ? n7239 : n7248;
  assign n7250 = pi07 ? n7239 : n7249;
  assign n7251 = pi06 ? n7244 : n7250;
  assign n7252 = pi14 ? n26 : ~n1832;
  assign n7253 = pi13 ? n7252 : ~n5431;
  assign n7254 = pi12 ? n26 : n7253;
  assign n7255 = pi13 ? n6233 : n26;
  assign n7256 = pi12 ? n26 : n7255;
  assign n7257 = pi11 ? n7254 : n7256;
  assign n7258 = pi10 ? n6193 : n7257;
  assign n7259 = pi14 ? n327 : ~n168;
  assign n7260 = pi13 ? n5886 : n7259;
  assign n7261 = pi12 ? n124 : n7260;
  assign n7262 = pi13 ? n3100 : n2904;
  assign n7263 = pi12 ? n26 : n7262;
  assign n7264 = pi11 ? n7261 : n7263;
  assign n7265 = pi12 ? n69 : n4534;
  assign n7266 = pi11 ? n4585 : n7265;
  assign n7267 = pi10 ? n7264 : n7266;
  assign n7268 = pi09 ? n7258 : n7267;
  assign n7269 = pi08 ? n7268 : n7265;
  assign n7270 = pi07 ? n6928 : n7269;
  assign n7271 = pi11 ? n7265 : n4585;
  assign n7272 = pi10 ? n7265 : n7271;
  assign n7273 = pi09 ? n7265 : n7272;
  assign n7274 = pi08 ? n7265 : n7273;
  assign n7275 = pi07 ? n7265 : n7274;
  assign n7276 = pi06 ? n7270 : n7275;
  assign n7277 = pi05 ? n7251 : n7276;
  assign n7278 = pi13 ? n1135 : ~n4341;
  assign n7279 = pi12 ? n26 : n7278;
  assign n7280 = pi13 ? n6771 : ~n415;
  assign n7281 = pi12 ? n26 : n7280;
  assign n7282 = pi11 ? n7279 : n7281;
  assign n7283 = pi10 ? n6222 : n7282;
  assign n7284 = pi09 ? n26 : n7283;
  assign n7285 = pi08 ? n26 : n7284;
  assign n7286 = pi13 ? n6208 : ~n126;
  assign n7287 = pi12 ? n26 : n7286;
  assign n7288 = pi11 ? n6265 : n7287;
  assign n7289 = pi13 ? n4325 : n125;
  assign n7290 = pi12 ? n26 : ~n7289;
  assign n7291 = pi11 ? n5468 : n7290;
  assign n7292 = pi10 ? n7288 : n7291;
  assign n7293 = pi14 ? n1872 : n168;
  assign n7294 = pi13 ? n351 : ~n7293;
  assign n7295 = pi12 ? n78 : n7294;
  assign n7296 = pi13 ? n6297 : n7293;
  assign n7297 = pi12 ? n78 : ~n7296;
  assign n7298 = pi11 ? n7295 : n7297;
  assign n7299 = pi13 ? n351 : ~n5479;
  assign n7300 = pi12 ? n78 : n7299;
  assign n7301 = pi12 ? n78 : n1894;
  assign n7302 = pi11 ? n7300 : n7301;
  assign n7303 = pi10 ? n7298 : n7302;
  assign n7304 = pi09 ? n7292 : n7303;
  assign n7305 = pi10 ? n5483 : n5205;
  assign n7306 = pi09 ? n7305 : n5205;
  assign n7307 = pi08 ? n7304 : n7306;
  assign n7308 = pi07 ? n7285 : n7307;
  assign n7309 = pi06 ? n7308 : n5205;
  assign n7310 = pi13 ? n6963 : ~n72;
  assign n7311 = pi12 ? n26 : n7310;
  assign n7312 = pi11 ? n4552 : n7311;
  assign n7313 = pi10 ? n6321 : n7312;
  assign n7314 = pi09 ? n26 : n7313;
  assign n7315 = pi08 ? n26 : n7314;
  assign n7316 = pi12 ? n26 : ~n6329;
  assign n7317 = pi11 ? n7316 : n6327;
  assign n7318 = pi12 ? n69 : ~n4602;
  assign n7319 = pi11 ? n5500 : n7318;
  assign n7320 = pi10 ? n7317 : n7319;
  assign n7321 = pi13 ? n4838 : n72;
  assign n7322 = pi12 ? n78 : ~n7321;
  assign n7323 = pi11 ? n7322 : n6336;
  assign n7324 = pi10 ? n7323 : n6336;
  assign n7325 = pi09 ? n7320 : n7324;
  assign n7326 = pi10 ? n6789 : n6340;
  assign n7327 = pi09 ? n7326 : n6340;
  assign n7328 = pi08 ? n7325 : n7327;
  assign n7329 = pi07 ? n7315 : n7328;
  assign n7330 = pi11 ? n6340 : n6301;
  assign n7331 = pi10 ? n6340 : n7330;
  assign n7332 = pi09 ? n6340 : n7331;
  assign n7333 = pi08 ? n6340 : n7332;
  assign n7334 = pi07 ? n6340 : n7333;
  assign n7335 = pi06 ? n7329 : n7334;
  assign n7336 = pi05 ? n7309 : n7335;
  assign n7337 = pi04 ? n7277 : n7336;
  assign n7338 = pi03 ? n7224 : n7337;
  assign n7339 = pi02 ? n7154 : n7338;
  assign n7340 = pi01 ? n6906 : n7339;
  assign n7341 = pi00 ? n6559 : n7340;
  assign n7342 = pi09 ? n26 : n2502;
  assign n7343 = pi08 ? n26 : n7342;
  assign n7344 = pi13 ? n26 : n3023;
  assign n7345 = pi12 ? n26 : n7344;
  assign n7346 = pi09 ? n2500 : n7345;
  assign n7347 = pi15 ? n291 : n60;
  assign n7348 = pi14 ? n26 : n7347;
  assign n7349 = pi13 ? n26 : n7348;
  assign n7350 = pi12 ? n26 : n7349;
  assign n7351 = pi12 ? n26 : n2857;
  assign n7352 = pi11 ? n7350 : n7351;
  assign n7353 = pi10 ? n7352 : n26;
  assign n7354 = pi09 ? n7353 : n2502;
  assign n7355 = pi08 ? n7346 : n7354;
  assign n7356 = pi07 ? n7343 : n7355;
  assign n7357 = pi09 ? n7345 : n7353;
  assign n7358 = pi09 ? n2502 : n7345;
  assign n7359 = pi08 ? n7357 : n7358;
  assign n7360 = pi12 ? n26 : n3023;
  assign n7361 = pi11 ? n26 : n7360;
  assign n7362 = pi14 ? n26 : n3250;
  assign n7363 = pi13 ? n7362 : n3023;
  assign n7364 = pi12 ? n26 : n7363;
  assign n7365 = pi11 ? n7360 : n7364;
  assign n7366 = pi10 ? n7361 : n7365;
  assign n7367 = pi09 ? n7353 : n7366;
  assign n7368 = pi13 ? n3023 : n3942;
  assign n7369 = pi12 ? n26 : n7368;
  assign n7370 = pi11 ? n7360 : n7369;
  assign n7371 = pi10 ? n7360 : n7370;
  assign n7372 = pi14 ? n26 : n4243;
  assign n7373 = pi13 ? n26 : n7372;
  assign n7374 = pi12 ? n26 : n7373;
  assign n7375 = pi11 ? n7360 : n7374;
  assign n7376 = pi13 ? n97 : n26;
  assign n7377 = pi12 ? n124 : n7376;
  assign n7378 = pi14 ? n291 : n26;
  assign n7379 = pi13 ? n2315 : n7378;
  assign n7380 = pi12 ? n69 : n7379;
  assign n7381 = pi11 ? n7377 : n7380;
  assign n7382 = pi10 ? n7375 : n7381;
  assign n7383 = pi09 ? n7371 : n7382;
  assign n7384 = pi08 ? n7367 : n7383;
  assign n7385 = pi07 ? n7359 : n7384;
  assign n7386 = pi06 ? n7356 : n7385;
  assign n7387 = pi05 ? n26 : n7386;
  assign n7388 = pi11 ? n26 : n2341;
  assign n7389 = pi13 ? n26 : n2319;
  assign n7390 = pi12 ? n26 : n7389;
  assign n7391 = pi10 ? n7388 : n7390;
  assign n7392 = pi09 ? n26 : n7391;
  assign n7393 = pi08 ? n26 : n7392;
  assign n7394 = pi10 ? n7390 : n2341;
  assign n7395 = pi12 ? n26 : n2891;
  assign n7396 = pi11 ? n7395 : n3028;
  assign n7397 = pi11 ? n7345 : n3191;
  assign n7398 = pi10 ? n7396 : n7397;
  assign n7399 = pi09 ? n7394 : n7398;
  assign n7400 = pi13 ? n26 : n2403;
  assign n7401 = pi12 ? n26 : n7400;
  assign n7402 = pi13 ? n97 : ~n507;
  assign n7403 = pi12 ? n26 : n7402;
  assign n7404 = pi11 ? n7401 : n7403;
  assign n7405 = pi10 ? n7404 : n26;
  assign n7406 = pi10 ? n7388 : n2341;
  assign n7407 = pi09 ? n7405 : n7406;
  assign n7408 = pi08 ? n7399 : n7407;
  assign n7409 = pi07 ? n7393 : n7408;
  assign n7410 = pi09 ? n7398 : n7405;
  assign n7411 = pi09 ? n7406 : n7398;
  assign n7412 = pi08 ? n7410 : n7411;
  assign n7413 = pi11 ? n26 : n7345;
  assign n7414 = pi14 ? n292 : n233;
  assign n7415 = pi13 ? n26 : n7414;
  assign n7416 = pi12 ? n26 : n7415;
  assign n7417 = pi11 ? n7345 : n7416;
  assign n7418 = pi10 ? n7413 : n7417;
  assign n7419 = pi09 ? n7405 : n7418;
  assign n7420 = pi14 ? n63 : ~n1437;
  assign n7421 = pi13 ? n7420 : n7414;
  assign n7422 = pi12 ? n26 : n7421;
  assign n7423 = pi14 ? n517 : n292;
  assign n7424 = pi13 ? n7423 : n7414;
  assign n7425 = pi12 ? n26 : n7424;
  assign n7426 = pi11 ? n7422 : n7425;
  assign n7427 = pi10 ? n7416 : n7426;
  assign n7428 = pi14 ? n292 : n1832;
  assign n7429 = pi13 ? n3023 : n7428;
  assign n7430 = pi12 ? n26 : n7429;
  assign n7431 = pi14 ? n292 : n147;
  assign n7432 = pi13 ? n26 : n7431;
  assign n7433 = pi12 ? n124 : n7432;
  assign n7434 = pi11 ? n7430 : n7433;
  assign n7435 = pi14 ? n1437 : ~n7347;
  assign n7436 = pi13 ? n2315 : ~n7435;
  assign n7437 = pi12 ? n69 : n7436;
  assign n7438 = pi13 ? n2315 : n2741;
  assign n7439 = pi12 ? n26 : n7438;
  assign n7440 = pi11 ? n7437 : n7439;
  assign n7441 = pi10 ? n7434 : n7440;
  assign n7442 = pi09 ? n7427 : n7441;
  assign n7443 = pi08 ? n7419 : n7442;
  assign n7444 = pi07 ? n7412 : n7443;
  assign n7445 = pi06 ? n7409 : n7444;
  assign n7446 = pi14 ? n5885 : n292;
  assign n7447 = pi13 ? n26 : n7446;
  assign n7448 = pi12 ? n26 : n7447;
  assign n7449 = pi11 ? n26 : n7448;
  assign n7450 = pi14 ? n5885 : n26;
  assign n7451 = pi13 ? n26 : n7450;
  assign n7452 = pi12 ? n26 : n7451;
  assign n7453 = pi10 ? n7449 : n7452;
  assign n7454 = pi09 ? n26 : n7453;
  assign n7455 = pi08 ? n26 : n7454;
  assign n7456 = pi13 ? n26 : n3942;
  assign n7457 = pi12 ? n26 : n7456;
  assign n7458 = pi11 ? n7345 : n7457;
  assign n7459 = pi10 ? n7452 : n7458;
  assign n7460 = pi09 ? n7452 : n7459;
  assign n7461 = pi14 ? n168 : ~n7347;
  assign n7462 = pi13 ? n68 : ~n7461;
  assign n7463 = pi12 ? n26 : n7462;
  assign n7464 = pi11 ? n7401 : n7463;
  assign n7465 = pi10 ? n7464 : n26;
  assign n7466 = pi09 ? n7465 : n7453;
  assign n7467 = pi08 ? n7460 : n7466;
  assign n7468 = pi07 ? n7455 : n7467;
  assign n7469 = pi09 ? n7459 : n7465;
  assign n7470 = pi09 ? n7453 : n7459;
  assign n7471 = pi08 ? n7469 : n7470;
  assign n7472 = pi10 ? n7413 : n7345;
  assign n7473 = pi09 ? n7465 : n7472;
  assign n7474 = pi13 ? n6109 : n3023;
  assign n7475 = pi12 ? n26 : n7474;
  assign n7476 = pi11 ? n7345 : n7475;
  assign n7477 = pi13 ? n1280 : n3023;
  assign n7478 = pi12 ? n26 : n7477;
  assign n7479 = pi13 ? n7423 : n2498;
  assign n7480 = pi12 ? n26 : n7479;
  assign n7481 = pi11 ? n7478 : n7480;
  assign n7482 = pi10 ? n7476 : n7481;
  assign n7483 = pi14 ? n2386 : n147;
  assign n7484 = pi13 ? n7483 : n130;
  assign n7485 = pi12 ? n69 : n7484;
  assign n7486 = pi11 ? n7360 : n7485;
  assign n7487 = pi15 ? n291 : n1200;
  assign n7488 = pi14 ? n26 : n7487;
  assign n7489 = pi13 ? n1252 : ~n7488;
  assign n7490 = pi12 ? n69 : ~n7489;
  assign n7491 = pi14 ? n233 : n517;
  assign n7492 = pi13 ? n7491 : n478;
  assign n7493 = pi12 ? n26 : n7492;
  assign n7494 = pi11 ? n7490 : n7493;
  assign n7495 = pi10 ? n7486 : n7494;
  assign n7496 = pi09 ? n7482 : n7495;
  assign n7497 = pi08 ? n7473 : n7496;
  assign n7498 = pi07 ? n7471 : n7497;
  assign n7499 = pi06 ? n7468 : n7498;
  assign n7500 = pi05 ? n7445 : n7499;
  assign n7501 = pi04 ? n7387 : n7500;
  assign n7502 = pi03 ? n26 : n7501;
  assign n7503 = pi02 ? n26 : n7502;
  assign n7504 = pi10 ? n3000 : n5908;
  assign n7505 = pi09 ? n26 : n7504;
  assign n7506 = pi08 ? n26 : n7505;
  assign n7507 = pi13 ? n97 : n478;
  assign n7508 = pi12 ? n26 : n7507;
  assign n7509 = pi10 ? n5908 : n7508;
  assign n7510 = pi13 ? n74 : n3023;
  assign n7511 = pi12 ? n26 : n7510;
  assign n7512 = pi11 ? n26 : n7511;
  assign n7513 = pi10 ? n26 : n7512;
  assign n7514 = pi09 ? n7509 : n7513;
  assign n7515 = pi13 ? n74 : n3942;
  assign n7516 = pi12 ? n26 : n7515;
  assign n7517 = pi14 ? n168 : ~n7487;
  assign n7518 = pi13 ? n68 : ~n7517;
  assign n7519 = pi12 ? n26 : n7518;
  assign n7520 = pi11 ? n7516 : n7519;
  assign n7521 = pi10 ? n7520 : n26;
  assign n7522 = pi14 ? n233 : n292;
  assign n7523 = pi13 ? n26 : n7522;
  assign n7524 = pi12 ? n26 : n7523;
  assign n7525 = pi11 ? n26 : n7524;
  assign n7526 = pi10 ? n7525 : n7508;
  assign n7527 = pi09 ? n7521 : n7526;
  assign n7528 = pi08 ? n7514 : n7527;
  assign n7529 = pi07 ? n7506 : n7528;
  assign n7530 = pi09 ? n7513 : n7521;
  assign n7531 = pi09 ? n7526 : n7513;
  assign n7532 = pi08 ? n7530 : n7531;
  assign n7533 = pi14 ? n327 : n73;
  assign n7534 = pi13 ? n26 : n7533;
  assign n7535 = pi12 ? n26 : n7534;
  assign n7536 = pi11 ? n26 : n7535;
  assign n7537 = pi14 ? n7347 : n73;
  assign n7538 = pi13 ? n26 : n7537;
  assign n7539 = pi12 ? n26 : n7538;
  assign n7540 = pi10 ? n7536 : n7539;
  assign n7541 = pi09 ? n7521 : n7540;
  assign n7542 = pi13 ? n198 : n7537;
  assign n7543 = pi12 ? n26 : n7542;
  assign n7544 = pi11 ? n7539 : n7543;
  assign n7545 = pi13 ? n1280 : n7537;
  assign n7546 = pi12 ? n26 : n7545;
  assign n7547 = pi14 ? n432 : ~n1437;
  assign n7548 = pi13 ? n7547 : n7537;
  assign n7549 = pi12 ? n26 : n7548;
  assign n7550 = pi11 ? n7546 : n7549;
  assign n7551 = pi10 ? n7544 : n7550;
  assign n7552 = pi14 ? n7347 : n233;
  assign n7553 = pi13 ? n2391 : n7552;
  assign n7554 = pi12 ? n26 : n7553;
  assign n7555 = pi13 ? n2391 : n3023;
  assign n7556 = pi12 ? n26 : n7555;
  assign n7557 = pi11 ? n7554 : n7556;
  assign n7558 = pi10 ? n7557 : n6162;
  assign n7559 = pi09 ? n7551 : n7558;
  assign n7560 = pi08 ? n7541 : n7559;
  assign n7561 = pi07 ? n7532 : n7560;
  assign n7562 = pi06 ? n7529 : n7561;
  assign n7563 = pi14 ? n147 : n517;
  assign n7564 = pi13 ? n26 : n7563;
  assign n7565 = pi12 ? n26 : n7564;
  assign n7566 = pi11 ? n26 : n7565;
  assign n7567 = pi13 ? n97 : n7522;
  assign n7568 = pi12 ? n26 : n7567;
  assign n7569 = pi11 ? n5908 : n7568;
  assign n7570 = pi10 ? n7566 : n7569;
  assign n7571 = pi09 ? n26 : n7570;
  assign n7572 = pi08 ? n26 : n7571;
  assign n7573 = pi11 ? n7568 : n7524;
  assign n7574 = pi14 ? n233 : n4950;
  assign n7575 = pi13 ? n68 : n7574;
  assign n7576 = pi12 ? n26 : n7575;
  assign n7577 = pi15 ? n28 : n70;
  assign n7578 = pi14 ? n26 : n7577;
  assign n7579 = pi15 ? n291 : ~n28;
  assign n7580 = pi14 ? n26 : n7579;
  assign n7581 = pi13 ? n7578 : n7580;
  assign n7582 = pi12 ? n26 : n7581;
  assign n7583 = pi11 ? n7576 : n7582;
  assign n7584 = pi10 ? n7573 : n7583;
  assign n7585 = pi10 ? n26 : n2501;
  assign n7586 = pi09 ? n7584 : n7585;
  assign n7587 = pi10 ? n7369 : n26;
  assign n7588 = pi13 ? n26 : n7491;
  assign n7589 = pi12 ? n26 : n7588;
  assign n7590 = pi11 ? n26 : n7589;
  assign n7591 = pi14 ? n233 : n63;
  assign n7592 = pi13 ? n68 : n7591;
  assign n7593 = pi12 ? n26 : n7592;
  assign n7594 = pi11 ? n7593 : n7582;
  assign n7595 = pi10 ? n7590 : n7594;
  assign n7596 = pi09 ? n7587 : n7595;
  assign n7597 = pi08 ? n7586 : n7596;
  assign n7598 = pi07 ? n7572 : n7597;
  assign n7599 = pi09 ? n7585 : n7587;
  assign n7600 = pi09 ? n7595 : n7585;
  assign n7601 = pi08 ? n7599 : n7600;
  assign n7602 = pi13 ? n26 : n3358;
  assign n7603 = pi12 ? n26 : n7602;
  assign n7604 = pi11 ? n26 : n7603;
  assign n7605 = pi10 ? n7604 : n7603;
  assign n7606 = pi09 ? n7587 : n7605;
  assign n7607 = pi13 ? n292 : n3358;
  assign n7608 = pi12 ? n26 : n7607;
  assign n7609 = pi11 ? n7603 : n7608;
  assign n7610 = pi10 ? n7603 : n7609;
  assign n7611 = pi11 ? n7603 : n4011;
  assign n7612 = pi13 ? n3918 : n1280;
  assign n7613 = pi12 ? n26 : n7612;
  assign n7614 = pi13 ? n6376 : n1280;
  assign n7615 = pi12 ? n26 : n7614;
  assign n7616 = pi11 ? n7613 : n7615;
  assign n7617 = pi10 ? n7611 : n7616;
  assign n7618 = pi09 ? n7610 : n7617;
  assign n7619 = pi08 ? n7606 : n7618;
  assign n7620 = pi07 ? n7601 : n7619;
  assign n7621 = pi06 ? n7598 : n7620;
  assign n7622 = pi05 ? n7562 : n7621;
  assign n7623 = pi14 ? n147 : n1400;
  assign n7624 = pi13 ? n97 : n7623;
  assign n7625 = pi12 ? n26 : n7624;
  assign n7626 = pi11 ? n26 : n7625;
  assign n7627 = pi13 ? n68 : n7491;
  assign n7628 = pi12 ? n26 : n7627;
  assign n7629 = pi13 ? n68 : n7522;
  assign n7630 = pi12 ? n26 : n7629;
  assign n7631 = pi11 ? n7628 : n7630;
  assign n7632 = pi10 ? n7626 : n7631;
  assign n7633 = pi09 ? n26 : n7632;
  assign n7634 = pi08 ? n26 : n7633;
  assign n7635 = pi13 ? n68 : n233;
  assign n7636 = pi12 ? n26 : n7635;
  assign n7637 = pi13 ? n68 : n3023;
  assign n7638 = pi12 ? n26 : n7637;
  assign n7639 = pi14 ? n63 : n5885;
  assign n7640 = pi14 ? n517 : n147;
  assign n7641 = pi13 ? n7639 : n7640;
  assign n7642 = pi12 ? n26 : n7641;
  assign n7643 = pi11 ? n7638 : n7642;
  assign n7644 = pi10 ? n7636 : n7643;
  assign n7645 = pi09 ? n7644 : n7585;
  assign n7646 = pi13 ? n26 : n292;
  assign n7647 = pi12 ? n26 : n7646;
  assign n7648 = pi11 ? n7647 : n2500;
  assign n7649 = pi14 ? n7347 : n292;
  assign n7650 = pi13 ? n26 : n7649;
  assign n7651 = pi12 ? n26 : n7650;
  assign n7652 = pi10 ? n7648 : n7651;
  assign n7653 = pi13 ? n26 : n2811;
  assign n7654 = pi12 ? n26 : n7653;
  assign n7655 = pi13 ? n68 : n2315;
  assign n7656 = pi12 ? n26 : n7655;
  assign n7657 = pi11 ? n7654 : n7656;
  assign n7658 = pi13 ? n68 : n773;
  assign n7659 = pi12 ? n26 : n7658;
  assign n7660 = pi13 ? n7578 : n2498;
  assign n7661 = pi12 ? n26 : n7660;
  assign n7662 = pi11 ? n7659 : n7661;
  assign n7663 = pi10 ? n7657 : n7662;
  assign n7664 = pi09 ? n7652 : n7663;
  assign n7665 = pi08 ? n7645 : n7664;
  assign n7666 = pi07 ? n7634 : n7665;
  assign n7667 = pi09 ? n7585 : n7652;
  assign n7668 = pi14 ? n327 : n292;
  assign n7669 = pi13 ? n26 : n7668;
  assign n7670 = pi12 ? n26 : n7669;
  assign n7671 = pi11 ? n26 : n7670;
  assign n7672 = pi10 ? n26 : n7671;
  assign n7673 = pi09 ? n7663 : n7672;
  assign n7674 = pi08 ? n7667 : n7673;
  assign n7675 = pi13 ? n2519 : n7649;
  assign n7676 = pi12 ? n26 : n7675;
  assign n7677 = pi11 ? n7651 : n7676;
  assign n7678 = pi14 ? n63 : ~n168;
  assign n7679 = pi13 ? n7678 : n7649;
  assign n7680 = pi12 ? n26 : n7679;
  assign n7681 = pi13 ? n2487 : n7649;
  assign n7682 = pi12 ? n26 : n7681;
  assign n7683 = pi11 ? n7680 : n7682;
  assign n7684 = pi10 ? n7677 : n7683;
  assign n7685 = pi13 ? n1280 : n1135;
  assign n7686 = pi12 ? n26 : n7685;
  assign n7687 = pi13 ? n1280 : n2759;
  assign n7688 = pi12 ? n26 : n7687;
  assign n7689 = pi11 ? n7686 : n7688;
  assign n7690 = pi10 ? n7689 : n5908;
  assign n7691 = pi09 ? n7684 : n7690;
  assign n7692 = pi13 ? n198 : n478;
  assign n7693 = pi12 ? n26 : n7692;
  assign n7694 = pi13 ? n6253 : n478;
  assign n7695 = pi12 ? n26 : n7694;
  assign n7696 = pi13 ? n6596 : n478;
  assign n7697 = pi12 ? n26 : n7696;
  assign n7698 = pi11 ? n7695 : n7697;
  assign n7699 = pi10 ? n7693 : n7698;
  assign n7700 = pi12 ? n26 : n478;
  assign n7701 = pi14 ? n125 : ~n1400;
  assign n7702 = pi13 ? n7701 : ~n2315;
  assign n7703 = pi12 ? n69 : ~n7702;
  assign n7704 = pi11 ? n7700 : n7703;
  assign n7705 = pi14 ? n292 : n1704;
  assign n7706 = pi13 ? n130 : n7705;
  assign n7707 = pi12 ? n26 : n7706;
  assign n7708 = pi13 ? n3942 : n3023;
  assign n7709 = pi12 ? n26 : n7708;
  assign n7710 = pi11 ? n7707 : n7709;
  assign n7711 = pi10 ? n7704 : n7710;
  assign n7712 = pi09 ? n7699 : n7711;
  assign n7713 = pi08 ? n7691 : n7712;
  assign n7714 = pi07 ? n7674 : n7713;
  assign n7715 = pi06 ? n7666 : n7714;
  assign n7716 = pi11 ? n26 : n7656;
  assign n7717 = pi10 ? n7716 : n7656;
  assign n7718 = pi09 ? n26 : n7717;
  assign n7719 = pi08 ? n26 : n7718;
  assign n7720 = pi13 ? n68 : n4125;
  assign n7721 = pi12 ? n26 : n7720;
  assign n7722 = pi11 ? n7636 : n7721;
  assign n7723 = pi13 ? n2312 : n4125;
  assign n7724 = pi12 ? n26 : n7723;
  assign n7725 = pi14 ? n73 : n5885;
  assign n7726 = pi13 ? n7725 : n4125;
  assign n7727 = pi12 ? n26 : n7726;
  assign n7728 = pi11 ? n7724 : n7727;
  assign n7729 = pi10 ? n7722 : n7728;
  assign n7730 = pi10 ? n26 : n7388;
  assign n7731 = pi09 ? n7729 : n7730;
  assign n7732 = pi11 ? n7395 : n2341;
  assign n7733 = pi13 ? n26 : n2762;
  assign n7734 = pi12 ? n26 : n7733;
  assign n7735 = pi11 ? n7734 : n5908;
  assign n7736 = pi10 ? n7732 : n7735;
  assign n7737 = pi13 ? n68 : n2698;
  assign n7738 = pi12 ? n26 : n7737;
  assign n7739 = pi11 ? n7654 : n7738;
  assign n7740 = pi14 ? n26 : n5885;
  assign n7741 = pi13 ? n7740 : n2387;
  assign n7742 = pi12 ? n26 : n7741;
  assign n7743 = pi11 ? n2911 : n7742;
  assign n7744 = pi10 ? n7739 : n7743;
  assign n7745 = pi09 ? n7736 : n7744;
  assign n7746 = pi08 ? n7731 : n7745;
  assign n7747 = pi07 ? n7719 : n7746;
  assign n7748 = pi09 ? n7730 : n7736;
  assign n7749 = pi11 ? n26 : n2372;
  assign n7750 = pi10 ? n26 : n7749;
  assign n7751 = pi09 ? n7744 : n7750;
  assign n7752 = pi08 ? n7748 : n7751;
  assign n7753 = pi11 ? n2372 : n4011;
  assign n7754 = pi10 ? n2372 : n7753;
  assign n7755 = pi14 ? n125 : n517;
  assign n7756 = pi13 ? n26 : n7755;
  assign n7757 = pi12 ? n26 : n7756;
  assign n7758 = pi11 ? n4011 : n7757;
  assign n7759 = pi11 ? n5908 : n7524;
  assign n7760 = pi10 ? n7758 : n7759;
  assign n7761 = pi09 ? n7754 : n7760;
  assign n7762 = pi13 ? n2332 : n7522;
  assign n7763 = pi12 ? n26 : n7762;
  assign n7764 = pi13 ? n2698 : n7522;
  assign n7765 = pi12 ? n26 : n7764;
  assign n7766 = pi11 ? n7763 : n7765;
  assign n7767 = pi10 ? n7524 : n7766;
  assign n7768 = pi14 ? n1437 : ~n1400;
  assign n7769 = pi14 ? n73 : n291;
  assign n7770 = pi13 ? n7768 : ~n7769;
  assign n7771 = pi12 ? n124 : ~n7770;
  assign n7772 = pi11 ? n7524 : n7771;
  assign n7773 = pi13 ? n176 : n292;
  assign n7774 = pi12 ? n26 : n7773;
  assign n7775 = pi13 ? n7414 : n26;
  assign n7776 = pi12 ? n26 : n7775;
  assign n7777 = pi11 ? n7774 : n7776;
  assign n7778 = pi10 ? n7772 : n7777;
  assign n7779 = pi09 ? n7767 : n7778;
  assign n7780 = pi08 ? n7761 : n7779;
  assign n7781 = pi07 ? n7752 : n7780;
  assign n7782 = pi06 ? n7747 : n7781;
  assign n7783 = pi05 ? n7715 : n7782;
  assign n7784 = pi04 ? n7622 : n7783;
  assign n7785 = pi14 ? n233 : n1400;
  assign n7786 = pi13 ? n68 : n7785;
  assign n7787 = pi12 ? n26 : n7786;
  assign n7788 = pi11 ? n7656 : n7787;
  assign n7789 = pi10 ? n7716 : n7788;
  assign n7790 = pi09 ? n26 : n7789;
  assign n7791 = pi08 ? n26 : n7790;
  assign n7792 = pi11 ? n7659 : n2911;
  assign n7793 = pi13 ? n336 : n3023;
  assign n7794 = pi12 ? n26 : n7793;
  assign n7795 = pi13 ? n7740 : n4125;
  assign n7796 = pi12 ? n26 : n7795;
  assign n7797 = pi11 ? n7794 : n7796;
  assign n7798 = pi10 ? n7792 : n7797;
  assign n7799 = pi11 ? n26 : n2761;
  assign n7800 = pi10 ? n26 : n7799;
  assign n7801 = pi09 ? n7798 : n7800;
  assign n7802 = pi11 ? n5908 : n2761;
  assign n7803 = pi11 ? n5908 : n7654;
  assign n7804 = pi10 ? n7802 : n7803;
  assign n7805 = pi11 ? n26 : n7738;
  assign n7806 = pi10 ? n7805 : n7743;
  assign n7807 = pi09 ? n7804 : n7806;
  assign n7808 = pi08 ? n7801 : n7807;
  assign n7809 = pi07 ? n7791 : n7808;
  assign n7810 = pi09 ? n7800 : n7804;
  assign n7811 = pi11 ? n26 : n4011;
  assign n7812 = pi10 ? n26 : n7811;
  assign n7813 = pi09 ? n7806 : n7812;
  assign n7814 = pi08 ? n7810 : n7813;
  assign n7815 = pi13 ? n26 : n4460;
  assign n7816 = pi12 ? n26 : n7815;
  assign n7817 = pi11 ? n4011 : n7816;
  assign n7818 = pi11 ? n7816 : n4011;
  assign n7819 = pi10 ? n7817 : n7818;
  assign n7820 = pi09 ? n4011 : n7819;
  assign n7821 = pi14 ? n147 : n233;
  assign n7822 = pi13 ? n26 : n7821;
  assign n7823 = pi12 ? n26 : n7822;
  assign n7824 = pi13 ? n26 : n233;
  assign n7825 = pi12 ? n26 : n7824;
  assign n7826 = pi10 ? n7823 : n7825;
  assign n7827 = pi14 ? n73 : n233;
  assign n7828 = pi13 ? n68 : n7827;
  assign n7829 = pi12 ? n26 : n7828;
  assign n7830 = pi11 ? n7825 : n7829;
  assign n7831 = pi13 ? n176 : n4125;
  assign n7832 = pi12 ? n26 : n7831;
  assign n7833 = pi14 ? n517 : n233;
  assign n7834 = pi13 ? n3023 : n7833;
  assign n7835 = pi12 ? n26 : n7834;
  assign n7836 = pi11 ? n7832 : n7835;
  assign n7837 = pi10 ? n7830 : n7836;
  assign n7838 = pi09 ? n7826 : n7837;
  assign n7839 = pi08 ? n7820 : n7838;
  assign n7840 = pi07 ? n7814 : n7839;
  assign n7841 = pi06 ? n7809 : n7840;
  assign n7842 = pi13 ? n1401 : n2315;
  assign n7843 = pi12 ? n26 : n7842;
  assign n7844 = pi11 ? n26 : n7843;
  assign n7845 = pi10 ? n7844 : n7656;
  assign n7846 = pi09 ? n26 : n7845;
  assign n7847 = pi08 ? n26 : n7846;
  assign n7848 = pi15 ? n44 : n291;
  assign n7849 = pi14 ? n26 : n7848;
  assign n7850 = pi13 ? n68 : n7849;
  assign n7851 = pi12 ? n26 : n7850;
  assign n7852 = pi13 ? n77 : n3023;
  assign n7853 = pi12 ? n26 : n7852;
  assign n7854 = pi11 ? n7851 : n7853;
  assign n7855 = pi10 ? n7854 : n7797;
  assign n7856 = pi09 ? n7855 : n26;
  assign n7857 = pi08 ? n7856 : n26;
  assign n7858 = pi07 ? n7847 : n7857;
  assign n7859 = pi06 ? n7858 : n26;
  assign n7860 = pi05 ? n7841 : n7859;
  assign n7861 = pi13 ? n1401 : n478;
  assign n7862 = pi12 ? n26 : n7861;
  assign n7863 = pi11 ? n26 : n7862;
  assign n7864 = pi10 ? n7863 : n7656;
  assign n7865 = pi09 ? n26 : n7864;
  assign n7866 = pi08 ? n26 : n7865;
  assign n7867 = pi12 ? n26 : n2929;
  assign n7868 = pi11 ? n7659 : n7867;
  assign n7869 = pi10 ? n7868 : n7797;
  assign n7870 = pi09 ? n7869 : n26;
  assign n7871 = pi08 ? n7870 : n26;
  assign n7872 = pi07 ? n7866 : n7871;
  assign n7873 = pi06 ? n7872 : n26;
  assign n7874 = pi13 ? n3996 : n2498;
  assign n7875 = pi12 ? n26 : n7874;
  assign n7876 = pi14 ? n2431 : n26;
  assign n7877 = pi13 ? n7450 : n7876;
  assign n7878 = pi12 ? n26 : n7877;
  assign n7879 = pi11 ? n7875 : n7878;
  assign n7880 = pi14 ? n7848 : n26;
  assign n7881 = pi13 ? n7450 : n7880;
  assign n7882 = pi12 ? n26 : n7881;
  assign n7883 = pi13 ? n7450 : n478;
  assign n7884 = pi12 ? n26 : n7883;
  assign n7885 = pi11 ? n7882 : n7884;
  assign n7886 = pi10 ? n7879 : n7885;
  assign n7887 = pi09 ? n7869 : n7886;
  assign n7888 = pi13 ? n7450 : n2631;
  assign n7889 = pi12 ? n26 : n7888;
  assign n7890 = pi08 ? n7887 : n7889;
  assign n7891 = pi07 ? n7847 : n7890;
  assign n7892 = pi06 ? n7891 : n7889;
  assign n7893 = pi05 ? n7873 : n7892;
  assign n7894 = pi04 ? n7860 : n7893;
  assign n7895 = pi03 ? n7784 : n7894;
  assign n7896 = pi14 ? n292 : n45;
  assign n7897 = pi13 ? n68 : n7896;
  assign n7898 = pi12 ? n26 : n7897;
  assign n7899 = pi11 ? n7656 : n7898;
  assign n7900 = pi10 ? n7844 : n7899;
  assign n7901 = pi09 ? n26 : n7900;
  assign n7902 = pi08 ? n26 : n7901;
  assign n7903 = pi13 ? n1280 : n2762;
  assign n7904 = pi12 ? n26 : n7903;
  assign n7905 = pi11 ? n2638 : n7904;
  assign n7906 = pi10 ? n7613 : n7905;
  assign n7907 = pi09 ? n7869 : n7906;
  assign n7908 = pi10 ? n2664 : n3143;
  assign n7909 = pi09 ? n7908 : n3143;
  assign n7910 = pi08 ? n7907 : n7909;
  assign n7911 = pi07 ? n7902 : n7910;
  assign n7912 = pi06 ? n7911 : n3143;
  assign n7913 = pi10 ? n7863 : n7899;
  assign n7914 = pi09 ? n26 : n7913;
  assign n7915 = pi08 ? n26 : n7914;
  assign n7916 = pi11 ? n2911 : n7867;
  assign n7917 = pi13 ? n336 : n4125;
  assign n7918 = pi12 ? n26 : n7917;
  assign n7919 = pi11 ? n7918 : n7796;
  assign n7920 = pi10 ? n7916 : n7919;
  assign n7921 = pi13 ? n4809 : n198;
  assign n7922 = pi12 ? n26 : n7921;
  assign n7923 = pi13 ? n1280 : n198;
  assign n7924 = pi12 ? n26 : n7923;
  assign n7925 = pi11 ? n7922 : n7924;
  assign n7926 = pi10 ? n7613 : n7925;
  assign n7927 = pi09 ? n7920 : n7926;
  assign n7928 = pi11 ? n2664 : n7904;
  assign n7929 = pi10 ? n7928 : n3143;
  assign n7930 = pi09 ? n7929 : n3143;
  assign n7931 = pi08 ? n7927 : n7930;
  assign n7932 = pi07 ? n7915 : n7931;
  assign n7933 = pi06 ? n7932 : n3143;
  assign n7934 = pi05 ? n7912 : n7933;
  assign n7935 = pi13 ? n68 : n478;
  assign n7936 = pi12 ? n26 : n7935;
  assign n7937 = pi11 ? n26 : n7936;
  assign n7938 = pi10 ? n7937 : n7899;
  assign n7939 = pi09 ? n26 : n7938;
  assign n7940 = pi08 ? n26 : n7939;
  assign n7941 = pi13 ? n336 : n26;
  assign n7942 = pi12 ? n26 : n7941;
  assign n7943 = pi11 ? n7942 : n7742;
  assign n7944 = pi10 ? n7868 : n7943;
  assign n7945 = pi13 ? n3023 : n1280;
  assign n7946 = pi12 ? n26 : n7945;
  assign n7947 = pi13 ? n1583 : n2762;
  assign n7948 = pi12 ? n26 : n7947;
  assign n7949 = pi11 ? n7948 : n4535;
  assign n7950 = pi10 ? n7946 : n7949;
  assign n7951 = pi09 ? n7944 : n7950;
  assign n7952 = pi10 ? n7613 : n4533;
  assign n7953 = pi09 ? n7952 : n4533;
  assign n7954 = pi08 ? n7951 : n7953;
  assign n7955 = pi07 ? n7940 : n7954;
  assign n7956 = pi13 ? n6376 : n26;
  assign n7957 = pi12 ? n26 : n7956;
  assign n7958 = pi11 ? n4533 : n7957;
  assign n7959 = pi10 ? n7958 : n7957;
  assign n7960 = pi09 ? n4533 : n7959;
  assign n7961 = pi08 ? n4533 : n7960;
  assign n7962 = pi07 ? n4533 : n7961;
  assign n7963 = pi06 ? n7955 : n7962;
  assign n7964 = pi13 ? n3023 : n26;
  assign n7965 = pi12 ? n26 : n7964;
  assign n7966 = pi11 ? n26 : n7965;
  assign n7967 = pi10 ? n26 : n7966;
  assign n7968 = pi11 ? n7965 : n2561;
  assign n7969 = pi13 ? n4737 : n26;
  assign n7970 = pi12 ? n26 : n7969;
  assign n7971 = pi11 ? n7970 : n7957;
  assign n7972 = pi10 ? n7968 : n7971;
  assign n7973 = pi09 ? n7967 : n7972;
  assign n7974 = pi08 ? n26 : n7973;
  assign n7975 = pi07 ? n26 : n7974;
  assign n7976 = pi06 ? n26 : n7975;
  assign n7977 = pi05 ? n7963 : n7976;
  assign n7978 = pi04 ? n7934 : n7977;
  assign n7979 = pi14 ? n292 : n1615;
  assign n7980 = pi13 ? n7979 : n26;
  assign n7981 = pi12 ? n69 : n7980;
  assign n7982 = pi11 ? n26 : n7981;
  assign n7983 = pi10 ? n26 : n7982;
  assign n7984 = pi14 ? n292 : n152;
  assign n7985 = pi13 ? n7984 : n26;
  assign n7986 = pi12 ? n26 : n7985;
  assign n7987 = pi11 ? n5293 : n7965;
  assign n7988 = pi10 ? n7986 : n7987;
  assign n7989 = pi09 ? n7983 : n7988;
  assign n7990 = pi08 ? n26 : n7989;
  assign n7991 = pi07 ? n26 : n7990;
  assign n7992 = pi06 ? n26 : n7991;
  assign n7993 = pi09 ? n26 : n7472;
  assign n7994 = pi08 ? n26 : n7993;
  assign n7995 = pi07 ? n7994 : n7345;
  assign n7996 = pi14 ? n63 : n292;
  assign n7997 = pi13 ? n7996 : n3023;
  assign n7998 = pi12 ? n26 : n7997;
  assign n7999 = pi11 ? n7345 : n7998;
  assign n8000 = pi10 ? n7345 : n7999;
  assign n8001 = pi09 ? n7345 : n8000;
  assign n8002 = pi13 ? n3031 : n3026;
  assign n8003 = pi12 ? n26 : n8002;
  assign n8004 = pi14 ? n45 : ~n1437;
  assign n8005 = pi13 ? n8004 : n7649;
  assign n8006 = pi12 ? n26 : n8005;
  assign n8007 = pi11 ? n8003 : n8006;
  assign n8008 = pi14 ? n26 : n1615;
  assign n8009 = pi13 ? n8008 : n2698;
  assign n8010 = pi12 ? n124 : n8009;
  assign n8011 = pi11 ? n7654 : n8010;
  assign n8012 = pi10 ? n8007 : n8011;
  assign n8013 = pi13 ? n7372 : n26;
  assign n8014 = pi12 ? n26 : n8013;
  assign n8015 = pi14 ? n292 : n168;
  assign n8016 = pi13 ? n8015 : n26;
  assign n8017 = pi12 ? n26 : n8016;
  assign n8018 = pi11 ? n8014 : n8017;
  assign n8019 = pi13 ? n7431 : n26;
  assign n8020 = pi12 ? n26 : n8019;
  assign n8021 = pi11 ? n5256 : n8020;
  assign n8022 = pi10 ? n8018 : n8021;
  assign n8023 = pi09 ? n8012 : n8022;
  assign n8024 = pi08 ? n8001 : n8023;
  assign n8025 = pi07 ? n7345 : n8024;
  assign n8026 = pi06 ? n7995 : n8025;
  assign n8027 = pi05 ? n7992 : n8026;
  assign n8028 = pi11 ? n26 : n2446;
  assign n8029 = pi13 ? n1280 : n2347;
  assign n8030 = pi12 ? n26 : n8029;
  assign n8031 = pi11 ? n26 : n8030;
  assign n8032 = pi10 ? n8028 : n8031;
  assign n8033 = pi09 ? n26 : n8032;
  assign n8034 = pi13 ? n2332 : n2811;
  assign n8035 = pi12 ? n26 : n8034;
  assign n8036 = pi11 ? n26 : n8035;
  assign n8037 = pi11 ? n5908 : n7738;
  assign n8038 = pi10 ? n8036 : n8037;
  assign n8039 = pi11 ? n2911 : n26;
  assign n8040 = pi13 ? n169 : n26;
  assign n8041 = pi12 ? n26 : n8040;
  assign n8042 = pi10 ? n8039 : n8041;
  assign n8043 = pi09 ? n8038 : n8042;
  assign n8044 = pi08 ? n8033 : n8043;
  assign n8045 = pi07 ? n26 : n8044;
  assign n8046 = pi06 ? n26 : n8045;
  assign n8047 = pi09 ? n26 : n7406;
  assign n8048 = pi08 ? n26 : n8047;
  assign n8049 = pi13 ? n2498 : n639;
  assign n8050 = pi12 ? n26 : n8049;
  assign n8051 = pi11 ? n2341 : n8050;
  assign n8052 = pi10 ? n2341 : n8051;
  assign n8053 = pi09 ? n8052 : n2341;
  assign n8054 = pi08 ? n2341 : n8053;
  assign n8055 = pi07 ? n8048 : n8054;
  assign n8056 = pi11 ? n2341 : n7395;
  assign n8057 = pi10 ? n8056 : n2384;
  assign n8058 = pi09 ? n2341 : n8057;
  assign n8059 = pi13 ? n2332 : n478;
  assign n8060 = pi12 ? n26 : n8059;
  assign n8061 = pi11 ? n5908 : n8060;
  assign n8062 = pi14 ? n4950 : n26;
  assign n8063 = pi13 ? n8062 : n478;
  assign n8064 = pi12 ? n26 : n8063;
  assign n8065 = pi11 ? n8064 : n7862;
  assign n8066 = pi10 ? n8061 : n8065;
  assign n8067 = pi12 ? n124 : n2929;
  assign n8068 = pi13 ? n7896 : n26;
  assign n8069 = pi12 ? n26 : n8068;
  assign n8070 = pi11 ? n8067 : n8069;
  assign n8071 = pi12 ? n26 : n5341;
  assign n8072 = pi10 ? n8070 : n8071;
  assign n8073 = pi09 ? n8066 : n8072;
  assign n8074 = pi08 ? n8058 : n8073;
  assign n8075 = pi07 ? n2341 : n8074;
  assign n8076 = pi06 ? n8055 : n8075;
  assign n8077 = pi05 ? n8046 : n8076;
  assign n8078 = pi04 ? n8027 : n8077;
  assign n8079 = pi03 ? n7978 : n8078;
  assign n8080 = pi02 ? n7895 : n8079;
  assign n8081 = pi01 ? n7503 : n8080;
  assign n8082 = pi10 ? n7811 : n4011;
  assign n8083 = pi09 ? n26 : n8082;
  assign n8084 = pi08 ? n26 : n8083;
  assign n8085 = pi07 ? n8084 : n4011;
  assign n8086 = pi11 ? n2761 : n5908;
  assign n8087 = pi10 ? n8086 : n4011;
  assign n8088 = pi09 ? n4011 : n8087;
  assign n8089 = pi13 ? n2698 : n591;
  assign n8090 = pi12 ? n26 : n8089;
  assign n8091 = pi11 ? n2483 : n8090;
  assign n8092 = pi13 ? n2698 : n478;
  assign n8093 = pi12 ? n26 : n8092;
  assign n8094 = pi11 ? n8093 : n7936;
  assign n8095 = pi10 ? n8091 : n8094;
  assign n8096 = pi10 ? n2911 : n8071;
  assign n8097 = pi09 ? n8095 : n8096;
  assign n8098 = pi08 ? n8088 : n8097;
  assign n8099 = pi07 ? n4011 : n8098;
  assign n8100 = pi06 ? n8085 : n8099;
  assign n8101 = pi11 ? n5908 : n7508;
  assign n8102 = pi10 ? n2484 : n8101;
  assign n8103 = pi09 ? n26 : n8102;
  assign n8104 = pi08 ? n26 : n8103;
  assign n8105 = pi07 ? n26 : n8104;
  assign n8106 = pi11 ? n7508 : n26;
  assign n8107 = pi10 ? n8106 : n26;
  assign n8108 = pi09 ? n8107 : n26;
  assign n8109 = pi08 ? n8108 : n26;
  assign n8110 = pi07 ? n8109 : n26;
  assign n8111 = pi06 ? n8105 : n8110;
  assign n8112 = pi05 ? n8100 : n8111;
  assign n8113 = pi11 ? n26 : n7630;
  assign n8114 = pi11 ? n7936 : n7656;
  assign n8115 = pi10 ? n8113 : n8114;
  assign n8116 = pi09 ? n26 : n8115;
  assign n8117 = pi08 ? n26 : n8116;
  assign n8118 = pi07 ? n26 : n8117;
  assign n8119 = pi13 ? n7578 : n2403;
  assign n8120 = pi12 ? n26 : n8119;
  assign n8121 = pi11 ? n8120 : n26;
  assign n8122 = pi10 ? n8121 : n26;
  assign n8123 = pi09 ? n8122 : n26;
  assign n8124 = pi08 ? n8123 : n26;
  assign n8125 = pi07 ? n8124 : n26;
  assign n8126 = pi06 ? n8118 : n8125;
  assign n8127 = pi10 ? n7413 : n7416;
  assign n8128 = pi09 ? n26 : n8127;
  assign n8129 = pi08 ? n26 : n8128;
  assign n8130 = pi12 ? n26 : n2498;
  assign n8131 = pi11 ? n7416 : n8130;
  assign n8132 = pi13 ? n7996 : n7649;
  assign n8133 = pi12 ? n26 : n8132;
  assign n8134 = pi14 ? n7347 : n26;
  assign n8135 = pi13 ? n3031 : n8134;
  assign n8136 = pi12 ? n26 : n8135;
  assign n8137 = pi11 ? n8133 : n8136;
  assign n8138 = pi10 ? n8131 : n8137;
  assign n8139 = pi11 ? n5908 : n7656;
  assign n8140 = pi11 ? n7936 : n7638;
  assign n8141 = pi10 ? n8139 : n8140;
  assign n8142 = pi09 ? n8138 : n8141;
  assign n8143 = pi08 ? n7416 : n8142;
  assign n8144 = pi07 ? n8129 : n8143;
  assign n8145 = pi13 ? n7740 : n321;
  assign n8146 = pi12 ? n26 : n8145;
  assign n8147 = pi14 ? n63 : n1832;
  assign n8148 = pi13 ? n8147 : n26;
  assign n8149 = pi12 ? n26 : n8148;
  assign n8150 = pi11 ? n8146 : n8149;
  assign n8151 = pi14 ? n7579 : n26;
  assign n8152 = pi13 ? n7450 : n8151;
  assign n8153 = pi12 ? n26 : n8152;
  assign n8154 = pi11 ? n8153 : n7882;
  assign n8155 = pi10 ? n8150 : n8154;
  assign n8156 = pi13 ? n7450 : n6596;
  assign n8157 = pi12 ? n26 : n8156;
  assign n8158 = pi11 ? n7884 : n8157;
  assign n8159 = pi10 ? n8158 : n7889;
  assign n8160 = pi09 ? n8155 : n8159;
  assign n8161 = pi08 ? n8160 : n7889;
  assign n8162 = pi07 ? n8161 : n7889;
  assign n8163 = pi06 ? n8144 : n8162;
  assign n8164 = pi05 ? n8126 : n8163;
  assign n8165 = pi04 ? n8112 : n8164;
  assign n8166 = pi13 ? n198 : n2347;
  assign n8167 = pi12 ? n26 : n8166;
  assign n8168 = pi11 ? n8167 : n26;
  assign n8169 = pi11 ? n2664 : n7654;
  assign n8170 = pi10 ? n8168 : n8169;
  assign n8171 = pi13 ? n68 : n2498;
  assign n8172 = pi12 ? n26 : n8171;
  assign n8173 = pi11 ? n7659 : n8172;
  assign n8174 = pi10 ? n8139 : n8173;
  assign n8175 = pi09 ? n8170 : n8174;
  assign n8176 = pi08 ? n26 : n8175;
  assign n8177 = pi07 ? n26 : n8176;
  assign n8178 = pi13 ? n3942 : n2498;
  assign n8179 = pi12 ? n26 : n8178;
  assign n8180 = pi11 ? n7796 : n8179;
  assign n8181 = pi14 ? n45 : n1832;
  assign n8182 = pi13 ? n8181 : n1280;
  assign n8183 = pi12 ? n26 : n8182;
  assign n8184 = pi11 ? n8183 : n2638;
  assign n8185 = pi10 ? n8180 : n8184;
  assign n8186 = pi11 ? n7904 : n2664;
  assign n8187 = pi10 ? n8186 : n2664;
  assign n8188 = pi09 ? n8185 : n8187;
  assign n8189 = pi08 ? n8188 : n2664;
  assign n8190 = pi07 ? n8189 : n2664;
  assign n8191 = pi06 ? n8177 : n8190;
  assign n8192 = pi11 ? n26 : n7395;
  assign n8193 = pi10 ? n8192 : n7395;
  assign n8194 = pi09 ? n26 : n8193;
  assign n8195 = pi08 ? n26 : n8194;
  assign n8196 = pi10 ? n7395 : n7732;
  assign n8197 = pi09 ? n7395 : n8196;
  assign n8198 = pi10 ? n5908 : n7654;
  assign n8199 = pi13 ? n26 : n2698;
  assign n8200 = pi12 ? n26 : n8199;
  assign n8201 = pi11 ? n8200 : n7843;
  assign n8202 = pi10 ? n8201 : n7792;
  assign n8203 = pi09 ? n8198 : n8202;
  assign n8204 = pi08 ? n8197 : n8203;
  assign n8205 = pi07 ? n8195 : n8204;
  assign n8206 = pi15 ? n44 : n60;
  assign n8207 = pi14 ? n26 : n8206;
  assign n8208 = pi13 ? n8207 : n4125;
  assign n8209 = pi12 ? n26 : n8208;
  assign n8210 = pi13 ? n3023 : n2498;
  assign n8211 = pi12 ? n26 : n8210;
  assign n8212 = pi11 ? n8209 : n8211;
  assign n8213 = pi13 ? n3996 : n1280;
  assign n8214 = pi12 ? n26 : n8213;
  assign n8215 = pi13 ? n3918 : n198;
  assign n8216 = pi12 ? n26 : n8215;
  assign n8217 = pi11 ? n8214 : n8216;
  assign n8218 = pi10 ? n8212 : n8217;
  assign n8219 = pi11 ? n7924 : n7904;
  assign n8220 = pi13 ? n2598 : n2762;
  assign n8221 = pi12 ? n26 : n8220;
  assign n8222 = pi11 ? n8221 : n2606;
  assign n8223 = pi10 ? n8219 : n8222;
  assign n8224 = pi09 ? n8218 : n8223;
  assign n8225 = pi08 ? n8224 : n2606;
  assign n8226 = pi07 ? n8225 : n2606;
  assign n8227 = pi06 ? n8205 : n8226;
  assign n8228 = pi05 ? n8191 : n8227;
  assign n8229 = pi11 ? n7654 : n5908;
  assign n8230 = pi10 ? n2761 : n8229;
  assign n8231 = pi11 ? n7738 : n7936;
  assign n8232 = pi11 ? n7867 : n2911;
  assign n8233 = pi10 ? n8231 : n8232;
  assign n8234 = pi09 ? n8230 : n8233;
  assign n8235 = pi08 ? n4011 : n8234;
  assign n8236 = pi07 ? n8084 : n8235;
  assign n8237 = pi13 ? n8207 : n2387;
  assign n8238 = pi12 ? n26 : n8237;
  assign n8239 = pi13 ? n3023 : n2762;
  assign n8240 = pi12 ? n26 : n8239;
  assign n8241 = pi11 ? n8238 : n8240;
  assign n8242 = pi13 ? n1583 : n1280;
  assign n8243 = pi12 ? n26 : n8242;
  assign n8244 = pi11 ? n8243 : n4925;
  assign n8245 = pi10 ? n8241 : n8244;
  assign n8246 = pi11 ? n4925 : n7613;
  assign n8247 = pi13 ? n4809 : n1280;
  assign n8248 = pi12 ? n26 : n8247;
  assign n8249 = pi11 ? n8248 : n2664;
  assign n8250 = pi10 ? n8246 : n8249;
  assign n8251 = pi09 ? n8245 : n8250;
  assign n8252 = pi13 ? n4809 : n26;
  assign n8253 = pi12 ? n26 : n8252;
  assign n8254 = pi08 ? n8251 : n8253;
  assign n8255 = pi14 ? n1400 : n233;
  assign n8256 = pi13 ? n8255 : n26;
  assign n8257 = pi12 ? n26 : n8256;
  assign n8258 = pi11 ? n8253 : n8257;
  assign n8259 = pi10 ? n8253 : n8258;
  assign n8260 = pi09 ? n8253 : n8259;
  assign n8261 = pi08 ? n8253 : n8260;
  assign n8262 = pi07 ? n8254 : n8261;
  assign n8263 = pi06 ? n8236 : n8262;
  assign n8264 = pi11 ? n2561 : n7776;
  assign n8265 = pi10 ? n7968 : n8264;
  assign n8266 = pi09 ? n7967 : n8265;
  assign n8267 = pi08 ? n26 : n8266;
  assign n8268 = pi07 ? n26 : n8267;
  assign n8269 = pi06 ? n26 : n8268;
  assign n8270 = pi05 ? n8263 : n8269;
  assign n8271 = pi04 ? n8228 : n8270;
  assign n8272 = pi03 ? n8165 : n8271;
  assign n8273 = pi13 ? n8008 : n26;
  assign n8274 = pi12 ? n69 : n8273;
  assign n8275 = pi11 ? n26 : n8274;
  assign n8276 = pi10 ? n26 : n8275;
  assign n8277 = pi11 ? n5256 : n7986;
  assign n8278 = pi10 ? n8277 : n7987;
  assign n8279 = pi09 ? n8276 : n8278;
  assign n8280 = pi08 ? n26 : n8279;
  assign n8281 = pi07 ? n26 : n8280;
  assign n8282 = pi06 ? n26 : n8281;
  assign n8283 = pi05 ? n8282 : n8026;
  assign n8284 = pi07 ? n8048 : n2341;
  assign n8285 = pi06 ? n8284 : n8075;
  assign n8286 = pi05 ? n8046 : n8285;
  assign n8287 = pi04 ? n8283 : n8286;
  assign n8288 = pi10 ? n7811 : n5908;
  assign n8289 = pi09 ? n26 : n8288;
  assign n8290 = pi08 ? n26 : n8289;
  assign n8291 = pi07 ? n8290 : n4011;
  assign n8292 = pi06 ? n8291 : n8099;
  assign n8293 = pi14 ? n147 : n292;
  assign n8294 = pi13 ? n26 : n8293;
  assign n8295 = pi12 ? n26 : n8294;
  assign n8296 = pi11 ? n26 : n8295;
  assign n8297 = pi10 ? n8296 : n5908;
  assign n8298 = pi09 ? n26 : n8297;
  assign n8299 = pi08 ? n26 : n8298;
  assign n8300 = pi10 ? n7508 : n26;
  assign n8301 = pi09 ? n8300 : n26;
  assign n8302 = pi08 ? n8301 : n26;
  assign n8303 = pi07 ? n8299 : n8302;
  assign n8304 = pi06 ? n8303 : n26;
  assign n8305 = pi05 ? n8292 : n8304;
  assign n8306 = pi13 ? n97 : n7491;
  assign n8307 = pi12 ? n26 : n8306;
  assign n8308 = pi11 ? n26 : n8307;
  assign n8309 = pi10 ? n8308 : n5132;
  assign n8310 = pi09 ? n26 : n8309;
  assign n8311 = pi08 ? n26 : n8310;
  assign n8312 = pi11 ? n7656 : n8120;
  assign n8313 = pi10 ? n8312 : n26;
  assign n8314 = pi09 ? n8313 : n26;
  assign n8315 = pi08 ? n8314 : n26;
  assign n8316 = pi07 ? n8311 : n8315;
  assign n8317 = pi06 ? n8316 : n26;
  assign n8318 = pi11 ? n26 : n7787;
  assign n8319 = pi14 ? n37 : ~n1400;
  assign n8320 = pi13 ? n68 : ~n8319;
  assign n8321 = pi12 ? n26 : n8320;
  assign n8322 = pi11 ? n5577 : n8321;
  assign n8323 = pi10 ? n8318 : n8322;
  assign n8324 = pi09 ? n26 : n8323;
  assign n8325 = pi08 ? n26 : n8324;
  assign n8326 = pi14 ? n517 : n320;
  assign n8327 = pi13 ? n7740 : n8326;
  assign n8328 = pi12 ? n26 : n8327;
  assign n8329 = pi11 ? n2911 : n8328;
  assign n8330 = pi13 ? n8147 : n1280;
  assign n8331 = pi12 ? n26 : n8330;
  assign n8332 = pi11 ? n8331 : n7878;
  assign n8333 = pi10 ? n8329 : n8332;
  assign n8334 = pi10 ? n7885 : n7889;
  assign n8335 = pi09 ? n8333 : n8334;
  assign n8336 = pi08 ? n8335 : n7889;
  assign n8337 = pi07 ? n8325 : n8336;
  assign n8338 = pi06 ? n8337 : n7889;
  assign n8339 = pi05 ? n8317 : n8338;
  assign n8340 = pi04 ? n8305 : n8339;
  assign n8341 = pi03 ? n8287 : n8340;
  assign n8342 = pi02 ? n8272 : n8341;
  assign n8343 = pi11 ? n7656 : n7659;
  assign n8344 = pi10 ? n7844 : n8343;
  assign n8345 = pi09 ? n26 : n8344;
  assign n8346 = pi08 ? n26 : n8345;
  assign n8347 = pi13 ? n3942 : n1280;
  assign n8348 = pi12 ? n26 : n8347;
  assign n8349 = pi11 ? n8348 : n8183;
  assign n8350 = pi10 ? n7797 : n8349;
  assign n8351 = pi10 ? n7905 : n2664;
  assign n8352 = pi09 ? n8350 : n8351;
  assign n8353 = pi08 ? n8352 : n2664;
  assign n8354 = pi07 ? n8346 : n8353;
  assign n8355 = pi06 ? n8354 : n2664;
  assign n8356 = pi14 ? n26 : n291;
  assign n8357 = pi13 ? n68 : n8356;
  assign n8358 = pi12 ? n26 : n8357;
  assign n8359 = pi11 ? n3565 : n8358;
  assign n8360 = pi10 ? n7844 : n8359;
  assign n8361 = pi09 ? n26 : n8360;
  assign n8362 = pi08 ? n26 : n8361;
  assign n8363 = pi11 ? n7946 : n8214;
  assign n8364 = pi10 ? n7797 : n8363;
  assign n8365 = pi13 ? n2391 : n198;
  assign n8366 = pi12 ? n26 : n8365;
  assign n8367 = pi11 ? n4533 : n8366;
  assign n8368 = pi11 ? n7904 : n8221;
  assign n8369 = pi10 ? n8367 : n8368;
  assign n8370 = pi09 ? n8364 : n8369;
  assign n8371 = pi08 ? n8370 : n2606;
  assign n8372 = pi07 ? n8362 : n8371;
  assign n8373 = pi06 ? n8372 : n2606;
  assign n8374 = pi05 ? n8355 : n8373;
  assign n8375 = pi10 ? n7716 : n7868;
  assign n8376 = pi09 ? n26 : n8375;
  assign n8377 = pi08 ? n26 : n8376;
  assign n8378 = pi13 ? n3023 : n7423;
  assign n8379 = pi12 ? n26 : n8378;
  assign n8380 = pi13 ? n3023 : n3031;
  assign n8381 = pi12 ? n26 : n8380;
  assign n8382 = pi11 ? n8379 : n8381;
  assign n8383 = pi10 ? n7797 : n8382;
  assign n8384 = pi10 ? n4925 : n7613;
  assign n8385 = pi09 ? n8383 : n8384;
  assign n8386 = pi11 ? n2664 : n8253;
  assign n8387 = pi10 ? n8386 : n8253;
  assign n8388 = pi09 ? n8387 : n8253;
  assign n8389 = pi08 ? n8385 : n8388;
  assign n8390 = pi07 ? n8377 : n8389;
  assign n8391 = pi13 ? n4809 : n2762;
  assign n8392 = pi12 ? n26 : n8391;
  assign n8393 = pi11 ? n8392 : n8253;
  assign n8394 = pi10 ? n8393 : n8253;
  assign n8395 = pi09 ? n8394 : n8253;
  assign n8396 = pi08 ? n8253 : n8395;
  assign n8397 = pi07 ? n8396 : n8253;
  assign n8398 = pi06 ? n8390 : n8397;
  assign n8399 = pi10 ? n26 : n7965;
  assign n8400 = pi10 ? n2561 : n26;
  assign n8401 = pi09 ? n8399 : n8400;
  assign n8402 = pi08 ? n8401 : n26;
  assign n8403 = pi07 ? n8402 : n26;
  assign n8404 = pi06 ? n26 : n8403;
  assign n8405 = pi05 ? n8398 : n8404;
  assign n8406 = pi04 ? n8374 : n8405;
  assign n8407 = pi11 ? n8274 : n5256;
  assign n8408 = pi10 ? n26 : n8407;
  assign n8409 = pi11 ? n5256 : n7776;
  assign n8410 = pi10 ? n8409 : n26;
  assign n8411 = pi09 ? n8408 : n8410;
  assign n8412 = pi08 ? n8411 : n26;
  assign n8413 = pi07 ? n8412 : n26;
  assign n8414 = pi06 ? n26 : n8413;
  assign n8415 = pi13 ? n3031 : n7649;
  assign n8416 = pi12 ? n26 : n8415;
  assign n8417 = pi11 ? n7998 : n8416;
  assign n8418 = pi10 ? n7416 : n8417;
  assign n8419 = pi09 ? n7416 : n8418;
  assign n8420 = pi08 ? n7416 : n8419;
  assign n8421 = pi07 ? n8129 : n8420;
  assign n8422 = pi13 ? n2631 : n2811;
  assign n8423 = pi12 ? n26 : n8422;
  assign n8424 = pi11 ? n8006 : n8423;
  assign n8425 = pi14 ? n292 : n4243;
  assign n8426 = pi13 ? n8425 : n26;
  assign n8427 = pi12 ? n26 : n8426;
  assign n8428 = pi11 ? n8010 : n8427;
  assign n8429 = pi10 ? n8424 : n8428;
  assign n8430 = pi14 ? n7577 : n26;
  assign n8431 = pi13 ? n8430 : n8151;
  assign n8432 = pi12 ? n26 : n8431;
  assign n8433 = pi11 ? n2446 : n8432;
  assign n8434 = pi10 ? n5256 : n8433;
  assign n8435 = pi09 ? n8429 : n8434;
  assign n8436 = pi09 ? n8159 : n7889;
  assign n8437 = pi08 ? n8435 : n8436;
  assign n8438 = pi07 ? n8437 : n7889;
  assign n8439 = pi06 ? n8421 : n8438;
  assign n8440 = pi05 ? n8414 : n8439;
  assign n8441 = pi11 ? n2446 : n7395;
  assign n8442 = pi11 ? n2664 : n7734;
  assign n8443 = pi10 ? n8441 : n8442;
  assign n8444 = pi09 ? n26 : n8443;
  assign n8445 = pi08 ? n26 : n8444;
  assign n8446 = pi07 ? n26 : n8445;
  assign n8447 = pi11 ? n8035 : n5908;
  assign n8448 = pi11 ? n7738 : n8069;
  assign n8449 = pi10 ? n8447 : n8448;
  assign n8450 = pi11 ? n8071 : n8041;
  assign n8451 = pi13 ? n3942 : n26;
  assign n8452 = pi12 ? n26 : n8451;
  assign n8453 = pi11 ? n8452 : n8183;
  assign n8454 = pi10 ? n8450 : n8453;
  assign n8455 = pi09 ? n8449 : n8454;
  assign n8456 = pi09 ? n8187 : n2664;
  assign n8457 = pi08 ? n8455 : n8456;
  assign n8458 = pi07 ? n8457 : n2664;
  assign n8459 = pi06 ? n8446 : n8458;
  assign n8460 = pi10 ? n8056 : n5908;
  assign n8461 = pi09 ? n7395 : n8460;
  assign n8462 = pi08 ? n7395 : n8461;
  assign n8463 = pi07 ? n8195 : n8462;
  assign n8464 = pi14 ? n4243 : n26;
  assign n8465 = pi13 ? n8464 : n478;
  assign n8466 = pi12 ? n26 : n8465;
  assign n8467 = pi11 ? n8466 : n8093;
  assign n8468 = pi11 ? n7862 : n8067;
  assign n8469 = pi10 ? n8467 : n8468;
  assign n8470 = pi13 ? n3996 : n2762;
  assign n8471 = pi12 ? n26 : n8470;
  assign n8472 = pi11 ? n7965 : n8471;
  assign n8473 = pi10 ? n8071 : n8472;
  assign n8474 = pi09 ? n8469 : n8473;
  assign n8475 = pi11 ? n7613 : n2393;
  assign n8476 = pi11 ? n7904 : n2606;
  assign n8477 = pi10 ? n8475 : n8476;
  assign n8478 = pi09 ? n8477 : n2606;
  assign n8479 = pi08 ? n8474 : n8478;
  assign n8480 = pi07 ? n8479 : n2606;
  assign n8481 = pi06 ? n8463 : n8480;
  assign n8482 = pi05 ? n8459 : n8481;
  assign n8483 = pi04 ? n8440 : n8482;
  assign n8484 = pi03 ? n8406 : n8483;
  assign n8485 = pi10 ? n7604 : n4011;
  assign n8486 = pi09 ? n26 : n8485;
  assign n8487 = pi08 ? n26 : n8486;
  assign n8488 = pi10 ? n8086 : n2483;
  assign n8489 = pi09 ? n4011 : n8488;
  assign n8490 = pi08 ? n4011 : n8489;
  assign n8491 = pi07 ? n8487 : n8490;
  assign n8492 = pi11 ? n7936 : n2911;
  assign n8493 = pi10 ? n5908 : n8492;
  assign n8494 = pi11 ? n2911 : n8071;
  assign n8495 = pi11 ? n8240 : n7946;
  assign n8496 = pi10 ? n8494 : n8495;
  assign n8497 = pi09 ? n8493 : n8496;
  assign n8498 = pi13 ? n8181 : n2762;
  assign n8499 = pi12 ? n26 : n8498;
  assign n8500 = pi11 ? n8183 : n4533;
  assign n8501 = pi10 ? n8499 : n8500;
  assign n8502 = pi09 ? n8501 : n8387;
  assign n8503 = pi08 ? n8497 : n8502;
  assign n8504 = pi07 ? n8503 : n8253;
  assign n8505 = pi06 ? n8491 : n8504;
  assign n8506 = pi10 ? n7525 : n5908;
  assign n8507 = pi09 ? n26 : n8506;
  assign n8508 = pi08 ? n26 : n8507;
  assign n8509 = pi07 ? n8508 : n8302;
  assign n8510 = pi06 ? n8509 : n26;
  assign n8511 = pi05 ? n8505 : n8510;
  assign n8512 = pi13 ? n97 : ~n38;
  assign n8513 = pi12 ? n26 : n8512;
  assign n8514 = pi14 ? n37 : ~n292;
  assign n8515 = pi13 ? n26 : ~n8514;
  assign n8516 = pi12 ? n26 : n8515;
  assign n8517 = pi11 ? n8513 : n8516;
  assign n8518 = pi10 ? n8308 : n8517;
  assign n8519 = pi09 ? n26 : n8518;
  assign n8520 = pi08 ? n26 : n8519;
  assign n8521 = pi07 ? n8520 : n8315;
  assign n8522 = pi06 ? n8521 : n26;
  assign n8523 = pi13 ? n7740 : n7640;
  assign n8524 = pi12 ? n26 : n8523;
  assign n8525 = pi11 ? n7638 : n8524;
  assign n8526 = pi10 ? n8525 : n8332;
  assign n8527 = pi13 ? n7450 : n6164;
  assign n8528 = pi12 ? n26 : n8527;
  assign n8529 = pi11 ? n7889 : n8528;
  assign n8530 = pi10 ? n7885 : n8529;
  assign n8531 = pi09 ? n8526 : n8530;
  assign n8532 = pi10 ? n8157 : n7889;
  assign n8533 = pi09 ? n8532 : n7889;
  assign n8534 = pi08 ? n8531 : n8533;
  assign n8535 = pi07 ? n8325 : n8534;
  assign n8536 = pi06 ? n8535 : n7889;
  assign n8537 = pi05 ? n8522 : n8536;
  assign n8538 = pi04 ? n8511 : n8537;
  assign n8539 = pi11 ? n7638 : n7796;
  assign n8540 = pi13 ? n8181 : n2741;
  assign n8541 = pi12 ? n26 : n8540;
  assign n8542 = pi11 ? n8348 : n8541;
  assign n8543 = pi10 ? n8539 : n8542;
  assign n8544 = pi13 ? n2598 : n7880;
  assign n8545 = pi12 ? n26 : n8544;
  assign n8546 = pi11 ? n7688 : n8545;
  assign n8547 = pi10 ? n8546 : n2606;
  assign n8548 = pi09 ? n8543 : n8547;
  assign n8549 = pi08 ? n8548 : n2606;
  assign n8550 = pi07 ? n8346 : n8549;
  assign n8551 = pi06 ? n8550 : n2606;
  assign n8552 = pi11 ? n7946 : n8183;
  assign n8553 = pi10 ? n7797 : n8552;
  assign n8554 = pi11 ? n8499 : n8366;
  assign n8555 = pi10 ? n8554 : n8186;
  assign n8556 = pi09 ? n8553 : n8555;
  assign n8557 = pi08 ? n8556 : n2664;
  assign n8558 = pi07 ? n8362 : n8557;
  assign n8559 = pi06 ? n8558 : n2664;
  assign n8560 = pi05 ? n8551 : n8559;
  assign n8561 = pi10 ? n7844 : n7868;
  assign n8562 = pi09 ? n26 : n8561;
  assign n8563 = pi08 ? n26 : n8562;
  assign n8564 = pi11 ? n8216 : n5258;
  assign n8565 = pi10 ? n4533 : n8564;
  assign n8566 = pi09 ? n8383 : n8565;
  assign n8567 = pi10 ? n8186 : n2393;
  assign n8568 = pi09 ? n8567 : n2393;
  assign n8569 = pi08 ? n8566 : n8568;
  assign n8570 = pi07 ? n8563 : n8569;
  assign n8571 = pi06 ? n8570 : n2393;
  assign n8572 = pi13 ? n3023 : n4809;
  assign n8573 = pi12 ? n26 : n8572;
  assign n8574 = pi11 ? n8573 : n7946;
  assign n8575 = pi10 ? n7943 : n8574;
  assign n8576 = pi10 ? n4926 : n8246;
  assign n8577 = pi09 ? n8575 : n8576;
  assign n8578 = pi10 ? n8248 : n4533;
  assign n8579 = pi09 ? n8578 : n4533;
  assign n8580 = pi08 ? n8577 : n8579;
  assign n8581 = pi07 ? n8377 : n8580;
  assign n8582 = pi06 ? n8581 : n4533;
  assign n8583 = pi05 ? n8571 : n8582;
  assign n8584 = pi04 ? n8560 : n8583;
  assign n8585 = pi03 ? n8538 : n8584;
  assign n8586 = pi02 ? n8484 : n8585;
  assign n8587 = pi01 ? n8342 : n8586;
  assign n8588 = pi00 ? n8081 : n8587;
  assign n8589 = pi13 ? n169 : n30;
  assign n8590 = pi12 ? n26 : n8589;
  assign n8591 = pi11 ? n26 : n8590;
  assign n8592 = pi13 ? n169 : ~n26;
  assign n8593 = pi12 ? n26 : n8592;
  assign n8594 = pi10 ? n8591 : n8593;
  assign n8595 = pi09 ? n26 : n8594;
  assign n8596 = pi08 ? n26 : n8595;
  assign n8597 = pi12 ? n26 : n135;
  assign n8598 = pi11 ? n8593 : n8597;
  assign n8599 = pi13 ? n176 : ~n26;
  assign n8600 = pi12 ? n26 : n8599;
  assign n8601 = pi11 ? n8597 : n8600;
  assign n8602 = pi10 ? n8598 : n8601;
  assign n8603 = pi12 ? n26 : n273;
  assign n8604 = pi11 ? n8600 : n8603;
  assign n8605 = pi12 ? n26 : n212;
  assign n8606 = pi11 ? n8603 : n8605;
  assign n8607 = pi10 ? n8604 : n8606;
  assign n8608 = pi09 ? n8602 : n8607;
  assign n8609 = pi11 ? n335 : n1373;
  assign n8610 = pi10 ? n8609 : n26;
  assign n8611 = pi13 ? n130 : n30;
  assign n8612 = pi12 ? n26 : n8611;
  assign n8613 = pi11 ? n26 : n8612;
  assign n8614 = pi10 ? n8613 : n8601;
  assign n8615 = pi09 ? n8610 : n8614;
  assign n8616 = pi08 ? n8608 : n8615;
  assign n8617 = pi07 ? n8596 : n8616;
  assign n8618 = pi09 ? n8607 : n8610;
  assign n8619 = pi09 ? n8614 : n8607;
  assign n8620 = pi08 ? n8618 : n8619;
  assign n8621 = pi09 ? n8610 : n8594;
  assign n8622 = pi14 ? n60 : n168;
  assign n8623 = pi13 ? n8622 : ~n97;
  assign n8624 = pi12 ? n26 : n8623;
  assign n8625 = pi11 ? n8593 : n8624;
  assign n8626 = pi14 ? n71 : ~n1615;
  assign n8627 = pi14 ? n26 : ~n73;
  assign n8628 = pi13 ? n8626 : n8627;
  assign n8629 = pi12 ? n69 : ~n8628;
  assign n8630 = pi13 ? n1344 : n240;
  assign n8631 = pi12 ? n78 : ~n8630;
  assign n8632 = pi11 ? n8629 : n8631;
  assign n8633 = pi10 ? n8625 : n8632;
  assign n8634 = pi09 ? n8593 : n8633;
  assign n8635 = pi08 ? n8621 : n8634;
  assign n8636 = pi07 ? n8620 : n8635;
  assign n8637 = pi06 ? n8617 : n8636;
  assign n8638 = pi05 ? n26 : n8637;
  assign n8639 = pi12 ? n26 : n3697;
  assign n8640 = pi11 ? n26 : n8639;
  assign n8641 = pi11 ? n8639 : n8593;
  assign n8642 = pi10 ? n8640 : n8641;
  assign n8643 = pi09 ? n26 : n8642;
  assign n8644 = pi08 ? n26 : n8643;
  assign n8645 = pi11 ? n99 : n731;
  assign n8646 = pi10 ? n8645 : n26;
  assign n8647 = pi11 ? n26 : n8597;
  assign n8648 = pi10 ? n8647 : n8601;
  assign n8649 = pi09 ? n8646 : n8648;
  assign n8650 = pi08 ? n8608 : n8649;
  assign n8651 = pi07 ? n8644 : n8650;
  assign n8652 = pi09 ? n8607 : n8646;
  assign n8653 = pi09 ? n8648 : n8607;
  assign n8654 = pi08 ? n8652 : n8653;
  assign n8655 = pi10 ? n8640 : n8639;
  assign n8656 = pi09 ? n8646 : n8655;
  assign n8657 = pi13 ? n240 : ~n26;
  assign n8658 = pi12 ? n26 : n8657;
  assign n8659 = pi12 ? n26 : n80;
  assign n8660 = pi11 ? n8658 : n8659;
  assign n8661 = pi10 ? n8639 : n8660;
  assign n8662 = pi12 ? n26 : n1268;
  assign n8663 = pi12 ? n124 : ~n26;
  assign n8664 = pi11 ? n8662 : n8663;
  assign n8665 = pi12 ? n78 : ~n69;
  assign n8666 = pi13 ? n4125 : n57;
  assign n8667 = pi12 ? n78 : ~n8666;
  assign n8668 = pi11 ? n8665 : n8667;
  assign n8669 = pi10 ? n8664 : n8668;
  assign n8670 = pi09 ? n8661 : n8669;
  assign n8671 = pi08 ? n8656 : n8670;
  assign n8672 = pi07 ? n8654 : n8671;
  assign n8673 = pi06 ? n8651 : n8672;
  assign n8674 = pi11 ? n8658 : n8639;
  assign n8675 = pi10 ? n8640 : n8674;
  assign n8676 = pi09 ? n26 : n8675;
  assign n8677 = pi08 ? n26 : n8676;
  assign n8678 = pi10 ? n8641 : n8598;
  assign n8679 = pi10 ? n8601 : n8603;
  assign n8680 = pi09 ? n8678 : n8679;
  assign n8681 = pi11 ? n8605 : n335;
  assign n8682 = pi10 ? n8681 : n26;
  assign n8683 = pi11 ? n26 : n8593;
  assign n8684 = pi10 ? n8683 : n8598;
  assign n8685 = pi09 ? n8682 : n8684;
  assign n8686 = pi08 ? n8680 : n8685;
  assign n8687 = pi07 ? n8677 : n8686;
  assign n8688 = pi09 ? n8679 : n8682;
  assign n8689 = pi09 ? n8684 : n8679;
  assign n8690 = pi08 ? n8688 : n8689;
  assign n8691 = pi11 ? n26 : n8658;
  assign n8692 = pi10 ? n8691 : n8658;
  assign n8693 = pi09 ? n8682 : n8692;
  assign n8694 = pi11 ? n8659 : n8662;
  assign n8695 = pi10 ? n8660 : n8694;
  assign n8696 = pi12 ? n26 : n3411;
  assign n8697 = pi12 ? n69 : ~n26;
  assign n8698 = pi11 ? n8696 : n8697;
  assign n8699 = pi12 ? n78 : ~n124;
  assign n8700 = pi13 ? n26 : n176;
  assign n8701 = pi12 ? n78 : ~n8700;
  assign n8702 = pi11 ? n8699 : n8701;
  assign n8703 = pi10 ? n8698 : n8702;
  assign n8704 = pi09 ? n8695 : n8703;
  assign n8705 = pi08 ? n8693 : n8704;
  assign n8706 = pi07 ? n8690 : n8705;
  assign n8707 = pi06 ? n8687 : n8706;
  assign n8708 = pi05 ? n8673 : n8707;
  assign n8709 = pi04 ? n8638 : n8708;
  assign n8710 = pi03 ? n26 : n8709;
  assign n8711 = pi02 ? n26 : n8710;
  assign n8712 = pi09 ? n26 : n8692;
  assign n8713 = pi08 ? n26 : n8712;
  assign n8714 = pi10 ? n8674 : n8598;
  assign n8715 = pi11 ? n26 : n8600;
  assign n8716 = pi10 ? n26 : n8715;
  assign n8717 = pi09 ? n8714 : n8716;
  assign n8718 = pi13 ? n77 : ~n97;
  assign n8719 = pi12 ? n26 : n8718;
  assign n8720 = pi11 ? n8600 : n8719;
  assign n8721 = pi10 ? n8720 : n26;
  assign n8722 = pi09 ? n8721 : n8684;
  assign n8723 = pi08 ? n8717 : n8722;
  assign n8724 = pi07 ? n8713 : n8723;
  assign n8725 = pi09 ? n8716 : n8721;
  assign n8726 = pi09 ? n8684 : n8716;
  assign n8727 = pi08 ? n8725 : n8726;
  assign n8728 = pi11 ? n26 : n8659;
  assign n8729 = pi10 ? n8728 : n8659;
  assign n8730 = pi09 ? n8721 : n8729;
  assign n8731 = pi13 ? n30 : ~n26;
  assign n8732 = pi12 ? n26 : n8731;
  assign n8733 = pi11 ? n8662 : n8732;
  assign n8734 = pi10 ? n8694 : n8733;
  assign n8735 = pi12 ? n26 : n2909;
  assign n8736 = pi12 ? n78 : ~n26;
  assign n8737 = pi11 ? n8735 : n8736;
  assign n8738 = pi13 ? n26 : n143;
  assign n8739 = pi12 ? n78 : ~n8738;
  assign n8740 = pi11 ? n8736 : n8739;
  assign n8741 = pi10 ? n8737 : n8740;
  assign n8742 = pi09 ? n8734 : n8741;
  assign n8743 = pi08 ? n8730 : n8742;
  assign n8744 = pi07 ? n8727 : n8743;
  assign n8745 = pi06 ? n8724 : n8744;
  assign n8746 = pi09 ? n26 : n8729;
  assign n8747 = pi08 ? n26 : n8746;
  assign n8748 = pi11 ? n8659 : n8658;
  assign n8749 = pi13 ? n169 : ~n97;
  assign n8750 = pi12 ? n26 : n8749;
  assign n8751 = pi11 ? n8639 : n8750;
  assign n8752 = pi10 ? n8748 : n8751;
  assign n8753 = pi10 ? n26 : n8683;
  assign n8754 = pi09 ? n8752 : n8753;
  assign n8755 = pi10 ? n8597 : n26;
  assign n8756 = pi10 ? n8683 : n8751;
  assign n8757 = pi09 ? n8755 : n8756;
  assign n8758 = pi08 ? n8754 : n8757;
  assign n8759 = pi07 ? n8747 : n8758;
  assign n8760 = pi09 ? n8753 : n8755;
  assign n8761 = pi09 ? n8756 : n8753;
  assign n8762 = pi08 ? n8760 : n8761;
  assign n8763 = pi11 ? n26 : n8662;
  assign n8764 = pi10 ? n8763 : n8662;
  assign n8765 = pi09 ? n8755 : n8764;
  assign n8766 = pi13 ? n38 : ~n26;
  assign n8767 = pi12 ? n26 : n8766;
  assign n8768 = pi11 ? n8662 : n8767;
  assign n8769 = pi11 ? n8767 : n8696;
  assign n8770 = pi10 ? n8768 : n8769;
  assign n8771 = pi09 ? n8770 : n8741;
  assign n8772 = pi08 ? n8765 : n8771;
  assign n8773 = pi07 ? n8762 : n8772;
  assign n8774 = pi06 ? n8759 : n8773;
  assign n8775 = pi05 ? n8745 : n8774;
  assign n8776 = pi09 ? n26 : n8764;
  assign n8777 = pi08 ? n26 : n8776;
  assign n8778 = pi13 ? n79 : ~n97;
  assign n8779 = pi12 ? n26 : n8778;
  assign n8780 = pi13 ? n240 : ~n68;
  assign n8781 = pi12 ? n26 : n8780;
  assign n8782 = pi11 ? n8779 : n8781;
  assign n8783 = pi10 ? n8662 : n8782;
  assign n8784 = pi10 ? n26 : n8640;
  assign n8785 = pi09 ? n8783 : n8784;
  assign n8786 = pi13 ? n57 : ~n97;
  assign n8787 = pi12 ? n26 : n8786;
  assign n8788 = pi13 ? n169 : ~n68;
  assign n8789 = pi12 ? n26 : n8788;
  assign n8790 = pi11 ? n8787 : n8789;
  assign n8791 = pi10 ? n8639 : n8790;
  assign n8792 = pi09 ? n8639 : n8791;
  assign n8793 = pi08 ? n8785 : n8792;
  assign n8794 = pi07 ? n8777 : n8793;
  assign n8795 = pi09 ? n8784 : n8639;
  assign n8796 = pi09 ? n8791 : n8784;
  assign n8797 = pi08 ? n8795 : n8796;
  assign n8798 = pi10 ? n8768 : n8767;
  assign n8799 = pi09 ? n8661 : n8798;
  assign n8800 = pi11 ? n8732 : n8696;
  assign n8801 = pi10 ? n8767 : n8800;
  assign n8802 = pi11 ? n8735 : n8697;
  assign n8803 = pi11 ? n8699 : n8739;
  assign n8804 = pi10 ? n8802 : n8803;
  assign n8805 = pi09 ? n8801 : n8804;
  assign n8806 = pi08 ? n8799 : n8805;
  assign n8807 = pi07 ? n8797 : n8806;
  assign n8808 = pi06 ? n8794 : n8807;
  assign n8809 = pi11 ? n26 : n8767;
  assign n8810 = pi10 ? n8809 : n8767;
  assign n8811 = pi09 ? n26 : n8810;
  assign n8812 = pi08 ? n26 : n8811;
  assign n8813 = pi13 ? n30 : ~n97;
  assign n8814 = pi12 ? n26 : n8813;
  assign n8815 = pi13 ? n30 : ~n77;
  assign n8816 = pi12 ? n26 : n8815;
  assign n8817 = pi11 ? n8814 : n8816;
  assign n8818 = pi10 ? n8767 : n8817;
  assign n8819 = pi10 ? n26 : n8691;
  assign n8820 = pi09 ? n8818 : n8819;
  assign n8821 = pi13 ? n240 : ~n97;
  assign n8822 = pi12 ? n26 : n8821;
  assign n8823 = pi13 ? n57 : ~n77;
  assign n8824 = pi12 ? n26 : n8823;
  assign n8825 = pi11 ? n8822 : n8824;
  assign n8826 = pi10 ? n8658 : n8825;
  assign n8827 = pi09 ? n8658 : n8826;
  assign n8828 = pi08 ? n8820 : n8827;
  assign n8829 = pi07 ? n8812 : n8828;
  assign n8830 = pi09 ? n8819 : n8658;
  assign n8831 = pi09 ? n8826 : n8819;
  assign n8832 = pi08 ? n8830 : n8831;
  assign n8833 = pi11 ? n8767 : n8732;
  assign n8834 = pi10 ? n8767 : n8833;
  assign n8835 = pi09 ? n8695 : n8834;
  assign n8836 = pi11 ? n8696 : n8735;
  assign n8837 = pi10 ? n8800 : n8836;
  assign n8838 = pi12 ? n124 : ~n124;
  assign n8839 = pi11 ? n8735 : n8838;
  assign n8840 = pi12 ? n69 : ~n69;
  assign n8841 = pi11 ? n8840 : n8739;
  assign n8842 = pi10 ? n8839 : n8841;
  assign n8843 = pi09 ? n8837 : n8842;
  assign n8844 = pi08 ? n8835 : n8843;
  assign n8845 = pi07 ? n8832 : n8844;
  assign n8846 = pi06 ? n8829 : n8845;
  assign n8847 = pi05 ? n8808 : n8846;
  assign n8848 = pi04 ? n8775 : n8847;
  assign n8849 = pi10 ? n8809 : n8833;
  assign n8850 = pi09 ? n26 : n8849;
  assign n8851 = pi08 ? n26 : n8850;
  assign n8852 = pi13 ? n126 : ~n97;
  assign n8853 = pi12 ? n26 : n8852;
  assign n8854 = pi11 ? n8732 : n8853;
  assign n8855 = pi13 ? n126 : ~n68;
  assign n8856 = pi12 ? n26 : n8855;
  assign n8857 = pi13 ? n507 : ~n77;
  assign n8858 = pi12 ? n26 : n8857;
  assign n8859 = pi11 ? n8856 : n8858;
  assign n8860 = pi10 ? n8854 : n8859;
  assign n8861 = pi13 ? n5528 : ~n4125;
  assign n8862 = pi12 ? n26 : n8861;
  assign n8863 = pi11 ? n26 : n8862;
  assign n8864 = pi10 ? n26 : n8863;
  assign n8865 = pi09 ? n8860 : n8864;
  assign n8866 = pi11 ? n8659 : n8779;
  assign n8867 = pi13 ? n79 : ~n68;
  assign n8868 = pi12 ? n26 : n8867;
  assign n8869 = pi14 ? n1355 : n71;
  assign n8870 = pi13 ? n240 : ~n8869;
  assign n8871 = pi12 ? n26 : n8870;
  assign n8872 = pi11 ? n8868 : n8871;
  assign n8873 = pi10 ? n8866 : n8872;
  assign n8874 = pi09 ? n8659 : n8873;
  assign n8875 = pi08 ? n8865 : n8874;
  assign n8876 = pi07 ? n8851 : n8875;
  assign n8877 = pi09 ? n8864 : n8659;
  assign n8878 = pi09 ? n8873 : n8864;
  assign n8879 = pi08 ? n8877 : n8878;
  assign n8880 = pi10 ? n8694 : n8768;
  assign n8881 = pi10 ? n8833 : n8732;
  assign n8882 = pi09 ? n8880 : n8881;
  assign n8883 = pi10 ? n8732 : n8836;
  assign n8884 = pi12 ? n26 : ~n124;
  assign n8885 = pi11 ? n8735 : n8884;
  assign n8886 = pi12 ? n69 : ~n78;
  assign n8887 = pi14 ? n1355 : n37;
  assign n8888 = pi13 ? n30 : ~n8887;
  assign n8889 = pi12 ? n78 : n8888;
  assign n8890 = pi11 ? n8886 : n8889;
  assign n8891 = pi10 ? n8885 : n8890;
  assign n8892 = pi09 ? n8883 : n8891;
  assign n8893 = pi08 ? n8882 : n8892;
  assign n8894 = pi07 ? n8879 : n8893;
  assign n8895 = pi06 ? n8876 : n8894;
  assign n8896 = pi11 ? n26 : n8732;
  assign n8897 = pi10 ? n8896 : n8800;
  assign n8898 = pi09 ? n26 : n8897;
  assign n8899 = pi08 ? n26 : n8898;
  assign n8900 = pi13 ? n507 : ~n97;
  assign n8901 = pi12 ? n26 : n8900;
  assign n8902 = pi11 ? n8696 : n8901;
  assign n8903 = pi13 ? n507 : ~n68;
  assign n8904 = pi12 ? n26 : n8903;
  assign n8905 = pi12 ? n26 : ~n78;
  assign n8906 = pi11 ? n8904 : n8905;
  assign n8907 = pi10 ? n8902 : n8906;
  assign n8908 = pi09 ? n8907 : n26;
  assign n8909 = pi08 ? n8908 : n26;
  assign n8910 = pi07 ? n8899 : n8909;
  assign n8911 = pi06 ? n8910 : n26;
  assign n8912 = pi05 ? n8895 : n8911;
  assign n8913 = pi12 ? n26 : ~n69;
  assign n8914 = pi12 ? n124 : ~n78;
  assign n8915 = pi11 ? n8913 : n8914;
  assign n8916 = pi10 ? n8902 : n8915;
  assign n8917 = pi09 ? n8916 : n26;
  assign n8918 = pi08 ? n8917 : n26;
  assign n8919 = pi07 ? n8899 : n8918;
  assign n8920 = pi06 ? n8919 : n26;
  assign n8921 = pi11 ? n26 : n8696;
  assign n8922 = pi10 ? n8921 : n8836;
  assign n8923 = pi09 ? n26 : n8922;
  assign n8924 = pi08 ? n26 : n8923;
  assign n8925 = pi12 ? n124 : ~n69;
  assign n8926 = pi11 ? n8925 : n8886;
  assign n8927 = pi10 ? n8885 : n8926;
  assign n8928 = pi12 ? n78 : ~n58;
  assign n8929 = pi11 ? n8701 : n8928;
  assign n8930 = pi12 ? n78 : ~n306;
  assign n8931 = pi12 ? n78 : ~n122;
  assign n8932 = pi11 ? n8930 : n8931;
  assign n8933 = pi10 ? n8929 : n8932;
  assign n8934 = pi09 ? n8927 : n8933;
  assign n8935 = pi13 ? n26 : n72;
  assign n8936 = pi12 ? n78 : ~n8935;
  assign n8937 = pi08 ? n8934 : n8936;
  assign n8938 = pi07 ? n8924 : n8937;
  assign n8939 = pi13 ? n4125 : n72;
  assign n8940 = pi12 ? n78 : ~n8939;
  assign n8941 = pi11 ? n8936 : n8940;
  assign n8942 = pi10 ? n8936 : n8941;
  assign n8943 = pi09 ? n8936 : n8942;
  assign n8944 = pi08 ? n8936 : n8943;
  assign n8945 = pi07 ? n8936 : n8944;
  assign n8946 = pi06 ? n8938 : n8945;
  assign n8947 = pi05 ? n8920 : n8946;
  assign n8948 = pi04 ? n8912 : n8947;
  assign n8949 = pi03 ? n8848 : n8948;
  assign n8950 = pi13 ? n26 : n130;
  assign n8951 = pi12 ? n78 : ~n8950;
  assign n8952 = pi11 ? n8701 : n8951;
  assign n8953 = pi11 ? n8928 : n8930;
  assign n8954 = pi10 ? n8952 : n8953;
  assign n8955 = pi09 ? n8927 : n8954;
  assign n8956 = pi10 ? n8932 : n8931;
  assign n8957 = pi09 ? n8956 : n8931;
  assign n8958 = pi08 ? n8955 : n8957;
  assign n8959 = pi07 ? n8924 : n8958;
  assign n8960 = pi06 ? n8959 : n8931;
  assign n8961 = pi11 ? n26 : n8735;
  assign n8962 = pi12 ? n26 : ~n26;
  assign n8963 = pi11 ? n8735 : n8962;
  assign n8964 = pi10 ? n8961 : n8963;
  assign n8965 = pi09 ? n26 : n8964;
  assign n8966 = pi08 ? n26 : n8965;
  assign n8967 = pi11 ? n8962 : n8838;
  assign n8968 = pi10 ? n8967 : n8926;
  assign n8969 = pi11 ? n8739 : n8951;
  assign n8970 = pi13 ? n26 : n169;
  assign n8971 = pi12 ? n78 : ~n8970;
  assign n8972 = pi11 ? n8971 : n8928;
  assign n8973 = pi10 ? n8969 : n8972;
  assign n8974 = pi09 ? n8968 : n8973;
  assign n8975 = pi10 ? n8953 : n8930;
  assign n8976 = pi09 ? n8975 : n8930;
  assign n8977 = pi08 ? n8974 : n8976;
  assign n8978 = pi07 ? n8966 : n8977;
  assign n8979 = pi06 ? n8978 : n8930;
  assign n8980 = pi05 ? n8960 : n8979;
  assign n8981 = pi14 ? n168 : n29;
  assign n8982 = pi13 ? n8981 : ~n4125;
  assign n8983 = pi12 ? n26 : n8982;
  assign n8984 = pi11 ? n26 : n8983;
  assign n8985 = pi10 ? n8984 : n8735;
  assign n8986 = pi09 ? n26 : n8985;
  assign n8987 = pi08 ? n26 : n8986;
  assign n8988 = pi11 ? n8962 : n8884;
  assign n8989 = pi10 ? n8988 : n8926;
  assign n8990 = pi11 ? n8739 : n8701;
  assign n8991 = pi10 ? n8990 : n8971;
  assign n8992 = pi09 ? n8989 : n8991;
  assign n8993 = pi10 ? n8972 : n8928;
  assign n8994 = pi09 ? n8993 : n8928;
  assign n8995 = pi08 ? n8992 : n8994;
  assign n8996 = pi07 ? n8987 : n8995;
  assign n8997 = pi06 ? n8996 : n8928;
  assign n8998 = pi11 ? n26 : n8971;
  assign n8999 = pi10 ? n26 : n8998;
  assign n9000 = pi09 ? n8999 : n8971;
  assign n9001 = pi08 ? n26 : n9000;
  assign n9002 = pi07 ? n26 : n9001;
  assign n9003 = pi06 ? n26 : n9002;
  assign n9004 = pi05 ? n8997 : n9003;
  assign n9005 = pi04 ? n8980 : n9004;
  assign n9006 = pi12 ? n69 : ~n8700;
  assign n9007 = pi11 ? n26 : n9006;
  assign n9008 = pi10 ? n26 : n9007;
  assign n9009 = pi10 ? n8951 : n8971;
  assign n9010 = pi09 ? n9008 : n9009;
  assign n9011 = pi08 ? n26 : n9010;
  assign n9012 = pi07 ? n26 : n9011;
  assign n9013 = pi06 ? n26 : n9012;
  assign n9014 = pi13 ? n57 : n30;
  assign n9015 = pi12 ? n26 : n9014;
  assign n9016 = pi11 ? n26 : n9015;
  assign n9017 = pi10 ? n9016 : n8639;
  assign n9018 = pi09 ? n26 : n9017;
  assign n9019 = pi08 ? n26 : n9018;
  assign n9020 = pi07 ? n9019 : n8639;
  assign n9021 = pi11 ? n8639 : n8822;
  assign n9022 = pi10 ? n8639 : n9021;
  assign n9023 = pi09 ? n8639 : n9022;
  assign n9024 = pi13 ? n72 : ~n77;
  assign n9025 = pi12 ? n26 : n9024;
  assign n9026 = pi11 ? n8868 : n9025;
  assign n9027 = pi13 ? n507 : ~n143;
  assign n9028 = pi12 ? n26 : n9027;
  assign n9029 = pi12 ? n124 : ~n8738;
  assign n9030 = pi11 ? n9028 : n9029;
  assign n9031 = pi10 ? n9026 : n9030;
  assign n9032 = pi11 ? n9006 : n8701;
  assign n9033 = pi10 ? n9032 : n8951;
  assign n9034 = pi09 ? n9031 : n9033;
  assign n9035 = pi08 ? n9023 : n9034;
  assign n9036 = pi07 ? n8639 : n9035;
  assign n9037 = pi06 ? n9020 : n9036;
  assign n9038 = pi05 ? n9013 : n9037;
  assign n9039 = pi07 ? n8713 : n8658;
  assign n9040 = pi10 ? n8658 : n8866;
  assign n9041 = pi09 ? n8658 : n9040;
  assign n9042 = pi13 ? n72 : ~n68;
  assign n9043 = pi12 ? n26 : n9042;
  assign n9044 = pi11 ? n9043 : n8816;
  assign n9045 = pi13 ? n126 : ~n143;
  assign n9046 = pi12 ? n26 : n9045;
  assign n9047 = pi12 ? n26 : ~n8738;
  assign n9048 = pi11 ? n9046 : n9047;
  assign n9049 = pi10 ? n9044 : n9048;
  assign n9050 = pi09 ? n9049 : n9033;
  assign n9051 = pi08 ? n9041 : n9050;
  assign n9052 = pi07 ? n8658 : n9051;
  assign n9053 = pi06 ? n9039 : n9052;
  assign n9054 = pi07 ? n8747 : n8659;
  assign n9055 = pi13 ? n72 : ~n97;
  assign n9056 = pi12 ? n26 : n9055;
  assign n9057 = pi11 ? n8662 : n9056;
  assign n9058 = pi10 ? n8659 : n9057;
  assign n9059 = pi09 ? n8659 : n9058;
  assign n9060 = pi13 ? n38 : ~n68;
  assign n9061 = pi12 ? n26 : n9060;
  assign n9062 = pi13 ? n30 : ~n68;
  assign n9063 = pi12 ? n26 : n9062;
  assign n9064 = pi11 ? n9061 : n9063;
  assign n9065 = pi11 ? n8858 : n8905;
  assign n9066 = pi10 ? n9064 : n9065;
  assign n9067 = pi12 ? n69 : ~n8738;
  assign n9068 = pi11 ? n9029 : n9067;
  assign n9069 = pi10 ? n9068 : n8701;
  assign n9070 = pi09 ? n9066 : n9069;
  assign n9071 = pi08 ? n9059 : n9070;
  assign n9072 = pi07 ? n8659 : n9071;
  assign n9073 = pi06 ? n9054 : n9072;
  assign n9074 = pi05 ? n9053 : n9073;
  assign n9075 = pi04 ? n9038 : n9074;
  assign n9076 = pi03 ? n9005 : n9075;
  assign n9077 = pi02 ? n8949 : n9076;
  assign n9078 = pi01 ? n8711 : n9077;
  assign n9079 = pi14 ? n71 : n29;
  assign n9080 = pi13 ? n9079 : ~n4125;
  assign n9081 = pi12 ? n26 : n9080;
  assign n9082 = pi11 ? n26 : n9081;
  assign n9083 = pi10 ? n9082 : n8662;
  assign n9084 = pi09 ? n26 : n9083;
  assign n9085 = pi08 ? n26 : n9084;
  assign n9086 = pi07 ? n9085 : n8662;
  assign n9087 = pi13 ? n38 : ~n97;
  assign n9088 = pi12 ? n26 : n9087;
  assign n9089 = pi11 ? n8767 : n9088;
  assign n9090 = pi10 ? n8662 : n9089;
  assign n9091 = pi09 ? n8662 : n9090;
  assign n9092 = pi13 ? n126 : ~n77;
  assign n9093 = pi12 ? n26 : n9092;
  assign n9094 = pi11 ? n9061 : n9093;
  assign n9095 = pi11 ? n8858 : n9047;
  assign n9096 = pi10 ? n9094 : n9095;
  assign n9097 = pi14 ? n1355 : n29;
  assign n9098 = pi13 ? n30 : ~n9097;
  assign n9099 = pi12 ? n78 : n9098;
  assign n9100 = pi11 ? n8701 : n9099;
  assign n9101 = pi10 ? n9068 : n9100;
  assign n9102 = pi09 ? n9096 : n9101;
  assign n9103 = pi08 ? n9091 : n9102;
  assign n9104 = pi07 ? n8662 : n9103;
  assign n9105 = pi06 ? n9086 : n9104;
  assign n9106 = pi07 ? n26 : n8812;
  assign n9107 = pi11 ? n8767 : n26;
  assign n9108 = pi10 ? n9107 : n26;
  assign n9109 = pi09 ? n9108 : n26;
  assign n9110 = pi08 ? n9109 : n26;
  assign n9111 = pi07 ? n9110 : n26;
  assign n9112 = pi06 ? n9106 : n9111;
  assign n9113 = pi05 ? n9105 : n9112;
  assign n9114 = pi07 ? n26 : n8851;
  assign n9115 = pi11 ? n8814 : n26;
  assign n9116 = pi10 ? n9115 : n26;
  assign n9117 = pi09 ? n9116 : n26;
  assign n9118 = pi08 ? n9117 : n26;
  assign n9119 = pi07 ? n9118 : n26;
  assign n9120 = pi06 ? n9114 : n9119;
  assign n9121 = pi10 ? n8833 : n8854;
  assign n9122 = pi09 ? n8661 : n9121;
  assign n9123 = pi08 ? n8639 : n9122;
  assign n9124 = pi07 ? n9019 : n9123;
  assign n9125 = pi11 ? n8856 : n9028;
  assign n9126 = pi13 ? n507 : ~n57;
  assign n9127 = pi12 ? n26 : n9126;
  assign n9128 = pi12 ? n26 : ~n306;
  assign n9129 = pi11 ? n9127 : n9128;
  assign n9130 = pi10 ? n9125 : n9129;
  assign n9131 = pi12 ? n124 : ~n122;
  assign n9132 = pi12 ? n69 : ~n8935;
  assign n9133 = pi11 ? n9131 : n9132;
  assign n9134 = pi10 ? n9133 : n8936;
  assign n9135 = pi09 ? n9130 : n9134;
  assign n9136 = pi08 ? n9135 : n8936;
  assign n9137 = pi07 ? n9136 : n8944;
  assign n9138 = pi06 ? n9124 : n9137;
  assign n9139 = pi05 ? n9120 : n9138;
  assign n9140 = pi04 ? n9113 : n9139;
  assign n9141 = pi11 ? n8659 : n8767;
  assign n9142 = pi10 ? n8660 : n9141;
  assign n9143 = pi09 ? n9142 : n9121;
  assign n9144 = pi08 ? n8658 : n9143;
  assign n9145 = pi07 ? n8713 : n9144;
  assign n9146 = pi13 ? n507 : ~n176;
  assign n9147 = pi12 ? n26 : n9146;
  assign n9148 = pi11 ? n9093 : n9147;
  assign n9149 = pi13 ? n507 : ~n130;
  assign n9150 = pi12 ? n26 : n9149;
  assign n9151 = pi12 ? n26 : ~n58;
  assign n9152 = pi11 ? n9150 : n9151;
  assign n9153 = pi10 ? n9148 : n9152;
  assign n9154 = pi12 ? n124 : ~n306;
  assign n9155 = pi12 ? n69 : ~n306;
  assign n9156 = pi11 ? n9154 : n9155;
  assign n9157 = pi10 ? n9156 : n8931;
  assign n9158 = pi09 ? n9153 : n9157;
  assign n9159 = pi08 ? n9158 : n8931;
  assign n9160 = pi07 ? n9159 : n8931;
  assign n9161 = pi06 ? n9145 : n9160;
  assign n9162 = pi10 ? n8694 : n8767;
  assign n9163 = pi11 ? n8853 : n8904;
  assign n9164 = pi10 ? n8800 : n9163;
  assign n9165 = pi09 ? n9162 : n9164;
  assign n9166 = pi08 ? n8659 : n9165;
  assign n9167 = pi07 ? n8747 : n9166;
  assign n9168 = pi12 ? n26 : ~n8950;
  assign n9169 = pi12 ? n124 : ~n8970;
  assign n9170 = pi11 ? n9168 : n9169;
  assign n9171 = pi10 ? n9095 : n9170;
  assign n9172 = pi12 ? n124 : ~n58;
  assign n9173 = pi12 ? n69 : ~n58;
  assign n9174 = pi11 ? n9172 : n9173;
  assign n9175 = pi10 ? n9174 : n8930;
  assign n9176 = pi09 ? n9171 : n9175;
  assign n9177 = pi08 ? n9176 : n8930;
  assign n9178 = pi07 ? n9177 : n8930;
  assign n9179 = pi06 ? n9167 : n9178;
  assign n9180 = pi05 ? n9161 : n9179;
  assign n9181 = pi10 ? n8768 : n8833;
  assign n9182 = pi09 ? n9181 : n9164;
  assign n9183 = pi08 ? n8662 : n9182;
  assign n9184 = pi07 ? n9085 : n9183;
  assign n9185 = pi11 ? n8858 : n9028;
  assign n9186 = pi12 ? n26 : ~n8700;
  assign n9187 = pi12 ? n26 : ~n8970;
  assign n9188 = pi11 ? n9186 : n9187;
  assign n9189 = pi10 ? n9185 : n9188;
  assign n9190 = pi12 ? n69 : ~n8970;
  assign n9191 = pi11 ? n9169 : n9190;
  assign n9192 = pi10 ? n9191 : n8928;
  assign n9193 = pi09 ? n9189 : n9192;
  assign n9194 = pi08 ? n9193 : n8928;
  assign n9195 = pi07 ? n9194 : n8928;
  assign n9196 = pi06 ? n9184 : n9195;
  assign n9197 = pi05 ? n9196 : n9003;
  assign n9198 = pi04 ? n9180 : n9197;
  assign n9199 = pi03 ? n9140 : n9198;
  assign n9200 = pi07 ? n8777 : n8662;
  assign n9201 = pi06 ? n9200 : n9104;
  assign n9202 = pi10 ? n8767 : n26;
  assign n9203 = pi09 ? n9202 : n26;
  assign n9204 = pi08 ? n9203 : n26;
  assign n9205 = pi07 ? n8812 : n9204;
  assign n9206 = pi06 ? n9205 : n26;
  assign n9207 = pi05 ? n9201 : n9206;
  assign n9208 = pi10 ? n8854 : n26;
  assign n9209 = pi09 ? n9208 : n26;
  assign n9210 = pi08 ? n9209 : n26;
  assign n9211 = pi07 ? n8851 : n9210;
  assign n9212 = pi06 ? n9211 : n26;
  assign n9213 = pi11 ? n9028 : n9151;
  assign n9214 = pi10 ? n9163 : n9213;
  assign n9215 = pi12 ? n69 : ~n122;
  assign n9216 = pi11 ? n9154 : n9215;
  assign n9217 = pi10 ? n9216 : n8936;
  assign n9218 = pi09 ? n9214 : n9217;
  assign n9219 = pi08 ? n9218 : n8936;
  assign n9220 = pi07 ? n8899 : n9219;
  assign n9221 = pi06 ? n9220 : n8945;
  assign n9222 = pi05 ? n9212 : n9221;
  assign n9223 = pi04 ? n9207 : n9222;
  assign n9224 = pi03 ? n9075 : n9223;
  assign n9225 = pi02 ? n9199 : n9224;
  assign n9226 = pi11 ? n8853 : n8858;
  assign n9227 = pi11 ? n9147 : n9168;
  assign n9228 = pi10 ? n9226 : n9227;
  assign n9229 = pi11 ? n9172 : n9155;
  assign n9230 = pi10 ? n9229 : n8932;
  assign n9231 = pi09 ? n9228 : n9230;
  assign n9232 = pi08 ? n9231 : n8931;
  assign n9233 = pi07 ? n8899 : n9232;
  assign n9234 = pi06 ? n9233 : n8931;
  assign n9235 = pi10 ? n8921 : n8902;
  assign n9236 = pi09 ? n26 : n9235;
  assign n9237 = pi08 ? n26 : n9236;
  assign n9238 = pi12 ? n124 : ~n8950;
  assign n9239 = pi11 ? n9047 : n9238;
  assign n9240 = pi10 ? n8906 : n9239;
  assign n9241 = pi11 ? n9169 : n9173;
  assign n9242 = pi10 ? n9241 : n8953;
  assign n9243 = pi09 ? n9240 : n9242;
  assign n9244 = pi08 ? n9243 : n8930;
  assign n9245 = pi07 ? n9237 : n9244;
  assign n9246 = pi06 ? n9245 : n8930;
  assign n9247 = pi05 ? n9234 : n9246;
  assign n9248 = pi14 ? n125 : n29;
  assign n9249 = pi13 ? n9248 : ~n4125;
  assign n9250 = pi12 ? n26 : n9249;
  assign n9251 = pi11 ? n26 : n9250;
  assign n9252 = pi10 ? n9251 : n8902;
  assign n9253 = pi09 ? n26 : n9252;
  assign n9254 = pi08 ? n26 : n9253;
  assign n9255 = pi11 ? n8904 : n8858;
  assign n9256 = pi11 ? n9047 : n9186;
  assign n9257 = pi10 ? n9255 : n9256;
  assign n9258 = pi10 ? n9191 : n8972;
  assign n9259 = pi09 ? n9257 : n9258;
  assign n9260 = pi08 ? n9259 : n8928;
  assign n9261 = pi07 ? n9254 : n9260;
  assign n9262 = pi14 ? n1355 : ~n26;
  assign n9263 = pi13 ? n30 : ~n9262;
  assign n9264 = pi12 ? n78 : n9263;
  assign n9265 = pi11 ? n8928 : n9264;
  assign n9266 = pi10 ? n8928 : n9265;
  assign n9267 = pi09 ? n8928 : n9266;
  assign n9268 = pi08 ? n8928 : n9267;
  assign n9269 = pi07 ? n8928 : n9268;
  assign n9270 = pi06 ? n9261 : n9269;
  assign n9271 = pi10 ? n26 : n8971;
  assign n9272 = pi10 ? n8971 : n26;
  assign n9273 = pi09 ? n9271 : n9272;
  assign n9274 = pi08 ? n9273 : n26;
  assign n9275 = pi07 ? n9274 : n26;
  assign n9276 = pi06 ? n26 : n9275;
  assign n9277 = pi05 ? n9270 : n9276;
  assign n9278 = pi04 ? n9247 : n9277;
  assign n9279 = pi12 ? n69 : ~n8950;
  assign n9280 = pi11 ? n9279 : n8951;
  assign n9281 = pi10 ? n26 : n9280;
  assign n9282 = pi09 ? n9281 : n9272;
  assign n9283 = pi08 ? n9282 : n26;
  assign n9284 = pi07 ? n9283 : n26;
  assign n9285 = pi06 ? n26 : n9284;
  assign n9286 = pi11 ? n8639 : n8787;
  assign n9287 = pi13 ? n79 : ~n77;
  assign n9288 = pi12 ? n26 : n9287;
  assign n9289 = pi11 ? n8781 : n9288;
  assign n9290 = pi10 ? n9286 : n9289;
  assign n9291 = pi09 ? n8639 : n9290;
  assign n9292 = pi08 ? n8639 : n9291;
  assign n9293 = pi07 ? n9019 : n9292;
  assign n9294 = pi13 ? n72 : ~n143;
  assign n9295 = pi12 ? n26 : n9294;
  assign n9296 = pi11 ? n9295 : n9028;
  assign n9297 = pi12 ? n124 : ~n8700;
  assign n9298 = pi11 ? n9297 : n9006;
  assign n9299 = pi10 ? n9296 : n9298;
  assign n9300 = pi11 ? n8971 : n8930;
  assign n9301 = pi10 ? n8951 : n9300;
  assign n9302 = pi09 ? n9299 : n9301;
  assign n9303 = pi11 ? n8931 : n8936;
  assign n9304 = pi10 ? n9303 : n8936;
  assign n9305 = pi09 ? n9304 : n8936;
  assign n9306 = pi08 ? n9302 : n9305;
  assign n9307 = pi07 ? n9306 : n8944;
  assign n9308 = pi06 ? n9293 : n9307;
  assign n9309 = pi05 ? n9285 : n9308;
  assign n9310 = pi11 ? n8658 : n8779;
  assign n9311 = pi10 ? n9310 : n9026;
  assign n9312 = pi09 ? n8658 : n9311;
  assign n9313 = pi08 ? n8658 : n9312;
  assign n9314 = pi07 ? n8713 : n9313;
  assign n9315 = pi13 ? n30 : ~n143;
  assign n9316 = pi12 ? n26 : n9315;
  assign n9317 = pi11 ? n9316 : n9046;
  assign n9318 = pi11 ? n9186 : n9006;
  assign n9319 = pi10 ? n9317 : n9318;
  assign n9320 = pi09 ? n9319 : n9009;
  assign n9321 = pi10 ? n8930 : n8931;
  assign n9322 = pi09 ? n9321 : n8931;
  assign n9323 = pi08 ? n9320 : n9322;
  assign n9324 = pi07 ? n9323 : n8931;
  assign n9325 = pi06 ? n9314 : n9324;
  assign n9326 = pi11 ? n8659 : n9056;
  assign n9327 = pi11 ? n9043 : n9061;
  assign n9328 = pi10 ? n9326 : n9327;
  assign n9329 = pi09 ? n8659 : n9328;
  assign n9330 = pi08 ? n8659 : n9329;
  assign n9331 = pi07 ? n8747 : n9330;
  assign n9332 = pi11 ? n8816 : n8858;
  assign n9333 = pi11 ? n9047 : n9029;
  assign n9334 = pi10 ? n9332 : n9333;
  assign n9335 = pi11 ? n8951 : n8971;
  assign n9336 = pi10 ? n9032 : n9335;
  assign n9337 = pi09 ? n9334 : n9336;
  assign n9338 = pi10 ? n8972 : n8930;
  assign n9339 = pi09 ? n9338 : n8930;
  assign n9340 = pi08 ? n9337 : n9339;
  assign n9341 = pi07 ? n9340 : n8930;
  assign n9342 = pi06 ? n9331 : n9341;
  assign n9343 = pi05 ? n9325 : n9342;
  assign n9344 = pi04 ? n9309 : n9343;
  assign n9345 = pi03 ? n9278 : n9344;
  assign n9346 = pi11 ? n8662 : n9088;
  assign n9347 = pi13 ? n38 : ~n77;
  assign n9348 = pi12 ? n26 : n9347;
  assign n9349 = pi11 ? n9061 : n9348;
  assign n9350 = pi10 ? n9346 : n9349;
  assign n9351 = pi09 ? n8662 : n9350;
  assign n9352 = pi08 ? n8662 : n9351;
  assign n9353 = pi07 ? n8777 : n9352;
  assign n9354 = pi11 ? n9093 : n9028;
  assign n9355 = pi10 ? n9354 : n9333;
  assign n9356 = pi09 ? n9355 : n9033;
  assign n9357 = pi10 ? n8971 : n8928;
  assign n9358 = pi09 ? n9357 : n8928;
  assign n9359 = pi08 ? n9356 : n9358;
  assign n9360 = pi07 ? n9359 : n9268;
  assign n9361 = pi06 ? n9353 : n9360;
  assign n9362 = pi05 ? n9361 : n9206;
  assign n9363 = pi11 ? n9155 : n8931;
  assign n9364 = pi10 ? n9363 : n8936;
  assign n9365 = pi09 ? n9214 : n9364;
  assign n9366 = pi08 ? n9365 : n8936;
  assign n9367 = pi07 ? n8899 : n9366;
  assign n9368 = pi06 ? n9367 : n8945;
  assign n9369 = pi05 ? n9212 : n9368;
  assign n9370 = pi04 ? n9362 : n9369;
  assign n9371 = pi11 ? n9186 : n9238;
  assign n9372 = pi10 ? n9226 : n9371;
  assign n9373 = pi10 ? n8953 : n8932;
  assign n9374 = pi09 ? n9372 : n9373;
  assign n9375 = pi08 ? n9374 : n8931;
  assign n9376 = pi07 ? n8899 : n9375;
  assign n9377 = pi06 ? n9376 : n8931;
  assign n9378 = pi11 ? n9029 : n9279;
  assign n9379 = pi10 ? n8906 : n9378;
  assign n9380 = pi10 ? n8972 : n8953;
  assign n9381 = pi09 ? n9379 : n9380;
  assign n9382 = pi08 ? n9381 : n8930;
  assign n9383 = pi07 ? n9237 : n9382;
  assign n9384 = pi06 ? n9383 : n8930;
  assign n9385 = pi05 ? n9377 : n9384;
  assign n9386 = pi11 ? n9029 : n9006;
  assign n9387 = pi10 ? n8906 : n9386;
  assign n9388 = pi10 ? n8971 : n8972;
  assign n9389 = pi09 ? n9387 : n9388;
  assign n9390 = pi08 ? n9389 : n8928;
  assign n9391 = pi07 ? n9237 : n9390;
  assign n9392 = pi06 ? n9391 : n8928;
  assign n9393 = pi11 ? n8735 : n8901;
  assign n9394 = pi10 ? n8984 : n9393;
  assign n9395 = pi09 ? n26 : n9394;
  assign n9396 = pi08 ? n26 : n9395;
  assign n9397 = pi11 ? n8913 : n8905;
  assign n9398 = pi10 ? n9397 : n9386;
  assign n9399 = pi10 ? n9335 : n8971;
  assign n9400 = pi09 ? n9398 : n9399;
  assign n9401 = pi08 ? n9400 : n8971;
  assign n9402 = pi07 ? n9396 : n9401;
  assign n9403 = pi14 ? n1355 : n168;
  assign n9404 = pi13 ? n30 : ~n9403;
  assign n9405 = pi12 ? n78 : n9404;
  assign n9406 = pi11 ? n8971 : n9405;
  assign n9407 = pi10 ? n8971 : n9406;
  assign n9408 = pi09 ? n8971 : n9407;
  assign n9409 = pi08 ? n8971 : n9408;
  assign n9410 = pi07 ? n8971 : n9409;
  assign n9411 = pi06 ? n9402 : n9410;
  assign n9412 = pi05 ? n9392 : n9411;
  assign n9413 = pi04 ? n9385 : n9412;
  assign n9414 = pi03 ? n9370 : n9413;
  assign n9415 = pi02 ? n9345 : n9414;
  assign n9416 = pi01 ? n9225 : n9415;
  assign n9417 = pi00 ? n9078 : n9416;
  assign po0 = ~n1247;
  assign po1 = ~n2306;
  assign po2 = ~n3763;
  assign po3 = ~n5527;
  assign po4 = ~n7341;
  assign po5 = ~n8588;
  assign po6 = ~n9417;
endmodule


