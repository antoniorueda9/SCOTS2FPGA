// Benchmark "DD" written by ABC on Wed Jun  5 14:52:31 2019

module DD ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24,
    po0, po1, po2, po3, po4, po5  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24;
  output po0, po1, po2, po3, po4, po5;
  wire n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
    n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
    n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
    n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
    n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
    n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
    n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
    n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
    n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
    n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
    n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
    n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
    n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
    n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
    n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
    n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
    n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
    n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
    n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
    n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
    n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
    n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
    n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
    n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
    n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
    n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
    n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
    n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
    n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
    n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
    n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
    n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
    n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
    n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
    n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
    n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
    n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
    n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
    n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
    n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
    n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
    n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
    n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
    n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
    n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
    n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
    n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
    n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
    n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
    n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
    n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
    n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
    n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
    n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
    n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
    n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
    n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
    n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
    n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
    n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
    n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
    n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
    n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
    n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
    n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
    n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
    n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
    n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
    n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
    n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
    n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
    n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
    n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
    n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
    n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
    n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
    n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
    n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
    n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
    n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
    n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
    n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
    n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
    n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
    n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
    n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
    n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
    n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
    n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
    n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
    n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
    n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
    n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
    n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
    n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
    n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
    n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
    n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
    n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
    n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
    n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
    n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
    n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
    n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
    n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
    n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
    n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
    n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
    n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
    n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
    n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
    n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
    n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
    n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
    n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
    n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
    n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
    n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
    n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
    n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
    n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
    n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
    n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
    n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
    n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
    n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
    n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
    n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
    n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
    n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
    n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
    n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
    n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
    n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
    n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
    n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
    n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
    n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
    n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
    n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
    n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
    n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
    n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
    n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
    n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
    n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
    n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
    n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
    n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
    n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
    n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
    n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
    n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
    n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
    n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
    n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
    n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
    n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
    n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
    n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
    n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
    n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
    n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
    n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
    n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
    n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
    n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
    n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
    n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
    n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
    n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
    n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
    n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
    n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
    n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
    n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
    n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
    n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
    n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
    n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
    n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
    n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
    n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
    n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
    n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
    n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
    n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
    n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
    n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
    n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
    n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
    n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
    n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
    n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
    n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
    n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
    n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
    n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
    n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
    n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
    n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
    n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
    n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
    n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
    n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
    n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
    n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
    n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
    n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
    n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
    n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
    n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
    n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
    n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
    n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
    n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
    n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
    n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
    n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
    n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
    n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
    n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
    n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
    n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
    n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
    n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
    n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
    n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
    n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
    n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
    n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
    n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
    n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
    n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
    n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
    n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
    n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
    n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
    n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
    n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
    n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
    n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
    n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
    n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
    n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
    n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
    n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
    n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
    n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
    n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
    n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
    n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
    n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
    n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
    n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
    n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
    n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
    n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
    n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
    n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
    n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
    n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
    n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
    n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
    n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
    n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
    n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
    n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
    n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
    n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
    n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
    n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
    n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
    n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
    n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
    n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
    n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
    n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
    n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
    n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
    n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
    n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
    n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
    n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
    n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
    n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
    n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
    n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
    n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
    n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
    n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
    n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
    n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
    n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
    n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
    n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
    n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
    n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
    n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
    n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
    n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
    n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
    n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
    n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
    n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
    n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
    n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
    n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
    n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
    n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
    n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
    n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
    n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
    n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
    n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
    n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
    n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
    n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
    n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
    n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
    n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
    n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
    n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
    n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
    n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
    n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
    n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
    n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
    n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
    n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
    n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
    n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
    n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
    n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
    n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
    n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
    n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
    n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
    n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
    n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
    n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
    n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
    n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
    n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
    n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
    n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
    n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
    n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
    n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
    n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
    n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
    n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
    n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
    n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
    n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
    n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
    n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
    n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
    n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
    n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
    n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
    n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
    n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
    n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
    n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
    n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
    n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
    n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
    n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
    n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
    n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
    n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
    n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
    n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
    n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
    n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
    n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
    n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
    n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
    n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
    n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
    n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
    n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
    n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
    n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
    n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
    n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
    n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
    n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
    n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
    n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
    n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
    n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
    n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
    n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
    n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
    n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
    n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
    n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
    n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
    n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
    n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
    n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
    n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
    n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
    n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
    n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
    n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
    n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
    n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
    n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
    n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
    n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
    n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
    n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
    n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
    n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
    n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
    n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
    n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
    n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
    n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
    n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
    n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
    n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
    n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
    n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
    n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
    n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
    n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
    n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
    n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
    n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
    n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
    n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
    n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
    n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
    n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
    n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
    n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
    n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
    n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
    n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
    n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
    n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
    n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
    n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
    n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
    n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
    n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
    n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
    n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
    n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
    n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
    n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
    n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
    n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
    n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
    n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
    n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
    n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
    n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
    n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
    n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
    n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
    n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
    n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
    n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
    n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
    n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
    n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
    n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
    n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
    n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
    n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
    n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
    n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
    n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
    n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
    n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
    n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
    n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
    n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
    n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
    n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
    n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
    n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
    n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
    n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
    n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
    n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
    n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
    n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
    n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
    n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
    n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
    n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
    n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
    n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
    n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
    n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
    n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
    n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
    n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
    n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
    n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
    n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
    n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
    n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
    n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
    n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
    n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
    n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
    n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
    n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
    n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
    n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
    n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
    n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
    n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
    n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
    n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
    n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
    n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
    n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
    n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
    n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
    n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
    n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
    n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
    n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
    n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
    n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
    n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
    n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
    n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
    n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
    n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
    n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
    n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
    n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
    n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
    n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
    n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
    n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
    n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
    n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
    n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
    n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
    n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
    n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
    n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
    n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
    n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
    n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
    n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
    n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
    n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
    n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
    n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
    n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
    n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
    n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
    n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
    n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
    n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
    n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
    n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
    n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
    n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
    n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
    n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
    n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
    n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
    n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
    n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
    n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
    n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
    n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
    n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
    n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
    n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
    n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
    n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
    n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
    n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
    n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
    n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
    n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
    n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
    n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
    n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
    n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
    n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
    n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
    n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
    n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
    n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
    n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
    n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
    n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
    n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
    n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
    n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
    n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
    n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
    n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
    n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
    n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
    n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
    n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
    n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
    n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
    n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
    n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
    n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
    n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
    n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
    n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
    n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
    n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
    n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
    n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
    n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
    n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
    n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
    n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
    n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
    n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
    n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
    n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
    n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
    n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
    n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
    n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
    n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
    n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
    n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
    n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
    n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
    n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
    n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
    n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
    n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
    n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
    n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
    n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
    n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
    n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
    n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
    n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
    n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
    n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
    n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
    n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
    n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
    n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
    n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
    n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
    n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
    n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
    n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
    n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
    n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
    n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
    n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
    n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
    n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
    n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
    n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
    n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
    n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
    n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
    n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
    n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
    n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
    n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
    n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
    n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
    n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
    n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
    n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
    n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
    n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
    n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
    n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
    n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
    n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
    n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
    n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
    n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
    n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
    n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
    n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
    n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
    n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
    n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
    n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429,
    n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
    n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
    n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
    n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
    n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
    n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
    n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
    n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
    n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
    n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
    n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
    n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
    n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
    n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
    n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
    n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
    n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
    n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
    n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
    n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726,
    n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
    n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
    n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
    n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798,
    n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
    n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
    n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852,
    n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870,
    n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
    n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
    n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
    n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942,
    n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
    n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
    n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
    n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
    n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
    n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014,
    n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
    n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
    n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
    n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
    n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
    n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
    n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
    n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086,
    n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
    n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
    n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
    n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
    n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
    n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
    n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
    n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
    n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
    n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
    n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212,
    n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230,
    n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
    n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
    n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
    n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
    n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
    n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
    n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
    n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
    n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
    n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
    n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
    n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
    n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
    n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
    n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
    n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
    n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
    n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
    n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
    n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
    n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
    n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
    n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
    n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
    n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
    n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
    n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
    n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
    n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716,
    n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
    n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
    n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
    n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
    n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
    n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
    n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
    n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788,
    n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
    n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
    n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
    n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
    n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
    n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
    n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
    n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
    n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
    n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
    n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
    n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
    n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
    n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
    n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932,
    n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950,
    n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
    n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
    n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
    n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
    n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
    n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
    n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
    n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
    n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
    n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
    n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
    n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
    n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
    n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
    n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
    n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
    n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
    n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
    n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
    n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
    n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
    n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
    n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
    n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238,
    n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
    n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
    n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292,
    n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310,
    n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
    n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
    n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
    n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
    n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
    n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364,
    n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
    n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382,
    n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
    n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
    n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
    n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
    n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
    n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
    n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
    n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454,
    n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
    n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
    n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
    n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
    n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
    n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
    n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
    n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
    n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
    n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
    n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
    n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
    n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
    n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
    n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598,
    n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
    n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
    n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
    n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
    n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
    n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
    n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
    n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
    n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
    n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
    n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
    n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
    n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
    n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
    n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
    n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
    n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
    n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
    n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
    n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
    n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
    n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
    n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
    n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
    n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
    n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
    n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
    n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
    n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
    n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
    n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
    n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
    n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
    n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
    n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102,
    n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
    n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
    n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
    n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
    n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
    n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
    n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
    n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
    n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
    n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
    n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
    n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
    n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
    n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
    n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
    n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
    n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
    n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
    n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
    n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
    n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
    n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
    n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
    n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
    n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
    n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
    n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
    n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
    n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
    n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
    n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
    n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
    n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
    n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
    n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
    n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
    n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
    n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
    n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
    n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
    n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
    n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
    n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
    n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
    n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
    n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
    n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
    n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
    n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
    n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
    n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
    n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
    n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
    n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
    n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
    n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
    n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
    n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
    n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
    n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
    n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
    n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
    n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
    n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
    n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
    n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
    n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
    n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
    n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
    n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
    n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
    n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
    n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
    n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
    n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
    n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
    n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
    n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
    n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
    n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542,
    n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
    n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
    n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
    n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614,
    n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
    n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
    n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
    n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686,
    n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
    n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
    n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
    n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758,
    n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
    n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
    n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
    n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
    n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
    n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
    n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
    n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
    n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
    n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
    n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
    n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
    n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
    n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
    n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
    n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
    n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
    n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
    n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
    n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
    n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
    n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
    n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
    n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
    n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
    n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
    n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
    n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
    n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
    n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
    n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
    n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
    n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
    n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
    n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
    n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
    n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
    n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
    n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334,
    n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
    n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
    n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
    n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
    n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
    n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
    n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
    n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406,
    n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
    n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
    n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
    n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
    n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
    n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
    n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
    n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
    n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550,
    n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559,
    n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
    n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
    n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
    n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
    n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
    n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
    n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
    n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
    n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
    n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
    n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
    n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
    n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
    n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
    n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784,
    n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
    n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
    n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838,
    n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856,
    n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
    n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
    n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
    n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928,
    n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
    n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
    n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
    n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000,
    n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
    n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
    n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054,
    n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072,
    n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
    n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
    n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
    n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
    n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
    n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
    n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198,
    n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216,
    n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
    n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
    n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
    n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
    n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
    n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
    n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
    n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
    n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
    n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
    n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
    n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
    n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
    n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
    n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
    n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486,
    n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
    n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504,
    n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
    n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
    n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558,
    n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
    n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
    n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
    n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
    n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630,
    n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
    n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648,
    n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
    n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
    n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
    n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
    n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
    n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
    n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720,
    n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
    n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
    n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
    n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
    n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
    n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
    n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846,
    n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864,
    n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
    n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
    n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
    n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936,
    n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
    n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
    n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990,
    n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
    n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
    n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
    n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
    n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
    n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
    n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
    n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
    n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
    n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
    n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
    n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
    n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
    n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
    n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
    n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
    n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
    n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
    n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
    n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
    n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
    n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
    n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764,
    n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
    n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
    n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
    n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
    n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
    n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
    n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
    n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980,
    n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989,
    n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
    n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
    n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
    n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
    n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
    n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
    n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
    n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061,
    n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
    n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
    n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
    n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
    n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
    n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
    n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
    n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
    n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
    n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
    n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
    n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
    n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
    n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
    n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
    n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412,
    n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
    n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
    n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
    n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
    n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
    n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
    n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
    n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
    n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
    n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
    n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
    n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
    n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
    n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
    n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
    n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
    n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
    n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
    n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
    n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628,
    n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637,
    n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
    n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
    n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
    n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
    n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
    n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
    n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709,
    n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
    n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
    n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
    n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
    n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
    n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
    n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
    n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
    n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
    n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
    n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
    n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
    n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
    n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853,
    n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
    n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
    n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
    n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916,
    n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925,
    n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
    n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
    n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
    n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
    n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
    n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
    n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997,
    n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
    n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
    n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
    n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
    n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
    n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
    n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060,
    n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
    n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
    n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
    n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
    n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114,
    n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
    n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132,
    n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141,
    n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
    n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
    n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
    n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
    n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204,
    n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213,
    n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
    n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
    n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
    n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
    n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258,
    n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
    n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
    n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285,
    n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
    n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
    n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
    n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
    n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
    n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
    n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348,
    n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357,
    n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
    n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
    n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
    n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
    n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
    n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
    n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
    n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
    n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
    n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
    n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
    n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
    n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
    n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
    n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501,
    n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
    n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
    n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
    n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
    n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
    n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
    n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564,
    n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573,
    n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
    n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
    n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
    n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
    n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
    n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
    n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
    n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
    n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
    n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
    n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
    n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
    n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
    n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
    n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
    n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789,
    n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
    n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
    n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816,
    n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
    n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
    n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
    n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
    n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861,
    n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
    n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
    n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888,
    n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
    n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906,
    n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
    n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
    n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933,
    n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
    n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
    n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960,
    n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
    n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
    n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
    n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
    n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005,
    n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
    n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023,
    n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
    n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
    n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
    n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077,
    n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
    n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095,
    n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
    n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
    n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
    n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
    n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
    n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149,
    n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
    n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167,
    n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176,
    n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
    n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
    n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
    n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
    n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221,
    n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
    n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239,
    n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248,
    n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
    n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
    n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
    n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
    n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293,
    n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
    n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320,
    n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
    n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
    n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
    n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
    n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
    n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
    n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
    n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
    n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437,
    n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
    n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455,
    n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
    n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
    n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
    n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
    n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
    n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509,
    n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
    n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
    n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
    n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
    n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
    n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
    n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
    n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581,
    n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
    n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599,
    n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608,
    n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
    n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
    n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
    n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644,
    n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653,
    n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
    n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
    n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680,
    n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
    n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
    n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
    n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
    n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725,
    n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
    n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743,
    n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752,
    n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
    n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
    n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
    n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788,
    n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797,
    n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
    n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815,
    n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824,
    n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
    n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
    n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
    n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
    n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
    n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887,
    n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
    n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
    n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
    n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
    n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
    n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941,
    n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
    n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959,
    n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968,
    n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
    n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
    n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
    n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013,
    n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
    n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040,
    n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
    n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
    n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
    n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076,
    n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085,
    n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
    n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103,
    n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
    n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
    n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
    n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
    n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148,
    n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157,
    n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
    n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
    n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184,
    n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
    n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202,
    n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
    n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
    n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229,
    n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
    n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
    n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
    n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
    n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
    n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328,
    n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
    n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
    n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
    n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400,
    n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
    n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
    n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
    n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
    n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445,
    n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
    n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463,
    n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472,
    n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
    n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
    n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
    n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
    n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535,
    n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544,
    n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
    n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562,
    n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
    n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
    n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589,
    n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
    n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616,
    n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
    n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634,
    n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
    n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652,
    n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661,
    n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
    n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679,
    n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688,
    n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
    n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
    n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
    n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
    n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
    n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
    n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
    n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805,
    n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
    n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823,
    n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832,
    n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
    n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850,
    n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
    n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868,
    n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877,
    n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
    n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895,
    n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904,
    n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
    n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922,
    n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
    n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940,
    n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949,
    n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
    n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
    n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976,
    n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
    n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994,
    n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
    n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
    n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021,
    n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
    n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039,
    n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048,
    n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
    n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
    n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
    n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084,
    n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093,
    n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
    n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111,
    n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120,
    n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
    n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
    n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156,
    n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165,
    n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
    n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183,
    n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192,
    n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
    n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
    n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
    n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228,
    n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237,
    n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
    n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255,
    n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264,
    n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
    n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282,
    n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
    n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300,
    n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309,
    n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
    n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
    n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
    n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
    n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
    n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
    n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
    n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381,
    n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
    n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
    n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
    n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
    n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426,
    n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
    n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444,
    n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453,
    n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
    n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
    n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
    n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
    n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
    n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
    n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516,
    n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525,
    n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
    n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
    n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552,
    n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
    n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
    n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
    n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588,
    n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597,
    n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
    n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
    n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624,
    n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
    n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642,
    n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
    n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660,
    n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669,
    n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
    n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
    n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696,
    n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
    n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714,
    n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
    n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732,
    n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741,
    n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
    n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
    n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
    n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786,
    n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
    n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804,
    n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813,
    n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
    n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831,
    n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840,
    n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
    n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
    n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
    n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876,
    n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885,
    n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
    n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903,
    n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912,
    n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
    n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
    n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
    n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948,
    n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957,
    n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
    n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975,
    n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984,
    n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
    n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002,
    n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
    n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020,
    n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029,
    n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
    n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047,
    n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056,
    n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
    n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
    n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092,
    n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101,
    n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
    n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119,
    n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
    n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173,
    n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191,
    n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200,
    n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
    n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
    n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236,
    n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
    n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
    n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
    n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308,
    n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317,
    n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
    n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
    n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
    n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
    n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
    n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
    n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
    n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389,
    n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
    n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
    n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
    n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
    n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452,
    n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
    n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
    n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
    n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524,
    n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
    n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
    n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
    n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
    n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
    n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632,
    n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650,
    n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
    n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668,
    n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677,
    n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
    n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704,
    n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
    n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722,
    n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740,
    n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749,
    n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
    n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776,
    n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
    n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794,
    n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
    n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812,
    n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821,
    n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
    n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839,
    n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
    n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
    n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866,
    n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
    n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884,
    n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893,
    n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
    n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911,
    n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920,
    n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
    n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938,
    n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956,
    n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965,
    n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
    n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983,
    n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992,
    n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
    n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010,
    n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
    n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028,
    n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037,
    n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
    n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
    n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064,
    n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
    n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082,
    n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
    n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100,
    n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109,
    n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
    n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127,
    n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
    n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
    n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
    n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
    n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172,
    n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181,
    n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
    n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199,
    n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
    n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
    n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226,
    n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
    n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244,
    n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253,
    n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
    n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271,
    n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280,
    n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
    n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298,
    n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
    n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316,
    n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325,
    n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
    n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
    n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
    n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
    n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388,
    n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397,
    n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
    n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415,
    n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424,
    n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
    n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442,
    n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
    n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460,
    n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
    n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487,
    n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496,
    n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
    n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514,
    n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
    n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532,
    n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541,
    n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
    n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568,
    n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
    n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
    n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
    n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604,
    n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613,
    n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
    n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
    n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640,
    n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
    n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
    n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
    n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676,
    n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685,
    n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
    n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703,
    n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712,
    n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
    n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
    n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
    n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748,
    n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757,
    n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
    n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775,
    n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784,
    n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
    n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
    n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829,
    n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847,
    n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
    n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
    n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
    n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892,
    n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901,
    n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
    n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919,
    n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
    n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
    n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
    n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
    n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964,
    n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973,
    n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
    n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991,
    n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
    n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
    n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
    n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
    n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036,
    n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045,
    n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
    n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063,
    n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
    n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
    n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
    n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117,
    n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
    n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
    n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
    n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
    n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
    n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
    n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180,
    n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189,
    n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
    n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207,
    n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
    n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
    n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
    n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
    n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252,
    n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261,
    n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
    n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
    n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
    n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
    n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
    n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
    n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324,
    n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333,
    n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
    n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351,
    n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
    n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
    n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
    n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
    n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396,
    n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405,
    n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
    n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423,
    n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
    n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
    n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
    n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
    n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468,
    n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477,
    n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
    n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495,
    n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
    n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
    n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
    n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531,
    n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540,
    n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549,
    n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
    n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567,
    n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
    n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
    n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594,
    n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603,
    n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612,
    n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621,
    n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
    n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639,
    n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
    n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
    n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666,
    n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675,
    n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684,
    n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693,
    n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
    n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711,
    n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720,
    n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
    n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738,
    n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747,
    n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756,
    n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765,
    n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
    n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783,
    n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
    n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
    n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
    n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819,
    n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828,
    n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837,
    n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
    n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
    n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
    n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
    n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
    n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
    n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900,
    n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909,
    n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
    n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927,
    n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936,
    n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
    n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954,
    n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963,
    n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972,
    n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981,
    n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
    n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999,
    n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008,
    n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
    n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026,
    n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035,
    n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044,
    n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053,
    n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
    n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071,
    n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080,
    n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
    n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
    n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
    n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116,
    n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125,
    n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
    n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143,
    n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
    n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
    n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170,
    n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179,
    n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188,
    n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197,
    n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
    n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215,
    n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
    n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
    n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242,
    n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251,
    n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260,
    n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269,
    n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
    n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287,
    n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
    n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
    n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
    n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
    n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332,
    n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341,
    n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
    n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359,
    n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368,
    n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
    n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
    n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395,
    n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404,
    n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413,
    n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
    n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431,
    n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
    n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
    n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
    n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467,
    n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476,
    n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485,
    n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
    n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
    n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
    n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
    n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
    n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
    n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
    n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
    n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
    n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
    n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
    n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
    n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620,
    n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629,
    n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
    n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647,
    n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
    n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
    n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
    n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683,
    n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692,
    n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701,
    n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
    n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
    n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
    n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
    n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
    n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
    n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764,
    n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773,
    n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
    n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
    n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
    n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
    n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
    n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
    n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836,
    n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845,
    n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
    n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863,
    n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
    n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
    n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
    n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
    n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908,
    n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917,
    n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
    n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
    n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
    n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
    n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980,
    n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989,
    n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
    n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
    n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
    n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
    n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
    n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
    n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052,
    n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061,
    n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
    n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079,
    n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
    n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
    n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
    n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124,
    n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133,
    n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
    n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151,
    n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160,
    n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
    n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
    n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196,
    n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
    n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223,
    n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
    n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
    n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
    n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259,
    n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268,
    n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277,
    n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
    n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295,
    n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
    n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
    n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
    n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331,
    n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340,
    n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349,
    n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
    n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367,
    n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
    n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
    n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
    n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403,
    n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412,
    n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421,
    n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
    n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439,
    n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
    n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
    n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
    n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475,
    n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484,
    n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493,
    n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502,
    n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511,
    n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
    n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
    n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
    n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
    n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556,
    n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565,
    n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574,
    n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583,
    n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
    n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
    n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
    n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
    n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628,
    n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637,
    n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646,
    n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
    n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
    n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700,
    n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
    n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727,
    n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
    n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
    n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
    n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763,
    n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772,
    n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, n39781,
    n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
    n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799,
    n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
    n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
    n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
    n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
    n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844,
    n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852, n39853,
    n39854, n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
    n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871,
    n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
    n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
    n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
    n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
    n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916,
    n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924, n39925,
    n39926, n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
    n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943,
    n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
    n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
    n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
    n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979,
    n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988,
    n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996, n39997,
    n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006,
    n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015,
    n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
    n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
    n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
    n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051,
    n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060,
    n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068, n40069,
    n40070, n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078,
    n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087,
    n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
    n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
    n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
    n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123,
    n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132,
    n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141,
    n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
    n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159,
    n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
    n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
    n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
    n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
    n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204,
    n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212, n40213,
    n40214, n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222,
    n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
    n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
    n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
    n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
    n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276,
    n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284, n40285,
    n40286, n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294,
    n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303,
    n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
    n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
    n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
    n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339,
    n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348,
    n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356, n40357,
    n40358, n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
    n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375,
    n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
    n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
    n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
    n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411,
    n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420,
    n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428, n40429,
    n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438,
    n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447,
    n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
    n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
    n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
    n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
    n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492,
    n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501,
    n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
    n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
    n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
    n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
    n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
    n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
    n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564,
    n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573,
    n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582,
    n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591,
    n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
    n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
    n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
    n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
    n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636,
    n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645,
    n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654,
    n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663,
    n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
    n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
    n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
    n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
    n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708,
    n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717,
    n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
    n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
    n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
    n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
    n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
    n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
    n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780,
    n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789,
    n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
    n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807,
    n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
    n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
    n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
    n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
    n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852,
    n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861,
    n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
    n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879,
    n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888,
    n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
    n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
    n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
    n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924,
    n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933,
    n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942,
    n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951,
    n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960,
    n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
    n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
    n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
    n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996,
    n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005,
    n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014,
    n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023,
    n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032,
    n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
    n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
    n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
    n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068,
    n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077,
    n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086,
    n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095,
    n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104,
    n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
    n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
    n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
    n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
    n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149,
    n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158,
    n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167,
    n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
    n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
    n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
    n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
    n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212,
    n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221,
    n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230,
    n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
    n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
    n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
    n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284,
    n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293,
    n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302,
    n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311,
    n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320,
    n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
    n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
    n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
    n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356,
    n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365,
    n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374,
    n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383,
    n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392,
    n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
    n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
    n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419,
    n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428,
    n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437,
    n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446,
    n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455,
    n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464,
    n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
    n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
    n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491,
    n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500,
    n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509,
    n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518,
    n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
    n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536,
    n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
    n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
    n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563,
    n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572,
    n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581,
    n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590,
    n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
    n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
    n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
    n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
    n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644,
    n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653,
    n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662,
    n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671,
    n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
    n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
    n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
    n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707,
    n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716,
    n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724, n41725,
    n41726, n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734,
    n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743,
    n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752,
    n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
    n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
    n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779,
    n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788,
    n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796, n41797,
    n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806,
    n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815,
    n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824,
    n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
    n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
    n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851,
    n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860,
    n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868, n41869,
    n41870, n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878,
    n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887,
    n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896,
    n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
    n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
    n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
    n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932,
    n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940, n41941,
    n41942, n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950,
    n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959,
    n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968,
    n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
    n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
    n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995,
    n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004,
    n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42013,
    n42014, n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022,
    n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031,
    n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
    n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
    n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
    n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
    n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076,
    n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085,
    n42086, n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
    n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103,
    n42104, n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112,
    n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
    n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
    n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139,
    n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148,
    n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157,
    n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
    n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174, n42175,
    n42176, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
    n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
    n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
    n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211,
    n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220,
    n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229,
    n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
    n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246, n42247,
    n42248, n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256,
    n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
    n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
    n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283,
    n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292,
    n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301,
    n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310,
    n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318, n42319,
    n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328,
    n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337,
    n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
    n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
    n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364,
    n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373,
    n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382,
    n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390, n42391,
    n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400,
    n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409,
    n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
    n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427,
    n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436,
    n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444, n42445,
    n42446, n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
    n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462, n42463,
    n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472,
    n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481,
    n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
    n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
    n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508,
    n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517,
    n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526,
    n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535,
    n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544,
    n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553,
    n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
    n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
    n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580,
    n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589,
    n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
    n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607,
    n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616,
    n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625,
    n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
    n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643,
    n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652,
    n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42661,
    n42662, n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
    n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679,
    n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688,
    n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697,
    n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
    n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715,
    n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724,
    n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732, n42733,
    n42734, n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
    n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751,
    n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760,
    n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769,
    n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
    n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787,
    n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796,
    n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804, n42805,
    n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814,
    n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823,
    n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
    n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
    n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
    n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859,
    n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868,
    n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876, n42877,
    n42878, n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886,
    n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895,
    n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904,
    n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
    n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
    n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931,
    n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940,
    n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949,
    n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
    n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967,
    n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976,
    n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985,
    n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
    n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
    n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012,
    n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020, n43021,
    n43022, n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030,
    n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039,
    n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048,
    n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057,
    n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
    n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
    n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084,
    n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092, n43093,
    n43094, n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
    n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111,
    n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120,
    n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
    n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
    n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156,
    n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165,
    n43166, n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174,
    n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182, n43183,
    n43184, n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192,
    n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201,
    n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
    n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
    n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228,
    n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237,
    n43238, n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246,
    n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255,
    n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264,
    n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273,
    n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
    n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
    n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300,
    n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308, n43309,
    n43310, n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318,
    n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326, n43327,
    n43328, n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336,
    n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
    n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
    n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
    n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372,
    n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381,
    n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
    n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399,
    n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
    n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
    n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
    n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
    n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444,
    n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453,
    n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
    n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471,
    n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
    n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
    n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
    n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
    n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516,
    n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525,
    n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
    n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543,
    n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552,
    n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
    n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
    n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588,
    n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597,
    n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
    n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615,
    n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624,
    n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
    n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
    n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
    n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660,
    n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669,
    n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
    n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687,
    n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
    n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
    n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
    n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
    n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732,
    n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741,
    n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
    n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759,
    n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768,
    n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
    n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
    n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
    n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804,
    n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813,
    n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
    n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831,
    n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840,
    n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
    n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
    n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
    n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876,
    n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885,
    n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
    n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903,
    n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
    n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
    n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
    n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
    n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948,
    n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957,
    n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
    n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975,
    n43976, n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984,
    n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993,
    n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
    n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
    n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020,
    n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029,
    n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038,
    n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047,
    n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056,
    n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065,
    n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
    n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
    n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092,
    n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100, n44101,
    n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110,
    n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119,
    n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128,
    n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137,
    n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
    n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
    n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164,
    n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173,
    n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
    n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191,
    n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200,
    n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209,
    n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
    n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
    n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236,
    n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245,
    n44246, n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254,
    n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263,
    n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272,
    n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281,
    n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
    n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
    n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308,
    n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316, n44317,
    n44318, n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326,
    n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335,
    n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344,
    n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353,
    n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
    n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
    n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380,
    n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388, n44389,
    n44390, n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398,
    n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406, n44407,
    n44408, n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416,
    n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425,
    n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
    n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
    n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452,
    n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460, n44461,
    n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
    n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478, n44479,
    n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488,
    n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497,
    n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
    n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
    n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524,
    n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532, n44533,
    n44534, n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542,
    n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551,
    n44552, n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560,
    n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
    n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
    n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
    n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596,
    n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604, n44605,
    n44606, n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614,
    n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622, n44623,
    n44624, n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632,
    n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
    n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
    n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
    n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668,
    n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676, n44677,
    n44678, n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686,
    n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694, n44695,
    n44696, n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704,
    n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713,
    n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
    n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
    n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740,
    n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748, n44749,
    n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758,
    n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766, n44767,
    n44768, n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776,
    n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785,
    n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
    n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
    n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812,
    n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821,
    n44822, n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
    n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838, n44839,
    n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848,
    n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857,
    n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
    n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
    n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884,
    n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892, n44893,
    n44894, n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
    n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910, n44911,
    n44912, n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920,
    n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929,
    n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
    n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
    n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956,
    n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965,
    n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
    n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983,
    n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
    n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
    n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
    n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
    n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028,
    n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037,
    n45038, n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046,
    n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055,
    n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064,
    n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073,
    n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
    n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
    n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100,
    n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109,
    n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118,
    n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127,
    n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136,
    n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145,
    n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
    n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
    n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172,
    n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180, n45181,
    n45182, n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190,
    n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199,
    n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208,
    n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217,
    n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
    n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
    n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244,
    n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252, n45253,
    n45254, n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262,
    n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271,
    n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280,
    n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289,
    n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
    n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307,
    n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316,
    n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324, n45325,
    n45326, n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334,
    n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343,
    n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
    n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361,
    n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
    n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379,
    n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388,
    n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397,
    n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
    n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415,
    n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424,
    n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
    n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
    n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
    n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460,
    n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469,
    n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
    n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487,
    n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496,
    n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505,
    n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
    n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523,
    n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532,
    n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541,
    n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550,
    n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559,
    n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568,
    n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577,
    n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
    n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595,
    n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604,
    n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613,
    n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622,
    n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631,
    n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640,
    n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649,
    n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
    n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667,
    n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676,
    n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685,
    n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
    n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703,
    n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712,
    n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721,
    n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
    n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739,
    n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748,
    n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756, n45757,
    n45758, n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
    n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775,
    n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784,
    n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793,
    n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
    n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811,
    n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820,
    n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828, n45829,
    n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838,
    n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847,
    n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
    n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865,
    n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
    n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883,
    n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892,
    n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900, n45901,
    n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910,
    n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919,
    n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928,
    n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
    n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
    n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955,
    n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964,
    n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973,
    n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
    n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991,
    n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000,
    n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009,
    n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
    n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027,
    n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036,
    n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045,
    n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054,
    n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063,
    n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072,
    n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081,
    n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
    n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099,
    n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108,
    n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116, n46117,
    n46118, n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
    n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135,
    n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144,
    n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153,
    n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
    n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171,
    n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180,
    n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188, n46189,
    n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198,
    n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207,
    n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216,
    n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225,
    n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
    n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243,
    n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252,
    n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261,
    n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270,
    n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279,
    n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288,
    n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297,
    n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
    n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315,
    n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324,
    n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333,
    n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342,
    n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351,
    n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360,
    n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369,
    n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
    n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387,
    n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396,
    n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405,
    n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414,
    n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423,
    n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432,
    n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441,
    n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
    n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459,
    n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468,
    n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477,
    n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486,
    n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495,
    n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504,
    n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513,
    n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
    n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531,
    n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540,
    n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549,
    n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558,
    n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567,
    n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576,
    n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585,
    n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
    n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603,
    n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612,
    n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621,
    n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630,
    n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639,
    n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648,
    n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657,
    n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
    n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675,
    n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684,
    n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693,
    n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702,
    n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711,
    n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720,
    n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729,
    n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
    n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747,
    n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756,
    n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765,
    n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774,
    n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783,
    n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792,
    n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801,
    n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
    n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
    n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828,
    n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837,
    n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846,
    n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855,
    n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864,
    n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873,
    n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
    n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891,
    n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900,
    n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909,
    n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918,
    n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927,
    n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936,
    n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945,
    n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
    n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
    n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972,
    n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981,
    n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990,
    n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999,
    n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008,
    n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017,
    n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
    n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035,
    n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044,
    n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052, n47053,
    n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062,
    n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071,
    n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080,
    n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
    n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
    n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107,
    n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116,
    n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125,
    n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
    n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143,
    n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152,
    n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
    n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
    n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179,
    n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188,
    n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197,
    n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206,
    n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215,
    n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224,
    n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233,
    n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
    n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251,
    n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260,
    n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269,
    n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
    n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287,
    n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296,
    n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305,
    n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
    n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323,
    n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332,
    n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340, n47341,
    n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350,
    n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359,
    n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
    n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
    n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
    n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395,
    n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404,
    n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413,
    n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422,
    n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431,
    n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440,
    n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449,
    n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
    n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467,
    n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476,
    n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484, n47485,
    n47486, n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494,
    n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503,
    n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512,
    n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521,
    n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
    n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539,
    n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548,
    n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557,
    n47558, n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566,
    n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575,
    n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584,
    n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593,
    n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
    n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611,
    n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620,
    n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629,
    n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638,
    n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647,
    n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656,
    n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
    n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
    n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683,
    n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692,
    n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701,
    n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710,
    n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719,
    n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728,
    n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737,
    n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
    n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755,
    n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764,
    n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773,
    n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782,
    n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791,
    n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800,
    n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809,
    n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
    n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827,
    n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836,
    n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845,
    n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
    n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863,
    n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872,
    n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881,
    n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
    n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899,
    n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908,
    n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917,
    n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926,
    n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935,
    n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944,
    n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953,
    n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
    n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971,
    n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980,
    n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989,
    n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998,
    n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007,
    n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016,
    n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025,
    n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
    n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043,
    n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052,
    n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061,
    n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070,
    n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079,
    n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088,
    n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097,
    n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
    n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115,
    n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124,
    n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133,
    n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
    n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151,
    n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
    n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169,
    n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
    n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187,
    n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196,
    n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205,
    n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214,
    n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223,
    n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232,
    n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241,
    n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
    n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259,
    n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268,
    n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277,
    n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286,
    n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295,
    n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304,
    n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313,
    n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
    n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331,
    n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340,
    n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349,
    n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358,
    n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367,
    n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376,
    n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385,
    n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
    n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403,
    n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412,
    n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421,
    n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430,
    n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439,
    n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448,
    n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457,
    n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
    n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475,
    n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484,
    n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493,
    n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502,
    n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511,
    n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520,
    n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529,
    n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
    n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547,
    n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556,
    n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565,
    n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574,
    n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583,
    n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592,
    n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601,
    n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
    n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619,
    n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628,
    n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637,
    n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646,
    n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655,
    n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664,
    n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673,
    n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
    n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691,
    n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700,
    n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709,
    n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718,
    n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727,
    n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
    n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745,
    n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
    n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763,
    n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772,
    n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781,
    n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790,
    n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799,
    n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808,
    n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817,
    n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
    n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835,
    n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844,
    n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853,
    n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862,
    n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871,
    n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880,
    n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889,
    n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
    n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907,
    n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916,
    n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925,
    n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934,
    n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943,
    n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952,
    n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961,
    n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
    n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979,
    n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988,
    n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997,
    n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006,
    n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015,
    n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024,
    n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033,
    n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
    n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051,
    n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060,
    n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069,
    n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078,
    n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087,
    n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096,
    n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105,
    n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
    n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123,
    n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132,
    n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141,
    n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150,
    n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159,
    n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168,
    n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177,
    n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
    n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195,
    n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204,
    n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213,
    n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222,
    n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231,
    n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240,
    n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249,
    n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
    n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267,
    n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276,
    n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285,
    n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294,
    n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303,
    n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312,
    n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321,
    n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
    n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339,
    n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348,
    n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357,
    n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366,
    n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375,
    n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384,
    n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393,
    n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
    n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411,
    n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420,
    n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429,
    n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438,
    n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447,
    n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456,
    n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465,
    n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
    n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483,
    n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492,
    n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500, n49501,
    n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510,
    n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519,
    n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528,
    n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537,
    n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
    n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555,
    n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564,
    n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573,
    n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582,
    n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591,
    n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600,
    n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609,
    n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
    n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627,
    n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636,
    n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645,
    n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654,
    n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663,
    n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672,
    n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681,
    n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
    n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699,
    n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708,
    n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716, n49717,
    n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726,
    n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735,
    n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744,
    n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753,
    n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
    n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771,
    n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780,
    n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789,
    n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
    n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807,
    n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816,
    n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825,
    n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
    n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843,
    n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852,
    n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860, n49861,
    n49862, n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870,
    n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879,
    n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888,
    n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897,
    n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
    n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915,
    n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924,
    n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933,
    n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942,
    n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951,
    n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960,
    n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969,
    n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
    n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987,
    n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996,
    n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004, n50005,
    n50006, n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
    n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023,
    n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032,
    n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041,
    n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
    n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059,
    n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068,
    n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076, n50077,
    n50078, n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086,
    n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095,
    n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104,
    n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113,
    n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
    n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131,
    n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140,
    n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148, n50149,
    n50150, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158,
    n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167,
    n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
    n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185,
    n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
    n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203,
    n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212,
    n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221,
    n50222, n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230,
    n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239,
    n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248,
    n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257,
    n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
    n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275,
    n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284,
    n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292, n50293,
    n50294, n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302,
    n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311,
    n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
    n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329,
    n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
    n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347,
    n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356,
    n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365,
    n50366, n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374,
    n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383,
    n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
    n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401,
    n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
    n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419,
    n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428,
    n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437,
    n50438, n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446,
    n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455,
    n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464,
    n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473,
    n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
    n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491,
    n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500,
    n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508, n50509,
    n50510, n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518,
    n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527,
    n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536,
    n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545,
    n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
    n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
    n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572,
    n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581,
    n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590,
    n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599,
    n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
    n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617,
    n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
    n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635,
    n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644,
    n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652, n50653,
    n50654, n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662,
    n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671,
    n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680,
    n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689,
    n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
    n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
    n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716,
    n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724, n50725,
    n50726, n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734,
    n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743,
    n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752,
    n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761,
    n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
    n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779,
    n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788,
    n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797,
    n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806,
    n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815,
    n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824,
    n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833,
    n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
    n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851,
    n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860,
    n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868, n50869,
    n50870, n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878,
    n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887,
    n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896,
    n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905,
    n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
    n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923,
    n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932,
    n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940, n50941,
    n50942, n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950,
    n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959,
    n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968,
    n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977,
    n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
    n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995,
    n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004,
    n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012, n51013,
    n51014, n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022,
    n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031,
    n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040,
    n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049,
    n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
    n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067,
    n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076,
    n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51085,
    n51086, n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094,
    n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103,
    n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112,
    n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121,
    n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
    n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139,
    n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148,
    n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157,
    n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166,
    n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175,
    n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184,
    n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193,
    n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
    n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211,
    n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220,
    n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228, n51229,
    n51230, n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238,
    n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247,
    n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256,
    n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265,
    n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
    n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283,
    n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292,
    n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301,
    n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310,
    n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319,
    n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328,
    n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337,
    n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
    n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355,
    n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364,
    n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373,
    n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382,
    n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391,
    n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400,
    n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409,
    n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
    n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427,
    n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436,
    n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445,
    n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454,
    n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463,
    n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472,
    n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481,
    n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
    n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499,
    n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508,
    n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517,
    n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526,
    n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535,
    n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544,
    n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553,
    n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
    n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571,
    n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580,
    n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589,
    n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598,
    n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607,
    n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616,
    n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625,
    n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
    n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643,
    n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652,
    n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661,
    n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670,
    n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679,
    n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688,
    n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697,
    n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
    n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715,
    n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724,
    n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733,
    n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742,
    n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751,
    n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760,
    n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769,
    n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
    n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787,
    n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796,
    n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805,
    n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814,
    n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823,
    n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832,
    n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841,
    n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
    n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859,
    n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868,
    n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877,
    n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886,
    n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895,
    n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904,
    n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913,
    n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
    n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931,
    n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940,
    n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949,
    n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958,
    n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967,
    n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976,
    n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985,
    n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
    n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003,
    n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012,
    n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021,
    n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030,
    n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039,
    n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048,
    n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057,
    n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
    n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075,
    n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084,
    n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093,
    n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102,
    n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111,
    n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120,
    n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129,
    n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
    n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147,
    n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156,
    n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165,
    n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174,
    n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183,
    n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192,
    n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201,
    n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
    n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219,
    n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228,
    n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237,
    n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246,
    n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255,
    n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264,
    n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273,
    n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
    n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291,
    n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
    n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309,
    n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318,
    n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327,
    n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336,
    n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345,
    n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
    n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363,
    n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372,
    n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381,
    n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390,
    n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399,
    n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408,
    n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417,
    n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
    n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435,
    n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444,
    n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453,
    n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462,
    n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471,
    n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480,
    n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489,
    n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
    n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507,
    n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
    n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525,
    n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534,
    n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543,
    n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552,
    n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561,
    n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
    n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579,
    n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
    n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597,
    n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606,
    n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615,
    n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624,
    n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633,
    n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
    n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651,
    n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660,
    n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669,
    n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678,
    n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687,
    n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696,
    n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705,
    n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
    n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723,
    n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732,
    n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741,
    n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750,
    n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759,
    n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768,
    n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777,
    n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
    n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795,
    n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804,
    n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813,
    n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822,
    n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831,
    n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840,
    n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849,
    n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
    n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867,
    n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876,
    n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885,
    n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894,
    n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903,
    n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912,
    n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921,
    n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
    n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939,
    n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948,
    n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957,
    n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966,
    n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975,
    n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984,
    n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993,
    n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
    n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011,
    n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020,
    n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029,
    n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038,
    n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047,
    n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056,
    n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065,
    n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
    n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083,
    n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
    n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101,
    n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110,
    n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119,
    n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128,
    n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137,
    n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
    n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155,
    n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164,
    n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173,
    n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182,
    n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191,
    n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200,
    n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
    n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
    n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227,
    n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
    n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245,
    n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254,
    n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263,
    n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272,
    n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281,
    n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
    n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299,
    n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308,
    n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317,
    n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326,
    n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335,
    n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344,
    n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353,
    n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
    n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371,
    n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380,
    n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389,
    n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398,
    n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407,
    n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416,
    n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425,
    n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
    n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443,
    n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452,
    n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461,
    n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470,
    n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479,
    n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488,
    n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497,
    n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
    n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515,
    n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524,
    n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533,
    n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542,
    n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550, n53551,
    n53552, n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560,
    n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569,
    n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
    n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587,
    n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596,
    n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605,
    n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614,
    n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623,
    n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632,
    n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641,
    n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
    n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659,
    n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668,
    n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677,
    n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686,
    n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695,
    n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704,
    n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713,
    n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
    n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731,
    n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740,
    n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749,
    n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758,
    n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766, n53767,
    n53768, n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776,
    n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785,
    n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
    n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803,
    n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812,
    n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821,
    n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830,
    n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838, n53839,
    n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848,
    n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857,
    n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
    n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875,
    n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884,
    n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893,
    n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902,
    n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911,
    n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920,
    n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929,
    n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
    n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947,
    n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956,
    n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965,
    n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974,
    n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983,
    n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992,
    n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001,
    n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
    n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019,
    n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028,
    n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037,
    n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046,
    n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055,
    n54056, n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064,
    n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073,
    n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
    n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091,
    n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100,
    n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108, n54109,
    n54110, n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118,
    n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127,
    n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136,
    n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145,
    n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
    n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163,
    n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172,
    n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181,
    n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190,
    n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199,
    n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208,
    n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217,
    n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
    n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235,
    n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244,
    n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, n54253,
    n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262,
    n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271,
    n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280,
    n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289,
    n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
    n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307,
    n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316,
    n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324, n54325,
    n54326, n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334,
    n54335, n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343,
    n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352,
    n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361,
    n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
    n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379,
    n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388,
    n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396, n54397,
    n54398, n54399, n54400, n54401, n54402, n54403, n54404, n54405, n54406,
    n54407, n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415,
    n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424,
    n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433,
    n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
    n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451,
    n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460,
    n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468, n54469,
    n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478,
    n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487,
    n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496,
    n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505,
    n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
    n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523,
    n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532,
    n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541,
    n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550,
    n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559,
    n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568,
    n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
    n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
    n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595,
    n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604,
    n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613,
    n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622,
    n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631,
    n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640,
    n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649,
    n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
    n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667,
    n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676,
    n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685,
    n54686, n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694,
    n54695, n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703,
    n54704, n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712,
    n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721,
    n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
    n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739,
    n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748,
    n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756, n54757,
    n54758, n54759, n54760, n54761, n54762, n54763, n54764, n54765, n54766,
    n54767, n54768, n54769, n54770, n54771, n54772, n54773, n54774, n54775,
    n54776, n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784,
    n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793,
    n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
    n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811,
    n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820,
    n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828, n54829,
    n54830, n54831, n54832, n54833, n54834, n54835, n54836, n54837, n54838,
    n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846, n54847,
    n54848, n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856,
    n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865,
    n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
    n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883,
    n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892,
    n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900, n54901,
    n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54910,
    n54911, n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919,
    n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928,
    n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937,
    n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
    n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955,
    n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964,
    n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972, n54973,
    n54974, n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982,
    n54983, n54984, n54985, n54986, n54987, n54988, n54989, n54990, n54991,
    n54992, n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000,
    n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009,
    n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
    n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027,
    n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036,
    n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044, n55045,
    n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053, n55054,
    n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062, n55063,
    n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072,
    n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081,
    n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090,
    n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099,
    n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108,
    n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116, n55117,
    n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125, n55126,
    n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135,
    n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144,
    n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153,
    n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162,
    n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171,
    n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180,
    n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189,
    n55190, n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198,
    n55199, n55200, n55201, n55202, n55203, n55204, n55205, n55206, n55207,
    n55208, n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216,
    n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225,
    n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234,
    n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243,
    n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252,
    n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261,
    n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269, n55270,
    n55271, n55272, n55273, n55274, n55275, n55276, n55277, n55278, n55279,
    n55280, n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288,
    n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297,
    n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
    n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315,
    n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324,
    n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333,
    n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342,
    n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351,
    n55352, n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360,
    n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369,
    n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
    n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387,
    n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396,
    n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404, n55405,
    n55406, n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414,
    n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422, n55423,
    n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432,
    n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441,
    n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450,
    n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459,
    n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468,
    n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476, n55477,
    n55478, n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486,
    n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494, n55495,
    n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504,
    n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513,
    n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522,
    n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531,
    n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540,
    n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549,
    n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558,
    n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567,
    n55568, n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576,
    n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585,
    n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594,
    n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603,
    n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612,
    n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620, n55621,
    n55622, n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630,
    n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639,
    n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648,
    n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657,
    n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666,
    n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675,
    n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684,
    n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692, n55693,
    n55694, n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702,
    n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711,
    n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720,
    n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729,
    n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738,
    n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747,
    n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756,
    n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764, n55765,
    n55766, n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774,
    n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782, n55783,
    n55784, n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792,
    n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801,
    n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810,
    n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819,
    n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828,
    n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836, n55837,
    n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845, n55846,
    n55847, n55848, n55849, n55850, n55851, n55852, n55853, n55854, n55855,
    n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864,
    n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873,
    n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
    n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891,
    n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900,
    n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909,
    n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918,
    n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927,
    n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936,
    n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945,
    n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954,
    n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963,
    n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972,
    n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981,
    n55982, n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990,
    n55991, n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999,
    n56000, n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008,
    n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017,
    n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026,
    n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035,
    n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044,
    n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053,
    n56054, n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062,
    n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071,
    n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080,
    n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089,
    n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098,
    n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107,
    n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116,
    n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125,
    n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134,
    n56135, n56136, n56137, n56138, n56139, n56140, n56141, n56142, n56143,
    n56144, n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152,
    n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161,
    n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170,
    n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179,
    n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188,
    n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196, n56197,
    n56198, n56199, n56200, n56201, n56202, n56203, n56204, n56205, n56206,
    n56207, n56208, n56209, n56210, n56211, n56212, n56213, n56214, n56215,
    n56216, n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224,
    n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233,
    n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
    n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251,
    n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260,
    n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268, n56269,
    n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277, n56278,
    n56279, n56280, n56281, n56282, n56283, n56284, n56285, n56286, n56287,
    n56288, n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296,
    n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305,
    n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314,
    n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323,
    n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332,
    n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340, n56341,
    n56342, n56343, n56344, n56345, n56346, n56347, n56348, n56349, n56350,
    n56351, n56352, n56353, n56354, n56355, n56356, n56357, n56358, n56359,
    n56360, n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368,
    n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377,
    n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386,
    n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394, n56395,
    n56396, n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404,
    n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412, n56413,
    n56414, n56415, n56416, n56417, n56418, n56419, n56420, n56421, n56422,
    n56423, n56424, n56425, n56426, n56427, n56428, n56429, n56430, n56431,
    n56432, n56433, n56434, n56435, n56436, n56437, n56438, n56439, n56440,
    n56441, n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449,
    n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458,
    n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466, n56467,
    n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476,
    n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484, n56485,
    n56486, n56487, n56488, n56489, n56490, n56491, n56492, n56493, n56494,
    n56495, n56496, n56497, n56498, n56499, n56500, n56501, n56502, n56503,
    n56504, n56505, n56506, n56507, n56508, n56509, n56510, n56511, n56512,
    n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521,
    n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
    n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539,
    n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548,
    n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556, n56557,
    n56558, n56559, n56560, n56561, n56562, n56563, n56564, n56565, n56566,
    n56567, n56568, n56569, n56570, n56571, n56572, n56573, n56574, n56575,
    n56576, n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584,
    n56585, n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593,
    n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
    n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611,
    n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620,
    n56621, n56622, n56623, n56624, n56625, n56626, n56627, n56628, n56629,
    n56630, n56631, n56632, n56633, n56634, n56635, n56636, n56637, n56638,
    n56639, n56640, n56641, n56642, n56643, n56644, n56645, n56646, n56647,
    n56648, n56649, n56650, n56651, n56652, n56653, n56654, n56655, n56656,
    n56657, n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665,
    n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674,
    n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683,
    n56684, n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692,
    n56693, n56694, n56695, n56696, n56697, n56698, n56699, n56700, n56701,
    n56702, n56703, n56704, n56705, n56706, n56707, n56708, n56709, n56710,
    n56711, n56712, n56713, n56714, n56715, n56716, n56717, n56718, n56719,
    n56720, n56721, n56722, n56723, n56724, n56725, n56726, n56727, n56728,
    n56729, n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737,
    n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746,
    n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754, n56755,
    n56756, n56757, n56758, n56759, n56760, n56761, n56762, n56763, n56764,
    n56765, n56766, n56767, n56768, n56769, n56770, n56771, n56772, n56773,
    n56774, n56775, n56776, n56777, n56778, n56779, n56780, n56781, n56782,
    n56783, n56784, n56785, n56786, n56787, n56788, n56789, n56790, n56791,
    n56792, n56793, n56794, n56795, n56796, n56797, n56798, n56799, n56800,
    n56801, n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809,
    n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818,
    n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826, n56827,
    n56828, n56829, n56830, n56831, n56832, n56833, n56834, n56835, n56836,
    n56837, n56838, n56839, n56840, n56841, n56842, n56843, n56844, n56845,
    n56846, n56847, n56848, n56849, n56850, n56851, n56852, n56853, n56854,
    n56855, n56856, n56857, n56858, n56859, n56860, n56861, n56862, n56863,
    n56864, n56865, n56866, n56867, n56868, n56869, n56870, n56871, n56872,
    n56873, n56874, n56875, n56876, n56877, n56878, n56879, n56880, n56881,
    n56882, n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890,
    n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898, n56899,
    n56900, n56901, n56902, n56903, n56904, n56905, n56906, n56907, n56908,
    n56909, n56910, n56911, n56912, n56913, n56914, n56915, n56916, n56917,
    n56918, n56919, n56920, n56921, n56922, n56923, n56924, n56925, n56926,
    n56927, n56928, n56929, n56930, n56931, n56932, n56933, n56934, n56935,
    n56936, n56937, n56938, n56939, n56940, n56941, n56942, n56943, n56944,
    n56945, n56946, n56947, n56948, n56949, n56950, n56951, n56952, n56953,
    n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962,
    n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970, n56971,
    n56972, n56973, n56974, n56975, n56976, n56977, n56978, n56979, n56980,
    n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988, n56989,
    n56990, n56991, n56992, n56993, n56994, n56995, n56996, n56997, n56998,
    n56999, n57000, n57001, n57002, n57003, n57004, n57005, n57006, n57007,
    n57008, n57009, n57010, n57011, n57012, n57013, n57014, n57015, n57016,
    n57017, n57018, n57019, n57020, n57021, n57022, n57023, n57024, n57025,
    n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034,
    n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042, n57043,
    n57044, n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052,
    n57053, n57054, n57055, n57056, n57057, n57058, n57059, n57060, n57061,
    n57062, n57063, n57064, n57065, n57066, n57067, n57068, n57069, n57070,
    n57071, n57072, n57073, n57074, n57075, n57076, n57077, n57078, n57079,
    n57080, n57081, n57082, n57083, n57084, n57085, n57086, n57087, n57088,
    n57089, n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097,
    n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
    n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115,
    n57116, n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124,
    n57125, n57126, n57127, n57128, n57129, n57130, n57131, n57132, n57133,
    n57134, n57135, n57136, n57137, n57138, n57139, n57140, n57141, n57142,
    n57143, n57144, n57145, n57146, n57147, n57148, n57149, n57150, n57151,
    n57152, n57153, n57154, n57155, n57156, n57157, n57158, n57159, n57160,
    n57161, n57162, n57163, n57164, n57165, n57166, n57167, n57168, n57169,
    n57170, n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178,
    n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186, n57187,
    n57188, n57189, n57190, n57191, n57192, n57193, n57194, n57195, n57196,
    n57197, n57198, n57199, n57200, n57201, n57202, n57203, n57204, n57205,
    n57206, n57207, n57208, n57209, n57210, n57211, n57212, n57213, n57214,
    n57215, n57216, n57217, n57218, n57219, n57220, n57221, n57222, n57223,
    n57224, n57225, n57226, n57227, n57228, n57229, n57230, n57231, n57232,
    n57233, n57234, n57235, n57236, n57237, n57238, n57239, n57240, n57241,
    n57242, n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250,
    n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258, n57259,
    n57260, n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268,
    n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276, n57277,
    n57278, n57279, n57280, n57281, n57282, n57283, n57284, n57285, n57286,
    n57287, n57288, n57289, n57290, n57291, n57292, n57293, n57294, n57295,
    n57296, n57297, n57298, n57299, n57300, n57301, n57302, n57303, n57304,
    n57305, n57306, n57307, n57308, n57309, n57310, n57311, n57312, n57313,
    n57314, n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322,
    n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330, n57331,
    n57332, n57333, n57334, n57335, n57336, n57337, n57338, n57339, n57340,
    n57341, n57342, n57343, n57344, n57345, n57346, n57347, n57348, n57349,
    n57350, n57351, n57352, n57353, n57354, n57355, n57356, n57357, n57358,
    n57359, n57360, n57361, n57362, n57363, n57364, n57365, n57366, n57367,
    n57368, n57369, n57370, n57371, n57372, n57373, n57374, n57375, n57376,
    n57377, n57378, n57379, n57380, n57381, n57382, n57383, n57384, n57385,
    n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394,
    n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402, n57403,
    n57404, n57405, n57406, n57407, n57408, n57409, n57410, n57411, n57412,
    n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420, n57421,
    n57422, n57423, n57424, n57425, n57426, n57427, n57428, n57429, n57430,
    n57431, n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439,
    n57440, n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448,
    n57449, n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457,
    n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
    n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474, n57475,
    n57476, n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484,
    n57485, n57486, n57487, n57488, n57489, n57490, n57491, n57492, n57493,
    n57494, n57495, n57496, n57497, n57498, n57499, n57500, n57501, n57502,
    n57503, n57504, n57505, n57506, n57507, n57508, n57509, n57510, n57511,
    n57512, n57513, n57514, n57515, n57516, n57517, n57518, n57519, n57520,
    n57521, n57522, n57523, n57524, n57525, n57526, n57527, n57528, n57529,
    n57530, n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538,
    n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546, n57547,
    n57548, n57549, n57550, n57551, n57552, n57553, n57554, n57555, n57556,
    n57557, n57558, n57559, n57560, n57561, n57562, n57563, n57564, n57565,
    n57566, n57567, n57568, n57569, n57570, n57571, n57572, n57573, n57574,
    n57575, n57576, n57577, n57578, n57579, n57580, n57581, n57582, n57583,
    n57584, n57585, n57586, n57587, n57588, n57589, n57590, n57591, n57592,
    n57593, n57594, n57595, n57596, n57597, n57598, n57599, n57600, n57601,
    n57602, n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610,
    n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618, n57619,
    n57620, n57621, n57622, n57623, n57624, n57625, n57626, n57627, n57628,
    n57629, n57630, n57631, n57632, n57633, n57634, n57635, n57636, n57637,
    n57638, n57639, n57640, n57641, n57642, n57643, n57644, n57645, n57646,
    n57647, n57648, n57649, n57650, n57651, n57652, n57653, n57654, n57655,
    n57656, n57657, n57658, n57659, n57660, n57661, n57662, n57663, n57664,
    n57665, n57666, n57667, n57668, n57669, n57670, n57671, n57672, n57673,
    n57674, n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682,
    n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690, n57691,
    n57692, n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700,
    n57701, n57702, n57703, n57704, n57705, n57706, n57707, n57708, n57709,
    n57710, n57711, n57712, n57713, n57714, n57715, n57716, n57717, n57718,
    n57719, n57720, n57721, n57722, n57723, n57724, n57725, n57726, n57727,
    n57728, n57729, n57730, n57731, n57732, n57733, n57734, n57735, n57736,
    n57737, n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745,
    n57746, n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
    n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762, n57763,
    n57764, n57765, n57766, n57767, n57768, n57769, n57770, n57771, n57772,
    n57773, n57774, n57775, n57776, n57777, n57778, n57779, n57780, n57781,
    n57782, n57783, n57784, n57785, n57786, n57787, n57788, n57789, n57790,
    n57791, n57792, n57793, n57794, n57795, n57796, n57797, n57798, n57799,
    n57800, n57801, n57802, n57803, n57804, n57805, n57806, n57807, n57808,
    n57809, n57810, n57811, n57812, n57813, n57814, n57815, n57816, n57817,
    n57818, n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826,
    n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834, n57835,
    n57836, n57837, n57838, n57839, n57840, n57841, n57842, n57843, n57844,
    n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852, n57853,
    n57854, n57855, n57856, n57857, n57858, n57859, n57860, n57861, n57862,
    n57863, n57864, n57865, n57866, n57867, n57868, n57869, n57870, n57871,
    n57872, n57873, n57874, n57875, n57876, n57877, n57878, n57879, n57880,
    n57881, n57882, n57883, n57884, n57885, n57886, n57887, n57888, n57889,
    n57890, n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
    n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906, n57907,
    n57908, n57909, n57910, n57911, n57912, n57913, n57914, n57915, n57916,
    n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924, n57925,
    n57926, n57927, n57928, n57929, n57930, n57931, n57932, n57933, n57934,
    n57935, n57936, n57937, n57938, n57939, n57940, n57941, n57942, n57943,
    n57944, n57945, n57946, n57947, n57948, n57949, n57950, n57951, n57952,
    n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961,
    n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
    n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978, n57979,
    n57980, n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988,
    n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997,
    n57998, n57999, n58000, n58001, n58002, n58003, n58004, n58005, n58006,
    n58007, n58008, n58009, n58010, n58011, n58012, n58013, n58014, n58015,
    n58016, n58017, n58018, n58019, n58020, n58021, n58022, n58023, n58024,
    n58025, n58026, n58027, n58028, n58029, n58030, n58031, n58032, n58033,
    n58034, n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042,
    n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050, n58051,
    n58052, n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060,
    n58061, n58062, n58063, n58064, n58065, n58066, n58067, n58068, n58069,
    n58070, n58071, n58072, n58073, n58074, n58075, n58076, n58077, n58078,
    n58079, n58080, n58081, n58082, n58083, n58084, n58085, n58086, n58087,
    n58088, n58089, n58090, n58091, n58092, n58093, n58094, n58095, n58096,
    n58097, n58098, n58099, n58100, n58101, n58102, n58103, n58104, n58105,
    n58106, n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114,
    n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122, n58123,
    n58124, n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132,
    n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140, n58141,
    n58142, n58143, n58144, n58145, n58146, n58147, n58148, n58149, n58150,
    n58151, n58152, n58153, n58154, n58155, n58156, n58157, n58158, n58159,
    n58160, n58161, n58162, n58163, n58164, n58165, n58166, n58167, n58168,
    n58169, n58170, n58171, n58172, n58173, n58174, n58175, n58176, n58177,
    n58178, n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186,
    n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194, n58195,
    n58196, n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204,
    n58205, n58206, n58207, n58208, n58209, n58210, n58211, n58212, n58213,
    n58214, n58215, n58216, n58217, n58218, n58219, n58220, n58221, n58222,
    n58223, n58224, n58225, n58226, n58227, n58228, n58229, n58230, n58231,
    n58232, n58233, n58234, n58235, n58236, n58237, n58238, n58239, n58240,
    n58241, n58242, n58243, n58244, n58245, n58246, n58247, n58248, n58249,
    n58250, n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258,
    n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266, n58267,
    n58268, n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276,
    n58277, n58278, n58279, n58280, n58281, n58282, n58283, n58284, n58285,
    n58286, n58287, n58288, n58289, n58290, n58291, n58292, n58293, n58294,
    n58295, n58296, n58297, n58298, n58299, n58300, n58301, n58302, n58303,
    n58304, n58305, n58306, n58307, n58308, n58309, n58310, n58311, n58312,
    n58313, n58314, n58315, n58316, n58317, n58318, n58319, n58320, n58321,
    n58322, n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330,
    n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338, n58339,
    n58340, n58341, n58342, n58343, n58344, n58345, n58346, n58347, n58348,
    n58349, n58350, n58351, n58352, n58353, n58354, n58355, n58356, n58357,
    n58358, n58359, n58360, n58361, n58362, n58363, n58364, n58365, n58366,
    n58367, n58368, n58369, n58370, n58371, n58372, n58373, n58374, n58375,
    n58376, n58377, n58378, n58379, n58380, n58381, n58382, n58383, n58384,
    n58385, n58386, n58387, n58388, n58389, n58390, n58391, n58392, n58393,
    n58394, n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402,
    n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410, n58411,
    n58412, n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420,
    n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428, n58429,
    n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437, n58438,
    n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446, n58447,
    n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455, n58456,
    n58457, n58458, n58459, n58460, n58461, n58462, n58463, n58464, n58465,
    n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
    n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482, n58483,
    n58484, n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492,
    n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500, n58501,
    n58502, n58503, n58504, n58505, n58506, n58507, n58508, n58509, n58510,
    n58511, n58512, n58513, n58514, n58515, n58516, n58517, n58518, n58519,
    n58520, n58521, n58522, n58523, n58524, n58525, n58526, n58527, n58528,
    n58529, n58530, n58531, n58532, n58533, n58534, n58535, n58536, n58537,
    n58538, n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
    n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554, n58555,
    n58556, n58557, n58558, n58559, n58560, n58561, n58562, n58563, n58564,
    n58565, n58566, n58567, n58568, n58569, n58570, n58571, n58572, n58573,
    n58574, n58575, n58576, n58577, n58578, n58579, n58580, n58581, n58582,
    n58583, n58584, n58585, n58586, n58587, n58588, n58589, n58590, n58591,
    n58592, n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600,
    n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608, n58609,
    n58610, n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618,
    n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626, n58627,
    n58628, n58629, n58630, n58631, n58632, n58633, n58634, n58635, n58636,
    n58637, n58638, n58639, n58640, n58641, n58642, n58643, n58644, n58645,
    n58646, n58647, n58648, n58649, n58650, n58651, n58652, n58653, n58654,
    n58655, n58656, n58657, n58658, n58659, n58660, n58661, n58662, n58663,
    n58664, n58665, n58666, n58667, n58668, n58669, n58670, n58671, n58672,
    n58673, n58674, n58675, n58676, n58677, n58678, n58679, n58680, n58681,
    n58682, n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690,
    n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698, n58699,
    n58700, n58701, n58702, n58703, n58704, n58705, n58706, n58707, n58708,
    n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716, n58717,
    n58718, n58719, n58720, n58721, n58722, n58723, n58724, n58725, n58726,
    n58727, n58728, n58729, n58730, n58731, n58732, n58733, n58734, n58735,
    n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58743, n58744,
    n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752, n58753,
    n58754, n58755, n58756, n58757, n58758, n58759, n58760, n58761, n58762,
    n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770, n58771,
    n58772, n58773, n58774, n58775, n58776, n58777, n58778, n58779, n58780,
    n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788, n58789,
    n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797, n58798,
    n58799, n58800, n58801, n58802, n58803, n58804, n58805, n58806, n58807,
    n58808, n58809, n58810, n58811, n58812, n58813, n58814, n58815, n58816,
    n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824, n58825,
    n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833, n58834,
    n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842, n58843,
    n58844, n58845, n58846, n58847, n58848, n58849, n58850, n58851, n58852,
    n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860, n58861,
    n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869, n58870,
    n58871, n58872, n58873, n58874, n58875, n58876, n58877, n58878, n58879,
    n58880, n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888,
    n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896, n58897,
    n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906,
    n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914, n58915,
    n58916, n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924,
    n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932, n58933,
    n58934, n58935, n58936, n58937, n58938, n58939, n58940, n58941, n58942,
    n58943, n58944, n58945, n58946, n58947, n58948, n58949, n58950, n58951,
    n58952, n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960,
    n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968, n58969,
    n58970, n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978,
    n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986, n58987,
    n58988, n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996,
    n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004, n59005,
    n59006, n59007, n59008, n59009, n59010, n59011, n59012, n59013, n59014,
    n59015, n59016, n59017, n59018, n59019, n59020, n59021, n59022, n59023,
    n59024, n59025, n59026, n59027, n59028, n59029, n59030, n59031, n59032,
    n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040, n59041,
    n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049, n59050,
    n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058, n59059,
    n59060, n59061, n59062, n59063, n59064, n59065, n59066, n59067, n59068,
    n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076, n59077,
    n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085, n59086,
    n59087, n59088, n59089, n59090, n59091, n59092, n59093, n59094, n59095,
    n59096, n59097, n59098, n59099, n59100, n59101, n59102, n59103, n59104,
    n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112, n59113,
    n59114, n59115, n59116, n59117, n59118, n59119, n59120, n59121, n59122,
    n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130, n59131,
    n59132, n59133, n59134, n59135, n59136, n59137, n59138, n59139, n59140,
    n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148, n59149,
    n59150, n59151, n59152, n59153, n59154, n59155, n59156, n59157, n59158,
    n59159, n59160, n59161, n59162, n59163, n59164, n59165, n59166, n59167,
    n59168, n59169, n59170, n59171, n59172, n59173, n59174, n59175, n59176,
    n59177, n59178, n59179, n59180, n59181, n59182, n59183, n59184, n59185,
    n59186, n59187, n59188, n59189, n59190, n59191, n59192, n59193, n59194,
    n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202, n59203,
    n59204, n59205, n59206, n59207, n59208, n59209, n59210, n59211, n59212,
    n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220, n59221,
    n59222, n59223, n59224, n59225, n59226, n59227, n59228, n59229, n59230,
    n59231, n59232, n59233, n59234, n59235, n59236, n59237, n59238, n59239,
    n59240, n59241, n59242, n59243, n59244, n59245, n59246, n59247, n59248,
    n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256, n59257,
    n59258, n59259, n59260, n59261, n59262, n59263, n59264, n59265, n59266,
    n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274, n59275,
    n59276, n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284,
    n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292, n59293,
    n59294, n59295, n59296, n59297, n59298, n59299, n59300, n59301, n59302,
    n59303, n59304, n59305, n59306, n59307, n59308, n59309, n59310, n59311,
    n59312, n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59320,
    n59321, n59322, n59323, n59324, n59325, n59326, n59327, n59328, n59329,
    n59330, n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338,
    n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346, n59347,
    n59348, n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356,
    n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364, n59365,
    n59366, n59367, n59368, n59369, n59370, n59371, n59372, n59373, n59374,
    n59375, n59376, n59377, n59378, n59379, n59380, n59381, n59382, n59383,
    n59384, n59385, n59386, n59387, n59388, n59389, n59390, n59391, n59392,
    n59393, n59394, n59395, n59396, n59397, n59398, n59399, n59400, n59401,
    n59402, n59403, n59404, n59405, n59406, n59407, n59408, n59409, n59410,
    n59411, n59412, n59413, n59414, n59415, n59416, n59417, n59418, n59419,
    n59420, n59421, n59422, n59423, n59424, n59425, n59426, n59427, n59428,
    n59429, n59430, n59431, n59432, n59433, n59434, n59435, n59436, n59437,
    n59438, n59439, n59440, n59441, n59442, n59443, n59444, n59445, n59446,
    n59447, n59448, n59449, n59450, n59451, n59452, n59453, n59454, n59455,
    n59456, n59457, n59458, n59459, n59460, n59461, n59462, n59463, n59464,
    n59465, n59466, n59467, n59468, n59469, n59470, n59471, n59472, n59473,
    n59474, n59475, n59476, n59477, n59478, n59479, n59480, n59481, n59482,
    n59483, n59484, n59485, n59486, n59487, n59488, n59489, n59490, n59491,
    n59492, n59493, n59494, n59495, n59496, n59497, n59498, n59499, n59500,
    n59501, n59502, n59503, n59504, n59505, n59506, n59507, n59508, n59509,
    n59510, n59511, n59512, n59513, n59514, n59515, n59516, n59517, n59518,
    n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526, n59527,
    n59528, n59529, n59530, n59531, n59532, n59533, n59534, n59535, n59536,
    n59537, n59538, n59539, n59540, n59541, n59542, n59543, n59544, n59545,
    n59546, n59547, n59548, n59549, n59550, n59551, n59552, n59553, n59554,
    n59555, n59556, n59557, n59558, n59559, n59560, n59561, n59562, n59563,
    n59564, n59565, n59566, n59567, n59568, n59569, n59570, n59571, n59572,
    n59573, n59574, n59575, n59576, n59577, n59578, n59579, n59580, n59581,
    n59582, n59583, n59584, n59585, n59586, n59587, n59588, n59589, n59590,
    n59591, n59592, n59593, n59594, n59595, n59596, n59597, n59598, n59599,
    n59600, n59601, n59602, n59603, n59604, n59605, n59606, n59607, n59608,
    n59609, n59610, n59611, n59612, n59613, n59614, n59615, n59616, n59617,
    n59618, n59619, n59620, n59621, n59622, n59623, n59624, n59625, n59626,
    n59627, n59628, n59629, n59630, n59631, n59632, n59633, n59634, n59635,
    n59636, n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644,
    n59645, n59646, n59647, n59648, n59649, n59650, n59651, n59652, n59653,
    n59654, n59655, n59656, n59657, n59658, n59659, n59660, n59661, n59662,
    n59663, n59664, n59665, n59666, n59667, n59668, n59669, n59670, n59671,
    n59672, n59673, n59674, n59675, n59676, n59677, n59678, n59679, n59680,
    n59681, n59682, n59683, n59684, n59685, n59686, n59687, n59688, n59689,
    n59690, n59691, n59692, n59693, n59694, n59695, n59696, n59697, n59698,
    n59699, n59700, n59701, n59702, n59703, n59704, n59705, n59706, n59707,
    n59708, n59709, n59710, n59711, n59712, n59713, n59714, n59715, n59716,
    n59717, n59718, n59719, n59720, n59721, n59722, n59723, n59724, n59725,
    n59726, n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734,
    n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742, n59743,
    n59744, n59745, n59746, n59747, n59748, n59749, n59750, n59751, n59752,
    n59753, n59754, n59755, n59756, n59757, n59758, n59759, n59760, n59761,
    n59762, n59763, n59764, n59765, n59766, n59767, n59768, n59769, n59770,
    n59771, n59772, n59773, n59774, n59775, n59776, n59777, n59778, n59779,
    n59780, n59781, n59782, n59783, n59784, n59785, n59786, n59787, n59788,
    n59789, n59790, n59791, n59792, n59793, n59794, n59795, n59796, n59797,
    n59798, n59799, n59800, n59801, n59802, n59803, n59804, n59805, n59806,
    n59807, n59808, n59809, n59810, n59811, n59812, n59813, n59814, n59815,
    n59816, n59817, n59818, n59819, n59820, n59821, n59822, n59823, n59824,
    n59825, n59826, n59827, n59828, n59829, n59830, n59831, n59832, n59833,
    n59834, n59835, n59836, n59837, n59838, n59839, n59840, n59841, n59842,
    n59843, n59844, n59845, n59846, n59847, n59848, n59849, n59850, n59851,
    n59852, n59853, n59854, n59855, n59856, n59857, n59858, n59859, n59860,
    n59861, n59862, n59863, n59864, n59865, n59866, n59867, n59868, n59869,
    n59870, n59871, n59872, n59873, n59874, n59875, n59876, n59877, n59878,
    n59879, n59880, n59881, n59882, n59883, n59884, n59885, n59886, n59887,
    n59888, n59889, n59890, n59891, n59892, n59893, n59894, n59895, n59896,
    n59897, n59898, n59899, n59900, n59901, n59902, n59903, n59904, n59905,
    n59906, n59907, n59908, n59909, n59910, n59911, n59912, n59913, n59914,
    n59915, n59916, n59917, n59918, n59919, n59920, n59921, n59922, n59923,
    n59924, n59925, n59926, n59927, n59928, n59929, n59930, n59931, n59932,
    n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59940, n59941,
    n59942, n59943, n59944, n59945, n59946, n59947, n59948, n59949, n59950,
    n59951, n59952, n59953, n59954, n59955, n59956, n59957, n59958, n59959,
    n59960, n59961, n59962, n59963, n59964, n59965, n59966, n59967, n59968,
    n59969, n59970, n59971, n59972, n59973, n59974, n59975, n59976, n59977,
    n59978, n59979, n59980, n59981, n59982, n59983, n59984, n59985, n59986,
    n59987, n59988, n59989, n59990, n59991, n59992, n59993, n59994, n59995,
    n59996, n59997, n59998, n59999, n60000, n60001, n60002, n60003, n60004,
    n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012, n60013,
    n60014, n60015, n60016, n60017, n60018, n60019, n60020, n60021, n60022,
    n60023, n60024, n60025, n60026, n60027, n60028, n60029, n60030, n60031,
    n60032, n60033, n60034, n60035, n60036, n60037, n60038, n60039, n60040,
    n60041, n60042, n60043, n60044, n60045, n60046, n60047, n60048, n60049,
    n60050, n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058,
    n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066, n60067,
    n60068, n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076,
    n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084, n60085,
    n60086, n60087, n60088, n60089, n60090, n60091, n60092, n60093, n60094,
    n60095, n60096, n60097, n60098, n60099, n60100, n60101, n60102, n60103,
    n60104, n60105, n60106, n60107, n60108, n60109, n60110, n60111, n60112,
    n60113, n60114, n60115, n60116, n60117, n60118, n60119, n60120, n60121,
    n60122, n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130,
    n60131, n60132, n60133, n60134, n60135, n60136, n60137, n60138, n60139,
    n60140, n60141, n60142, n60143, n60144, n60145, n60146, n60147, n60148,
    n60149, n60150, n60151, n60152, n60153, n60154, n60155, n60156, n60157,
    n60158, n60159, n60160, n60161, n60162, n60163, n60164, n60165, n60166,
    n60167, n60168, n60169, n60170, n60171, n60172, n60173, n60174, n60175,
    n60176, n60177, n60178, n60179, n60180, n60181, n60182, n60183, n60184,
    n60185, n60186, n60187, n60188, n60189, n60190, n60191, n60192, n60193,
    n60194, n60195, n60196, n60197, n60198, n60199, n60200, n60201, n60202,
    n60203, n60204, n60205, n60206, n60207, n60208, n60209, n60210, n60211,
    n60212, n60213, n60214, n60215, n60216, n60217, n60218, n60219, n60220,
    n60221, n60222, n60223, n60224, n60225, n60226, n60227, n60228, n60229,
    n60230, n60231, n60232, n60233, n60234, n60235, n60236, n60237, n60238,
    n60239, n60240, n60241, n60242, n60243, n60244, n60245, n60246, n60247,
    n60248, n60249, n60250, n60251, n60252, n60253, n60254, n60255, n60256,
    n60257, n60258, n60259, n60260, n60261, n60262, n60263, n60264, n60265,
    n60266, n60267, n60268, n60269, n60270, n60271, n60272, n60273, n60274,
    n60275, n60276, n60277, n60278, n60279, n60280, n60281, n60282, n60283,
    n60284, n60285, n60286, n60287, n60288, n60289, n60290, n60291, n60292,
    n60293, n60294, n60295, n60296, n60297, n60298, n60299, n60300, n60301,
    n60302, n60303, n60304, n60305, n60306, n60307, n60308, n60309, n60310,
    n60311, n60312, n60313, n60314, n60315, n60316, n60317, n60318, n60319,
    n60320, n60321, n60322, n60323, n60324, n60325, n60326, n60327, n60328,
    n60329, n60330, n60331, n60332, n60333, n60334, n60335, n60336, n60337,
    n60338, n60339, n60340, n60341, n60342, n60343, n60344, n60345, n60346,
    n60347, n60348, n60349, n60350, n60351, n60352, n60353, n60354, n60355,
    n60356, n60357, n60358, n60359, n60360, n60361, n60362, n60363, n60364,
    n60365, n60366, n60367, n60368, n60369, n60370, n60371, n60372, n60373,
    n60374, n60375, n60376, n60377, n60378, n60379, n60380, n60381, n60382,
    n60383, n60384, n60385, n60386, n60387, n60388, n60389, n60390, n60391,
    n60392, n60393, n60394, n60395, n60396, n60397, n60398, n60399, n60400,
    n60401, n60402, n60403, n60404, n60405, n60406, n60407, n60408, n60409,
    n60410, n60411, n60412, n60413, n60414, n60415, n60416, n60417, n60418,
    n60419, n60420, n60421, n60422, n60423, n60424, n60425, n60426, n60427,
    n60428, n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60436,
    n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444, n60445,
    n60446, n60447, n60448, n60449, n60450, n60451, n60452, n60453, n60454,
    n60455, n60456, n60457, n60458, n60459, n60460, n60461, n60462, n60463,
    n60464, n60465, n60466, n60467, n60468, n60469, n60470, n60471, n60472,
    n60473, n60474, n60475, n60476, n60477, n60478, n60479, n60480, n60481,
    n60482, n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490,
    n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498, n60499,
    n60500, n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508,
    n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516, n60517,
    n60518, n60519, n60520, n60521, n60522, n60523, n60524, n60525, n60526,
    n60527, n60528, n60529, n60530, n60531, n60532, n60533, n60534, n60535,
    n60536, n60537, n60538, n60539, n60540, n60541, n60542, n60543, n60544,
    n60545, n60546, n60547, n60548, n60549, n60550, n60551, n60552, n60553,
    n60554, n60555, n60556, n60557, n60558, n60559, n60560, n60561, n60562,
    n60563, n60564, n60565, n60566, n60567, n60568, n60569, n60570, n60571,
    n60572, n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580,
    n60581, n60582, n60583, n60584, n60585, n60586, n60587, n60588, n60589,
    n60590, n60591, n60592, n60593, n60594, n60595, n60596, n60597, n60598,
    n60599, n60600, n60601, n60602, n60603, n60604, n60605, n60606, n60607,
    n60608, n60609, n60610, n60611, n60612, n60613, n60614, n60615, n60616,
    n60617, n60618, n60619, n60620, n60621, n60622, n60623, n60624, n60625,
    n60626, n60627, n60628, n60629, n60630, n60631, n60632, n60633, n60634,
    n60635, n60636, n60637, n60638, n60639, n60640, n60641, n60642, n60643,
    n60644, n60645, n60646, n60647, n60648, n60649, n60650, n60651, n60652,
    n60653, n60654, n60655, n60656, n60657, n60658, n60659, n60660, n60661,
    n60662, n60663, n60664, n60665, n60666, n60667, n60668, n60669, n60670,
    n60671, n60672, n60673, n60674, n60675, n60676, n60677, n60678, n60679,
    n60680, n60681, n60682, n60683, n60684, n60685, n60686, n60687, n60688,
    n60689, n60690, n60691, n60692, n60693, n60694, n60695, n60696, n60697,
    n60698, n60699, n60700, n60701, n60702, n60703, n60704, n60705, n60706,
    n60707, n60708, n60709, n60710, n60711, n60712, n60713, n60714, n60715,
    n60716, n60717, n60718, n60719, n60720, n60721, n60722, n60723, n60724,
    n60725, n60726, n60727, n60728, n60729, n60730, n60731, n60732, n60733,
    n60734, n60735, n60736, n60737, n60738, n60739, n60740, n60741, n60742,
    n60743, n60744, n60745, n60746, n60747, n60748, n60749, n60750, n60751,
    n60752, n60753, n60754, n60755, n60756, n60757, n60758, n60759, n60760,
    n60761, n60762, n60763, n60764, n60765, n60766, n60767, n60768, n60769,
    n60770, n60771, n60772, n60773, n60774, n60775, n60776, n60777, n60778,
    n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786, n60787,
    n60788, n60789, n60790, n60791, n60792, n60793, n60794, n60795, n60796,
    n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60804, n60805,
    n60806, n60807, n60808, n60809, n60810, n60811, n60812, n60813, n60814,
    n60815, n60816, n60817, n60818, n60819, n60820, n60821, n60822, n60823,
    n60824, n60825, n60826, n60827, n60828, n60829, n60830, n60831, n60832,
    n60833, n60834, n60835, n60836, n60837, n60838, n60839, n60840, n60841,
    n60842, n60843, n60844, n60845, n60846, n60847, n60848, n60849, n60850,
    n60851, n60852, n60853, n60854, n60855, n60856, n60857, n60858, n60859,
    n60860, n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868,
    n60869, n60870, n60871, n60872, n60873, n60874, n60875, n60876, n60877,
    n60878, n60879, n60880, n60881, n60882, n60883, n60884, n60885, n60886,
    n60887, n60888, n60889, n60890, n60891, n60892, n60893, n60894, n60895,
    n60896, n60897, n60898, n60899, n60900, n60901, n60902, n60903, n60904,
    n60905, n60906, n60907, n60908, n60909, n60910, n60911, n60912, n60913,
    n60914, n60915, n60916, n60917, n60918, n60919, n60920, n60921, n60922,
    n60923, n60924, n60925, n60926, n60927, n60928, n60929, n60930, n60931,
    n60932, n60933, n60934, n60935, n60936, n60937, n60938, n60939, n60940,
    n60941, n60942, n60943, n60944, n60945, n60946, n60947, n60948, n60949,
    n60950, n60951, n60952, n60953, n60954, n60955, n60956, n60957, n60958,
    n60959, n60960, n60961, n60962, n60963, n60964, n60965, n60966, n60967,
    n60968, n60969, n60970, n60971, n60972, n60973, n60974, n60975, n60976,
    n60977, n60978, n60979, n60980, n60981, n60982, n60983, n60984, n60985,
    n60986, n60987, n60988, n60989, n60990, n60991, n60992, n60993, n60994,
    n60995, n60996, n60997, n60998, n60999, n61000, n61001, n61002, n61003,
    n61004, n61005, n61006, n61007, n61008, n61009, n61010, n61011, n61012,
    n61013, n61014, n61015, n61016, n61017, n61018, n61019, n61020, n61021,
    n61022, n61023, n61024, n61025, n61026, n61027, n61028, n61029, n61030,
    n61031, n61032, n61033, n61034, n61035, n61036, n61037, n61038, n61039,
    n61040, n61041, n61042, n61043, n61044, n61045, n61046, n61047, n61048,
    n61049, n61050, n61051, n61052, n61053, n61054, n61055, n61056, n61057,
    n61058, n61059, n61060, n61061, n61062, n61063, n61064, n61065, n61066,
    n61067, n61068, n61069, n61070, n61071, n61072, n61073, n61074, n61075,
    n61076, n61077, n61078, n61079, n61080, n61081, n61082, n61083, n61084,
    n61085, n61086, n61087, n61088, n61089, n61090, n61091, n61092, n61093,
    n61094, n61095, n61096, n61097, n61098, n61099, n61100, n61101, n61102,
    n61103, n61104, n61105, n61106, n61107, n61108, n61109, n61110, n61111,
    n61112, n61113, n61114, n61115, n61116, n61117, n61118, n61119, n61120,
    n61121, n61122, n61123, n61124, n61125, n61126, n61127, n61128, n61129,
    n61130, n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138,
    n61139, n61140, n61141, n61142, n61143, n61144, n61145, n61146, n61147,
    n61148, n61149, n61150, n61151, n61152, n61153, n61154, n61155, n61156,
    n61157, n61158, n61159, n61160, n61161, n61162, n61163, n61164, n61165,
    n61166, n61167, n61168, n61169, n61170, n61171, n61172, n61173, n61174,
    n61175, n61176, n61177, n61178, n61179, n61180, n61181, n61182, n61183,
    n61184, n61185, n61186, n61187, n61188, n61189, n61190, n61191, n61192,
    n61193, n61194, n61195, n61196, n61197, n61198, n61199, n61200, n61201,
    n61202, n61203, n61204, n61205, n61206, n61207, n61208, n61209, n61210,
    n61211, n61212, n61213, n61214, n61215, n61216, n61217, n61218, n61219,
    n61220, n61221, n61222, n61223, n61224, n61225, n61226, n61227, n61228,
    n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236, n61237,
    n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61245, n61246,
    n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61254, n61255,
    n61256, n61257, n61258, n61259, n61260, n61261, n61262, n61263, n61264,
    n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272, n61273,
    n61274, n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282,
    n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290, n61291,
    n61292, n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300,
    n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308, n61309,
    n61310, n61311, n61312, n61313, n61314, n61315, n61316, n61317, n61318,
    n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326, n61327,
    n61328, n61329, n61330, n61331, n61332, n61333, n61334, n61335, n61336,
    n61337, n61338, n61339, n61340, n61341, n61342, n61343, n61344, n61345,
    n61346, n61347, n61348, n61349, n61350, n61351, n61352, n61353, n61354,
    n61355, n61356, n61357, n61358, n61359, n61360, n61361, n61362, n61363,
    n61364, n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372,
    n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380, n61381,
    n61382, n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390,
    n61391, n61392, n61393, n61394, n61395, n61396, n61397, n61398, n61399,
    n61400, n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408,
    n61409, n61410, n61411, n61412, n61413, n61414, n61415, n61416, n61417,
    n61418, n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426,
    n61427, n61428, n61429, n61430, n61431, n61432, n61433, n61434, n61435,
    n61436, n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444,
    n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452, n61453,
    n61454, n61455, n61456, n61457, n61458, n61459, n61460, n61461, n61462,
    n61463, n61464, n61465, n61466, n61467, n61468, n61469, n61470, n61471,
    n61472, n61473, n61474, n61475, n61476, n61477, n61478, n61479, n61480,
    n61481, n61482, n61483, n61484, n61485, n61486, n61487, n61488, n61489,
    n61490, n61491, n61492, n61493, n61494, n61495, n61496, n61497, n61498,
    n61499, n61500, n61501, n61502, n61503, n61504, n61505, n61506, n61507,
    n61508, n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516,
    n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524, n61525,
    n61526, n61527, n61528, n61529, n61530, n61531, n61532, n61533, n61534,
    n61535, n61536, n61537, n61538, n61539, n61540, n61541, n61542, n61543,
    n61544, n61545, n61546, n61547, n61548, n61549, n61550, n61551, n61552,
    n61553, n61554, n61555, n61556, n61557, n61558, n61559, n61560, n61561,
    n61562, n61563, n61564, n61565, n61566, n61567, n61568, n61569, n61570,
    n61571, n61572, n61573, n61574, n61575, n61576, n61577, n61578, n61579,
    n61580, n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588,
    n61589, n61590, n61591, n61592, n61593, n61594, n61595, n61596, n61597,
    n61598, n61599, n61600, n61601, n61602, n61603, n61604, n61605, n61606,
    n61607, n61608, n61609, n61610, n61611, n61612, n61613, n61614, n61615,
    n61616, n61617, n61618, n61619, n61620, n61621, n61622, n61623, n61624,
    n61625, n61626, n61627, n61628, n61629, n61630, n61631, n61632, n61633,
    n61634, n61635, n61636, n61637, n61638, n61639, n61640, n61641, n61642,
    n61643, n61644, n61645, n61646, n61647, n61648, n61649, n61650, n61651,
    n61652, n61653, n61654, n61655, n61656, n61657, n61658, n61659, n61660,
    n61661, n61662, n61663, n61664, n61665, n61666, n61667, n61668, n61669,
    n61670, n61671, n61672, n61673, n61674, n61675, n61676, n61677, n61678,
    n61679, n61680, n61681, n61682, n61683, n61684, n61685, n61686, n61687,
    n61688, n61689, n61690, n61691, n61692, n61693, n61694, n61695, n61696,
    n61697, n61698, n61699, n61700, n61701, n61702, n61703, n61704, n61705,
    n61706, n61707, n61708, n61709, n61710, n61711, n61712, n61713, n61714,
    n61715, n61716, n61717, n61718, n61719, n61720, n61721, n61722, n61723,
    n61724, n61725, n61726, n61727, n61728, n61729, n61730, n61731, n61732,
    n61733, n61734, n61735, n61736, n61737, n61738, n61739, n61740, n61741,
    n61742, n61743, n61744, n61745, n61746, n61747, n61748, n61749, n61750,
    n61751, n61752, n61753, n61754, n61755, n61756, n61757, n61758, n61759,
    n61760, n61761, n61762, n61763, n61764, n61765, n61766, n61767, n61768,
    n61769, n61770, n61771, n61772, n61773, n61774, n61775, n61776, n61777,
    n61778, n61779, n61780, n61781, n61782, n61783, n61784, n61785, n61786,
    n61787, n61788, n61789, n61790, n61791, n61792, n61793, n61794, n61795,
    n61796, n61797, n61798, n61799, n61800, n61801, n61802, n61803, n61804,
    n61805, n61806, n61807, n61808, n61809, n61810, n61811, n61812, n61813,
    n61814, n61815, n61816, n61817, n61818, n61819, n61820, n61821, n61822,
    n61823, n61824, n61825, n61826, n61827, n61828, n61829, n61830, n61831,
    n61832, n61833, n61834, n61835, n61836, n61837, n61838, n61839, n61840,
    n61841, n61842, n61843, n61844, n61845, n61846, n61847, n61848, n61849,
    n61850, n61851, n61852, n61853, n61854, n61855, n61856, n61857, n61858,
    n61859, n61860, n61861, n61862, n61863, n61864, n61865, n61866, n61867,
    n61868, n61869, n61870, n61871, n61872, n61873, n61874, n61875, n61876,
    n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884, n61885,
    n61886, n61887, n61888, n61889, n61890, n61891, n61892, n61893, n61894,
    n61895, n61896, n61897, n61898, n61899, n61900, n61901, n61902, n61903,
    n61904, n61905, n61906, n61907, n61908, n61909, n61910, n61911, n61912,
    n61913, n61914, n61915, n61916, n61917, n61918, n61919, n61920, n61921,
    n61922, n61923, n61924, n61925, n61926, n61927, n61928, n61929, n61930,
    n61931, n61932, n61933, n61934, n61935, n61936, n61937, n61938, n61939,
    n61940, n61941, n61942, n61943, n61944, n61945, n61946, n61947, n61948,
    n61949, n61950, n61951, n61952, n61953, n61954, n61955, n61956, n61957,
    n61958, n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966,
    n61967, n61968, n61969, n61970, n61971, n61972, n61973, n61974, n61975,
    n61976, n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984,
    n61985, n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993,
    n61994, n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62002,
    n62003, n62004, n62005, n62006, n62007, n62008, n62009, n62010, n62011,
    n62012, n62013, n62014, n62015, n62016, n62017, n62018, n62019, n62020,
    n62021, n62022, n62023, n62024, n62025, n62026, n62027, n62028, n62029,
    n62030, n62031, n62032, n62033, n62034, n62035, n62036, n62037, n62038,
    n62039, n62040, n62041, n62042, n62043, n62044, n62045, n62046, n62047,
    n62048, n62049, n62050, n62051, n62052, n62053, n62054, n62055, n62056,
    n62057, n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065,
    n62066, n62067, n62068, n62069, n62070, n62071, n62072, n62073, n62074,
    n62075, n62076, n62077, n62078, n62079, n62080, n62081, n62082, n62083,
    n62084, n62085, n62086, n62087, n62088, n62089, n62090, n62091, n62092,
    n62093, n62094, n62095, n62096, n62097, n62098, n62099, n62100, n62101,
    n62102, n62103, n62104, n62105, n62106, n62107, n62108, n62109, n62110,
    n62111, n62112, n62113, n62114, n62115, n62116, n62117, n62118, n62119,
    n62120, n62121, n62122, n62123, n62124, n62125, n62126, n62127, n62128,
    n62129, n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137,
    n62138, n62139, n62140, n62141, n62142, n62143, n62144, n62145, n62146,
    n62147, n62148, n62149, n62150, n62151, n62152, n62153, n62154, n62155,
    n62156, n62157, n62158, n62159, n62160, n62161, n62162, n62163, n62164,
    n62165, n62166, n62167, n62168, n62169, n62170, n62171, n62172, n62173,
    n62174, n62175, n62176, n62177, n62178, n62179, n62180, n62181, n62182,
    n62183, n62184, n62185, n62186, n62187, n62188, n62189, n62190, n62191,
    n62192, n62193, n62194, n62195, n62196, n62197, n62198, n62199, n62200,
    n62201, n62202, n62203, n62204, n62205, n62206, n62207, n62208, n62209,
    n62210, n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218,
    n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226, n62227,
    n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235, n62236,
    n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244, n62245,
    n62246, n62247, n62248, n62249, n62250, n62251, n62252, n62253, n62254,
    n62255, n62256, n62257, n62258, n62259, n62260, n62261, n62262, n62263,
    n62264, n62265, n62266, n62267, n62268, n62269, n62270, n62271, n62272,
    n62273, n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281,
    n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290,
    n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299,
    n62300, n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308,
    n62309, n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317,
    n62318, n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326,
    n62327, n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335,
    n62336, n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344,
    n62345, n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353,
    n62354, n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362,
    n62363, n62364, n62365, n62366, n62367, n62368, n62369, n62370, n62371,
    n62372, n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380,
    n62381, n62382, n62383, n62384, n62385, n62386, n62387, n62388, n62389,
    n62390, n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398,
    n62399, n62400, n62401, n62402, n62403, n62404, n62405, n62406, n62407,
    n62408, n62409, n62410, n62411, n62412, n62413, n62414, n62415, n62416,
    n62417, n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425,
    n62426, n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434,
    n62435, n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443,
    n62444, n62445, n62446, n62447, n62448, n62449, n62450, n62451, n62452,
    n62453, n62454, n62455, n62456, n62457, n62458, n62459, n62460, n62461,
    n62462, n62463, n62464, n62465, n62466, n62467, n62468, n62469, n62470,
    n62471, n62472, n62473, n62474, n62475, n62476, n62477, n62478, n62479,
    n62480, n62481, n62482, n62483, n62484, n62485, n62486, n62487, n62488,
    n62489, n62490, n62491, n62492, n62493, n62494, n62495, n62496, n62497,
    n62498, n62499, n62500, n62501, n62502, n62503, n62504, n62505, n62506,
    n62507, n62508, n62509, n62510, n62511, n62512, n62513, n62514, n62515,
    n62516, n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524,
    n62525, n62526, n62527, n62528, n62529, n62530, n62531, n62532, n62533,
    n62534, n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542,
    n62543, n62544, n62545, n62546, n62547, n62548, n62549, n62550, n62551,
    n62552, n62553, n62554, n62555, n62556, n62557, n62558, n62559, n62560,
    n62561, n62562, n62563, n62564, n62565, n62566, n62567, n62568, n62569,
    n62570, n62571, n62572, n62573, n62574, n62575, n62576, n62577, n62578,
    n62579, n62580, n62581, n62582, n62583, n62584, n62585, n62586, n62587,
    n62588, n62589, n62590, n62591, n62592, n62593, n62594, n62595, n62596,
    n62597, n62598, n62599, n62600, n62601, n62602, n62603, n62604, n62605,
    n62606, n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614,
    n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622, n62623,
    n62624, n62625, n62626, n62627, n62628, n62629, n62630, n62631, n62632,
    n62633, n62634, n62635, n62636, n62637, n62638, n62639, n62640, n62641,
    n62642, n62643, n62644, n62645, n62646, n62647, n62648, n62649, n62650,
    n62651, n62652, n62653, n62654, n62655, n62656, n62657, n62658, n62659,
    n62660, n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668,
    n62669, n62670, n62671, n62672, n62673, n62674, n62675, n62676, n62677,
    n62678, n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686,
    n62687, n62688, n62689, n62690, n62691, n62692, n62693, n62694, n62695,
    n62696, n62697, n62698, n62699, n62700, n62701, n62702, n62703, n62704,
    n62705, n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713,
    n62714, n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722,
    n62723, n62724, n62725, n62726, n62727, n62728, n62729, n62730, n62731,
    n62732, n62733, n62734, n62735, n62736, n62737, n62738, n62739, n62740,
    n62741, n62742, n62743, n62744, n62745, n62746, n62747, n62748, n62749,
    n62750, n62751, n62752, n62753, n62754, n62755, n62756, n62757, n62758,
    n62759, n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767,
    n62768, n62769, n62770, n62771, n62772, n62773, n62774, n62775, n62776,
    n62777, n62778, n62779, n62780, n62781, n62782, n62783, n62784, n62785,
    n62786, n62787, n62788, n62789, n62790, n62791, n62792, n62793, n62794,
    n62795, n62796, n62797, n62798, n62799, n62800, n62801, n62802, n62803,
    n62804, n62805, n62806, n62807, n62808, n62809, n62810, n62811, n62812,
    n62813, n62814, n62815, n62816, n62817, n62818, n62819, n62820, n62821,
    n62822, n62823, n62824, n62825, n62826, n62827, n62828, n62829, n62830,
    n62831, n62832, n62833, n62834, n62835, n62836, n62837, n62838, n62839,
    n62840, n62841, n62842, n62843, n62844, n62845, n62846, n62847, n62848,
    n62849, n62850, n62851, n62852, n62853, n62854, n62855, n62856, n62857,
    n62858, n62859, n62860, n62861, n62862, n62863, n62864, n62865, n62866,
    n62867, n62868, n62869, n62870, n62871, n62872, n62873, n62874, n62875,
    n62876, n62877, n62878, n62879, n62880, n62881, n62882, n62883, n62884,
    n62885, n62886, n62887, n62888, n62889, n62890, n62891, n62892, n62893,
    n62894, n62895, n62896, n62897, n62898, n62899, n62900, n62901, n62902,
    n62903, n62904, n62905, n62906, n62907, n62908, n62909, n62910, n62911,
    n62912, n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920,
    n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928, n62929,
    n62930, n62931, n62932, n62933, n62934, n62935, n62936, n62937, n62938,
    n62939, n62940, n62941, n62942, n62943, n62944, n62945, n62946, n62947,
    n62948, n62949, n62950, n62951, n62952, n62953, n62954, n62955, n62956,
    n62957, n62958, n62959, n62960, n62961, n62962, n62963, n62964, n62965,
    n62966, n62967, n62968, n62969, n62970, n62971, n62972, n62973, n62974,
    n62975, n62976, n62977, n62978, n62979, n62980, n62981, n62982, n62983,
    n62984, n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992,
    n62993, n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001,
    n63002, n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010,
    n63011, n63012, n63013, n63014, n63015, n63016, n63017, n63018, n63019,
    n63020, n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028,
    n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036, n63037,
    n63038, n63039, n63040, n63041, n63042, n63043, n63044, n63045, n63046,
    n63047, n63048, n63049, n63050, n63051, n63052, n63053, n63054, n63055,
    n63056, n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064,
    n63065, n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073,
    n63074, n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082,
    n63083, n63084, n63085, n63086, n63087, n63088, n63089, n63090, n63091,
    n63092, n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100,
    n63101, n63102, n63103, n63104, n63105, n63106, n63107, n63108, n63109,
    n63110, n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63118,
    n63119, n63120, n63121, n63122, n63123, n63124, n63125, n63126, n63127,
    n63128, n63129, n63130, n63131, n63132, n63133, n63134, n63135, n63136,
    n63137, n63138, n63139, n63140, n63141, n63142, n63143, n63144, n63145,
    n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153, n63154,
    n63155, n63156, n63157, n63158, n63159, n63160, n63161, n63162, n63163,
    n63164, n63165, n63166, n63167, n63168, n63169, n63170, n63171, n63172,
    n63173, n63174, n63175, n63176, n63177, n63178, n63179, n63180, n63181,
    n63182, n63183, n63184, n63185, n63186, n63187, n63188, n63189, n63190,
    n63191, n63192, n63193, n63194, n63195, n63196, n63197, n63198, n63199,
    n63200, n63201, n63202, n63203, n63204, n63205, n63206, n63207, n63208,
    n63209, n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217,
    n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225, n63226,
    n63227, n63228, n63229, n63230, n63231, n63232, n63233, n63234, n63235,
    n63236, n63237, n63238, n63239, n63240, n63241, n63242, n63243, n63244,
    n63245, n63246, n63247, n63248, n63249, n63250, n63251, n63252, n63253,
    n63254, n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262,
    n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270, n63271,
    n63272, n63273, n63274, n63275, n63276, n63277, n63278, n63279, n63280,
    n63281, n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289,
    n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298,
    n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306, n63307,
    n63308, n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316,
    n63317, n63318, n63319, n63320, n63321, n63322, n63323, n63324, n63325,
    n63326, n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63334,
    n63335, n63336, n63337, n63338, n63339, n63340, n63341, n63342, n63343,
    n63344, n63345, n63346, n63347, n63348, n63349, n63350, n63351, n63352,
    n63353, n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361,
    n63362, n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370,
    n63371, n63372, n63373, n63374, n63375, n63376, n63377, n63378, n63379,
    n63380, n63381, n63382, n63383, n63384, n63385, n63386, n63387, n63388,
    n63389, n63390, n63391, n63392, n63393, n63394, n63395, n63396, n63397,
    n63398, n63399, n63400, n63401, n63402, n63403, n63404, n63405, n63406,
    n63407, n63408, n63409, n63410, n63411, n63412, n63413, n63414, n63415,
    n63416, n63417, n63418, n63419, n63420, n63421, n63422, n63423, n63424,
    n63425, n63426, n63427, n63428, n63429, n63430, n63431, n63432, n63433,
    n63434, n63435, n63436, n63437, n63438, n63439, n63440, n63441, n63442,
    n63443, n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451,
    n63452, n63453, n63454, n63455, n63456, n63457, n63458, n63459, n63460,
    n63461, n63462, n63463, n63464, n63465, n63466, n63467, n63468, n63469,
    n63470, n63471, n63472, n63473, n63474, n63475, n63476, n63477, n63478,
    n63479, n63480, n63481, n63482, n63483, n63484, n63485, n63486, n63487,
    n63488, n63489, n63490, n63491, n63492, n63493, n63494, n63495, n63496,
    n63497, n63498, n63499, n63500, n63501, n63502, n63503, n63504, n63505,
    n63506, n63507, n63508, n63509, n63510, n63511, n63512, n63513, n63514,
    n63515, n63516, n63517, n63518, n63519, n63520, n63521, n63522, n63523,
    n63524, n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532,
    n63533, n63534, n63535, n63536, n63537, n63538, n63539, n63540, n63541,
    n63542, n63543, n63544, n63545, n63546, n63547, n63548, n63549, n63550,
    n63551, n63552, n63553, n63554, n63555, n63556, n63557, n63558, n63559,
    n63560, n63561, n63562, n63563, n63564, n63565, n63566, n63567, n63568,
    n63569, n63570, n63571, n63572, n63573, n63574, n63575, n63576, n63577,
    n63578, n63579, n63580, n63581, n63582, n63583, n63584, n63585, n63586,
    n63587, n63588, n63589, n63590, n63591, n63592, n63593, n63594, n63595,
    n63596, n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604,
    n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612, n63613,
    n63614, n63615, n63616, n63617, n63618, n63619, n63620, n63621, n63622,
    n63623, n63624, n63625, n63626, n63627, n63628, n63629, n63630, n63631,
    n63632, n63633, n63634, n63635, n63636, n63637, n63638, n63639, n63640,
    n63641, n63642, n63643, n63644, n63645, n63646, n63647, n63648, n63649,
    n63650, n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658,
    n63659, n63660, n63661, n63662, n63663, n63664, n63665, n63666, n63667,
    n63668, n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676,
    n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684, n63685,
    n63686, n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694,
    n63695, n63696, n63697, n63698, n63699, n63700, n63701, n63702, n63703,
    n63704, n63705, n63706, n63707, n63708, n63709, n63710, n63711, n63712,
    n63713, n63714, n63715, n63716, n63717, n63718, n63719, n63720, n63721,
    n63722, n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730,
    n63731, n63732, n63733, n63734, n63735, n63736, n63737, n63738, n63739,
    n63740, n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748,
    n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756, n63757,
    n63758, n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766,
    n63767, n63768, n63769, n63770, n63771, n63772, n63773, n63774, n63775,
    n63776, n63777, n63778, n63779, n63780, n63781, n63782, n63783, n63784,
    n63785, n63786, n63787, n63788, n63789, n63790, n63791, n63792, n63793,
    n63794, n63795, n63796, n63797, n63798, n63799, n63800, n63801, n63802,
    n63803, n63804, n63805, n63806, n63807, n63808, n63809, n63810, n63811,
    n63812, n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
    n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828, n63829,
    n63830, n63831, n63832, n63833, n63834, n63835, n63836, n63837, n63838,
    n63839, n63840, n63841, n63842, n63843, n63844, n63845, n63846, n63847,
    n63848, n63849, n63850, n63851, n63852, n63853, n63854, n63855, n63856,
    n63857, n63858, n63859, n63860, n63861, n63862, n63863, n63864, n63865,
    n63866, n63867, n63868, n63869, n63870, n63871, n63872, n63873, n63874,
    n63875, n63876, n63877, n63878, n63879, n63880, n63881, n63882, n63883,
    n63884, n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892,
    n63893, n63894, n63895, n63896, n63897, n63898, n63899, n63900, n63901,
    n63902, n63903, n63904, n63905, n63906, n63907, n63908, n63909, n63910,
    n63911, n63912, n63913, n63914, n63915, n63916, n63917, n63918, n63919,
    n63920, n63921, n63922, n63923, n63924, n63925, n63926, n63927, n63928,
    n63929, n63930, n63931, n63932, n63933, n63934, n63935, n63936, n63937,
    n63938, n63939, n63940, n63941, n63942, n63943, n63944, n63945, n63946,
    n63947, n63948, n63949, n63950, n63951, n63952, n63953, n63954, n63955,
    n63956, n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964,
    n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972, n63973,
    n63974, n63975, n63976, n63977, n63978, n63979, n63980, n63981, n63982,
    n63983, n63984, n63985, n63986, n63987, n63988, n63989, n63990, n63991,
    n63992, n63993, n63994, n63995, n63996, n63997, n63998, n63999, n64000,
    n64001, n64002, n64003, n64004, n64005, n64006, n64007, n64008, n64009,
    n64010, n64011, n64012, n64013, n64014, n64015, n64016, n64017, n64018,
    n64019, n64020, n64021, n64022, n64023, n64024, n64025, n64026, n64027,
    n64028, n64029, n64030, n64031, n64032, n64033, n64034, n64035, n64036,
    n64037, n64038, n64039, n64040, n64041, n64042, n64043, n64044, n64045,
    n64046, n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054,
    n64055, n64056, n64057, n64058, n64059, n64060, n64061, n64062, n64063,
    n64064, n64065, n64066, n64067, n64068, n64069, n64070, n64071, n64072,
    n64073, n64074, n64075, n64076, n64077, n64078, n64079, n64080, n64081,
    n64082, n64083, n64084, n64085, n64086, n64087, n64088, n64089, n64090,
    n64091, n64092, n64093, n64094, n64095, n64096, n64097, n64098, n64099,
    n64100, n64101, n64102, n64103, n64104, n64105, n64106, n64107, n64108,
    n64109, n64110, n64111, n64112, n64113, n64114, n64115, n64116, n64117,
    n64118, n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64126,
    n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134, n64135,
    n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143, n64144,
    n64145, n64146, n64147, n64148, n64149, n64150, n64151, n64152, n64153,
    n64154, n64155, n64156, n64157, n64158, n64159, n64160, n64161, n64162,
    n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170, n64171,
    n64172, n64173, n64174, n64175, n64176, n64177, n64178, n64179, n64180,
    n64181, n64182, n64183, n64184, n64185, n64186, n64187, n64188, n64189,
    n64190, n64191, n64192, n64193, n64194, n64195, n64196, n64197, n64198,
    n64199, n64200, n64201, n64202, n64203, n64204, n64205, n64206, n64207,
    n64208, n64209, n64210, n64211, n64212, n64213, n64214, n64215, n64216,
    n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224, n64225,
    n64226, n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234,
    n64235, n64236, n64237, n64238, n64239, n64240, n64241, n64242, n64243,
    n64244, n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252,
    n64253, n64254, n64255, n64256, n64257, n64258, n64259, n64260, n64261,
    n64262, n64263, n64264, n64265, n64266, n64267, n64268, n64269, n64270,
    n64271, n64272, n64273, n64274, n64275, n64276, n64277, n64278, n64279,
    n64280, n64281, n64282, n64283, n64284, n64285, n64286, n64287, n64288,
    n64289, n64290, n64291, n64292, n64293, n64294, n64295, n64296, n64297,
    n64298, n64299, n64300, n64301, n64302, n64303, n64304, n64305, n64306,
    n64307, n64308, n64309, n64310, n64311, n64312, n64313, n64314, n64315,
    n64316, n64317, n64318, n64319, n64320, n64321, n64322, n64323, n64324,
    n64325, n64326, n64327, n64328, n64329, n64330, n64331, n64332, n64333,
    n64334, n64335, n64336, n64337, n64338, n64339, n64340, n64341, n64342,
    n64343, n64344, n64345, n64346, n64347, n64348, n64349, n64350, n64351,
    n64352, n64353, n64354, n64355, n64356, n64357, n64358, n64359, n64360,
    n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368, n64369,
    n64370, n64371, n64372, n64373, n64374, n64375, n64376, n64377, n64378,
    n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386, n64387,
    n64388, n64389, n64390, n64391, n64392, n64393, n64394, n64395, n64396,
    n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404, n64405,
    n64406, n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414,
    n64415, n64416, n64417, n64418, n64419, n64420, n64421, n64422, n64423,
    n64424, n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432,
    n64433, n64434, n64435, n64436, n64437, n64438, n64439, n64440, n64441,
    n64442, n64443, n64444, n64445, n64446, n64447, n64448, n64449, n64450,
    n64451, n64452, n64453, n64454, n64455, n64456, n64457, n64458, n64459,
    n64460, n64461, n64462, n64463, n64464, n64465, n64466, n64467, n64468,
    n64469, n64470, n64471, n64472, n64473, n64474, n64475, n64476, n64477,
    n64478, n64479, n64480, n64481, n64482, n64483, n64484, n64485, n64486,
    n64487, n64488, n64489, n64490, n64491, n64492, n64493, n64494, n64495,
    n64496, n64497, n64498, n64499, n64500, n64501, n64502, n64503, n64504,
    n64505, n64506, n64507, n64508, n64509, n64510, n64511, n64512, n64513,
    n64514, n64515, n64516, n64517, n64518, n64519, n64520, n64521, n64522,
    n64523, n64524, n64525, n64526, n64527, n64528, n64529, n64530, n64531,
    n64532, n64533, n64534, n64535, n64536, n64537, n64538, n64539, n64540,
    n64541, n64542, n64543, n64544, n64545, n64546, n64547, n64548, n64549,
    n64550, n64551, n64552, n64553, n64554, n64555, n64556, n64557, n64558,
    n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566, n64567,
    n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64575, n64576,
    n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64584, n64585,
    n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593, n64594,
    n64595, n64596, n64597, n64598, n64599, n64600, n64601, n64602, n64603,
    n64604, n64605, n64606, n64607, n64608, n64609, n64610, n64611, n64612,
    n64613, n64614, n64615, n64616, n64617, n64618, n64619, n64620, n64621,
    n64622, n64623, n64624, n64625, n64626, n64627, n64628, n64629, n64630,
    n64631, n64632, n64633, n64634, n64635, n64636, n64637, n64638, n64639,
    n64640, n64641, n64642, n64643, n64644, n64645, n64646, n64647, n64648,
    n64649, n64650, n64651, n64652, n64653, n64654, n64655, n64656, n64657,
    n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665, n64666,
    n64667, n64668, n64669, n64670, n64671, n64672, n64673, n64674, n64675,
    n64676, n64677, n64678, n64679, n64680, n64681, n64682, n64683, n64684,
    n64685, n64686, n64687, n64688, n64689, n64690, n64691, n64692, n64693,
    n64694, n64695, n64696, n64697, n64698, n64699, n64700, n64701, n64702,
    n64703, n64704, n64705, n64706, n64707, n64708, n64709, n64710, n64711,
    n64712, n64713, n64714, n64715, n64716, n64717, n64718, n64719, n64720,
    n64721, n64722, n64723, n64724, n64725, n64726, n64727, n64728, n64729,
    n64730, n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738,
    n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746, n64747,
    n64748, n64749, n64750, n64751, n64752, n64753, n64754, n64755, n64756,
    n64757, n64758, n64759, n64760, n64761, n64762, n64763, n64764, n64765,
    n64766, n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774,
    n64775, n64776, n64777, n64778, n64779, n64780, n64781, n64782, n64783,
    n64784, n64785, n64786, n64787, n64788, n64789, n64790, n64791, n64792,
    n64793, n64794, n64795, n64796, n64797, n64798, n64799, n64800, n64801,
    n64802, n64803, n64804, n64805, n64806, n64807, n64808, n64809, n64810,
    n64811, n64812, n64813, n64814, n64815, n64816, n64817, n64818, n64819,
    n64820, n64821, n64822, n64823, n64824, n64825, n64826, n64827, n64828,
    n64829, n64830, n64831, n64832, n64833, n64834, n64835, n64836, n64837,
    n64838, n64839, n64840, n64841, n64842, n64843, n64844, n64845, n64846,
    n64847, n64848, n64849, n64850, n64851, n64852, n64853, n64854, n64855,
    n64856, n64857, n64858, n64859, n64860, n64861, n64862, n64863, n64864,
    n64865, n64866, n64867, n64868, n64869, n64870, n64871, n64872, n64873,
    n64874, n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882,
    n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890, n64891,
    n64892, n64893, n64894, n64895, n64896, n64897, n64898, n64899, n64900,
    n64901, n64902, n64903, n64904, n64905, n64906, n64907, n64908, n64909,
    n64910, n64911, n64912, n64913, n64914, n64915, n64916, n64917, n64918,
    n64919, n64920, n64921, n64922, n64923, n64924, n64925, n64926, n64927,
    n64928, n64929, n64930, n64931, n64932, n64933, n64934, n64935, n64936,
    n64937, n64938, n64939, n64940, n64941, n64942, n64943, n64944, n64945,
    n64946, n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954,
    n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962, n64963,
    n64964, n64965, n64966, n64967, n64968, n64969, n64970, n64971, n64972,
    n64973, n64974, n64975, n64976, n64977, n64978, n64979, n64980, n64981,
    n64982, n64983, n64984, n64985, n64986, n64987, n64988, n64989, n64990,
    n64991, n64992, n64993, n64994, n64995, n64996, n64997, n64998, n64999,
    n65000, n65001, n65002, n65003, n65004, n65005, n65006, n65007, n65008,
    n65009, n65010, n65011, n65012, n65013, n65014, n65015, n65016, n65017,
    n65018, n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026,
    n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034, n65035,
    n65036, n65037, n65038, n65039, n65040, n65041, n65042, n65043, n65044,
    n65045, n65046, n65047, n65048, n65049, n65050, n65051, n65052, n65053,
    n65054, n65055, n65056, n65057, n65058, n65059, n65060, n65061, n65062,
    n65063, n65064, n65065, n65066, n65067, n65068, n65069, n65070, n65071,
    n65072, n65073, n65074, n65075, n65076, n65077, n65078, n65079, n65080,
    n65081, n65082, n65083, n65084, n65085, n65086, n65087, n65088, n65089,
    n65090, n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098,
    n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106, n65107,
    n65108, n65109, n65110, n65111, n65112, n65113, n65114, n65115, n65116,
    n65117, n65118, n65119, n65120, n65121, n65122, n65123, n65124, n65125,
    n65126, n65127, n65128, n65129, n65130, n65131, n65132, n65133, n65134,
    n65135, n65136, n65137, n65138, n65139, n65140, n65141, n65142, n65143,
    n65144, n65145, n65146, n65147, n65148, n65149, n65150, n65151, n65152,
    n65153, n65154, n65155, n65156, n65157, n65158, n65159, n65160, n65161,
    n65162, n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170,
    n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178, n65179,
    n65180, n65181, n65182, n65183, n65184, n65185, n65186, n65187, n65188,
    n65189, n65190, n65191, n65192, n65193, n65194, n65195, n65196, n65197,
    n65198, n65199, n65200, n65201, n65202, n65203, n65204, n65205, n65206,
    n65207, n65208, n65209, n65210, n65211, n65212, n65213, n65214, n65215,
    n65216, n65217, n65218, n65219, n65220, n65221, n65222, n65223, n65224,
    n65225, n65226, n65227, n65228, n65229, n65230, n65231, n65232, n65233,
    n65234, n65235, n65236, n65237, n65238, n65239, n65240, n65241, n65242,
    n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250, n65251,
    n65252, n65253, n65254, n65255, n65256, n65257, n65258, n65259, n65260,
    n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268, n65269,
    n65270, n65271, n65272, n65273, n65274, n65275, n65276, n65277, n65278,
    n65279, n65280, n65281, n65282, n65283, n65284, n65285, n65286, n65287,
    n65288, n65289, n65290, n65291, n65292, n65293, n65294, n65295, n65296,
    n65297, n65298, n65299, n65300, n65301, n65302, n65303, n65304, n65305,
    n65306, n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314,
    n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322, n65323,
    n65324, n65325, n65326, n65327, n65328, n65329, n65330, n65331, n65332,
    n65333, n65334, n65335, n65336, n65337, n65338, n65339, n65340, n65341,
    n65342, n65343, n65344, n65345, n65346, n65347, n65348, n65349, n65350,
    n65351, n65352, n65353, n65354, n65355, n65356, n65357, n65358, n65359,
    n65360, n65361, n65362, n65363, n65364, n65365, n65366, n65367, n65368,
    n65369, n65370, n65371, n65372, n65373, n65374, n65375, n65376, n65377,
    n65378, n65379, n65380, n65381, n65382, n65383, n65384, n65385, n65386,
    n65387, n65388, n65389, n65390, n65391, n65392, n65393, n65394, n65395,
    n65396, n65397, n65398, n65399, n65400, n65401, n65402, n65403, n65404,
    n65405, n65406, n65407, n65408, n65409, n65410, n65411, n65412, n65413,
    n65414, n65415, n65416, n65417, n65418, n65419, n65420, n65421, n65422,
    n65423, n65424, n65425, n65426, n65427, n65428, n65429, n65430, n65431,
    n65432, n65433, n65434, n65435, n65436, n65437, n65438, n65439, n65440,
    n65441, n65442, n65443, n65444, n65445, n65446, n65447, n65448, n65449,
    n65450, n65451, n65452, n65453, n65454, n65455, n65456, n65457, n65458,
    n65459, n65460, n65461, n65462, n65463, n65464, n65465, n65466, n65467,
    n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475, n65476,
    n65477, n65478, n65479, n65480, n65481, n65482, n65483, n65484, n65485,
    n65486, n65487, n65488, n65489, n65490, n65491, n65492, n65493, n65494,
    n65495, n65496, n65497, n65498, n65499, n65500, n65501, n65502, n65503,
    n65504, n65505, n65506, n65507, n65508, n65509, n65510, n65511, n65512,
    n65513, n65514, n65515, n65516, n65517, n65518, n65519, n65520, n65521,
    n65522, n65523, n65524, n65525, n65526, n65527, n65528, n65529, n65530,
    n65531, n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539,
    n65540, n65541, n65542, n65543, n65544, n65545, n65546, n65547, n65548,
    n65549, n65550, n65551, n65552, n65553, n65554, n65555, n65556, n65557,
    n65558, n65559, n65560, n65561, n65562, n65563, n65564, n65565, n65566,
    n65567, n65568, n65569, n65570, n65571, n65572, n65573, n65574, n65575,
    n65576, n65577, n65578, n65579, n65580, n65581, n65582, n65583, n65584,
    n65585, n65586, n65587, n65588, n65589, n65590, n65591, n65592, n65593,
    n65594, n65595, n65596, n65597, n65598, n65599, n65600, n65601, n65602,
    n65603, n65604, n65605, n65606, n65607, n65608, n65609, n65610, n65611,
    n65612, n65613, n65614, n65615, n65616, n65617, n65618, n65619, n65620,
    n65621, n65622, n65623, n65624, n65625, n65626, n65627, n65628, n65629,
    n65630, n65631, n65632, n65633, n65634, n65635, n65636, n65637, n65638,
    n65639, n65640, n65641, n65642, n65643, n65644, n65645, n65646, n65647,
    n65648, n65649, n65650, n65651, n65652, n65653, n65654, n65655, n65656,
    n65657, n65658, n65659, n65660, n65661, n65662, n65663, n65664, n65665,
    n65666, n65667, n65668, n65669, n65670, n65671, n65672, n65673, n65674,
    n65675, n65676, n65677, n65678, n65679, n65680, n65681, n65682, n65683,
    n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691, n65692,
    n65693, n65694, n65695, n65696, n65697, n65698, n65699, n65700, n65701,
    n65702, n65703, n65704, n65705, n65706, n65707, n65708, n65709, n65710,
    n65711, n65712, n65713, n65714, n65715, n65716, n65717, n65718, n65719,
    n65720, n65721, n65722, n65723, n65724, n65725, n65726, n65727, n65728,
    n65729, n65730, n65731, n65732, n65733, n65734, n65735, n65736, n65737,
    n65738, n65739, n65740, n65741, n65742, n65743, n65744, n65745, n65746,
    n65747, n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755,
    n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763, n65764,
    n65765, n65766, n65767, n65768, n65769, n65770, n65771, n65772, n65773,
    n65774, n65775, n65776, n65777, n65778, n65779, n65780, n65781, n65782,
    n65783, n65784, n65785, n65786, n65787, n65788, n65789, n65790, n65791,
    n65792, n65793, n65794, n65795, n65796, n65797, n65798, n65799, n65800,
    n65801, n65802, n65803, n65804, n65805, n65806, n65807, n65808, n65809,
    n65810, n65811, n65812, n65813, n65814, n65815, n65816, n65817, n65818,
    n65819, n65820, n65821, n65822, n65823, n65824, n65825, n65826, n65827,
    n65828, n65829, n65830, n65831, n65832, n65833, n65834, n65835, n65836,
    n65837, n65838, n65839, n65840, n65841, n65842, n65843, n65844, n65845,
    n65846, n65847, n65848, n65849, n65850, n65851, n65852, n65853, n65854,
    n65855, n65856, n65857, n65858, n65859, n65860, n65861, n65862, n65863,
    n65864, n65865, n65866, n65867, n65868, n65869, n65870, n65871, n65872,
    n65873, n65874, n65875, n65876, n65877, n65878, n65879, n65880, n65881,
    n65882, n65883, n65884, n65885, n65886, n65887, n65888, n65889, n65890,
    n65891, n65892, n65893, n65894, n65895, n65896, n65897, n65898, n65899,
    n65900, n65901, n65902, n65903, n65904, n65905, n65906, n65907, n65908,
    n65909, n65910, n65911, n65912, n65913, n65914, n65915, n65916, n65917,
    n65918, n65919, n65920, n65921, n65922, n65923, n65924, n65925, n65926,
    n65927, n65928, n65929, n65930, n65931, n65932, n65933, n65934, n65935,
    n65936, n65937, n65938, n65939, n65940, n65941, n65942, n65943, n65944,
    n65945, n65946, n65947, n65948, n65949, n65950, n65951, n65952, n65953,
    n65954, n65955, n65956, n65957, n65958, n65959, n65960, n65961, n65962,
    n65963, n65964, n65965, n65966, n65967, n65968, n65969, n65970, n65971,
    n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979, n65980,
    n65981, n65982, n65983, n65984, n65985, n65986, n65987, n65988, n65989,
    n65990, n65991, n65992, n65993, n65994, n65995, n65996, n65997, n65998,
    n65999, n66000, n66001, n66002, n66003, n66004, n66005, n66006, n66007,
    n66008, n66009, n66010, n66011, n66012, n66013, n66014, n66015, n66016,
    n66017, n66018, n66019, n66020, n66021, n66022, n66023, n66024, n66025,
    n66026, n66027, n66028, n66029, n66030, n66031, n66032, n66033, n66034,
    n66035, n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043,
    n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051, n66052,
    n66053, n66054, n66055, n66056, n66057, n66058, n66059, n66060, n66061,
    n66062, n66063, n66064, n66065, n66066, n66067, n66068, n66069, n66070,
    n66071, n66072, n66073, n66074, n66075, n66076, n66077, n66078, n66079,
    n66080, n66081, n66082, n66083, n66084, n66085, n66086, n66087, n66088,
    n66089, n66090, n66091, n66092, n66093, n66094, n66095, n66096, n66097,
    n66098, n66099, n66100, n66101, n66102, n66103, n66104, n66105, n66106,
    n66107, n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115,
    n66116, n66117, n66118, n66119, n66120, n66121, n66122, n66123, n66124,
    n66125, n66126, n66127, n66128, n66129, n66130, n66131, n66132, n66133,
    n66134, n66135, n66136, n66137, n66138, n66139, n66140, n66141, n66142,
    n66143, n66144, n66145, n66146, n66147, n66148, n66149, n66150, n66151,
    n66152, n66153, n66154, n66155, n66156, n66157, n66158, n66159, n66160,
    n66161, n66162, n66163, n66164, n66165, n66166, n66167, n66168, n66169,
    n66170, n66171, n66172, n66173, n66174, n66175, n66176, n66177, n66178,
    n66179, n66180, n66181, n66182, n66183, n66184, n66185, n66186, n66187,
    n66188, n66189, n66190, n66191, n66192, n66193, n66194, n66195, n66196,
    n66197, n66198, n66199, n66200, n66201, n66202, n66203, n66204, n66205,
    n66206, n66207, n66208, n66209, n66210, n66211, n66212, n66213, n66214,
    n66215, n66216, n66217, n66218, n66219, n66220, n66221, n66222, n66223,
    n66224, n66225, n66226, n66227, n66228, n66229, n66230, n66231, n66232,
    n66233, n66234, n66235, n66236, n66237, n66238, n66239, n66240, n66241,
    n66242, n66243, n66244, n66245, n66246, n66247, n66248, n66249, n66250,
    n66251, n66252, n66253, n66254, n66255, n66256, n66257, n66258, n66259,
    n66260, n66261, n66262, n66263, n66264, n66265, n66266, n66267, n66268,
    n66269, n66270, n66271, n66272, n66273, n66274, n66275, n66276, n66277,
    n66278, n66279, n66280, n66281, n66282, n66283, n66284, n66285, n66286,
    n66287, n66288, n66289, n66290, n66291, n66292, n66293, n66294, n66295,
    n66296, n66297, n66298, n66299, n66300, n66301, n66302, n66303, n66304,
    n66305, n66306, n66307, n66308, n66309, n66310, n66311, n66312, n66313,
    n66314, n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66322,
    n66323, n66324, n66325, n66326, n66327, n66328, n66329, n66330, n66331,
    n66332, n66333, n66334, n66335, n66336, n66337, n66338, n66339, n66340,
    n66341, n66342, n66343, n66344, n66345, n66346, n66347, n66348, n66349,
    n66350, n66351, n66352, n66353, n66354, n66355, n66356, n66357, n66358,
    n66359, n66360, n66361, n66362, n66363, n66364, n66365, n66366, n66367,
    n66368, n66369, n66370, n66371, n66372, n66373, n66374, n66375, n66376,
    n66377, n66378, n66379, n66380, n66381, n66382, n66383, n66384, n66385,
    n66386, n66387, n66388, n66389, n66390, n66391, n66392, n66393, n66394,
    n66395, n66396, n66397, n66398, n66399, n66400, n66401, n66402, n66403,
    n66404, n66405, n66406, n66407, n66408, n66409, n66410, n66411, n66412,
    n66413, n66414, n66415, n66416, n66417, n66418, n66419, n66420, n66421,
    n66422, n66423, n66424, n66425, n66426, n66427, n66428, n66429, n66430,
    n66431, n66432, n66433, n66434, n66435, n66436, n66437, n66438, n66439,
    n66440, n66441, n66442, n66443, n66444, n66445, n66446, n66447, n66448,
    n66449, n66450, n66451, n66452, n66453, n66454, n66455, n66456, n66457,
    n66458, n66459, n66460, n66461, n66462, n66463, n66464, n66465, n66466,
    n66467, n66468, n66469, n66470, n66471, n66472, n66473, n66474, n66475,
    n66476, n66477, n66478, n66479, n66480, n66481, n66482, n66483, n66484,
    n66485, n66486, n66487, n66488, n66489, n66490, n66491, n66492, n66493,
    n66494, n66495, n66496, n66497, n66498, n66499, n66500, n66501, n66502,
    n66503, n66504, n66505, n66506, n66507, n66508, n66509, n66510, n66511,
    n66512, n66513, n66514, n66515, n66516, n66517, n66518, n66519, n66520,
    n66521, n66522, n66523, n66524, n66525, n66526, n66527, n66528, n66529,
    n66530, n66531, n66532, n66533, n66534, n66535, n66536, n66537, n66538,
    n66539, n66540, n66541, n66542, n66543, n66544, n66545, n66546, n66547,
    n66548, n66549, n66550, n66551, n66552, n66553, n66554, n66555, n66556,
    n66557, n66558, n66559, n66560, n66561, n66562, n66563, n66564, n66565,
    n66566, n66567, n66568, n66569, n66570, n66571, n66572, n66573, n66574,
    n66575, n66576, n66577, n66578, n66579, n66580, n66581, n66582, n66583,
    n66584, n66585, n66586, n66587, n66588, n66589, n66590, n66591, n66592,
    n66593, n66594, n66595, n66596, n66597, n66598, n66599, n66600, n66601,
    n66602, n66603, n66604, n66605, n66606, n66607, n66608, n66609, n66610,
    n66611, n66612, n66613, n66614, n66615, n66616, n66617, n66618, n66619,
    n66620, n66621, n66622, n66623, n66624, n66625, n66626, n66627, n66628,
    n66629, n66630, n66631, n66632, n66633, n66634, n66635, n66636, n66637,
    n66638, n66639, n66640, n66641, n66642, n66643, n66644, n66645, n66646,
    n66647, n66648, n66649, n66650, n66651, n66652, n66653, n66654, n66655,
    n66656, n66657, n66658, n66659, n66660, n66661, n66662, n66663, n66664,
    n66665, n66666, n66667, n66668, n66669, n66670, n66671, n66672, n66673,
    n66674, n66675, n66676, n66677, n66678, n66679, n66680, n66681, n66682,
    n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690, n66691,
    n66692, n66693, n66694, n66695, n66696, n66697, n66698, n66699, n66700,
    n66701, n66702, n66703, n66704, n66705, n66706, n66707, n66708, n66709,
    n66710, n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718,
    n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726, n66727,
    n66728, n66729, n66730, n66731, n66732, n66733, n66734, n66735, n66736,
    n66737, n66738, n66739, n66740, n66741, n66742, n66743, n66744, n66745,
    n66746, n66747, n66748, n66749, n66750, n66751, n66752, n66753, n66754,
    n66755, n66756, n66757, n66758, n66759, n66760, n66761, n66762, n66763,
    n66764, n66765, n66766, n66767, n66768, n66769, n66770, n66771, n66772,
    n66773, n66774, n66775, n66776, n66777, n66778, n66779, n66780, n66781,
    n66782, n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790,
    n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798, n66799,
    n66800, n66801, n66802, n66803, n66804, n66805, n66806, n66807, n66808,
    n66809, n66810, n66811, n66812, n66813, n66814, n66815, n66816, n66817,
    n66818, n66819, n66820, n66821, n66822, n66823, n66824, n66825, n66826,
    n66827, n66828, n66829, n66830, n66831, n66832, n66833, n66834, n66835,
    n66836, n66837, n66838, n66839, n66840, n66841, n66842, n66843, n66844,
    n66845, n66846, n66847, n66848, n66849, n66850, n66851, n66852, n66853,
    n66854, n66855, n66856, n66857, n66858, n66859, n66860, n66861, n66862,
    n66863, n66864, n66865, n66866, n66867, n66868, n66869, n66870, n66871,
    n66872, n66873, n66874, n66875, n66876, n66877, n66878, n66879, n66880,
    n66881, n66882, n66883, n66884, n66885, n66886, n66887, n66888, n66889,
    n66890, n66891, n66892, n66893, n66894, n66895, n66896, n66897, n66898,
    n66899, n66900, n66901, n66902, n66903, n66904, n66905, n66906, n66907,
    n66908, n66909, n66910, n66911, n66912, n66913, n66914, n66915, n66916,
    n66917, n66918, n66919, n66920, n66921, n66922, n66923, n66924, n66925,
    n66926, n66927, n66928, n66929, n66930, n66931, n66932, n66933, n66934,
    n66935, n66936, n66937, n66938, n66939, n66940, n66941, n66942, n66943,
    n66944, n66945, n66946, n66947, n66948, n66949, n66950, n66951, n66952,
    n66953, n66954, n66955, n66956, n66957, n66958, n66959, n66960, n66961,
    n66962, n66963, n66964, n66965, n66966, n66967, n66968, n66969, n66970,
    n66971, n66972, n66973, n66974, n66975, n66976, n66977, n66978, n66979,
    n66980, n66981, n66982, n66983, n66984, n66985, n66986, n66987, n66988,
    n66989, n66990, n66991, n66992, n66993, n66994, n66995, n66996, n66997,
    n66998, n66999, n67000, n67001, n67002, n67003, n67004, n67005, n67006,
    n67007, n67008, n67009, n67010, n67011, n67012, n67013, n67014, n67015,
    n67016, n67017, n67018, n67019, n67020, n67021, n67022, n67023, n67024,
    n67025, n67026, n67027, n67028, n67029, n67030, n67031, n67032, n67033,
    n67034, n67035, n67036, n67037, n67038, n67039, n67040, n67041, n67042,
    n67043, n67044, n67045, n67046, n67047, n67048, n67049, n67050, n67051,
    n67052, n67053, n67054, n67055, n67056, n67057, n67058, n67059, n67060,
    n67061, n67062, n67063, n67064, n67065, n67066, n67067, n67068, n67069,
    n67070, n67071, n67072, n67073, n67074, n67075, n67076, n67077, n67078,
    n67079, n67080, n67081, n67082, n67083, n67084, n67085, n67086, n67087,
    n67088, n67089, n67090, n67091, n67092, n67093, n67094, n67095, n67096,
    n67097, n67098, n67099, n67100, n67101, n67102, n67103, n67104, n67105,
    n67106, n67107, n67108, n67109, n67110, n67111, n67112, n67113, n67114,
    n67115, n67116, n67117, n67118, n67119, n67120, n67121, n67122, n67123,
    n67124, n67125, n67126, n67127, n67128, n67129, n67130, n67131, n67132,
    n67133, n67134, n67135, n67136, n67137, n67138, n67139, n67140, n67141,
    n67142, n67143, n67144, n67145, n67146, n67147, n67148, n67149, n67150,
    n67151, n67152, n67153, n67154, n67155, n67156, n67157, n67158, n67159,
    n67160, n67161, n67162, n67163, n67164, n67165, n67166, n67167, n67168,
    n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176, n67177,
    n67178, n67179, n67180, n67181, n67182, n67183, n67184, n67185, n67186,
    n67187, n67188, n67189, n67190, n67191, n67192, n67193, n67194, n67195,
    n67196, n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204,
    n67205, n67206, n67207, n67208, n67209, n67210, n67211, n67212, n67213,
    n67214, n67215, n67216, n67217, n67218, n67219, n67220, n67221, n67222,
    n67223, n67224, n67225, n67226, n67227, n67228, n67229, n67230, n67231,
    n67232, n67233, n67234, n67235, n67236, n67237, n67238, n67239, n67240,
    n67241, n67242, n67243, n67244, n67245, n67246, n67247, n67248, n67249,
    n67250, n67251, n67252, n67253, n67254, n67255, n67256, n67257, n67258,
    n67259, n67260, n67261, n67262, n67263, n67264, n67265, n67266, n67267,
    n67268, n67269, n67270, n67271, n67272, n67273, n67274, n67275, n67276,
    n67277, n67278, n67279, n67280, n67281, n67282, n67283, n67284, n67285,
    n67286, n67287, n67288, n67289, n67290, n67291, n67292, n67293, n67294,
    n67295, n67296, n67297, n67298, n67299, n67300, n67301, n67302, n67303,
    n67304, n67305, n67306, n67307, n67308, n67309, n67310, n67311, n67312,
    n67313, n67314, n67315, n67316, n67317, n67318, n67319, n67320, n67321,
    n67322, n67323, n67324, n67325, n67326, n67327, n67328, n67329, n67330,
    n67331, n67332, n67333, n67334, n67335, n67336, n67337, n67338, n67339,
    n67340, n67341, n67342, n67343, n67344, n67345, n67346, n67347, n67348,
    n67349, n67350, n67351, n67352, n67353, n67354, n67355, n67356, n67357,
    n67358, n67359, n67360, n67361, n67362, n67363, n67364, n67365, n67366,
    n67367, n67368, n67369, n67370, n67371, n67372, n67373, n67374, n67375,
    n67376, n67377, n67378, n67379, n67380, n67381, n67382, n67383, n67384,
    n67385, n67386, n67387, n67388, n67389, n67390, n67391, n67392, n67393,
    n67394, n67395, n67396, n67397, n67398, n67399, n67400, n67401, n67402,
    n67403, n67404, n67405, n67406, n67407, n67408, n67409, n67410, n67411,
    n67412, n67413, n67414, n67415, n67416, n67417, n67418, n67419, n67420,
    n67421, n67422, n67423, n67424, n67425, n67426, n67427, n67428, n67429,
    n67430, n67431, n67432, n67433, n67434, n67435, n67436, n67437, n67438,
    n67439, n67440, n67441, n67442, n67443, n67444, n67445, n67446, n67447,
    n67448, n67449, n67450, n67451, n67452, n67453, n67454, n67455, n67456,
    n67457, n67458, n67459, n67460, n67461, n67462, n67463, n67464, n67465,
    n67466, n67467, n67468, n67469, n67470, n67471, n67472, n67473, n67474,
    n67475, n67476, n67477, n67478, n67479, n67480, n67481, n67482, n67483,
    n67484, n67485, n67486, n67487, n67488, n67489, n67490, n67491, n67492,
    n67493, n67494, n67495, n67496, n67497, n67498, n67499, n67500, n67501,
    n67502, n67503, n67504, n67505, n67506, n67507, n67508, n67509, n67510,
    n67511, n67512, n67513, n67514, n67515, n67516, n67517, n67518, n67519,
    n67520, n67521, n67522, n67523, n67524, n67525, n67526, n67527, n67528,
    n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536, n67537,
    n67538, n67539, n67540, n67541, n67542, n67543, n67544, n67545, n67546,
    n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554, n67555,
    n67556, n67557, n67558, n67559, n67560, n67561, n67562, n67563, n67564,
    n67565, n67566, n67567, n67568, n67569, n67570, n67571, n67572, n67573,
    n67574, n67575, n67576, n67577, n67578, n67579, n67580, n67581, n67582,
    n67583, n67584, n67585, n67586, n67587, n67588, n67589, n67590, n67591,
    n67592, n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600,
    n67601, n67602, n67603, n67604, n67605, n67606, n67607, n67608, n67609,
    n67610, n67611, n67612, n67613, n67614, n67615, n67616, n67617, n67618,
    n67619, n67620, n67621, n67622, n67623, n67624, n67625, n67626, n67627,
    n67628, n67629, n67630, n67631, n67632, n67633, n67634, n67635, n67636,
    n67637, n67638, n67639, n67640, n67641, n67642, n67643, n67644, n67645,
    n67646, n67647, n67648, n67649, n67650, n67651, n67652, n67653, n67654,
    n67655, n67656, n67657, n67658, n67659, n67660, n67661, n67662, n67663,
    n67664, n67665, n67666, n67667, n67668, n67669, n67670, n67671, n67672,
    n67673, n67674, n67675, n67676, n67677, n67678, n67679, n67680, n67681,
    n67682, n67683, n67684, n67685, n67686, n67687, n67688, n67689, n67690,
    n67691, n67692, n67693, n67694, n67695, n67696, n67697, n67698, n67699,
    n67700, n67701, n67702, n67703, n67704, n67705, n67706, n67707, n67708,
    n67709, n67710, n67711, n67712, n67713, n67714, n67715, n67716, n67717,
    n67718, n67719, n67720, n67721, n67722, n67723, n67724, n67725, n67726,
    n67727, n67728, n67729, n67730, n67731, n67732, n67733, n67734, n67735,
    n67736, n67737, n67738, n67739, n67740, n67741, n67742, n67743, n67744,
    n67745, n67746, n67747, n67748, n67749, n67750, n67751, n67752, n67753,
    n67754, n67755, n67756, n67757, n67758, n67759, n67760, n67761, n67762,
    n67763, n67764, n67765, n67766, n67767, n67768, n67769, n67770, n67771,
    n67772, n67773, n67774, n67775, n67776, n67777, n67778, n67779, n67780,
    n67781, n67782, n67783, n67784, n67785, n67786, n67787, n67788, n67789,
    n67790, n67791, n67792, n67793, n67794, n67795, n67796, n67797, n67798,
    n67799, n67800, n67801, n67802, n67803, n67804, n67805, n67806, n67807,
    n67808, n67809, n67810, n67811, n67812, n67813, n67814, n67815, n67816,
    n67817, n67818, n67819, n67820, n67821, n67822, n67823, n67824, n67825,
    n67826, n67827, n67828, n67829, n67830, n67831, n67832, n67833, n67834,
    n67835, n67836, n67837, n67838, n67839, n67840, n67841, n67842, n67843,
    n67844, n67845, n67846, n67847, n67848, n67849, n67850, n67851, n67852,
    n67853, n67854, n67855, n67856, n67857, n67858, n67859, n67860, n67861,
    n67862, n67863, n67864, n67865, n67866, n67867, n67868, n67869, n67870,
    n67871, n67872, n67873, n67874, n67875, n67876, n67877, n67878, n67879,
    n67880, n67881, n67882, n67883, n67884, n67885, n67886, n67887, n67888,
    n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896, n67897,
    n67898, n67899, n67900, n67901, n67902, n67903, n67904, n67905, n67906,
    n67907, n67908, n67909, n67910, n67911, n67912, n67913, n67914, n67915,
    n67916, n67917, n67918, n67919, n67920, n67921, n67922, n67923, n67924,
    n67925, n67926, n67927, n67928, n67929, n67930, n67931, n67932, n67933,
    n67934, n67935, n67936, n67937, n67938, n67939, n67940, n67941, n67942,
    n67943, n67944, n67945, n67946, n67947, n67948, n67949, n67950, n67951,
    n67952, n67953, n67954, n67955, n67956, n67957, n67958, n67959, n67960,
    n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968, n67969,
    n67970, n67971, n67972, n67973, n67974, n67975, n67976, n67977, n67978,
    n67979, n67980, n67981, n67982, n67983, n67984, n67985, n67986, n67987,
    n67988, n67989, n67990, n67991, n67992, n67993, n67994, n67995, n67996,
    n67997, n67998, n67999, n68000, n68001, n68002, n68003, n68004, n68005,
    n68006, n68007, n68008, n68009, n68010, n68011, n68012, n68013, n68014,
    n68015, n68016, n68017, n68018, n68019, n68020, n68021, n68022, n68023,
    n68024, n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032,
    n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040, n68041,
    n68042, n68043, n68044, n68045, n68046, n68047, n68048, n68049, n68050,
    n68051, n68052, n68053, n68054, n68055, n68056, n68057, n68058, n68059,
    n68060, n68061, n68062, n68063, n68064, n68065, n68066, n68067, n68068,
    n68069, n68070, n68071, n68072, n68073, n68074, n68075, n68076, n68077,
    n68078, n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086,
    n68087, n68088, n68089, n68090, n68091, n68092, n68093, n68094, n68095,
    n68096, n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104,
    n68105, n68106, n68107, n68108, n68109, n68110, n68111, n68112, n68113,
    n68114, n68115, n68116, n68117, n68118, n68119, n68120, n68121, n68122,
    n68123, n68124, n68125, n68126, n68127, n68128, n68129, n68130, n68131,
    n68132, n68133, n68134, n68135, n68136, n68137, n68138, n68139, n68140,
    n68141, n68142, n68143, n68144, n68145, n68146, n68147, n68148, n68149,
    n68150, n68151, n68152, n68153, n68154, n68155, n68156, n68157, n68158,
    n68159, n68160, n68161, n68162, n68163, n68164, n68165, n68166, n68167,
    n68168, n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176,
    n68177, n68178, n68179, n68180, n68181, n68182, n68183, n68184, n68185,
    n68186, n68187, n68188, n68189, n68190, n68191, n68192, n68193, n68194,
    n68195, n68196, n68197, n68198, n68199, n68200, n68201, n68202, n68203,
    n68204, n68205, n68206, n68207, n68208, n68209, n68210, n68211, n68212,
    n68213, n68214, n68215, n68216, n68217, n68218, n68219, n68220, n68221,
    n68222, n68223, n68224, n68225, n68226, n68227, n68228, n68229, n68230,
    n68231, n68232, n68233, n68234, n68235, n68236, n68237, n68238, n68239,
    n68240, n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248,
    n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256, n68257,
    n68258, n68259, n68260, n68261, n68262, n68263, n68264, n68265, n68266,
    n68267, n68268, n68269, n68270, n68271, n68272, n68273, n68274, n68275,
    n68276, n68277, n68278, n68279, n68280, n68281, n68282, n68283, n68284,
    n68285, n68286, n68287, n68288, n68289, n68290, n68291, n68292, n68293,
    n68294, n68295, n68296, n68297, n68298, n68299, n68300, n68301, n68302,
    n68303, n68304, n68305, n68306, n68307, n68308, n68309, n68310, n68311,
    n68312, n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320,
    n68321, n68322, n68323, n68324, n68325, n68326, n68327, n68328, n68329,
    n68330, n68331, n68332, n68333, n68334, n68335, n68336, n68337, n68338,
    n68339, n68340, n68341, n68342, n68343, n68344, n68345, n68346, n68347,
    n68348, n68349, n68350, n68351, n68352, n68353, n68354, n68355, n68356,
    n68357, n68358, n68359, n68360, n68361, n68362, n68363, n68364, n68365,
    n68366, n68367, n68368, n68369, n68370, n68371, n68372, n68373, n68374,
    n68375, n68376, n68377, n68378, n68379, n68380, n68381, n68382, n68383,
    n68384, n68385, n68386, n68387, n68388, n68389, n68390, n68391, n68392,
    n68393, n68394, n68395, n68396, n68397, n68398, n68399, n68400, n68401,
    n68402, n68403, n68404, n68405, n68406, n68407, n68408, n68409, n68410,
    n68411, n68412, n68413, n68414, n68415, n68416, n68417, n68418, n68419,
    n68420, n68421, n68422, n68423, n68424, n68425, n68426, n68427, n68428,
    n68429, n68430, n68431, n68432, n68433, n68434, n68435, n68436, n68437,
    n68438, n68439, n68440, n68441, n68442, n68443, n68444, n68445, n68446,
    n68447, n68448, n68449, n68450, n68451, n68452, n68453, n68454, n68455,
    n68456, n68457, n68458, n68459, n68460, n68461, n68462, n68463, n68464,
    n68465, n68466, n68467, n68468, n68469, n68470, n68471, n68472, n68473,
    n68474, n68475, n68476, n68477, n68478, n68479, n68480, n68481, n68482,
    n68483, n68484, n68485, n68486, n68487, n68488, n68489, n68490, n68491,
    n68492, n68493, n68494, n68495, n68496, n68497, n68498, n68499, n68500,
    n68501, n68502, n68503, n68504, n68505, n68506, n68507, n68508, n68509,
    n68510, n68511, n68512, n68513, n68514, n68515, n68516, n68517, n68518,
    n68519, n68520, n68521, n68522, n68523, n68524, n68525, n68526, n68527,
    n68528, n68529, n68530, n68531, n68532, n68533, n68534, n68535, n68536,
    n68537, n68538, n68539, n68540, n68541, n68542, n68543, n68544, n68545,
    n68546, n68547, n68548, n68549, n68550, n68551, n68552, n68553, n68554,
    n68555, n68556, n68557, n68558, n68559, n68560, n68561, n68562, n68563,
    n68564, n68565, n68566, n68567, n68568, n68569, n68570, n68571, n68572,
    n68573, n68574, n68575, n68576, n68577, n68578, n68579, n68580, n68581,
    n68582, n68583, n68584, n68585, n68586, n68587, n68588, n68589, n68590,
    n68591, n68592, n68593, n68594, n68595, n68596, n68597, n68598, n68599,
    n68600, n68601, n68602, n68603, n68604, n68605, n68606, n68607, n68608,
    n68609, n68610, n68611, n68612, n68613, n68614, n68615, n68616, n68617,
    n68618, n68619, n68620, n68621, n68622, n68623, n68624, n68625, n68626,
    n68627, n68628, n68629, n68630, n68631, n68632, n68633, n68634, n68635,
    n68636, n68637, n68638, n68639, n68640, n68641, n68642, n68643, n68644,
    n68645, n68646, n68647, n68648, n68649, n68650, n68651, n68652, n68653,
    n68654, n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662,
    n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671,
    n68672, n68673, n68674, n68675, n68676, n68677, n68678, n68679, n68680,
    n68681, n68682, n68683, n68684, n68685, n68686, n68687, n68688, n68689,
    n68690, n68691, n68692, n68693, n68694, n68695, n68696, n68697, n68698,
    n68699, n68700, n68701, n68702, n68703, n68704, n68705, n68706, n68707,
    n68708, n68709, n68710, n68711, n68712, n68713, n68714, n68715, n68716,
    n68717, n68718, n68719, n68720, n68721, n68722, n68723, n68724, n68725,
    n68726, n68727, n68728, n68729, n68730, n68731, n68732, n68733, n68734,
    n68735, n68736, n68737, n68738, n68739, n68740, n68741, n68742, n68743,
    n68744, n68745, n68746, n68747, n68748, n68749, n68750, n68751, n68752,
    n68753, n68754, n68755, n68756, n68757, n68758, n68759, n68760, n68761,
    n68762, n68763, n68764, n68765, n68766, n68767, n68768, n68769, n68770,
    n68771, n68772, n68773, n68774, n68775, n68776, n68777, n68778, n68779,
    n68780, n68781, n68782, n68783, n68784, n68785, n68786, n68787, n68788,
    n68789, n68790, n68791, n68792, n68793, n68794, n68795, n68796, n68797,
    n68798, n68799, n68800, n68801, n68802, n68803, n68804, n68805, n68806,
    n68807, n68808, n68809, n68810, n68811, n68812, n68813, n68814, n68815,
    n68816, n68817, n68818, n68819, n68820, n68821, n68822, n68823, n68824,
    n68825, n68826, n68827, n68828, n68829, n68830, n68831, n68832, n68833,
    n68834, n68835, n68836, n68837, n68838, n68839, n68840, n68841, n68842,
    n68843, n68844, n68845, n68846, n68847, n68848, n68849, n68850, n68851,
    n68852, n68853, n68854, n68855, n68856, n68857, n68858, n68859, n68860,
    n68861, n68862, n68863, n68864, n68865, n68866, n68867, n68868, n68869,
    n68870, n68871, n68872, n68873, n68874, n68875, n68876, n68877, n68878,
    n68879, n68880, n68881, n68882, n68883, n68884, n68885, n68886, n68887,
    n68888, n68889, n68890, n68891, n68892, n68893, n68894, n68895, n68896,
    n68897, n68898, n68899, n68900, n68901, n68902, n68903, n68904, n68905,
    n68906, n68907, n68908, n68909, n68910, n68911, n68912, n68913, n68914,
    n68915, n68916, n68917, n68918, n68919, n68920, n68921, n68922, n68923,
    n68924, n68925, n68926, n68927, n68928, n68929, n68930, n68931, n68932,
    n68933, n68934, n68935, n68936, n68937, n68938, n68939, n68940, n68941,
    n68942, n68943, n68944, n68945, n68946, n68947, n68948, n68949, n68950,
    n68951, n68952, n68953, n68954, n68955, n68956, n68957, n68958, n68959,
    n68960, n68961, n68962, n68963, n68964, n68965, n68966, n68967, n68968,
    n68969, n68970, n68971, n68972, n68973, n68974, n68975, n68976, n68977,
    n68978, n68979, n68980, n68981, n68982, n68983, n68984, n68985, n68986,
    n68987, n68988, n68989, n68990, n68991, n68992, n68993, n68994, n68995,
    n68996, n68997, n68998, n68999, n69000, n69001, n69002, n69003, n69004,
    n69005, n69006, n69007, n69008, n69009, n69010, n69011, n69012, n69013,
    n69014, n69015, n69016, n69017, n69018, n69019, n69020, n69021, n69022,
    n69023, n69024, n69025, n69026, n69027, n69028, n69029, n69030, n69031,
    n69032, n69033, n69034, n69035, n69036, n69037, n69038, n69039, n69040,
    n69041, n69042, n69043, n69044, n69045, n69046, n69047, n69048, n69049,
    n69050, n69051, n69052, n69053, n69054, n69055, n69056, n69057, n69058,
    n69059, n69060, n69061, n69062, n69063, n69064, n69065, n69066, n69067,
    n69068, n69069, n69070, n69071, n69072, n69073, n69074, n69075, n69076,
    n69077, n69078, n69079, n69080, n69081, n69082, n69083, n69084, n69085,
    n69086, n69087, n69088, n69089, n69090, n69091, n69092, n69093, n69094,
    n69095, n69096, n69097, n69098, n69099, n69100, n69101, n69102, n69103,
    n69104, n69105, n69106, n69107, n69108, n69109, n69110, n69111, n69112,
    n69113, n69114, n69115, n69116, n69117, n69118, n69119, n69120, n69121,
    n69122, n69123, n69124, n69125, n69126, n69127, n69128, n69129, n69130,
    n69131, n69132, n69133, n69134, n69135, n69136, n69137, n69138, n69139,
    n69140, n69141, n69142, n69143, n69144, n69145, n69146, n69147, n69148,
    n69149, n69150, n69151, n69152, n69153, n69154, n69155, n69156, n69157,
    n69158, n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69166,
    n69167, n69168, n69169, n69170, n69171, n69172, n69173, n69174, n69175,
    n69176, n69177, n69178, n69179, n69180, n69181, n69182, n69183, n69184,
    n69185, n69186, n69187, n69188, n69189, n69190, n69191, n69192, n69193,
    n69194, n69195, n69196, n69197, n69198, n69199, n69200, n69201, n69202,
    n69203, n69204, n69205, n69206, n69207, n69208, n69209, n69210, n69211,
    n69212, n69213, n69214, n69215, n69216, n69217, n69218, n69219, n69220,
    n69221, n69222, n69223, n69224, n69225, n69226, n69227, n69228, n69229,
    n69230, n69231, n69232, n69233, n69234, n69235, n69236, n69237, n69238,
    n69239, n69240, n69241, n69242, n69243, n69244, n69245, n69246, n69247,
    n69248, n69249, n69250, n69251, n69252, n69253, n69254, n69255, n69256,
    n69257, n69258, n69259, n69260, n69261, n69262, n69263, n69264, n69265,
    n69266, n69267, n69268, n69269, n69270, n69271, n69272, n69273, n69274,
    n69275, n69276, n69277, n69278, n69279, n69280, n69281, n69282, n69283,
    n69284, n69285, n69286, n69287, n69288, n69289, n69290, n69291, n69292,
    n69293, n69294, n69295, n69296, n69297, n69298, n69299, n69300, n69301,
    n69302, n69303, n69304, n69305, n69306, n69307, n69308, n69309, n69310,
    n69311, n69312, n69313, n69314, n69315, n69316, n69317, n69318, n69319,
    n69320, n69321, n69322, n69323, n69324, n69325, n69326, n69327, n69328,
    n69329, n69330, n69331, n69332, n69333, n69334, n69335, n69336, n69337,
    n69338, n69339, n69340, n69341, n69342, n69343, n69344, n69345, n69346,
    n69347, n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355,
    n69356, n69357, n69358, n69359, n69360, n69361, n69362, n69363, n69364,
    n69365, n69366, n69367, n69368, n69369, n69370, n69371, n69372, n69373,
    n69374, n69375, n69376, n69377, n69378, n69379, n69380, n69381, n69382,
    n69383, n69384, n69385, n69386, n69387, n69388, n69389, n69390, n69391,
    n69392, n69393, n69394, n69395, n69396, n69397, n69398, n69399, n69400,
    n69401, n69402, n69403, n69404, n69405, n69406, n69407, n69408, n69409,
    n69410, n69411, n69412, n69413, n69414, n69415, n69416, n69417, n69418,
    n69419, n69420, n69421, n69422, n69423, n69424, n69425, n69426, n69427,
    n69428, n69429, n69430, n69431, n69432, n69433, n69434, n69435, n69436,
    n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444, n69445,
    n69446, n69447, n69448, n69449, n69450, n69451, n69452, n69453, n69454,
    n69455, n69456, n69457, n69458, n69459, n69460, n69461, n69462, n69463,
    n69464, n69465, n69466, n69467, n69468, n69469, n69470, n69471, n69472,
    n69473, n69474, n69475, n69476, n69477, n69478, n69479, n69480, n69481,
    n69482, n69483, n69484, n69485, n69486, n69487, n69488, n69489, n69490,
    n69491, n69492, n69493, n69494, n69495, n69496, n69497, n69498, n69499,
    n69500, n69501, n69502, n69503, n69504, n69505, n69506, n69507, n69508,
    n69509, n69510, n69511, n69512, n69513, n69514, n69515, n69516, n69517,
    n69518, n69519, n69520, n69521, n69522, n69523, n69524, n69525, n69526,
    n69527, n69528, n69529, n69530, n69531, n69532, n69533, n69534, n69535,
    n69536, n69537, n69538, n69539, n69540, n69541, n69542, n69543, n69544,
    n69545, n69546, n69547, n69548, n69549, n69550, n69551, n69552, n69553,
    n69554, n69555, n69556, n69557, n69558, n69559, n69560, n69561, n69562,
    n69563, n69564, n69565, n69566, n69567, n69568, n69569, n69570, n69571,
    n69572, n69573, n69574, n69575, n69576, n69577, n69578, n69579, n69580,
    n69581, n69582, n69583, n69584, n69585, n69586, n69587, n69588, n69589,
    n69590, n69591, n69592, n69593, n69594, n69595, n69596, n69597, n69598,
    n69599, n69600, n69601, n69602, n69603, n69604, n69605, n69606, n69607,
    n69608, n69609, n69610, n69611, n69612, n69613, n69614, n69615, n69616,
    n69617, n69618, n69619, n69620, n69621, n69622, n69623, n69624, n69625,
    n69626, n69627, n69628, n69629, n69630, n69631, n69632, n69633, n69634,
    n69635, n69636, n69637, n69638, n69639, n69640, n69641, n69642, n69643,
    n69644, n69645, n69646, n69647, n69648, n69649, n69650, n69651, n69652,
    n69653, n69654, n69655, n69656, n69657, n69658, n69659, n69660, n69661,
    n69662, n69663, n69664, n69665, n69666, n69667, n69668, n69669, n69670,
    n69671, n69672, n69673, n69674, n69675, n69676, n69677, n69678, n69679,
    n69680, n69681, n69682, n69683, n69684, n69685, n69686, n69687, n69688,
    n69689, n69690, n69691, n69692, n69693, n69694, n69695, n69696, n69697,
    n69698, n69699, n69700, n69701, n69702, n69703, n69704, n69705, n69706,
    n69707, n69708, n69709, n69710, n69711, n69712, n69713, n69714, n69715,
    n69716, n69717, n69718, n69719, n69720, n69721, n69722, n69723, n69724,
    n69725, n69726, n69727, n69728, n69729, n69730, n69731, n69732, n69733,
    n69734, n69735, n69736, n69737, n69738, n69739, n69740, n69741, n69742,
    n69743, n69744, n69745, n69746, n69747, n69748, n69749, n69750, n69751,
    n69752, n69753, n69754, n69755, n69756, n69757, n69758, n69759, n69760,
    n69761, n69762, n69763, n69764, n69765, n69766, n69767, n69768, n69769,
    n69770, n69771, n69772, n69773, n69774, n69775, n69776, n69777, n69778,
    n69779, n69780, n69781, n69782, n69783, n69784, n69785, n69786, n69787,
    n69788, n69789, n69790, n69791, n69792, n69793, n69794, n69795, n69796,
    n69797, n69798, n69799, n69800, n69801, n69802, n69803, n69804, n69805,
    n69806, n69807, n69808, n69809, n69810, n69811, n69812, n69813, n69814,
    n69815, n69816, n69817, n69818, n69819, n69820, n69821, n69822, n69823,
    n69824, n69825, n69826, n69827, n69828, n69829, n69830, n69831, n69832,
    n69833, n69834, n69835, n69836, n69837, n69838, n69839, n69840, n69841,
    n69842, n69843, n69844, n69845, n69846, n69847, n69848, n69849, n69850,
    n69851, n69852, n69853, n69854, n69855, n69856, n69857, n69858, n69859,
    n69860, n69861, n69862, n69863, n69864, n69865, n69866, n69867, n69868,
    n69869, n69870, n69871, n69872, n69873, n69874, n69875, n69876, n69877,
    n69878, n69879, n69880, n69881, n69882, n69883, n69884, n69885, n69886,
    n69887, n69888, n69889, n69890, n69891, n69892, n69893, n69894, n69895,
    n69896, n69897, n69898, n69899, n69900, n69901, n69902, n69903, n69904,
    n69905, n69906, n69907, n69908, n69909, n69910, n69911, n69912, n69913,
    n69914, n69915, n69916, n69917, n69918, n69919, n69920, n69921, n69922,
    n69923, n69924, n69925, n69926, n69927, n69928, n69929, n69930, n69931,
    n69932, n69933, n69934, n69935, n69936, n69937, n69938, n69939, n69940,
    n69941, n69942, n69943, n69944, n69945, n69946, n69947, n69948, n69949,
    n69950, n69951, n69952, n69953, n69954, n69955, n69956, n69957, n69958,
    n69959, n69960, n69961, n69962, n69963, n69964, n69965, n69966, n69967,
    n69968, n69969, n69970, n69971, n69972, n69973, n69974, n69975, n69976,
    n69977, n69978, n69979, n69980, n69981, n69982, n69983, n69984, n69985,
    n69986, n69987, n69988, n69989, n69990, n69991, n69992, n69993, n69994,
    n69995, n69996, n69997, n69998, n69999, n70000, n70001, n70002, n70003,
    n70004, n70005, n70006, n70007, n70008, n70009, n70010, n70011, n70012,
    n70013, n70014, n70015, n70016, n70017, n70018, n70019, n70020, n70021,
    n70022, n70023, n70024, n70025, n70026, n70027, n70028, n70029, n70030,
    n70031, n70032, n70033, n70034, n70035, n70036, n70037, n70038, n70039,
    n70040, n70041, n70042, n70043, n70044, n70045, n70046, n70047, n70048,
    n70049, n70050, n70051, n70052, n70053, n70054, n70055, n70056, n70057,
    n70058, n70059, n70060, n70061, n70062, n70063, n70064, n70065, n70066,
    n70067, n70068, n70069, n70070, n70071, n70072, n70073, n70074, n70075,
    n70076, n70077, n70078, n70079, n70080, n70081, n70082, n70083, n70084,
    n70085, n70086, n70087, n70088, n70089, n70090, n70091, n70092, n70093,
    n70094, n70095, n70096, n70097, n70098, n70099, n70100, n70101, n70102,
    n70103, n70104, n70105, n70106, n70107, n70108, n70109, n70110, n70111,
    n70112, n70113, n70114, n70115, n70116, n70117, n70118, n70119, n70120,
    n70121, n70122, n70123, n70124, n70125, n70126, n70127, n70128, n70129,
    n70130, n70131, n70132, n70133, n70134, n70135, n70136, n70137, n70138,
    n70139, n70140, n70141, n70142, n70143, n70144, n70145, n70146, n70147,
    n70148, n70149, n70150, n70151, n70152, n70153, n70154, n70155, n70156,
    n70157, n70158, n70159, n70160, n70161, n70162, n70163, n70164, n70165,
    n70166, n70167, n70168, n70169, n70170, n70171, n70172, n70173, n70174,
    n70175, n70176, n70177, n70178, n70179, n70180, n70181, n70182, n70183,
    n70184, n70185, n70186, n70187, n70188, n70189, n70190, n70191, n70192,
    n70193, n70194, n70195, n70196, n70197, n70198, n70199, n70200, n70201,
    n70202, n70203, n70204, n70205, n70206, n70207, n70208, n70209, n70210,
    n70211, n70212, n70213, n70214, n70215, n70216, n70217, n70218, n70219,
    n70220, n70221, n70222, n70223, n70224, n70225, n70226, n70227, n70228,
    n70229, n70230, n70231, n70232, n70233, n70234, n70235, n70236, n70237,
    n70238, n70239, n70240, n70241, n70242, n70243, n70244, n70245, n70246,
    n70247, n70248, n70249, n70250, n70251, n70252, n70253, n70254, n70255,
    n70256, n70257, n70258, n70259, n70260, n70261, n70262, n70263, n70264,
    n70265, n70266, n70267, n70268, n70269, n70270, n70271, n70272, n70273,
    n70274, n70275, n70276, n70277, n70278, n70279, n70280, n70281, n70282,
    n70283, n70284, n70285, n70286, n70287, n70288, n70289, n70290, n70291,
    n70292, n70293, n70294, n70295, n70296, n70297, n70298, n70299, n70300,
    n70301, n70302, n70303, n70304, n70305, n70306, n70307, n70308, n70309,
    n70310, n70311, n70312, n70313, n70314, n70315, n70316, n70317, n70318,
    n70319, n70320, n70321, n70322, n70323, n70324, n70325, n70326, n70327,
    n70328, n70329, n70330, n70331, n70332, n70333, n70334, n70335, n70336,
    n70337, n70338, n70339, n70340, n70341, n70342, n70343, n70344, n70345,
    n70346, n70347, n70348, n70349, n70350, n70351, n70352, n70353, n70354,
    n70355, n70356, n70357, n70358, n70359, n70360, n70361, n70362, n70363,
    n70364, n70365, n70366, n70367, n70368, n70369, n70370, n70371, n70372,
    n70373, n70374, n70375, n70376, n70377, n70378, n70379, n70380, n70381,
    n70382, n70383, n70384, n70385, n70386, n70387, n70388, n70389, n70390,
    n70391, n70392, n70393, n70394, n70395, n70396, n70397, n70398, n70399,
    n70400, n70401, n70402, n70403, n70404, n70405, n70406, n70407, n70408,
    n70409, n70410, n70411, n70412, n70413, n70414, n70415, n70416, n70417,
    n70418, n70419, n70420, n70421, n70422, n70423, n70424, n70425, n70426,
    n70427, n70428, n70429, n70430, n70431, n70432, n70433, n70434, n70435,
    n70436, n70437, n70438, n70439, n70440, n70441, n70442, n70443, n70444,
    n70445, n70446, n70447, n70448, n70449, n70450, n70451, n70452, n70453,
    n70454, n70455, n70456, n70457, n70458, n70459, n70460, n70461, n70462,
    n70463, n70464, n70465, n70466, n70467, n70468, n70469, n70470, n70471,
    n70472, n70473, n70474, n70475, n70476, n70477, n70478, n70479, n70480,
    n70481, n70482, n70483, n70484, n70485, n70486, n70487, n70488, n70489,
    n70490, n70491, n70492, n70493, n70494, n70495, n70496, n70497, n70498,
    n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507,
    n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516,
    n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524, n70525,
    n70526, n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534,
    n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542, n70543,
    n70544, n70545, n70546, n70547, n70548, n70549, n70550, n70551, n70552,
    n70553, n70554, n70555, n70556, n70557, n70558, n70559, n70560, n70561,
    n70562, n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570,
    n70571, n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579,
    n70580, n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588,
    n70589, n70590, n70591, n70592, n70593, n70594, n70595, n70596, n70597,
    n70598, n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606,
    n70607, n70608, n70609, n70610, n70611, n70612, n70613, n70614, n70615,
    n70616, n70617, n70618, n70619, n70620, n70621, n70622, n70623, n70624,
    n70625, n70626, n70627, n70628, n70629, n70630, n70631, n70632, n70633,
    n70634, n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642,
    n70643, n70644, n70645, n70646, n70647, n70648, n70649, n70650, n70651,
    n70652, n70653, n70654, n70655, n70656, n70657, n70658, n70659, n70660,
    n70661, n70662, n70663, n70664, n70665, n70666, n70667, n70668, n70669,
    n70670, n70671, n70672, n70673, n70674, n70675, n70676, n70677, n70678,
    n70679, n70680, n70681, n70682, n70683, n70684, n70685, n70686, n70687,
    n70688, n70689, n70690, n70691, n70692, n70693, n70694, n70695, n70696,
    n70697, n70698, n70699, n70700, n70701, n70702, n70703, n70704, n70705,
    n70706, n70707, n70708, n70709, n70710, n70711, n70712, n70713, n70714,
    n70715, n70716, n70717, n70718, n70719, n70720, n70721, n70722, n70723,
    n70724, n70725, n70726, n70727, n70728, n70729, n70730, n70731, n70732,
    n70733, n70734, n70735, n70736, n70737, n70738, n70739, n70740, n70741,
    n70742, n70743, n70744, n70745, n70746, n70747, n70748, n70749, n70750,
    n70751, n70752, n70753, n70754, n70755, n70756, n70757, n70758, n70759,
    n70760, n70761, n70762, n70763, n70764, n70765, n70766, n70767, n70768,
    n70769, n70770, n70771, n70772, n70773, n70774, n70775, n70776, n70777,
    n70778, n70779, n70780, n70781, n70782, n70783, n70784, n70785, n70786,
    n70787, n70788, n70789, n70790, n70791, n70792, n70793, n70794, n70795,
    n70796, n70797, n70798, n70799, n70800, n70801, n70802, n70803, n70804,
    n70805, n70806, n70807, n70808, n70809, n70810, n70811, n70812, n70813,
    n70814, n70815, n70816, n70817, n70818, n70819, n70820, n70821, n70822,
    n70823, n70824, n70825, n70826, n70827, n70828, n70829, n70830, n70831,
    n70832, n70833, n70834, n70835, n70836, n70837, n70838, n70839, n70840,
    n70841, n70842, n70843, n70844, n70845, n70846, n70847, n70848, n70849,
    n70850, n70851, n70852, n70853, n70854, n70855, n70856, n70857, n70858,
    n70859, n70860, n70861, n70862, n70863, n70864, n70865, n70866, n70867,
    n70868, n70869, n70870, n70871, n70872, n70873, n70874, n70875, n70876,
    n70877, n70878, n70879, n70880, n70881, n70882, n70883, n70884, n70885,
    n70886, n70887, n70888, n70889, n70890, n70891, n70892, n70893, n70894,
    n70895, n70896, n70897, n70898, n70899, n70900, n70901, n70902, n70903,
    n70904, n70905, n70906, n70907, n70908, n70909, n70910, n70911, n70912,
    n70913, n70914, n70915, n70916, n70917, n70918, n70919, n70920, n70921,
    n70922, n70923, n70924, n70925, n70926, n70927, n70928, n70929, n70930,
    n70931, n70932, n70933, n70934, n70935, n70936, n70937, n70938, n70939,
    n70940, n70941, n70942, n70943, n70944, n70945, n70946, n70947, n70948,
    n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956, n70957,
    n70958, n70959, n70960, n70961, n70962, n70963, n70964, n70965, n70966,
    n70967, n70968, n70969, n70970, n70971, n70972, n70973, n70974, n70975,
    n70976, n70977, n70978, n70979, n70980, n70981, n70982, n70983, n70984,
    n70985, n70986, n70987, n70988, n70989, n70990, n70991, n70992, n70993,
    n70994, n70995, n70996, n70997, n70998, n70999, n71000, n71001, n71002,
    n71003, n71004, n71005, n71006, n71007, n71008, n71009, n71010, n71011,
    n71012, n71013, n71014, n71015, n71016, n71017, n71018, n71019, n71020,
    n71021, n71022, n71023, n71024, n71025, n71026, n71027, n71028, n71029,
    n71030, n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038,
    n71039, n71040, n71041, n71042, n71043, n71044, n71045, n71046, n71047,
    n71048, n71049, n71050, n71051, n71052, n71053, n71054, n71055, n71056,
    n71057, n71058, n71059, n71060, n71061, n71062, n71063, n71064, n71065,
    n71066, n71067, n71068, n71069, n71070, n71071, n71072, n71073, n71074,
    n71075, n71076, n71077, n71078, n71079, n71080, n71081, n71082, n71083,
    n71084, n71085, n71086, n71087, n71088, n71089, n71090, n71091, n71092,
    n71093, n71094, n71095, n71096, n71097, n71098, n71099, n71100, n71101,
    n71102, n71103, n71104, n71105, n71106, n71107, n71108, n71109, n71110,
    n71111, n71112, n71113, n71114, n71115, n71116, n71117, n71118, n71119,
    n71120, n71121, n71122, n71123, n71124, n71125, n71126, n71127, n71128,
    n71129, n71130, n71131, n71132, n71133, n71134, n71135, n71136, n71137,
    n71138, n71139, n71140, n71141, n71142, n71143, n71144, n71145, n71146,
    n71147, n71148, n71149, n71150, n71151, n71152, n71153, n71154, n71155,
    n71156, n71157, n71158, n71159, n71160, n71161, n71162, n71163, n71164,
    n71165, n71166, n71167, n71168, n71169, n71170, n71171, n71172, n71173,
    n71174, n71175, n71176, n71177, n71178, n71179, n71180, n71181, n71182,
    n71183, n71184, n71185, n71186, n71187, n71188, n71189, n71190, n71191,
    n71192, n71193, n71194, n71195, n71196, n71197, n71198, n71199, n71200,
    n71201, n71202, n71203, n71204, n71205, n71206, n71207, n71208, n71209,
    n71210, n71211, n71212, n71213, n71214, n71215, n71216, n71217, n71218,
    n71219, n71220, n71221, n71222, n71223, n71224, n71225, n71226, n71227,
    n71228, n71229, n71230, n71231, n71232, n71233, n71234, n71235, n71236,
    n71237, n71238, n71239, n71240, n71241, n71242, n71243, n71244, n71245,
    n71246, n71247, n71248, n71249, n71250, n71251, n71252, n71253, n71254,
    n71255, n71256, n71257, n71258, n71259, n71260, n71261, n71262, n71263,
    n71264, n71265, n71266, n71267, n71268, n71269, n71270, n71271, n71272,
    n71273, n71274, n71275, n71276, n71277, n71278, n71279, n71280, n71281,
    n71282, n71283, n71284, n71285, n71286, n71287, n71288, n71289, n71290,
    n71291, n71292, n71293, n71294, n71295, n71296, n71297, n71298, n71299,
    n71300, n71301, n71302, n71303, n71304, n71305, n71306, n71307, n71308,
    n71309, n71310, n71311, n71312, n71313, n71314, n71315, n71316, n71317,
    n71318, n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326,
    n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334, n71335,
    n71336, n71337, n71338, n71339, n71340, n71341, n71342, n71343, n71344,
    n71345, n71346, n71347, n71348, n71349, n71350, n71351, n71352, n71353,
    n71354, n71355, n71356, n71357, n71358, n71359, n71360, n71361, n71362,
    n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370, n71371,
    n71372, n71373, n71374, n71375, n71376, n71377, n71378, n71379, n71380,
    n71381, n71382, n71383, n71384, n71385, n71386, n71387, n71388, n71389,
    n71390, n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398,
    n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406, n71407,
    n71408, n71409, n71410, n71411, n71412, n71413, n71414, n71415, n71416,
    n71417, n71418, n71419, n71420, n71421, n71422, n71423, n71424, n71425,
    n71426, n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434,
    n71435, n71436, n71437, n71438, n71439, n71440, n71441, n71442, n71443,
    n71444, n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452,
    n71453, n71454, n71455, n71456, n71457, n71458, n71459, n71460, n71461,
    n71462, n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470,
    n71471, n71472, n71473, n71474, n71475, n71476, n71477, n71478, n71479,
    n71480, n71481, n71482, n71483, n71484, n71485, n71486, n71487, n71488,
    n71489, n71490, n71491, n71492, n71493, n71494, n71495, n71496, n71497,
    n71498, n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506,
    n71507, n71508, n71509, n71510, n71511, n71512, n71513, n71514, n71515,
    n71516, n71517, n71518, n71519, n71520, n71521, n71522, n71523, n71524,
    n71525, n71526, n71527, n71528, n71529, n71530, n71531, n71532, n71533,
    n71534, n71535, n71536, n71537, n71538, n71539, n71540, n71541, n71542,
    n71543, n71544, n71545, n71546, n71547, n71548, n71549, n71550, n71551,
    n71552, n71553, n71554, n71555, n71556, n71557, n71558, n71559, n71560,
    n71561, n71562, n71563, n71564, n71565, n71566, n71567, n71568, n71569,
    n71570, n71571, n71572, n71573, n71574, n71575, n71576, n71577, n71578,
    n71579, n71580, n71581, n71582, n71583, n71584, n71585, n71586, n71587,
    n71588, n71589, n71590, n71591, n71592, n71593, n71594, n71595, n71596,
    n71597, n71598, n71599, n71600, n71601, n71602, n71603, n71604, n71605,
    n71606, n71607, n71608, n71609, n71610, n71611, n71612, n71613, n71614,
    n71615, n71616, n71617, n71618, n71619, n71620, n71621, n71622, n71623,
    n71624, n71625, n71626, n71627, n71628, n71629, n71630, n71631, n71632,
    n71633, n71634, n71635, n71636, n71637, n71638, n71639, n71640, n71641,
    n71642, n71643, n71644, n71645, n71646, n71647, n71648, n71649, n71650,
    n71651, n71652, n71653, n71654, n71655, n71656, n71657, n71658, n71659,
    n71660, n71661, n71662, n71663, n71664, n71665, n71666, n71667, n71668,
    n71669, n71670, n71671, n71672, n71673, n71674, n71675, n71676, n71677,
    n71678, n71679, n71680, n71681, n71682, n71683, n71684, n71685, n71686,
    n71687, n71688, n71689, n71690, n71691, n71692, n71693, n71694, n71695,
    n71696, n71697, n71698, n71699, n71700, n71701, n71702, n71703, n71704,
    n71705, n71706, n71707, n71708, n71709, n71710, n71711, n71712, n71713,
    n71714, n71715, n71716, n71717, n71718, n71719, n71720, n71721, n71722,
    n71723, n71724, n71725, n71726, n71727, n71728, n71729, n71730, n71731,
    n71732, n71733, n71734, n71735, n71736, n71737, n71738, n71739, n71740,
    n71741, n71742, n71743, n71744, n71745, n71746, n71747, n71748, n71749,
    n71750, n71751, n71752, n71753, n71754, n71755, n71756, n71757, n71758,
    n71759, n71760, n71761, n71762, n71763, n71764, n71765, n71766, n71767,
    n71768, n71769, n71770, n71771, n71772, n71773, n71774, n71775, n71776,
    n71777, n71778, n71779, n71780, n71781, n71782, n71783, n71784, n71785,
    n71786, n71787, n71788, n71789, n71790, n71791, n71792, n71793, n71794,
    n71795, n71796, n71797, n71798, n71799, n71800, n71801, n71802, n71803,
    n71804, n71805, n71806, n71807, n71808, n71809, n71810, n71811, n71812,
    n71813, n71814, n71815, n71816, n71817, n71818, n71819, n71820, n71821,
    n71822, n71823, n71824, n71825, n71826, n71827, n71828, n71829, n71830,
    n71831, n71832, n71833, n71834, n71835, n71836, n71837, n71838, n71839,
    n71840, n71841, n71842, n71843, n71844, n71845, n71846, n71847, n71848,
    n71849, n71850, n71851, n71852, n71853, n71854, n71855, n71856, n71857,
    n71858, n71859, n71860, n71861, n71862, n71863, n71864, n71865, n71866,
    n71867, n71868, n71869, n71870, n71871, n71872, n71873, n71874, n71875,
    n71876, n71877, n71878, n71879, n71880, n71881, n71882, n71883, n71884,
    n71885, n71886, n71887, n71888, n71889, n71890, n71891, n71892, n71893,
    n71894, n71895, n71896, n71897, n71898, n71899, n71900, n71901, n71902,
    n71903, n71904, n71905, n71906, n71907, n71908, n71909, n71910, n71911,
    n71912, n71913, n71914, n71915, n71916, n71917, n71918, n71919, n71920,
    n71921, n71922, n71923, n71924, n71925, n71926, n71927, n71928, n71929,
    n71930, n71931, n71932, n71933, n71934, n71935, n71936, n71937, n71938,
    n71939, n71940, n71941, n71942, n71943, n71944, n71945, n71946, n71947,
    n71948, n71949, n71950, n71951, n71952, n71953, n71954, n71955, n71956,
    n71957, n71958, n71959, n71960, n71961, n71962, n71963, n71964, n71965,
    n71966, n71967, n71968, n71969, n71970, n71971, n71972, n71973, n71974,
    n71975, n71976, n71977, n71978, n71979, n71980, n71981, n71982, n71983,
    n71984, n71985, n71986, n71987, n71988, n71989, n71990, n71991, n71992,
    n71993, n71994, n71995, n71996, n71997, n71998, n71999, n72000, n72001,
    n72002, n72003, n72004, n72005, n72006, n72007, n72008, n72009, n72010,
    n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018, n72019,
    n72020, n72021, n72022, n72023, n72024, n72025, n72026, n72027, n72028,
    n72029, n72030, n72031, n72032, n72033, n72034, n72035, n72036, n72037,
    n72038, n72039, n72040, n72041, n72042, n72043, n72044, n72045, n72046,
    n72047, n72048, n72049, n72050, n72051, n72052, n72053, n72054, n72055,
    n72056, n72057, n72058, n72059, n72060, n72061, n72062, n72063, n72064,
    n72065, n72066, n72067, n72068, n72069, n72070, n72071, n72072, n72073,
    n72074, n72075, n72076, n72077, n72078, n72079, n72080, n72081, n72082,
    n72083, n72084, n72085, n72086, n72087, n72088, n72089, n72090, n72091,
    n72092, n72093, n72094, n72095, n72096, n72097, n72098, n72099, n72100,
    n72101, n72102, n72103, n72104, n72105, n72106, n72107, n72108, n72109,
    n72110, n72111, n72112, n72113, n72114, n72115, n72116, n72117, n72118,
    n72119, n72120, n72121, n72122, n72123, n72124, n72125, n72126, n72127,
    n72128, n72129, n72130, n72131, n72132, n72133, n72134, n72135, n72136,
    n72137, n72138, n72139, n72140, n72141, n72142, n72143, n72144, n72145,
    n72146, n72147, n72148, n72149, n72150, n72151, n72152, n72153, n72154,
    n72155, n72156, n72157, n72158, n72159, n72160, n72161, n72162, n72163,
    n72164, n72165, n72166, n72167, n72168, n72169, n72170, n72171, n72172,
    n72173, n72174, n72175, n72176, n72177, n72178, n72179, n72180, n72181,
    n72182, n72183, n72184, n72185, n72186, n72187, n72188, n72189, n72190,
    n72191, n72192, n72193, n72194, n72195, n72196, n72197, n72198, n72199,
    n72200, n72201, n72202, n72203, n72204, n72205, n72206, n72207, n72208,
    n72209, n72210, n72211, n72212, n72213, n72214, n72215, n72216, n72217,
    n72218, n72219, n72220, n72221, n72222, n72223, n72224, n72225, n72226,
    n72227, n72228, n72229, n72230, n72231, n72232, n72233, n72234, n72235,
    n72236, n72237, n72238, n72239, n72240, n72241, n72242, n72243, n72244,
    n72245, n72246, n72247, n72248, n72249, n72250, n72251, n72252, n72253,
    n72254, n72255, n72256, n72257, n72258, n72259, n72260, n72261, n72262,
    n72263, n72264, n72265, n72266, n72267, n72268, n72269, n72270, n72271,
    n72272, n72273, n72274, n72275, n72276, n72277, n72278, n72279, n72280,
    n72281, n72282, n72283, n72284, n72285, n72286, n72287, n72288, n72289,
    n72290, n72291, n72292, n72293, n72294, n72295, n72296, n72297, n72298,
    n72299, n72300, n72301, n72302, n72303, n72304, n72305, n72306, n72307,
    n72308, n72309, n72310, n72311, n72312, n72313, n72314, n72315, n72316,
    n72317, n72318, n72319, n72320, n72321, n72322, n72323, n72324, n72325,
    n72326, n72327, n72328, n72329, n72330, n72331, n72332, n72333, n72334,
    n72335, n72336, n72337, n72338, n72339, n72340, n72341, n72342, n72343,
    n72344, n72345, n72346, n72347, n72348, n72349, n72350, n72351, n72352,
    n72353, n72354, n72355, n72356, n72357, n72358, n72359, n72360, n72361,
    n72362, n72363, n72364, n72365, n72366, n72367, n72368, n72369, n72370,
    n72371, n72372, n72373, n72374, n72375, n72376, n72377, n72378, n72379,
    n72380, n72381, n72382, n72383, n72384, n72385, n72386, n72387, n72388,
    n72389, n72390, n72391, n72392, n72393, n72394, n72395, n72396, n72397,
    n72398, n72399, n72400, n72401, n72402, n72403, n72404, n72405, n72406,
    n72407, n72408, n72409, n72410, n72411, n72412, n72413, n72414, n72415,
    n72416, n72417, n72418, n72419, n72420, n72421, n72422, n72423, n72424,
    n72425, n72426, n72427, n72428, n72429, n72430, n72431, n72432, n72433,
    n72434, n72435, n72436, n72437, n72438, n72439, n72440, n72441, n72442,
    n72443, n72444, n72445, n72446, n72447, n72448, n72449, n72450, n72451,
    n72452, n72453, n72454, n72455, n72456, n72457, n72458, n72459, n72460,
    n72461, n72462, n72463, n72464, n72465, n72466, n72467, n72468, n72469,
    n72470, n72471, n72472, n72473, n72474, n72475, n72476, n72477, n72478,
    n72479, n72480, n72481, n72482, n72483, n72484, n72485, n72486, n72487,
    n72488, n72489, n72490, n72491, n72492, n72493, n72494, n72495, n72496,
    n72497, n72498, n72499, n72500, n72501, n72502, n72503, n72504, n72505,
    n72506, n72507, n72508, n72509, n72510, n72511, n72512, n72513, n72514,
    n72515, n72516, n72517, n72518, n72519, n72520, n72521, n72522, n72523,
    n72524, n72525, n72526, n72527, n72528, n72529, n72530, n72531, n72532,
    n72533, n72534, n72535, n72536, n72537, n72538, n72539, n72540, n72541,
    n72542, n72543, n72544, n72545, n72546, n72547, n72548, n72549, n72550,
    n72551, n72552, n72553, n72554, n72555, n72556, n72557, n72558, n72559,
    n72560, n72561, n72562, n72563, n72564, n72565, n72566, n72567, n72568,
    n72569, n72570, n72571, n72572, n72573, n72574, n72575, n72576, n72577,
    n72578, n72579, n72580, n72581, n72582, n72583, n72584, n72585, n72586,
    n72587, n72588, n72589, n72590, n72591, n72592, n72593, n72594, n72595,
    n72596, n72597, n72598, n72599, n72600, n72601, n72602, n72603, n72604,
    n72605, n72606, n72607, n72608, n72609, n72610, n72611, n72612, n72613,
    n72614, n72615, n72616, n72617, n72618, n72619, n72620, n72621, n72622,
    n72623, n72624, n72625, n72626, n72627, n72628, n72629, n72630, n72631,
    n72632, n72633, n72634, n72635, n72636, n72637, n72638, n72639, n72640,
    n72641, n72642, n72643, n72644, n72645, n72646, n72647, n72648, n72649,
    n72650, n72651, n72652, n72653, n72654, n72655, n72656, n72657, n72658,
    n72659, n72660, n72661, n72662, n72663, n72664, n72665, n72666, n72667,
    n72668, n72669, n72670, n72671, n72672, n72673, n72674, n72675, n72676,
    n72677, n72678, n72679, n72680, n72681, n72682, n72683, n72684, n72685,
    n72686, n72687, n72688, n72689, n72690, n72691, n72692, n72693, n72694,
    n72695, n72696, n72697, n72698, n72699, n72700, n72701, n72702, n72703,
    n72704, n72705, n72706, n72707, n72708, n72709, n72710, n72711, n72712,
    n72713, n72714, n72715, n72716, n72717, n72718, n72719, n72720, n72721,
    n72722, n72723, n72724, n72725, n72726, n72727, n72728, n72729, n72730,
    n72731, n72732, n72733, n72734, n72735, n72736, n72737, n72738, n72739,
    n72740, n72741, n72742, n72743, n72744, n72745, n72746, n72747, n72748,
    n72749, n72750, n72751, n72752, n72753, n72754, n72755, n72756, n72757,
    n72758, n72759, n72760, n72761, n72762, n72763, n72764, n72765, n72766,
    n72767, n72768, n72769, n72770, n72771, n72772, n72773, n72774, n72775,
    n72776, n72777, n72778, n72779, n72780, n72781, n72782, n72783, n72784,
    n72785, n72786, n72787, n72788, n72789, n72790, n72791, n72792, n72793,
    n72794, n72795, n72796, n72797, n72798, n72799, n72800, n72801, n72802,
    n72803, n72804, n72805, n72806, n72807, n72808, n72809, n72810, n72811,
    n72812, n72813, n72814, n72815, n72816, n72817, n72818, n72819, n72820,
    n72821, n72822, n72823, n72824, n72825, n72826, n72827, n72828, n72829,
    n72830, n72831, n72832, n72833, n72834, n72835, n72836, n72837, n72838,
    n72839, n72840, n72841, n72842, n72843, n72844, n72845, n72846, n72847,
    n72848, n72849, n72850, n72851, n72852, n72853, n72854, n72855, n72856,
    n72857, n72858, n72859, n72860, n72861, n72862, n72863, n72864, n72865,
    n72866, n72867, n72868, n72869, n72870, n72871, n72872, n72873, n72874,
    n72875, n72876, n72877, n72878, n72879, n72880, n72881, n72882, n72883,
    n72884, n72885, n72886, n72887, n72888, n72889, n72890, n72891, n72892,
    n72893, n72894, n72895, n72896, n72897, n72898, n72899, n72900, n72901,
    n72902, n72903, n72904, n72905, n72906, n72907, n72908, n72909, n72910,
    n72911, n72912, n72913, n72914, n72915, n72916, n72917, n72918, n72919,
    n72920, n72921, n72922, n72923, n72924, n72925, n72926, n72927, n72928,
    n72929, n72930, n72931, n72932, n72933, n72934, n72935, n72936, n72937,
    n72938, n72939, n72940, n72941, n72942, n72943, n72944, n72945, n72946,
    n72947, n72948, n72949, n72950, n72951, n72952, n72953, n72954, n72955,
    n72956, n72957, n72958, n72959, n72960, n72961, n72962, n72963, n72964,
    n72965, n72966, n72967, n72968, n72969, n72970, n72971, n72972, n72973,
    n72974, n72975, n72976, n72977, n72978, n72979, n72980, n72981, n72982,
    n72983, n72984, n72985, n72986, n72987, n72988, n72989, n72990, n72991,
    n72992, n72993, n72994, n72995, n72996, n72997, n72998, n72999, n73000,
    n73001, n73002, n73003, n73004, n73005, n73006, n73007, n73008, n73009,
    n73010, n73011, n73012, n73013, n73014, n73015, n73016, n73017, n73018,
    n73019, n73020, n73021, n73022, n73023, n73024, n73025, n73026, n73027,
    n73028, n73029, n73030, n73031, n73032, n73033, n73034, n73035, n73036,
    n73037, n73038, n73039, n73040, n73041, n73042, n73043, n73044, n73045,
    n73046, n73047, n73048, n73049, n73050, n73051, n73052, n73053, n73054,
    n73055, n73056, n73057, n73058, n73059, n73060, n73061, n73062, n73063,
    n73064, n73065, n73066, n73067, n73068, n73069, n73070, n73071, n73072,
    n73073, n73074, n73075, n73076, n73077, n73078, n73079, n73080, n73081,
    n73082, n73083, n73084, n73085, n73086, n73087, n73088, n73089, n73090,
    n73091, n73092, n73093, n73094, n73095, n73096, n73097, n73098, n73099,
    n73100, n73101, n73102, n73103, n73104, n73105, n73106, n73107, n73108,
    n73109, n73110, n73111, n73112, n73113, n73114, n73115, n73116, n73117,
    n73118, n73119, n73120, n73121, n73122, n73123, n73124, n73125, n73126,
    n73127, n73128, n73129, n73130, n73131, n73132, n73133, n73134, n73135,
    n73136, n73137, n73138, n73139, n73140, n73141, n73142, n73143, n73144,
    n73145, n73146, n73147, n73148, n73149, n73150, n73151, n73152, n73153,
    n73154, n73155, n73156, n73157, n73158, n73159, n73160, n73161, n73162,
    n73163, n73164, n73165, n73166, n73167, n73168, n73169, n73170, n73171,
    n73172, n73173, n73174, n73175, n73176, n73177, n73178, n73179, n73180,
    n73181, n73182, n73183, n73184, n73185, n73186, n73187, n73188, n73189,
    n73190, n73191, n73192, n73193, n73194, n73195, n73196, n73197, n73198,
    n73199, n73200, n73201, n73202, n73203, n73204, n73205, n73206, n73207,
    n73208, n73209, n73210, n73211, n73212, n73213, n73214, n73215, n73216,
    n73217, n73218, n73219, n73220, n73221, n73222, n73223, n73224, n73225,
    n73226, n73227, n73228, n73229, n73230, n73231, n73232, n73233, n73234,
    n73235, n73236, n73237, n73238, n73239, n73240, n73241, n73242, n73243,
    n73244, n73245, n73246, n73247, n73248, n73249, n73250, n73251, n73252,
    n73253, n73254, n73255, n73256, n73257, n73258, n73259, n73260, n73261,
    n73262, n73263, n73264, n73265, n73266, n73267, n73268, n73269, n73270,
    n73271, n73272, n73273, n73274, n73275, n73276, n73277, n73278, n73279,
    n73280, n73281, n73282, n73283, n73284, n73285, n73286, n73287, n73288,
    n73289, n73290, n73291, n73292, n73293, n73294, n73295, n73296, n73297,
    n73298, n73299, n73300, n73301, n73302, n73303, n73304, n73305, n73306,
    n73307, n73308, n73309, n73310, n73311, n73312, n73313, n73314, n73315,
    n73316, n73317, n73318, n73319, n73320, n73321, n73322, n73323, n73324,
    n73325, n73326, n73327, n73328, n73329, n73330, n73331, n73332, n73333,
    n73334, n73335, n73336, n73337, n73338, n73339, n73340, n73341, n73342,
    n73343, n73344, n73345, n73346, n73347, n73348, n73349, n73350, n73351,
    n73352, n73353, n73354, n73355, n73356, n73357, n73358, n73359, n73360,
    n73361, n73362, n73363, n73364, n73365, n73366, n73367, n73368, n73369,
    n73370, n73371, n73372, n73373, n73374, n73375, n73376, n73377, n73378,
    n73379, n73380, n73381, n73382, n73383, n73384, n73385, n73386, n73387,
    n73388, n73389, n73390, n73391, n73392, n73393, n73394, n73395, n73396,
    n73397, n73398, n73399, n73400, n73401, n73402, n73403, n73404, n73405,
    n73406, n73407, n73408, n73409, n73410, n73411, n73412, n73413, n73414,
    n73415, n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423,
    n73424, n73425, n73426, n73427, n73428, n73429, n73430, n73431, n73432,
    n73433, n73434, n73435, n73436, n73437, n73438, n73439, n73440, n73441,
    n73442, n73443, n73444, n73445, n73446, n73447, n73448, n73449, n73450,
    n73451, n73452, n73453, n73454, n73455, n73456, n73457, n73458, n73459,
    n73460, n73461, n73462, n73463, n73464, n73465, n73466, n73467, n73468,
    n73469, n73470, n73471, n73472, n73473, n73474, n73475, n73476, n73477,
    n73478, n73479, n73480, n73481, n73482, n73483, n73484, n73485, n73486,
    n73487, n73488, n73489, n73490, n73491, n73492, n73493, n73494, n73495,
    n73496, n73497, n73498, n73499, n73500, n73501, n73502, n73503, n73504,
    n73505, n73506, n73507, n73508, n73509, n73510, n73511, n73512, n73513,
    n73514, n73515, n73516, n73517, n73518, n73519, n73520, n73521, n73522,
    n73523, n73524, n73525, n73526, n73527, n73528, n73529, n73530, n73531,
    n73532, n73533, n73534, n73535, n73536, n73537, n73538, n73539, n73540,
    n73541, n73542, n73543, n73544, n73545, n73546, n73547, n73548, n73549,
    n73550, n73551, n73552, n73553, n73554, n73555, n73556, n73557, n73558,
    n73559, n73560, n73561, n73562, n73563, n73564, n73565, n73566, n73567,
    n73568, n73569, n73570, n73571, n73572, n73573, n73574, n73575, n73576,
    n73577, n73578, n73579, n73580, n73581, n73582, n73583, n73584, n73585,
    n73586, n73587, n73588, n73589, n73590, n73591, n73592, n73593, n73594,
    n73595, n73596, n73597, n73598, n73599, n73600, n73601, n73602, n73603,
    n73604, n73605, n73606, n73607, n73608, n73609, n73610, n73611, n73612,
    n73613, n73614, n73615, n73616, n73617, n73618, n73619, n73620, n73621,
    n73622, n73623, n73624, n73625, n73626, n73627, n73628, n73629, n73630,
    n73631, n73632, n73633, n73634, n73635, n73636, n73637, n73638, n73639,
    n73640, n73641, n73642, n73643, n73644, n73645, n73646, n73647, n73648,
    n73649, n73650, n73651, n73652, n73653, n73654, n73655, n73656, n73657,
    n73658, n73659, n73660, n73661, n73662, n73663, n73664, n73665, n73666,
    n73667, n73668, n73669, n73670, n73671, n73672, n73673, n73674, n73675,
    n73676, n73677, n73678, n73679, n73680, n73681, n73682, n73683, n73684,
    n73685, n73686, n73687, n73688, n73689, n73690, n73691, n73692, n73693,
    n73694, n73695, n73696, n73697, n73698, n73699, n73700, n73701, n73702,
    n73703, n73704, n73705, n73706, n73707, n73708, n73709, n73710, n73711,
    n73712, n73713, n73714, n73715, n73716, n73717, n73718, n73719, n73720,
    n73721, n73722, n73723, n73724, n73725, n73726, n73727, n73728, n73729,
    n73730, n73731, n73732, n73733, n73734, n73735, n73736, n73737, n73738,
    n73739, n73740, n73741, n73742, n73743, n73744, n73745, n73746, n73747,
    n73748, n73749, n73750, n73751, n73752, n73753, n73754, n73755, n73756,
    n73757, n73758, n73759, n73760, n73761, n73762, n73763, n73764, n73765,
    n73766, n73767, n73768, n73769, n73770, n73771, n73772, n73773, n73774,
    n73775, n73776, n73777, n73778, n73779, n73780, n73781, n73782, n73783,
    n73784, n73785, n73786, n73787, n73788, n73789, n73790, n73791, n73792,
    n73793, n73794, n73795, n73796, n73797, n73798, n73799, n73800, n73801,
    n73802, n73803, n73804, n73805, n73806, n73807, n73808, n73809, n73810,
    n73811, n73812, n73813, n73814, n73815, n73816, n73817, n73818, n73819,
    n73820, n73821, n73822, n73823, n73824, n73825, n73826, n73827, n73828,
    n73829, n73830, n73831, n73832, n73833, n73834, n73835, n73836, n73837,
    n73838, n73839, n73840, n73841, n73842, n73843, n73844, n73845, n73846,
    n73847, n73848, n73849, n73850, n73851, n73852, n73853, n73854, n73855,
    n73856, n73857, n73858, n73859, n73860, n73861, n73862, n73863, n73864,
    n73865, n73866, n73867, n73868, n73869, n73870, n73871, n73872, n73873,
    n73874, n73875, n73876, n73877, n73878, n73879, n73880, n73881, n73882,
    n73883, n73884, n73885, n73886, n73887, n73888, n73889, n73890, n73891,
    n73892, n73893, n73894, n73895, n73896, n73897, n73898, n73899, n73900,
    n73901, n73902, n73903, n73904, n73905, n73906, n73907, n73908, n73909,
    n73910, n73911, n73912, n73913, n73914, n73915, n73916, n73917, n73918,
    n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927,
    n73928, n73929, n73930, n73931, n73932, n73933, n73934, n73935, n73936,
    n73937, n73938, n73939, n73940, n73941, n73942, n73943, n73944, n73945,
    n73946, n73947, n73948, n73949, n73950, n73951, n73952, n73953, n73954,
    n73955, n73956, n73957, n73958, n73959, n73960, n73961, n73962, n73963,
    n73964, n73965, n73966, n73967, n73968, n73969, n73970, n73971, n73972,
    n73973, n73974, n73975, n73976, n73977, n73978, n73979, n73980, n73981,
    n73982, n73983, n73984, n73985, n73986, n73987, n73988, n73989, n73990,
    n73991, n73992, n73993, n73994, n73995, n73996, n73997, n73998, n73999,
    n74000, n74001, n74002, n74003, n74004, n74005, n74006, n74007, n74008,
    n74009, n74010, n74011, n74012, n74013, n74014, n74015, n74016, n74017,
    n74018, n74019, n74020, n74021, n74022, n74023, n74024, n74025, n74026,
    n74027, n74028, n74029, n74030, n74031, n74032, n74033, n74034, n74035,
    n74036, n74037, n74038, n74039, n74040, n74041, n74042, n74043, n74044,
    n74045, n74046, n74047, n74048, n74049, n74050, n74051, n74052, n74053,
    n74054, n74055, n74056, n74057, n74058, n74059, n74060, n74061, n74062,
    n74063, n74064, n74065, n74066, n74067, n74068, n74069, n74070, n74071,
    n74072, n74073, n74074, n74075, n74076, n74077, n74078, n74079, n74080,
    n74081, n74082, n74083, n74084, n74085, n74086, n74087, n74088, n74089,
    n74090, n74091, n74092, n74093, n74094, n74095, n74096, n74097, n74098,
    n74099, n74100, n74101, n74102, n74103, n74104, n74105, n74106, n74107,
    n74108, n74109, n74110, n74111, n74112, n74113, n74114, n74115, n74116,
    n74117, n74118, n74119, n74120, n74121, n74122, n74123, n74124, n74125,
    n74126, n74127, n74128, n74129, n74130, n74131, n74132, n74133, n74134,
    n74135, n74136, n74137, n74138, n74139, n74140, n74141, n74142, n74143,
    n74144, n74145, n74146, n74147, n74148, n74149, n74150, n74151, n74152,
    n74153, n74154, n74155, n74156, n74157, n74158, n74159, n74160, n74161,
    n74162, n74163, n74164, n74165, n74166, n74167, n74168, n74169, n74170,
    n74171, n74172, n74173, n74174, n74175, n74176, n74177, n74178, n74179,
    n74180, n74181, n74182, n74183, n74184, n74185, n74186, n74187, n74188,
    n74189, n74190, n74191, n74192, n74193, n74194, n74195, n74196, n74197,
    n74198, n74199, n74200, n74201, n74202, n74203, n74204, n74205, n74206,
    n74207, n74208, n74209, n74210, n74211, n74212, n74213, n74214, n74215,
    n74216, n74217, n74218, n74219, n74220, n74221, n74222, n74223, n74224,
    n74225, n74226, n74227, n74228, n74229, n74230, n74231, n74232, n74233,
    n74234, n74235, n74236, n74237, n74238, n74239, n74240, n74241, n74242,
    n74243, n74244, n74245, n74246, n74247, n74248, n74249, n74250, n74251,
    n74252, n74253, n74254, n74255, n74256, n74257, n74258, n74259, n74260,
    n74261, n74262, n74263, n74264, n74265, n74266, n74267, n74268, n74269,
    n74270, n74271, n74272, n74273, n74274, n74275, n74276, n74277, n74278,
    n74279, n74280, n74281, n74282, n74283, n74284, n74285, n74286, n74287,
    n74288, n74289, n74290, n74291, n74292, n74293, n74294, n74295, n74296,
    n74297, n74298, n74299, n74300, n74301, n74302, n74303, n74304, n74305,
    n74306, n74307, n74308, n74309, n74310, n74311, n74312, n74313, n74314,
    n74315, n74316, n74317, n74318, n74319, n74320, n74321, n74322, n74323,
    n74324, n74325, n74326, n74327, n74328, n74329, n74330, n74331, n74332,
    n74333, n74334, n74335, n74336, n74337, n74338, n74339, n74340, n74341,
    n74342, n74343, n74344, n74345, n74346, n74347, n74348, n74349, n74350,
    n74351, n74352, n74353, n74354, n74355, n74356, n74357, n74358, n74359,
    n74360, n74361, n74362, n74363, n74364, n74365, n74366, n74367, n74368,
    n74369, n74370, n74371, n74372, n74373, n74374, n74375, n74376, n74377,
    n74378, n74379, n74380, n74381, n74382, n74383, n74384, n74385, n74386,
    n74387, n74388, n74389, n74390, n74391, n74392, n74393, n74394, n74395,
    n74396, n74397, n74398, n74399, n74400, n74401, n74402, n74403, n74404,
    n74405, n74406, n74407, n74408, n74409, n74410, n74411, n74412, n74413,
    n74414, n74415, n74416, n74417, n74418, n74419, n74420, n74421, n74422,
    n74423, n74424, n74425, n74426, n74427, n74428, n74429, n74430, n74431,
    n74432, n74433, n74434, n74435, n74436, n74437, n74438, n74439, n74440,
    n74441, n74442, n74443, n74444, n74445, n74446, n74447, n74448, n74449,
    n74450, n74451, n74452, n74453, n74454, n74455, n74456, n74457, n74458,
    n74459, n74460, n74461, n74462, n74463, n74464, n74465, n74466, n74467,
    n74468, n74469, n74470, n74471, n74472, n74473, n74474, n74475, n74476,
    n74477, n74478, n74479, n74480, n74481, n74482, n74483, n74484, n74485,
    n74486, n74487, n74488, n74489, n74490, n74491, n74492, n74493, n74494,
    n74495, n74496, n74497, n74498, n74499, n74500, n74501, n74502, n74503,
    n74504, n74505, n74506, n74507, n74508, n74509, n74510, n74511, n74512,
    n74513, n74514, n74515, n74516, n74517, n74518, n74519, n74520, n74521,
    n74522, n74523, n74524, n74525, n74526, n74527, n74528, n74529, n74530,
    n74531, n74532, n74533, n74534, n74535, n74536, n74537, n74538, n74539,
    n74540, n74541, n74542, n74543, n74544, n74545, n74546, n74547, n74548,
    n74549, n74550, n74551, n74552, n74553, n74554, n74555, n74556, n74557,
    n74558, n74559, n74560, n74561, n74562, n74563, n74564, n74565, n74566,
    n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574, n74575,
    n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583, n74584,
    n74585, n74586, n74587, n74588, n74589, n74590, n74591, n74592, n74593,
    n74594, n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602,
    n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610, n74611,
    n74612, n74613, n74614, n74615, n74616, n74617, n74618, n74619, n74620,
    n74621, n74622, n74623, n74624, n74625, n74626, n74627, n74628, n74629,
    n74630, n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638,
    n74639, n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647,
    n74648, n74649, n74650, n74651, n74652, n74653, n74654, n74655, n74656,
    n74657, n74658, n74659, n74660, n74661, n74662, n74663, n74664, n74665,
    n74666, n74667, n74668, n74669, n74670, n74671, n74672, n74673, n74674,
    n74675, n74676, n74677, n74678, n74679, n74680, n74681, n74682, n74683,
    n74684, n74685, n74686, n74687, n74688, n74689, n74690, n74691, n74692,
    n74693, n74694, n74695, n74696, n74697, n74698, n74699, n74700, n74701,
    n74702, n74703, n74704, n74705, n74706, n74707, n74708, n74709, n74710,
    n74711, n74712, n74713, n74714, n74715, n74716, n74717, n74718, n74719,
    n74720, n74721, n74722, n74723, n74724, n74725, n74726, n74727, n74728,
    n74729, n74730, n74731, n74732, n74733, n74734, n74735, n74736, n74737,
    n74738, n74739, n74740, n74741, n74742, n74743, n74744, n74745, n74746,
    n74747, n74748, n74749, n74750, n74751, n74752, n74753, n74754, n74755,
    n74756, n74757, n74758, n74759, n74760, n74761, n74762, n74763, n74764,
    n74765, n74766, n74767, n74768, n74769, n74770, n74771, n74772, n74773,
    n74774, n74775, n74776, n74777, n74778, n74779, n74780, n74781, n74782,
    n74783, n74784, n74785, n74786, n74787, n74788, n74789, n74790, n74791,
    n74792, n74793, n74794, n74795, n74796, n74797, n74798, n74799, n74800,
    n74801, n74802, n74803, n74804, n74805, n74806, n74807, n74808, n74809,
    n74810, n74811, n74812, n74813, n74814, n74815, n74816, n74817, n74818,
    n74819, n74820, n74821, n74822, n74823, n74824, n74825, n74826, n74827,
    n74828, n74829, n74830, n74831, n74832, n74833, n74834, n74835, n74836,
    n74837, n74838, n74839, n74840, n74841, n74842, n74843, n74844, n74845,
    n74846, n74847, n74848, n74849, n74850, n74851, n74852, n74853, n74854,
    n74855, n74856, n74857, n74858, n74859, n74860, n74861, n74862, n74863,
    n74864, n74865, n74866, n74867, n74868, n74869, n74870, n74871, n74872,
    n74873, n74874, n74875, n74876, n74877, n74878, n74879, n74880, n74881,
    n74882, n74883, n74884, n74885, n74886, n74887, n74888, n74889, n74890,
    n74891, n74892, n74893, n74894, n74895, n74896, n74897, n74898, n74899,
    n74900, n74901, n74902, n74903, n74904, n74905, n74906, n74907, n74908,
    n74909, n74910, n74911, n74912, n74913, n74914, n74915, n74916, n74917,
    n74918, n74919, n74920, n74921, n74922, n74923, n74924, n74925, n74926,
    n74927, n74928, n74929, n74930, n74931, n74932, n74933, n74934, n74935,
    n74936, n74937, n74938, n74939, n74940, n74941, n74942, n74943, n74944,
    n74945, n74946, n74947, n74948, n74949, n74950, n74951, n74952, n74953,
    n74954, n74955, n74956, n74957, n74958, n74959, n74960, n74961, n74962,
    n74963, n74964, n74965, n74966, n74967, n74968, n74969, n74970, n74971,
    n74972, n74973, n74974, n74975, n74976, n74977, n74978, n74979, n74980,
    n74981, n74982, n74983, n74984, n74985, n74986, n74987, n74988, n74989,
    n74990, n74991, n74992, n74993, n74994, n74995, n74996, n74997, n74998,
    n74999, n75000, n75001, n75002, n75003, n75004, n75005, n75006, n75007,
    n75008, n75009, n75010, n75011, n75012, n75013, n75014, n75015, n75016,
    n75017, n75018, n75019, n75020, n75021, n75022, n75023, n75024, n75025,
    n75026, n75027, n75028, n75029, n75030, n75031, n75032, n75033, n75034,
    n75035, n75036, n75037, n75038, n75039, n75040, n75041, n75042, n75043,
    n75044, n75045, n75046, n75047, n75048, n75049, n75050, n75051, n75052,
    n75053, n75054, n75055, n75056, n75057, n75058, n75059, n75060, n75061,
    n75062, n75063, n75064, n75065, n75066, n75067, n75068, n75069, n75070,
    n75071, n75072, n75073, n75074, n75075, n75076, n75077, n75078, n75079,
    n75080, n75081, n75082, n75083, n75084, n75085, n75086, n75087, n75088,
    n75089, n75090, n75091, n75092, n75093, n75094, n75095, n75096, n75097,
    n75098, n75099, n75100, n75101, n75102, n75103, n75104, n75105, n75106,
    n75107, n75108, n75109, n75110, n75111, n75112, n75113, n75114, n75115,
    n75116, n75117, n75118, n75119, n75120, n75121, n75122, n75123, n75124,
    n75125, n75126, n75127, n75128, n75129, n75130, n75131, n75132, n75133,
    n75134, n75135, n75136, n75137, n75138, n75139, n75140, n75141, n75142,
    n75143, n75144, n75145, n75146, n75147, n75148, n75149, n75150, n75151,
    n75152, n75153, n75154, n75155, n75156, n75157, n75158, n75159, n75160,
    n75161, n75162, n75163, n75164, n75165, n75166, n75167, n75168, n75169,
    n75170, n75171, n75172, n75173, n75174, n75175, n75176, n75177, n75178,
    n75179, n75180, n75181, n75182, n75183, n75184, n75185, n75186, n75187,
    n75188, n75189, n75190, n75191, n75192, n75193, n75194, n75195, n75196,
    n75197, n75198, n75199, n75200, n75201, n75202, n75203, n75204, n75205,
    n75206, n75207, n75208, n75209, n75210, n75211, n75212, n75213, n75214,
    n75215, n75216, n75217, n75218, n75219, n75220, n75221, n75222, n75223,
    n75224, n75225, n75226, n75227, n75228, n75229, n75230, n75231, n75232,
    n75233, n75234, n75235, n75236, n75237, n75238, n75239, n75240, n75241,
    n75242, n75243, n75244, n75245, n75246, n75247, n75248, n75249, n75250,
    n75251, n75252, n75253, n75254, n75255, n75256, n75257, n75258, n75259,
    n75260, n75261, n75262, n75263, n75264, n75265, n75266, n75267, n75268,
    n75269, n75270, n75271, n75272, n75273, n75274, n75275, n75276, n75277,
    n75278, n75279, n75280, n75281, n75282, n75283, n75284, n75285, n75286,
    n75287, n75288, n75289, n75290, n75291, n75292, n75293, n75294, n75295,
    n75296, n75297, n75298, n75299, n75300, n75301, n75302, n75303, n75304,
    n75305, n75306, n75307, n75308, n75309, n75310, n75311, n75312, n75313,
    n75314, n75315, n75316, n75317, n75318, n75319, n75320, n75321, n75322,
    n75323, n75324, n75325, n75326, n75327, n75328, n75329, n75330, n75331,
    n75332, n75333, n75334, n75335, n75336, n75337, n75338, n75339, n75340,
    n75341, n75342, n75343, n75344, n75345, n75346, n75347, n75348, n75349,
    n75350, n75351, n75352, n75353, n75354, n75355, n75356, n75357, n75358,
    n75359, n75360, n75361, n75362, n75363, n75364, n75365, n75366, n75367,
    n75368, n75369, n75370, n75371, n75372, n75373, n75374, n75375, n75376,
    n75377, n75378, n75379, n75380, n75381, n75382, n75383, n75384, n75385,
    n75386, n75387, n75388, n75389, n75390, n75391, n75392, n75393, n75394,
    n75395, n75396, n75397, n75398, n75399, n75400, n75401, n75402, n75403,
    n75404, n75405, n75406, n75407, n75408, n75409, n75410, n75411, n75412,
    n75413, n75414, n75415, n75416, n75417, n75418, n75419, n75420, n75421,
    n75422, n75423, n75424, n75425, n75426, n75427, n75428, n75429, n75430,
    n75431, n75432, n75433, n75434, n75435, n75436, n75437, n75438, n75439,
    n75440, n75441, n75442, n75443, n75444, n75445, n75446, n75447, n75448,
    n75449, n75450, n75451, n75452, n75453, n75454, n75455, n75456, n75457,
    n75458, n75459, n75460, n75461, n75462, n75463, n75464, n75465, n75466,
    n75467, n75468, n75469, n75470, n75471, n75472, n75473, n75474, n75475,
    n75476, n75477, n75478, n75479, n75480, n75481, n75482, n75483, n75484,
    n75485, n75486, n75487, n75488, n75489, n75490, n75491, n75492, n75493,
    n75494, n75495, n75496, n75497, n75498, n75499, n75500, n75501, n75502,
    n75503, n75504, n75505, n75506, n75507, n75508, n75509, n75510, n75511,
    n75512, n75513, n75514, n75515, n75516, n75517, n75518, n75519, n75520,
    n75521, n75522, n75523, n75524, n75525, n75526, n75527, n75528, n75529,
    n75530, n75531, n75532, n75533, n75534, n75535, n75536, n75537, n75538,
    n75539, n75540, n75541, n75542, n75543, n75544, n75545, n75546, n75547,
    n75548, n75549, n75550, n75551, n75552, n75553, n75554, n75555, n75556,
    n75557, n75558, n75559, n75560, n75561, n75562, n75563, n75564, n75565,
    n75566, n75567, n75568, n75569, n75570, n75571, n75572, n75573, n75574,
    n75575, n75576, n75577, n75578, n75579, n75580, n75581, n75582, n75583,
    n75584, n75585, n75586, n75587, n75588, n75589, n75590, n75591, n75592,
    n75593, n75594, n75595, n75596, n75597, n75598, n75599, n75600, n75601,
    n75602, n75603, n75604, n75605, n75606, n75607, n75608, n75609, n75610,
    n75611, n75612, n75613, n75614, n75615, n75616, n75617, n75618, n75619,
    n75620, n75621, n75622, n75623, n75624, n75625, n75626, n75627, n75628,
    n75629, n75630, n75631, n75632, n75633, n75634, n75635, n75636, n75637,
    n75638, n75639, n75640, n75641, n75642, n75643, n75644, n75645, n75646,
    n75647, n75648, n75649, n75650, n75651, n75652, n75653, n75654, n75655,
    n75656, n75657, n75658, n75659, n75660, n75661, n75662, n75663, n75664,
    n75665, n75666, n75667, n75668, n75669, n75670, n75671, n75672, n75673,
    n75674, n75675, n75676, n75677, n75678, n75679, n75680, n75681, n75682,
    n75683, n75684, n75685, n75686, n75687, n75688, n75689, n75690, n75691,
    n75692, n75693, n75694, n75695, n75696, n75697, n75698, n75699, n75700,
    n75701, n75702, n75703, n75704, n75705, n75706, n75707, n75708, n75709,
    n75710, n75711, n75712, n75713, n75714, n75715, n75716, n75717, n75718,
    n75719, n75720, n75721, n75722, n75723, n75724, n75725, n75726, n75727,
    n75728, n75729, n75730, n75731, n75732, n75733, n75734, n75735, n75736,
    n75737, n75738, n75739, n75740, n75741, n75742, n75743, n75744, n75745,
    n75746, n75747, n75748, n75749, n75750, n75751, n75752, n75753, n75754,
    n75755, n75756, n75757, n75758, n75759, n75760, n75761, n75762, n75763,
    n75764, n75765, n75766, n75767, n75768, n75769, n75770, n75771, n75772,
    n75773, n75774, n75775, n75776, n75777, n75778, n75779, n75780, n75781,
    n75782, n75783, n75784, n75785, n75786, n75787, n75788, n75789, n75790,
    n75791, n75792, n75793, n75794, n75795, n75796, n75797, n75798, n75799,
    n75800, n75801, n75802, n75803, n75804, n75805, n75806, n75807, n75808,
    n75809, n75810, n75811, n75812, n75813, n75814, n75815, n75816, n75817,
    n75818, n75819, n75820, n75821, n75822, n75823, n75824, n75825, n75826,
    n75827, n75828, n75829, n75830, n75831, n75832, n75833, n75834, n75835,
    n75836, n75837, n75838, n75839, n75840, n75841, n75842, n75843, n75844,
    n75845, n75846, n75847, n75848, n75849, n75850, n75851, n75852, n75853,
    n75854, n75855, n75856, n75857, n75858, n75859, n75860, n75861, n75862,
    n75863, n75864, n75865, n75866, n75867, n75868, n75869, n75870, n75871,
    n75872, n75873, n75874, n75875, n75876, n75877, n75878, n75879, n75880,
    n75881, n75882, n75883, n75884, n75885, n75886, n75887, n75888, n75889,
    n75890, n75891, n75892, n75893, n75894, n75895, n75896, n75897, n75898,
    n75899, n75900, n75901, n75902, n75903, n75904, n75905, n75906, n75907,
    n75908, n75909, n75910, n75911, n75912, n75913, n75914, n75915, n75916,
    n75917, n75918, n75919, n75920, n75921, n75922, n75923, n75924, n75925,
    n75926, n75927, n75928, n75929, n75930, n75931, n75932, n75933, n75934,
    n75935, n75936, n75937, n75938, n75939, n75940, n75941, n75942, n75943,
    n75944, n75945, n75946, n75947, n75948, n75949, n75950, n75951, n75952,
    n75953, n75954, n75955, n75956, n75957, n75958, n75959, n75960, n75961,
    n75962, n75963, n75964, n75965, n75966, n75967, n75968, n75969, n75970,
    n75971, n75972, n75973, n75974, n75975, n75976, n75977, n75978, n75979,
    n75980, n75981, n75982, n75983, n75984, n75985, n75986, n75987, n75988,
    n75989, n75990, n75991, n75992, n75993, n75994, n75995, n75996, n75997,
    n75998, n75999, n76000, n76001, n76002, n76003, n76004, n76005, n76006,
    n76007, n76008, n76009, n76010, n76011, n76012, n76013, n76014, n76015,
    n76016, n76017, n76018, n76019, n76020, n76021, n76022, n76023, n76024,
    n76025, n76026, n76027, n76028, n76029, n76030, n76031, n76032, n76033,
    n76034, n76035, n76036, n76037, n76038, n76039, n76040, n76041, n76042,
    n76043, n76044, n76045, n76046, n76047, n76048, n76049, n76050, n76051,
    n76052, n76053, n76054, n76055, n76056, n76057, n76058, n76059, n76060,
    n76061, n76062, n76063, n76064, n76065, n76066, n76067, n76068, n76069,
    n76070, n76071, n76072, n76073, n76074, n76075, n76076, n76077, n76078,
    n76079, n76080, n76081, n76082, n76083, n76084, n76085, n76086, n76087,
    n76088, n76089, n76090, n76091, n76092, n76093, n76094, n76095, n76096,
    n76097, n76098, n76099, n76100, n76101, n76102, n76103, n76104, n76105,
    n76106, n76107, n76108, n76109, n76110, n76111, n76112, n76113, n76114,
    n76115, n76116, n76117, n76118, n76119, n76120, n76121, n76122, n76123,
    n76124, n76125, n76126, n76127, n76128, n76129, n76130, n76131, n76132,
    n76133, n76134, n76135, n76136, n76137, n76138, n76139, n76140, n76141,
    n76142, n76143, n76144, n76145, n76146, n76147, n76148, n76149, n76150,
    n76151, n76152, n76153, n76154, n76155, n76156, n76157, n76158, n76159,
    n76160, n76161, n76162, n76163, n76164, n76165, n76166, n76167, n76168,
    n76169, n76170, n76171, n76172, n76173, n76174, n76175, n76176, n76177,
    n76178, n76179, n76180, n76181, n76182, n76183, n76184, n76185, n76186,
    n76187, n76188, n76189, n76190, n76191, n76192, n76193, n76194, n76195,
    n76196, n76197, n76198, n76199, n76200, n76201, n76202, n76203, n76204,
    n76205, n76206, n76207, n76208, n76209, n76210, n76211, n76212, n76213,
    n76214, n76215, n76216, n76217, n76218, n76219, n76220, n76221, n76222,
    n76223, n76224, n76225, n76226, n76227, n76228, n76229, n76230, n76231,
    n76232, n76233, n76234, n76235, n76236, n76237, n76238, n76239, n76240,
    n76241, n76242, n76243, n76244, n76245, n76246, n76247, n76248, n76249,
    n76250, n76251, n76252, n76253, n76254, n76255, n76256, n76257, n76258,
    n76259, n76260, n76261, n76262, n76263, n76264, n76265, n76266, n76267,
    n76268, n76269, n76270, n76271, n76272, n76273, n76274, n76275, n76276,
    n76277, n76278, n76279, n76280, n76281, n76282, n76283, n76284, n76285,
    n76286, n76287, n76288, n76289, n76290, n76291, n76292, n76293, n76294,
    n76295, n76296, n76297, n76298, n76299, n76300, n76301, n76302, n76303,
    n76304, n76305, n76306, n76307, n76308, n76309, n76310, n76311, n76312,
    n76313, n76314, n76315, n76316, n76317, n76318, n76319, n76320, n76321,
    n76322, n76323, n76324, n76325, n76326, n76327, n76328, n76329, n76330,
    n76331, n76332, n76333, n76334, n76335, n76336, n76337, n76338, n76339,
    n76340, n76341, n76342, n76343, n76344, n76345, n76346, n76347, n76348,
    n76349, n76350, n76351, n76352, n76353, n76354, n76355, n76356, n76357,
    n76358, n76359, n76360, n76361, n76362, n76363, n76364, n76365, n76366,
    n76367, n76368, n76369, n76370, n76371, n76372, n76373, n76374, n76375,
    n76376, n76377, n76378, n76379, n76380, n76381, n76382, n76383, n76384,
    n76385, n76386, n76387, n76388, n76389, n76390, n76391, n76392, n76393,
    n76394, n76395, n76396, n76397, n76398, n76399, n76400, n76401, n76402,
    n76403, n76404, n76405, n76406, n76407, n76408, n76409, n76410, n76411,
    n76412, n76413, n76414, n76415, n76416, n76417, n76418, n76419, n76420,
    n76421, n76422, n76423, n76424, n76425, n76426, n76427, n76428, n76429,
    n76430, n76431, n76432, n76433, n76434, n76435, n76436, n76437, n76438,
    n76439, n76440, n76441, n76442, n76443, n76444, n76445, n76446, n76447,
    n76448, n76449, n76450, n76451, n76452, n76453, n76454, n76455, n76456,
    n76457, n76458, n76459, n76460, n76461, n76462, n76463, n76464, n76465,
    n76466, n76467, n76468, n76469, n76470, n76471, n76472, n76473, n76474,
    n76475, n76476, n76477, n76478, n76479, n76480, n76481, n76482, n76483,
    n76484, n76485, n76486, n76487, n76488, n76489, n76490, n76491, n76492,
    n76493, n76494, n76495, n76496, n76497, n76498, n76499, n76500, n76501,
    n76502, n76503, n76504, n76505, n76506, n76507, n76508, n76509, n76510,
    n76511, n76512, n76513, n76514, n76515, n76516, n76517, n76518, n76519,
    n76520, n76521, n76522, n76523, n76524, n76525, n76526, n76527, n76528,
    n76529, n76530, n76531, n76532, n76533, n76534, n76535, n76536, n76537,
    n76538, n76539, n76540, n76541, n76542, n76543, n76544, n76545, n76546,
    n76547, n76548, n76549, n76550, n76551, n76552, n76553, n76554, n76555,
    n76556, n76557, n76558, n76559, n76560, n76561, n76562, n76563, n76564,
    n76565, n76566, n76567, n76568, n76569, n76570, n76571, n76572, n76573,
    n76574, n76575, n76576, n76577, n76578, n76579, n76580, n76581, n76582,
    n76583, n76584, n76585, n76586, n76587, n76588, n76589, n76590, n76591,
    n76592, n76593, n76594, n76595, n76596, n76597, n76598, n76599, n76600,
    n76601, n76602, n76603, n76604, n76605, n76606, n76607, n76608, n76609,
    n76610, n76611, n76612, n76613, n76614, n76615, n76616, n76617, n76618,
    n76619, n76620, n76621, n76622, n76623, n76624, n76625, n76626, n76627,
    n76628, n76629, n76630, n76631, n76632, n76633, n76634, n76635, n76636,
    n76637, n76638, n76639, n76640, n76641, n76642, n76643, n76644, n76645,
    n76646, n76647, n76648, n76649, n76650, n76651, n76652, n76653, n76654,
    n76655, n76656, n76657, n76658, n76659, n76660, n76661, n76662, n76663,
    n76664, n76665, n76666, n76667, n76668, n76669, n76670, n76671, n76672,
    n76673, n76674, n76675, n76676, n76677, n76678, n76679, n76680, n76681,
    n76682, n76683, n76684, n76685, n76686, n76687, n76688, n76689, n76690,
    n76691, n76692, n76693, n76694, n76695, n76696, n76697, n76698, n76699,
    n76700, n76701, n76702, n76703, n76704, n76705, n76706, n76707, n76708,
    n76709, n76710, n76711, n76712, n76713, n76714, n76715, n76716, n76717,
    n76718, n76719, n76720, n76721, n76722, n76723, n76724, n76725, n76726,
    n76727, n76728, n76729, n76730, n76731, n76732, n76733, n76734, n76735,
    n76736, n76737, n76738, n76739, n76740, n76741, n76742, n76743, n76744,
    n76745, n76746, n76747, n76748, n76749, n76750, n76751, n76752, n76753,
    n76754, n76755, n76756, n76757, n76758, n76759, n76760, n76761, n76762,
    n76763, n76764, n76765, n76766, n76767, n76768, n76769, n76770, n76771,
    n76772, n76773, n76774, n76775, n76776, n76777, n76778, n76779, n76780,
    n76781, n76782, n76783, n76784, n76785, n76786, n76787, n76788, n76789,
    n76790, n76791, n76792, n76793, n76794, n76795, n76796, n76797, n76798,
    n76799, n76800, n76801, n76802, n76803, n76804, n76805, n76806, n76807,
    n76808, n76809, n76810, n76811, n76812, n76813, n76814, n76815, n76816,
    n76817, n76818, n76819, n76820, n76821, n76822, n76823, n76824, n76825,
    n76826, n76827, n76828, n76829, n76830, n76831, n76832, n76833, n76834,
    n76835, n76836, n76837, n76838, n76839, n76840, n76841, n76842, n76843,
    n76844, n76845, n76846, n76847, n76848, n76849, n76850, n76851, n76852,
    n76853, n76854, n76855, n76856, n76857, n76858, n76859, n76860, n76861,
    n76862, n76863, n76864, n76865, n76866, n76867, n76868, n76869, n76870,
    n76871, n76872, n76873, n76874, n76875, n76876, n76877, n76878, n76879,
    n76880, n76881, n76882, n76883, n76884, n76885, n76886, n76887, n76888,
    n76889, n76890, n76891, n76892, n76893, n76894, n76895, n76896, n76897,
    n76898, n76899, n76900, n76901, n76902, n76903, n76904, n76905, n76906,
    n76907, n76908, n76909, n76910, n76911, n76912, n76913, n76914, n76915,
    n76916, n76917, n76918, n76919, n76920, n76921, n76922, n76923, n76924,
    n76925, n76926, n76927, n76928, n76929, n76930, n76931, n76932, n76933,
    n76934, n76935, n76936, n76937, n76938, n76939, n76940, n76941, n76942,
    n76943, n76944, n76945, n76946, n76947, n76948, n76949, n76950, n76951,
    n76952, n76953, n76954, n76955, n76956, n76957, n76958, n76959, n76960,
    n76961, n76962, n76963, n76964, n76965, n76966, n76967, n76968, n76969,
    n76970, n76971, n76972, n76973, n76974, n76975, n76976, n76977, n76978,
    n76979, n76980, n76981, n76982, n76983, n76984, n76985, n76986, n76987,
    n76988, n76989, n76990, n76991, n76992, n76993, n76994, n76995, n76996,
    n76997, n76998, n76999, n77000, n77001, n77002, n77003, n77004, n77005,
    n77006, n77007, n77008, n77009, n77010, n77011, n77012, n77013, n77014,
    n77015, n77016, n77017, n77018, n77019, n77020, n77021, n77022, n77023,
    n77024, n77025, n77026, n77027, n77028, n77029, n77030, n77031, n77032,
    n77033, n77034, n77035, n77036, n77037, n77038, n77039, n77040, n77041,
    n77042, n77043, n77044, n77045, n77046, n77047, n77048, n77049, n77050,
    n77051, n77052, n77053, n77054, n77055, n77056, n77057, n77058, n77059,
    n77060, n77061, n77062, n77063, n77064, n77065, n77066, n77067, n77068,
    n77069, n77070, n77071, n77072, n77073, n77074, n77075, n77076, n77077,
    n77078, n77079, n77080, n77081, n77082, n77083, n77084, n77085, n77086,
    n77087, n77088, n77089, n77090, n77091, n77092, n77093, n77094, n77095,
    n77096, n77097, n77098, n77099, n77100, n77101, n77102, n77103, n77104,
    n77105, n77106, n77107, n77108, n77109, n77110, n77111, n77112, n77113,
    n77114, n77115, n77116, n77117, n77118, n77119, n77120, n77121, n77122,
    n77123, n77124, n77125, n77126, n77127, n77128, n77129, n77130, n77131,
    n77132, n77133, n77134, n77135, n77136, n77137, n77138, n77139, n77140,
    n77141, n77142, n77143, n77144, n77145, n77146, n77147, n77148, n77149,
    n77150, n77151, n77152, n77153, n77154, n77155, n77156, n77157, n77158,
    n77159, n77160, n77161, n77162, n77163, n77164, n77165, n77166, n77167,
    n77168, n77169, n77170, n77171, n77172, n77173, n77174, n77175, n77176,
    n77177, n77178, n77179, n77180, n77181, n77182, n77183, n77184, n77185,
    n77186, n77187, n77188, n77189, n77190, n77191, n77192, n77193, n77194,
    n77195, n77196, n77197, n77198, n77199, n77200, n77201, n77202, n77203,
    n77204, n77205, n77206, n77207, n77208, n77209, n77210, n77211, n77212,
    n77213, n77214, n77215, n77216, n77217, n77218, n77219, n77220, n77221,
    n77222, n77223, n77224, n77225, n77226, n77227, n77228, n77229, n77230,
    n77231, n77232, n77233, n77234, n77235, n77236, n77237, n77238, n77239,
    n77240, n77241, n77242, n77243, n77244, n77245, n77246, n77247, n77248,
    n77249, n77250, n77251, n77252, n77253, n77254, n77255, n77256, n77257,
    n77258, n77259, n77260, n77261, n77262, n77263, n77264, n77265, n77266,
    n77267, n77268, n77269, n77270, n77271, n77272, n77273, n77274, n77275,
    n77276, n77277, n77278, n77279, n77280, n77281, n77282, n77283, n77284,
    n77285, n77286, n77287, n77288, n77289, n77290, n77291, n77292, n77293,
    n77294, n77295, n77296, n77297, n77298, n77299, n77300, n77301, n77302,
    n77303, n77304, n77305, n77306, n77307, n77308, n77309, n77310, n77311,
    n77312, n77313, n77314, n77315, n77316, n77317, n77318, n77319, n77320,
    n77321, n77322, n77323, n77324, n77325, n77326, n77327, n77328, n77329,
    n77330, n77331, n77332, n77333, n77334, n77335, n77336, n77337, n77338,
    n77339, n77340, n77341, n77342, n77343, n77344, n77345, n77346, n77347,
    n77348, n77349, n77350, n77351, n77352, n77353, n77354, n77355, n77356,
    n77357, n77358, n77359, n77360, n77361, n77362, n77363, n77364, n77365,
    n77366, n77367, n77368, n77369, n77370, n77371, n77372, n77373, n77374,
    n77375, n77376, n77377, n77378, n77379, n77380, n77381, n77382, n77383,
    n77384, n77385, n77386, n77387, n77388, n77389, n77390, n77391, n77392,
    n77393, n77394, n77395, n77396, n77397, n77398, n77399, n77400, n77401,
    n77402, n77403, n77404, n77405, n77406, n77407, n77408, n77409, n77410,
    n77411, n77412, n77413, n77414, n77415, n77416, n77417, n77418, n77419,
    n77420, n77421, n77422, n77423, n77424, n77425, n77426, n77427, n77428,
    n77429, n77430, n77431, n77432, n77433, n77434, n77435, n77436, n77437,
    n77438, n77439, n77440, n77441, n77442, n77443, n77444, n77445, n77446,
    n77447, n77448, n77449, n77450, n77451, n77452, n77453, n77454, n77455,
    n77456, n77457, n77458, n77459, n77460, n77461, n77462, n77463, n77464,
    n77465, n77466, n77467, n77468, n77469, n77470, n77471, n77472, n77473,
    n77474, n77475, n77476, n77477, n77478, n77479, n77480, n77481, n77482,
    n77483, n77484, n77485, n77486, n77487, n77488, n77489, n77490, n77491,
    n77492, n77493, n77494, n77495, n77496, n77497, n77498, n77499, n77500,
    n77501, n77502, n77503, n77504, n77505, n77506, n77507, n77508, n77509,
    n77510, n77511, n77512, n77513, n77514, n77515, n77516, n77517, n77518,
    n77519, n77520, n77521, n77522, n77523, n77524, n77525, n77526, n77527,
    n77528, n77529, n77530, n77531, n77532, n77533, n77534, n77535, n77536,
    n77537, n77538, n77539, n77540, n77541, n77542, n77543, n77544, n77545,
    n77546, n77547, n77548, n77549, n77550, n77551, n77552, n77553, n77554,
    n77555, n77556, n77557, n77558, n77559, n77560, n77561, n77562, n77563,
    n77564, n77565, n77566, n77567, n77568, n77569, n77570, n77571, n77572,
    n77573, n77574, n77575, n77576, n77577, n77578, n77579, n77580, n77581,
    n77582, n77583, n77584, n77585, n77586, n77587, n77588, n77589, n77590,
    n77591, n77592, n77593, n77594, n77595, n77596, n77597, n77598, n77599,
    n77600, n77601, n77602, n77603, n77604, n77605, n77606, n77607, n77608,
    n77609, n77610, n77611, n77612, n77613, n77614, n77615, n77616, n77617,
    n77618, n77619, n77620, n77621, n77622, n77623, n77624, n77625, n77626,
    n77627, n77628, n77629, n77630, n77631, n77632, n77633, n77634, n77635,
    n77636, n77637, n77638, n77639, n77640, n77641, n77642, n77643, n77644,
    n77645, n77646, n77647, n77648, n77649, n77650, n77651, n77652, n77653,
    n77654, n77655, n77656, n77657, n77658, n77659, n77660, n77661, n77662,
    n77663, n77664, n77665, n77666, n77667, n77668, n77669, n77670, n77671,
    n77672, n77673, n77674, n77675, n77676, n77677, n77678, n77679, n77680,
    n77681, n77682, n77683, n77684, n77685, n77686, n77687, n77688, n77689,
    n77690, n77691, n77692, n77693, n77694, n77695, n77696, n77697, n77698,
    n77699, n77700, n77701, n77702, n77703, n77704, n77705, n77706, n77707,
    n77708, n77709, n77710, n77711, n77712, n77713, n77714, n77715, n77716,
    n77717, n77718, n77719, n77720, n77721, n77722, n77723, n77724, n77725,
    n77726, n77727, n77728, n77729, n77730, n77731, n77732, n77733, n77734,
    n77735, n77736, n77737, n77738, n77739, n77740, n77741, n77742, n77743,
    n77744, n77745, n77746, n77747, n77748, n77749, n77750, n77751, n77752,
    n77753, n77754, n77755, n77756, n77757, n77758, n77759, n77760, n77761,
    n77762, n77763, n77764, n77765, n77766, n77767, n77768, n77769, n77770,
    n77771, n77772, n77773, n77774, n77775, n77776, n77777, n77778, n77779,
    n77780, n77781, n77782, n77783, n77784, n77785, n77786, n77787, n77788,
    n77789, n77790, n77791, n77792, n77793, n77794, n77795, n77796, n77797,
    n77798, n77799, n77800, n77801, n77802, n77803, n77804, n77805, n77806,
    n77807, n77808, n77809, n77810, n77811, n77812, n77813, n77814, n77815,
    n77816, n77817, n77818, n77819, n77820, n77821, n77822, n77823, n77824,
    n77825, n77826, n77827, n77828, n77829, n77830, n77831, n77832, n77833,
    n77834, n77835, n77836, n77837, n77838, n77839, n77840, n77841, n77842,
    n77843, n77844, n77845, n77846, n77847, n77848, n77849, n77850, n77851,
    n77852, n77853, n77854, n77855, n77856, n77857, n77858, n77859, n77860,
    n77861, n77862, n77863, n77864, n77865, n77866, n77867, n77868, n77869,
    n77870, n77871, n77872, n77873, n77874, n77875, n77876, n77877, n77878,
    n77879, n77880, n77881, n77882, n77883, n77884, n77885, n77886, n77887,
    n77888, n77889, n77890, n77891, n77892, n77893, n77894, n77895, n77896,
    n77897, n77898, n77899, n77900, n77901, n77902, n77903, n77904, n77905,
    n77906, n77907, n77908, n77909, n77910, n77911, n77912, n77913, n77914,
    n77915, n77916, n77917, n77918, n77919, n77920, n77921, n77922, n77923,
    n77924, n77925, n77926, n77927, n77928, n77929, n77930, n77931, n77932,
    n77933, n77934, n77935, n77936, n77937, n77938, n77939, n77940, n77941,
    n77942, n77943, n77944, n77945, n77946, n77947, n77948, n77949, n77950,
    n77951, n77952, n77953, n77954, n77955, n77956, n77957, n77958, n77959,
    n77960, n77961, n77962, n77963, n77964, n77965, n77966, n77967, n77968,
    n77969, n77970, n77971, n77972, n77973, n77974, n77975, n77976, n77977,
    n77978, n77979, n77980, n77981, n77982, n77983, n77984, n77985, n77986,
    n77987, n77988, n77989, n77990, n77991, n77992, n77993, n77994, n77995,
    n77996, n77997, n77998, n77999, n78000, n78001, n78002, n78003, n78004,
    n78005, n78006, n78007, n78008, n78009, n78010, n78011, n78012, n78013,
    n78014, n78015, n78016, n78017, n78018, n78019, n78020, n78021, n78022,
    n78023, n78024, n78025, n78026, n78027, n78028, n78029, n78030, n78031,
    n78032, n78033, n78034, n78035, n78036, n78037, n78038, n78039, n78040,
    n78041, n78042, n78043, n78044, n78045, n78046, n78047, n78048, n78049,
    n78050, n78051, n78052, n78053, n78054, n78055, n78056, n78057, n78058,
    n78059, n78060, n78061, n78062, n78063, n78064, n78065, n78066, n78067,
    n78068, n78069, n78070, n78071, n78072, n78073, n78074, n78075, n78076,
    n78077, n78078, n78079, n78080, n78081, n78082, n78083, n78084, n78085,
    n78086, n78087, n78088, n78089, n78090, n78091, n78092, n78093, n78094,
    n78095, n78096, n78097, n78098, n78099, n78100, n78101, n78102, n78103,
    n78104, n78105, n78106, n78107, n78108, n78109, n78110, n78111, n78112,
    n78113, n78114, n78115, n78116, n78117, n78118, n78119, n78120, n78121,
    n78122, n78123, n78124, n78125, n78126, n78127, n78128, n78129, n78130,
    n78131, n78132, n78133, n78134, n78135, n78136, n78137, n78138, n78139,
    n78140, n78141, n78142, n78143, n78144, n78145, n78146, n78147, n78148,
    n78149, n78150, n78151, n78152, n78153, n78154, n78155, n78156, n78157,
    n78158, n78159, n78160, n78161, n78162, n78163, n78164, n78165, n78166,
    n78167, n78168, n78169, n78170, n78171, n78172, n78173, n78174, n78175,
    n78176, n78177, n78178, n78179, n78180, n78181, n78182, n78183, n78184,
    n78185, n78186, n78187, n78188, n78189, n78190, n78191, n78192, n78193,
    n78194, n78195, n78196, n78197, n78198, n78199, n78200, n78201, n78202,
    n78203, n78204, n78205, n78206, n78207, n78208, n78209, n78210, n78211,
    n78212, n78213, n78214, n78215, n78216, n78217, n78218, n78219, n78220,
    n78221, n78222, n78223, n78224, n78225, n78226, n78227, n78228, n78229,
    n78230, n78231, n78232, n78233, n78234, n78235, n78236, n78237, n78238,
    n78239, n78240, n78241, n78242, n78243, n78244, n78245, n78246, n78247,
    n78248, n78249, n78250, n78251, n78252, n78253, n78254, n78255, n78256,
    n78257, n78258, n78259, n78260, n78261, n78262, n78263, n78264, n78265,
    n78266, n78267, n78268, n78269, n78270, n78271, n78272, n78273, n78274,
    n78275, n78276, n78277, n78278, n78279, n78280, n78281, n78282, n78283,
    n78284, n78285, n78286, n78287, n78288, n78289, n78290, n78291, n78292,
    n78293, n78294, n78295, n78296, n78297, n78298, n78299, n78300, n78301,
    n78302, n78303, n78304, n78305, n78306, n78307, n78308, n78309, n78310,
    n78311, n78312, n78313, n78314, n78315, n78316, n78317, n78318, n78319,
    n78320, n78321, n78322, n78323, n78324, n78325, n78326, n78327, n78328,
    n78329, n78330, n78331, n78332, n78333, n78334, n78335, n78336, n78337,
    n78338, n78339, n78340, n78341, n78342, n78343, n78344, n78345, n78346,
    n78347, n78348, n78349, n78350, n78351, n78352, n78353, n78354, n78355,
    n78356, n78357, n78358, n78359, n78360, n78361, n78362, n78363, n78364,
    n78365, n78366, n78367, n78368, n78369, n78370, n78371, n78372, n78373,
    n78374, n78375, n78376, n78377, n78378, n78379, n78380, n78381, n78382,
    n78383, n78384, n78385, n78386, n78387, n78388, n78389, n78390, n78391,
    n78392, n78393, n78394, n78395, n78396, n78397, n78398, n78399, n78400,
    n78401, n78402, n78403, n78404, n78405, n78406, n78407, n78408, n78409,
    n78410, n78411, n78412, n78413, n78414, n78415, n78416, n78417, n78418,
    n78419, n78420, n78421, n78422, n78423, n78424, n78425, n78426, n78427,
    n78428, n78429, n78430, n78431, n78432, n78433, n78434, n78435, n78436,
    n78437, n78438, n78439, n78440, n78441, n78442, n78443, n78444, n78445,
    n78446, n78447, n78448, n78449, n78450, n78451, n78452, n78453, n78454,
    n78455, n78456, n78457, n78458, n78459, n78460, n78461, n78462, n78463,
    n78464, n78465, n78466, n78467, n78468, n78469, n78470, n78471, n78472,
    n78473, n78474, n78475, n78476, n78477, n78478, n78479, n78480, n78481,
    n78482, n78483, n78484, n78485, n78486, n78487, n78488, n78489, n78490,
    n78491, n78492, n78493, n78494, n78495, n78496, n78497, n78498, n78499,
    n78500, n78501, n78502, n78503, n78504, n78505, n78506, n78507, n78508,
    n78509, n78510, n78511, n78512, n78513, n78514, n78515, n78516, n78517,
    n78518, n78519, n78520, n78521, n78522, n78523, n78524, n78525, n78526,
    n78527, n78528, n78529, n78530, n78531, n78532, n78533, n78534, n78535,
    n78536, n78537, n78538, n78539, n78540, n78541, n78542, n78543, n78544,
    n78545, n78546, n78547, n78548, n78549, n78550, n78551, n78552, n78553,
    n78554, n78555, n78556, n78557, n78558, n78559, n78560, n78561, n78562,
    n78563, n78564, n78565, n78566, n78567, n78568, n78569, n78570, n78571,
    n78572, n78573, n78574, n78575, n78576, n78577, n78578, n78579, n78580,
    n78581, n78582, n78583, n78584, n78585, n78586, n78587, n78588, n78589,
    n78590, n78591, n78592, n78593, n78594, n78595, n78596, n78597, n78598,
    n78599, n78600, n78601, n78602, n78603, n78604, n78605, n78606, n78607,
    n78608, n78609, n78610, n78611, n78612, n78613, n78614, n78615, n78616,
    n78617, n78618, n78619, n78620, n78621, n78622, n78623, n78624, n78625,
    n78626, n78627, n78628, n78629, n78630, n78631, n78632, n78633, n78634,
    n78635, n78636, n78637, n78638, n78639, n78640, n78641, n78642, n78643,
    n78644, n78645, n78646, n78647, n78648, n78649, n78650, n78651, n78652,
    n78653, n78654, n78655, n78656, n78657, n78658, n78659, n78660, n78661,
    n78662, n78663, n78664, n78665, n78666, n78667, n78668, n78669, n78670,
    n78671, n78672, n78673, n78674, n78675, n78676, n78677, n78678, n78679,
    n78680, n78681, n78682, n78683, n78684, n78685, n78686, n78687, n78688,
    n78689, n78690, n78691, n78692, n78693, n78694, n78695, n78696, n78697,
    n78698, n78699, n78700, n78701, n78702, n78703, n78704, n78705, n78706,
    n78707, n78708, n78709, n78710, n78711, n78712, n78713, n78714, n78715,
    n78716, n78717, n78718, n78719, n78720, n78721, n78722, n78723, n78724,
    n78725, n78726, n78727, n78728, n78729, n78730, n78731, n78732, n78733,
    n78734, n78735, n78736, n78737, n78738, n78739, n78740, n78741, n78742,
    n78743, n78744, n78745, n78746, n78747, n78748, n78749, n78750, n78751,
    n78752, n78753, n78754, n78755, n78756, n78757, n78758, n78759, n78760,
    n78761, n78762, n78763, n78764, n78765, n78766, n78767, n78768, n78769,
    n78770, n78771, n78772, n78773, n78774, n78775, n78776, n78777, n78778,
    n78779, n78780, n78781, n78782, n78783, n78784, n78785, n78786, n78787,
    n78788, n78789, n78790, n78791, n78792, n78793, n78794, n78795, n78796,
    n78797, n78798, n78799, n78800, n78801, n78802, n78803, n78804, n78805,
    n78806, n78807, n78808, n78809, n78810, n78811, n78812, n78813, n78814,
    n78815, n78816, n78817, n78818, n78819, n78820, n78821, n78822, n78823,
    n78824, n78825, n78826, n78827, n78828, n78829, n78830, n78831, n78832,
    n78833, n78834, n78835, n78836, n78837, n78838, n78839, n78840, n78841,
    n78842, n78843, n78844, n78845, n78846, n78847, n78848, n78849, n78850,
    n78851, n78852, n78853, n78854, n78855, n78856, n78857, n78858, n78859,
    n78860, n78861, n78862, n78863, n78864, n78865, n78866, n78867, n78868,
    n78869, n78870, n78871, n78872, n78873, n78874, n78875, n78876, n78877,
    n78878, n78879, n78880, n78881, n78882, n78883, n78884, n78885, n78886,
    n78887, n78888, n78889, n78890, n78891, n78892, n78893, n78894, n78895,
    n78896, n78897, n78898, n78899, n78900, n78901, n78902, n78903, n78904,
    n78905, n78906, n78907, n78908, n78909, n78910, n78911, n78912, n78913,
    n78914, n78915, n78916, n78917, n78918, n78919, n78920, n78921, n78922,
    n78923, n78924, n78925, n78926, n78927, n78928, n78929, n78930, n78931,
    n78932, n78933, n78934, n78935, n78936, n78937, n78938, n78939, n78940,
    n78941, n78942, n78943, n78944, n78945, n78946, n78947, n78948, n78949,
    n78950, n78951, n78952, n78953, n78954, n78955, n78956, n78957, n78958,
    n78959, n78960, n78961, n78962, n78963, n78964, n78965, n78966, n78967,
    n78968, n78969, n78970, n78971, n78972, n78973, n78974, n78975, n78976,
    n78977, n78978, n78979, n78980, n78981, n78982, n78983, n78984, n78985,
    n78986, n78987, n78988, n78989, n78990, n78991, n78992, n78993, n78994,
    n78995, n78996, n78997, n78998, n78999, n79000, n79001, n79002, n79003,
    n79004, n79005, n79006, n79007, n79008, n79009, n79010, n79011, n79012,
    n79013, n79014, n79015, n79016, n79017, n79018, n79019, n79020, n79021,
    n79022, n79023, n79024, n79025, n79026, n79027, n79028, n79029, n79030,
    n79031, n79032, n79033, n79034, n79035, n79036, n79037, n79038, n79039,
    n79040, n79041, n79042, n79043, n79044, n79045, n79046, n79047, n79048,
    n79049, n79050, n79051, n79052, n79053, n79054, n79055, n79056, n79057,
    n79058, n79059, n79060, n79061, n79062, n79063, n79064, n79065, n79066,
    n79067, n79068, n79069, n79070, n79071, n79072, n79073, n79074, n79075,
    n79076, n79077, n79078, n79079, n79080, n79081, n79082, n79083, n79084,
    n79085, n79086, n79087, n79088, n79089, n79090, n79091, n79092, n79093,
    n79094, n79095, n79096, n79097, n79098, n79099, n79100, n79101, n79102,
    n79103, n79104, n79105, n79106, n79107, n79108, n79109, n79110, n79111,
    n79112, n79113, n79114, n79115, n79116, n79117, n79118, n79119, n79120,
    n79121, n79122, n79123, n79124, n79125, n79126, n79127, n79128, n79129,
    n79130, n79131, n79132, n79133, n79134, n79135, n79136, n79137, n79138,
    n79139, n79140, n79141, n79142, n79143, n79144, n79145, n79146, n79147,
    n79148, n79149, n79150, n79151, n79152, n79153, n79154, n79155, n79156,
    n79157, n79158, n79159, n79160, n79161, n79162, n79163, n79164, n79165,
    n79166, n79167, n79168, n79169, n79170, n79171, n79172, n79173, n79174,
    n79175, n79176, n79177, n79178, n79179, n79180, n79181, n79182, n79183,
    n79184, n79185, n79186, n79187, n79188, n79189, n79190, n79191, n79192,
    n79193, n79194, n79195, n79196, n79197, n79198, n79199, n79200, n79201,
    n79202, n79203, n79204, n79205, n79206, n79207, n79208, n79209, n79210,
    n79211, n79212, n79213, n79214, n79215, n79216, n79217, n79218, n79219,
    n79220, n79221, n79222, n79223, n79224, n79225, n79226, n79227, n79228,
    n79229, n79230, n79231, n79232, n79233, n79234, n79235, n79236, n79237,
    n79238, n79239, n79240, n79241, n79242, n79243, n79244, n79245, n79246,
    n79247, n79248, n79249, n79250, n79251, n79252, n79253, n79254, n79255,
    n79256, n79257, n79258, n79259, n79260, n79261, n79262, n79263, n79264,
    n79265, n79266, n79267, n79268, n79269, n79270, n79271, n79272, n79273,
    n79274, n79275, n79276, n79277, n79278, n79279, n79280, n79281, n79282,
    n79283, n79284, n79285, n79286, n79287, n79288, n79289, n79290, n79291,
    n79292, n79293, n79294, n79295, n79296, n79297, n79298, n79299, n79300,
    n79301, n79302, n79303, n79304, n79305, n79306, n79307, n79308, n79309,
    n79310, n79311, n79312, n79313, n79314, n79315, n79316, n79317, n79318,
    n79319, n79320, n79321, n79322, n79323, n79324, n79325, n79326, n79327,
    n79328, n79329, n79330, n79331, n79332, n79333, n79334, n79335, n79336,
    n79337, n79338, n79339, n79340, n79341, n79342, n79343, n79344, n79345,
    n79346, n79347, n79348, n79349, n79350, n79351, n79352, n79353, n79354,
    n79355, n79356, n79357, n79358, n79359, n79360, n79361, n79362, n79363,
    n79364, n79365, n79366, n79367, n79368, n79369, n79370, n79371, n79372,
    n79373, n79374, n79375, n79376, n79377, n79378, n79379, n79380, n79381,
    n79382, n79383, n79384, n79385, n79386, n79387, n79388, n79389, n79390,
    n79391, n79392, n79393, n79394, n79395, n79396, n79397, n79398, n79399,
    n79400, n79401, n79402, n79403, n79404, n79405, n79406, n79407, n79408,
    n79409, n79410, n79411, n79412, n79413, n79414, n79415, n79416, n79417,
    n79418, n79419, n79420, n79421, n79422, n79423, n79424, n79425, n79426,
    n79427, n79428, n79429, n79430, n79431, n79432, n79433, n79434, n79435,
    n79436, n79437, n79438, n79439, n79440, n79441, n79442, n79443, n79444,
    n79445, n79446, n79447, n79448, n79449, n79450, n79451, n79452, n79453,
    n79454, n79455, n79456, n79457, n79458, n79459, n79460, n79461, n79462,
    n79463, n79464, n79465, n79466, n79467, n79468, n79469, n79470, n79471,
    n79472, n79473, n79474, n79475, n79476, n79477, n79478, n79479, n79480,
    n79481, n79482, n79483, n79484, n79485, n79486, n79487, n79488, n79489,
    n79490, n79491, n79492, n79493, n79494, n79495, n79496, n79497, n79498,
    n79499, n79500, n79501, n79502, n79503, n79504, n79505, n79506, n79507,
    n79508, n79509, n79510, n79511, n79512, n79513, n79514, n79515, n79516,
    n79517, n79518, n79519, n79520, n79521, n79522, n79523, n79524, n79525,
    n79526, n79527, n79528, n79529, n79530, n79531, n79532, n79533, n79534,
    n79535, n79536, n79537, n79538, n79539, n79540, n79541, n79542, n79543,
    n79544, n79545, n79546, n79547, n79548, n79549, n79550, n79551, n79552,
    n79553, n79554, n79555, n79556, n79557, n79558, n79559, n79560, n79561,
    n79562, n79563, n79564, n79565, n79566, n79567, n79568, n79569, n79570,
    n79571, n79572, n79573, n79574, n79575, n79576, n79577, n79578, n79579,
    n79580, n79581, n79582, n79583, n79584, n79585, n79586, n79587, n79588,
    n79589, n79590, n79591, n79592, n79593, n79594, n79595, n79596, n79597,
    n79598, n79599, n79600, n79601, n79602, n79603, n79604, n79605, n79606,
    n79607, n79608, n79609, n79610, n79611, n79612, n79613, n79614, n79615,
    n79616, n79617, n79618, n79619, n79620, n79621, n79622, n79623, n79624,
    n79625, n79626, n79627, n79628, n79629, n79630, n79631, n79632, n79633,
    n79634, n79635, n79636, n79637, n79638, n79639, n79640, n79641, n79642,
    n79643, n79644, n79645, n79646, n79647, n79648, n79649, n79650, n79651,
    n79652, n79653, n79654, n79655, n79656, n79657, n79658, n79659, n79660,
    n79661, n79662, n79663, n79664, n79665, n79666, n79667, n79668, n79669,
    n79670, n79671, n79672, n79673, n79674, n79675, n79676, n79677, n79678,
    n79679, n79680, n79681, n79682, n79683, n79684, n79685, n79686, n79687,
    n79688, n79689, n79690, n79691, n79692, n79693, n79694, n79695, n79696,
    n79697, n79698, n79699, n79700, n79701, n79702, n79703, n79704, n79705,
    n79706, n79707, n79708, n79709, n79710, n79711, n79712, n79713, n79714,
    n79715, n79716, n79717, n79718, n79719, n79720, n79721, n79722, n79723,
    n79724, n79725, n79726, n79727, n79728, n79729, n79730, n79731, n79732,
    n79733, n79734, n79735, n79736, n79737, n79738, n79739, n79740, n79741,
    n79742, n79743, n79744, n79745, n79746, n79747, n79748, n79749, n79750,
    n79751, n79752, n79753, n79754, n79755, n79756, n79757, n79758, n79759,
    n79760, n79761, n79762, n79763, n79764, n79765, n79766, n79767, n79768,
    n79769, n79770, n79771, n79772, n79773, n79774, n79775, n79776, n79777,
    n79778, n79779, n79780, n79781, n79782, n79783, n79784, n79785, n79786,
    n79787, n79788, n79789, n79790, n79791, n79792, n79793, n79794, n79795,
    n79796, n79797, n79798, n79799, n79800, n79801, n79802, n79803, n79804,
    n79805, n79806, n79807, n79808, n79809, n79810, n79811, n79812, n79813,
    n79814, n79815, n79816, n79817, n79818, n79819, n79820, n79821, n79822,
    n79823, n79824, n79825, n79826, n79827, n79828, n79829, n79830, n79831,
    n79832, n79833, n79834, n79835, n79836, n79837, n79838, n79839, n79840,
    n79841, n79842, n79843, n79844, n79845, n79846, n79847, n79848, n79849,
    n79850, n79851, n79852, n79853, n79854, n79855, n79856, n79857, n79858,
    n79859, n79860, n79861, n79862, n79863, n79864, n79865, n79866, n79867,
    n79868, n79869, n79870, n79871, n79872, n79873, n79874, n79875, n79876,
    n79877, n79878, n79879, n79880, n79881, n79882, n79883, n79884, n79885,
    n79886, n79887, n79888, n79889, n79890, n79891, n79892, n79893, n79894,
    n79895, n79896, n79897, n79898, n79899, n79900, n79901, n79902, n79903,
    n79904, n79905, n79906, n79907, n79908, n79909, n79910, n79911, n79912,
    n79913, n79914, n79915, n79916, n79917, n79918, n79919, n79920, n79921,
    n79922, n79923, n79924, n79925, n79926, n79927, n79928, n79929, n79930,
    n79931, n79932, n79933, n79934, n79935, n79936, n79937, n79938, n79939,
    n79940, n79941, n79942, n79943, n79944, n79945, n79946, n79947, n79948,
    n79949, n79950, n79951, n79952, n79953, n79954, n79955, n79956, n79957,
    n79958, n79959, n79960, n79961, n79962, n79963, n79964, n79965, n79966,
    n79967, n79968, n79969, n79970, n79971, n79972, n79973, n79974, n79975,
    n79976, n79977, n79978, n79979, n79980, n79981, n79982, n79983, n79984,
    n79985, n79986, n79987, n79988, n79989, n79990, n79991, n79992, n79993,
    n79994, n79995, n79996, n79997, n79998, n79999, n80000, n80001, n80002,
    n80003, n80004, n80005, n80006, n80007, n80008, n80009, n80010, n80011,
    n80012, n80013, n80014, n80015, n80016, n80017, n80018, n80019, n80020,
    n80021, n80022, n80023, n80024, n80025, n80026, n80027, n80028, n80029,
    n80030, n80031, n80032, n80033, n80034, n80035, n80036, n80037, n80038,
    n80039, n80040, n80041, n80042, n80043, n80044, n80045, n80046, n80047,
    n80048, n80049, n80050, n80051, n80052, n80053, n80054, n80055, n80056,
    n80057, n80058, n80059, n80060, n80061, n80062, n80063, n80064, n80065,
    n80066, n80067, n80068, n80069, n80070, n80071, n80072, n80073, n80074,
    n80075, n80076, n80077, n80078, n80079, n80080, n80081, n80082, n80083,
    n80084, n80085, n80086, n80087, n80088, n80089, n80090, n80091, n80092,
    n80093, n80094, n80095, n80096, n80097, n80098, n80099, n80100, n80101,
    n80102, n80103, n80104, n80105, n80106, n80107, n80108, n80109, n80110,
    n80111, n80112, n80113, n80114, n80115, n80116, n80117, n80118, n80119,
    n80120, n80121, n80122, n80123, n80124, n80125, n80126, n80127, n80128,
    n80129, n80130, n80131, n80132, n80133, n80134, n80135, n80136, n80137,
    n80138, n80139, n80140, n80141, n80142, n80143, n80144, n80145, n80146,
    n80147, n80148, n80149, n80150, n80151, n80152, n80153, n80154, n80155,
    n80156, n80157, n80158, n80159, n80160, n80161, n80162, n80163, n80164,
    n80165, n80166, n80167, n80168, n80169, n80170, n80171, n80172, n80173,
    n80174, n80175, n80176, n80177, n80178, n80179, n80180, n80181, n80182,
    n80183, n80184, n80185, n80186, n80187, n80188, n80189, n80190, n80191,
    n80192, n80193, n80194, n80195, n80196, n80197, n80198, n80199, n80200,
    n80201, n80202, n80203, n80204, n80205, n80206, n80207, n80208, n80209,
    n80210, n80211, n80212, n80213, n80214, n80215, n80216, n80217, n80218,
    n80219, n80220, n80221, n80222, n80223, n80224, n80225, n80226, n80227,
    n80228, n80229, n80230, n80231, n80232, n80233, n80234, n80235, n80236,
    n80237, n80238, n80239, n80240, n80241, n80242, n80243, n80244, n80245,
    n80246, n80247, n80248, n80249, n80250, n80251, n80252, n80253, n80254,
    n80255, n80256, n80257, n80258, n80259, n80260, n80261, n80262, n80263,
    n80264, n80265, n80266, n80267, n80268, n80269, n80270, n80271, n80272,
    n80273, n80274, n80275, n80276, n80277, n80278, n80279, n80280, n80281,
    n80282, n80283, n80284, n80285, n80286, n80287, n80288, n80289, n80290,
    n80291, n80292, n80293, n80294, n80295, n80296, n80297, n80298, n80299,
    n80300, n80301, n80302, n80303, n80304, n80305, n80306, n80307, n80308,
    n80309, n80310, n80311, n80312, n80313, n80314, n80315, n80316, n80317,
    n80318, n80319, n80320, n80321, n80322, n80323, n80324, n80325, n80326,
    n80327, n80328, n80329, n80330, n80331, n80332, n80333, n80334, n80335,
    n80336, n80337, n80338, n80339, n80340, n80341, n80342, n80343, n80344,
    n80345, n80346, n80347, n80348, n80349, n80350, n80351, n80352, n80353,
    n80354, n80355, n80356, n80357, n80358, n80359, n80360, n80361, n80362,
    n80363, n80364, n80365, n80366, n80367, n80368, n80369, n80370, n80371,
    n80372, n80373, n80374, n80375, n80376, n80377, n80378, n80379, n80380,
    n80381, n80382, n80383, n80384, n80385, n80386, n80387, n80388, n80389,
    n80390, n80391, n80392, n80393, n80394, n80395, n80396, n80397, n80398,
    n80399, n80400, n80401, n80402, n80403, n80404, n80405, n80406, n80407,
    n80408, n80409, n80410, n80411, n80412, n80413, n80414, n80415, n80416,
    n80417, n80418, n80419, n80420, n80421, n80422, n80423, n80424, n80425,
    n80426, n80427, n80428, n80429, n80430, n80431, n80432, n80433, n80434,
    n80435, n80436, n80437, n80438, n80439, n80440, n80441, n80442, n80443,
    n80444, n80445, n80446, n80447, n80448, n80449, n80450, n80451, n80452,
    n80453, n80454, n80455, n80456, n80457, n80458, n80459, n80460, n80461,
    n80462, n80463, n80464, n80465, n80466, n80467, n80468, n80469, n80470,
    n80471, n80472, n80473, n80474, n80475, n80476, n80477, n80478, n80479,
    n80480, n80481, n80482, n80483, n80484, n80485, n80486, n80487, n80488,
    n80489, n80490, n80491, n80492, n80493, n80494, n80495, n80496, n80497,
    n80498, n80499, n80500, n80501, n80502, n80503, n80504, n80505, n80506,
    n80507, n80508, n80509, n80510, n80511, n80512, n80513, n80514, n80515,
    n80516, n80517, n80518, n80519, n80520, n80521, n80522, n80523, n80524,
    n80525, n80526, n80527, n80528, n80529, n80530, n80531, n80532, n80533,
    n80534, n80535, n80536, n80537, n80538, n80539, n80540, n80541, n80542,
    n80543, n80544, n80545, n80546, n80547, n80548, n80549, n80550, n80551,
    n80552, n80553, n80554, n80555, n80556, n80557, n80558, n80559, n80560,
    n80561, n80562, n80563, n80564, n80565, n80566, n80567, n80568, n80569,
    n80570, n80571, n80572, n80573, n80574, n80575, n80576, n80577, n80578,
    n80579, n80580, n80581, n80582, n80583, n80584, n80585, n80586, n80587,
    n80588, n80589, n80590, n80591, n80592, n80593, n80594, n80595, n80596,
    n80597, n80598, n80599, n80600, n80601, n80602, n80603, n80604, n80605,
    n80606, n80607, n80608, n80609, n80610, n80611, n80612, n80613, n80614,
    n80615, n80616, n80617, n80618, n80619, n80620, n80621, n80622, n80623,
    n80624, n80625, n80626, n80627, n80628, n80629, n80630, n80631, n80632,
    n80633, n80634, n80635, n80636, n80637, n80638, n80639, n80640, n80641,
    n80642, n80643, n80644, n80645, n80646, n80647, n80648, n80649, n80650,
    n80651, n80652, n80653, n80654, n80655, n80656, n80657, n80658, n80659,
    n80660, n80661, n80662, n80663, n80664, n80665, n80666, n80667, n80668,
    n80669, n80670, n80671, n80672, n80673, n80674, n80675, n80676, n80677,
    n80678, n80679, n80680, n80681, n80682, n80683, n80684, n80685, n80686,
    n80687, n80688, n80689, n80690, n80691, n80692, n80693, n80694, n80695,
    n80696, n80697, n80698, n80699, n80700, n80701, n80702, n80703, n80704,
    n80705, n80706, n80707, n80708, n80709, n80710, n80711, n80712, n80713,
    n80714, n80715, n80716, n80717, n80718, n80719, n80720, n80721, n80722,
    n80723, n80724, n80725, n80726, n80727, n80728, n80729, n80730, n80731,
    n80732, n80733, n80734, n80735, n80736, n80737, n80738, n80739, n80740,
    n80741, n80742, n80743, n80744, n80745, n80746, n80747, n80748, n80749,
    n80750, n80751, n80752, n80753, n80754, n80755, n80756, n80757, n80758,
    n80759, n80760, n80761, n80762, n80763, n80764, n80765, n80766, n80767,
    n80768, n80769, n80770, n80771, n80772, n80773, n80774, n80775, n80776,
    n80777, n80778, n80779, n80780, n80781, n80782, n80783, n80784, n80785,
    n80786, n80787, n80788, n80789, n80790, n80791, n80792, n80793, n80794,
    n80795, n80796, n80797, n80798, n80799, n80800, n80801, n80802, n80803,
    n80804, n80805, n80806, n80807, n80808, n80809, n80810, n80811, n80812,
    n80813, n80814, n80815, n80816, n80817, n80818, n80819, n80820, n80821,
    n80822, n80823, n80824, n80825, n80826, n80827, n80828, n80829, n80830,
    n80831, n80832, n80833, n80834, n80835, n80836, n80837, n80838, n80839,
    n80840, n80841, n80842, n80843, n80844, n80845, n80846, n80847, n80848,
    n80849, n80850, n80851, n80852, n80853, n80854, n80855, n80856, n80857,
    n80858, n80859, n80860, n80861, n80862, n80863, n80864, n80865, n80866,
    n80867, n80868, n80869, n80870, n80871, n80872, n80873, n80874, n80875,
    n80876, n80877, n80878, n80879, n80880, n80881, n80882, n80883, n80884,
    n80885, n80886, n80887, n80888, n80889, n80890, n80891, n80892, n80893,
    n80894, n80895, n80896, n80897, n80898, n80899, n80900, n80901, n80902,
    n80903, n80904, n80905, n80906, n80907, n80908, n80909, n80910, n80911,
    n80912, n80913, n80914, n80915, n80916, n80917, n80918, n80919, n80920,
    n80921, n80922, n80923, n80924, n80925, n80926, n80927, n80928, n80929,
    n80930, n80931, n80932, n80933, n80934, n80935, n80936, n80937, n80938,
    n80939, n80940, n80941, n80942, n80943, n80944, n80945, n80946, n80947,
    n80948, n80949, n80950, n80951, n80952, n80953, n80954, n80955, n80956,
    n80957, n80958, n80959, n80960, n80961, n80962, n80963, n80964, n80965,
    n80966, n80967, n80968, n80969, n80970, n80971, n80972, n80973, n80974,
    n80975, n80976, n80977, n80978, n80979, n80980, n80981, n80982, n80983,
    n80984, n80985, n80986, n80987, n80988, n80989, n80990, n80991, n80992,
    n80993, n80994, n80995, n80996, n80997, n80998, n80999, n81000, n81001,
    n81002, n81003, n81004, n81005, n81006, n81007, n81008, n81009, n81010,
    n81011, n81012, n81013, n81014, n81015, n81016, n81017, n81018, n81019,
    n81020, n81021, n81022, n81023, n81024, n81025, n81026, n81027, n81028,
    n81029, n81030, n81031, n81032, n81033, n81034, n81035, n81036, n81037,
    n81038, n81039, n81040, n81041, n81042, n81043, n81044, n81045, n81046,
    n81047, n81048, n81049, n81050, n81051, n81052, n81053, n81054, n81055,
    n81056, n81057, n81058, n81059, n81060, n81061, n81062, n81063, n81064,
    n81065, n81066, n81067, n81068, n81069, n81070, n81071, n81072, n81073,
    n81074, n81075, n81076, n81077, n81078, n81079, n81080, n81081, n81082,
    n81083, n81084, n81085, n81086, n81087, n81088, n81089, n81090, n81091,
    n81092, n81093, n81094, n81095, n81096, n81097, n81098, n81099, n81100,
    n81101, n81102, n81103, n81104, n81105, n81106, n81107, n81108, n81109,
    n81110, n81111, n81112, n81113, n81114, n81115, n81116, n81117, n81118,
    n81119, n81120, n81121, n81122, n81123, n81124, n81125, n81126, n81127,
    n81128, n81129, n81130, n81131, n81132, n81133, n81134, n81135, n81136,
    n81137, n81138, n81139, n81140, n81141, n81142, n81143, n81144, n81145,
    n81146, n81147, n81148, n81149, n81150, n81151, n81152, n81153, n81154,
    n81155, n81156, n81157, n81158, n81159, n81160, n81161, n81162, n81163,
    n81164, n81165, n81166, n81167, n81168, n81169, n81170, n81171, n81172,
    n81173, n81174, n81175, n81176, n81177, n81178, n81179, n81180, n81181,
    n81182, n81183, n81184, n81185, n81186, n81187, n81188, n81189, n81190,
    n81191, n81192, n81193, n81194, n81195, n81196, n81197, n81198, n81199,
    n81200, n81201, n81202, n81203, n81204, n81205, n81206, n81207, n81208,
    n81209, n81210, n81211, n81212, n81213, n81214, n81215, n81216, n81217,
    n81218, n81219, n81220, n81221, n81222, n81223, n81224, n81225, n81226,
    n81227, n81228, n81229, n81230, n81231, n81232, n81233, n81234, n81235,
    n81236, n81237, n81238, n81239, n81240, n81241, n81242, n81243, n81244,
    n81245, n81246, n81247, n81248, n81249, n81250, n81251, n81252, n81253,
    n81254, n81255, n81256, n81257, n81258, n81259, n81260, n81261, n81262,
    n81263, n81264, n81265, n81266, n81267, n81268, n81269, n81270, n81271,
    n81272, n81273, n81274, n81275, n81276, n81277, n81278, n81279, n81280,
    n81281, n81282, n81283, n81284, n81285, n81286, n81287, n81288, n81289,
    n81290, n81291, n81292, n81293, n81294, n81295, n81296, n81297, n81298,
    n81299, n81300, n81301, n81302, n81303, n81304, n81305, n81306, n81307,
    n81308, n81309, n81310, n81311, n81312, n81313, n81314, n81315, n81316,
    n81317, n81318, n81319, n81320, n81321, n81322, n81323, n81324, n81325,
    n81326, n81327, n81328, n81329, n81330, n81331, n81332, n81333, n81334,
    n81335, n81336, n81337, n81338, n81339, n81340, n81341, n81342, n81343,
    n81344, n81345, n81346, n81347, n81348, n81349, n81350, n81351, n81352,
    n81353, n81354, n81355, n81356, n81357, n81358, n81359, n81360, n81361,
    n81362, n81363, n81364, n81365, n81366, n81367, n81368, n81369, n81370,
    n81371, n81372, n81373, n81374, n81375, n81376, n81377, n81378, n81379,
    n81380, n81381, n81382, n81383, n81384, n81385, n81386, n81387, n81388,
    n81389, n81390, n81391, n81392, n81393, n81394, n81395, n81396, n81397,
    n81398, n81399, n81400, n81401, n81402, n81403, n81404, n81405, n81406,
    n81407, n81408, n81409, n81410, n81411, n81412, n81413, n81414, n81415,
    n81416, n81417, n81418, n81419, n81420, n81421, n81422, n81423, n81424,
    n81425, n81426, n81427, n81428, n81429, n81430, n81431, n81432, n81433,
    n81434, n81435, n81436, n81437, n81438, n81439, n81440, n81441, n81442,
    n81443, n81444, n81445, n81446, n81447, n81448, n81449, n81450, n81451,
    n81452, n81453, n81454, n81455, n81456, n81457, n81458, n81459, n81460,
    n81461, n81462, n81463, n81464, n81465, n81466, n81467, n81468, n81469,
    n81470, n81471, n81472, n81473, n81474, n81475, n81476, n81477, n81478,
    n81479, n81480, n81481, n81482, n81483, n81484, n81485, n81486, n81487,
    n81488, n81489, n81490, n81491, n81492, n81493, n81494, n81495, n81496,
    n81497, n81498, n81499, n81500, n81501, n81502, n81503, n81504, n81505,
    n81506, n81507, n81508, n81509, n81510, n81511, n81512, n81513, n81514,
    n81515, n81516, n81517, n81518, n81519, n81520, n81521, n81522, n81523,
    n81524, n81525, n81526, n81527, n81528, n81529, n81530, n81531, n81532,
    n81533, n81534, n81535, n81536, n81537, n81538, n81539, n81540, n81541,
    n81542, n81543, n81544, n81545, n81546, n81547, n81548, n81549, n81550,
    n81551, n81552, n81553, n81554, n81555, n81556, n81557, n81558, n81559,
    n81560, n81561, n81562, n81563, n81564, n81565, n81566, n81567, n81568,
    n81569, n81570, n81571, n81572, n81573, n81574, n81575, n81576, n81577,
    n81578, n81579, n81580, n81581, n81582, n81583, n81584, n81585, n81586,
    n81587, n81588, n81589, n81590, n81591, n81592, n81593, n81594, n81595,
    n81596, n81597, n81598, n81599, n81600, n81601, n81602, n81603, n81604,
    n81605, n81606, n81607, n81608, n81609, n81610, n81611, n81612, n81613,
    n81614, n81615, n81616, n81617, n81618, n81619, n81620, n81621, n81622,
    n81623, n81624, n81625, n81626, n81627, n81628, n81629, n81630, n81631,
    n81632, n81633, n81634, n81635, n81636, n81637, n81638, n81639, n81640,
    n81641, n81642, n81643, n81644, n81645, n81646, n81647, n81648, n81649,
    n81650, n81651, n81652, n81653, n81654, n81655, n81656, n81657, n81658,
    n81659, n81660, n81661, n81662, n81663, n81664, n81665, n81666, n81667,
    n81668, n81669, n81670, n81671, n81672, n81673, n81674, n81675, n81676,
    n81677, n81678, n81679, n81680, n81681, n81682, n81683, n81684, n81685,
    n81686, n81687, n81688, n81689, n81690, n81691, n81692, n81693, n81694,
    n81695, n81696, n81697, n81698, n81699, n81700, n81701, n81702, n81703,
    n81704, n81705, n81706, n81707, n81708, n81709, n81710, n81711, n81712,
    n81713, n81714, n81715, n81716, n81717, n81718, n81719, n81720, n81721,
    n81722, n81723, n81724, n81725, n81726, n81727, n81728, n81729, n81730,
    n81731, n81732, n81733, n81734, n81735, n81736, n81737, n81738, n81739,
    n81740, n81741, n81742, n81743, n81744, n81745, n81746, n81747, n81748,
    n81749, n81750, n81751, n81752, n81753, n81754, n81755, n81756, n81757,
    n81758, n81759, n81760, n81761, n81762, n81763, n81764, n81765, n81766,
    n81767, n81768, n81769, n81770, n81771, n81772, n81773, n81774, n81775,
    n81776, n81777, n81778, n81779, n81780, n81781, n81782, n81783, n81784,
    n81785, n81786, n81787, n81788, n81789, n81790, n81791, n81792, n81793,
    n81794, n81795, n81796, n81797, n81798, n81799, n81800, n81801, n81802,
    n81803, n81804, n81805, n81806, n81807, n81808, n81809, n81810, n81811,
    n81812, n81813, n81814, n81815, n81816, n81817, n81818, n81819, n81820,
    n81821, n81822, n81823, n81824, n81825, n81826, n81827, n81828, n81829,
    n81830, n81831, n81832, n81833, n81834, n81835, n81836, n81837, n81838,
    n81839, n81840, n81841, n81842, n81843, n81844, n81845, n81846, n81847,
    n81848, n81849, n81850, n81851, n81852, n81853, n81854, n81855, n81856,
    n81857, n81858, n81859, n81860, n81861, n81862, n81863, n81864, n81865,
    n81866, n81867, n81868, n81869, n81870, n81871, n81872, n81873, n81874,
    n81875, n81876, n81877, n81878, n81879, n81880, n81881, n81882, n81883,
    n81884, n81885, n81886, n81887, n81888, n81889, n81890, n81891, n81892,
    n81893, n81894, n81895, n81896, n81897, n81898, n81899, n81900, n81901,
    n81902, n81903, n81904, n81905, n81906, n81907, n81908, n81909, n81910,
    n81911, n81912, n81913, n81914, n81915, n81916, n81917, n81918, n81919,
    n81920, n81921, n81922, n81923, n81924, n81925, n81926, n81927, n81928,
    n81929, n81930, n81931, n81932, n81933, n81934, n81935, n81936, n81937,
    n81938, n81939, n81940, n81941, n81942, n81943, n81944, n81945, n81946,
    n81947, n81948, n81949, n81950, n81951, n81952, n81953, n81954, n81955,
    n81956, n81957, n81958, n81959, n81960, n81961, n81962, n81963, n81964,
    n81965, n81966, n81967, n81968, n81969, n81970, n81971, n81972, n81973,
    n81974, n81975, n81976, n81977, n81978, n81979, n81980, n81981, n81982,
    n81983, n81984, n81985, n81986, n81987, n81988, n81989, n81990, n81991,
    n81992, n81993, n81994, n81995, n81996, n81997, n81998, n81999, n82000,
    n82001, n82002, n82003, n82004, n82005, n82006, n82007, n82008, n82009,
    n82010, n82011, n82012, n82013, n82014, n82015, n82016, n82017, n82018,
    n82019, n82020, n82021, n82022, n82023, n82024, n82025, n82026, n82027,
    n82028, n82029, n82030, n82031, n82032, n82033, n82034, n82035, n82036,
    n82037, n82038, n82039, n82040, n82041, n82042, n82043, n82044, n82045,
    n82046, n82047, n82048, n82049, n82050, n82051, n82052, n82053, n82054,
    n82055, n82056, n82057, n82058, n82059, n82060, n82061, n82062, n82063,
    n82064, n82065, n82066, n82067, n82068, n82069, n82070, n82071, n82072,
    n82073, n82074, n82075, n82076, n82077, n82078, n82079, n82080, n82081,
    n82082, n82083, n82084, n82085, n82086, n82087, n82088, n82089, n82090,
    n82091, n82092, n82093, n82094, n82095, n82096, n82097, n82098, n82099,
    n82100, n82101, n82102, n82103, n82104, n82105, n82106, n82107, n82108,
    n82109, n82110, n82111, n82112, n82113, n82114, n82115, n82116, n82117,
    n82118, n82119, n82120, n82121, n82122, n82123, n82124, n82125, n82126,
    n82127, n82128, n82129, n82130, n82131, n82132, n82133, n82134, n82135,
    n82136, n82137, n82138, n82139, n82140, n82141, n82142, n82143, n82144,
    n82145, n82146, n82147, n82148, n82149, n82150, n82151, n82152, n82153,
    n82154, n82155, n82156, n82157, n82158, n82159, n82160, n82161, n82162,
    n82163, n82164, n82165, n82166, n82167, n82168, n82169, n82170, n82171,
    n82172, n82173, n82174, n82175, n82176, n82177, n82178, n82179, n82180,
    n82181, n82182, n82183, n82184, n82185, n82186, n82187, n82188, n82189,
    n82190, n82191, n82192, n82193, n82194, n82195, n82196, n82197, n82198,
    n82199, n82200, n82201, n82202, n82203, n82204, n82205, n82206, n82207,
    n82208, n82209, n82210, n82211, n82212, n82213, n82214, n82215, n82216,
    n82217, n82218, n82219, n82220, n82221, n82222, n82223, n82224, n82225,
    n82226, n82227, n82228, n82229, n82230, n82231, n82232, n82233, n82234,
    n82235, n82236, n82237, n82238, n82239, n82240, n82241, n82242, n82243,
    n82244, n82245, n82246, n82247, n82248, n82249, n82250, n82251, n82252,
    n82253, n82254, n82255, n82256, n82257, n82258, n82259, n82260, n82261,
    n82262, n82263, n82264, n82265, n82266, n82267, n82268, n82269, n82270,
    n82271, n82272, n82273, n82274, n82275, n82276, n82277, n82278, n82279,
    n82280, n82281, n82282, n82283, n82284, n82285, n82286, n82287, n82288,
    n82289, n82290, n82291, n82292, n82293, n82294, n82295, n82296, n82297,
    n82298, n82299, n82300, n82301, n82302, n82303, n82304, n82305, n82306,
    n82307, n82308, n82309, n82310, n82311, n82312, n82313, n82314, n82315,
    n82316, n82317, n82318, n82319, n82320, n82321, n82322, n82323, n82324,
    n82325, n82326, n82327, n82328, n82329, n82330, n82331, n82332, n82333,
    n82334, n82335, n82336, n82337, n82338, n82339, n82340, n82341, n82342,
    n82343, n82344, n82345, n82346, n82347, n82348, n82349, n82350, n82351,
    n82352, n82353, n82354, n82355, n82356, n82357, n82358, n82359, n82360,
    n82361, n82362, n82363, n82364, n82365, n82366, n82367, n82368, n82369,
    n82370, n82371, n82372, n82373, n82374, n82375, n82376, n82377, n82378,
    n82379, n82380, n82381, n82382, n82383, n82384, n82385, n82386, n82387,
    n82388, n82389, n82390, n82391, n82392, n82393, n82394, n82395, n82396,
    n82397, n82398, n82399, n82400, n82401, n82402, n82403, n82404, n82405,
    n82406, n82407, n82408, n82409, n82410, n82411, n82412, n82413, n82414,
    n82415, n82416, n82417, n82418, n82419, n82420, n82421, n82422, n82423,
    n82424, n82425, n82426, n82427, n82428, n82429, n82430, n82431, n82432,
    n82433, n82434, n82435, n82436, n82437, n82438, n82439, n82440, n82441,
    n82442, n82443, n82444, n82445, n82446, n82447, n82448, n82449, n82450,
    n82451, n82452, n82453, n82454, n82455, n82456, n82457, n82458, n82459,
    n82460, n82461, n82462, n82463, n82464, n82465, n82466, n82467, n82468,
    n82469, n82470, n82471, n82472, n82473, n82474, n82475, n82476, n82477,
    n82478, n82479, n82480, n82481, n82482, n82483, n82484, n82485, n82486,
    n82487, n82488, n82489, n82490, n82491, n82492, n82493, n82494, n82495,
    n82496, n82497, n82498, n82499, n82500, n82501, n82502, n82503, n82504,
    n82505, n82506, n82507, n82508, n82509, n82510, n82511, n82512, n82513,
    n82514, n82515, n82516, n82517, n82518, n82519, n82520, n82521, n82522,
    n82523, n82524, n82525, n82526, n82527, n82528, n82529, n82530, n82531,
    n82532, n82533, n82534, n82535, n82536, n82537, n82538, n82539, n82540,
    n82541, n82542, n82543, n82544, n82545, n82546, n82547, n82548, n82549,
    n82550, n82551, n82552, n82553, n82554, n82555, n82556, n82557, n82558,
    n82559, n82560, n82561, n82562, n82563, n82564, n82565, n82566, n82567,
    n82568, n82569, n82570, n82571, n82572, n82573, n82574, n82575, n82576,
    n82577, n82578, n82579, n82580, n82581, n82582, n82583, n82584, n82585,
    n82586, n82587, n82588, n82589, n82590, n82591, n82592, n82593, n82594,
    n82595, n82596, n82597, n82598, n82599, n82600, n82601, n82602, n82603,
    n82604, n82605, n82606, n82607, n82608, n82609, n82610, n82611, n82612,
    n82613, n82614, n82615, n82616, n82617, n82618, n82619, n82620, n82621,
    n82622, n82623, n82624, n82625, n82626, n82627, n82628, n82629, n82630,
    n82631, n82632, n82633, n82634, n82635, n82636, n82637, n82638, n82639,
    n82640, n82641, n82642, n82643, n82644, n82645, n82646, n82647, n82648,
    n82649, n82650, n82651, n82652, n82653, n82654, n82655, n82656, n82657,
    n82658, n82659, n82660, n82661, n82662, n82663, n82664, n82665, n82666,
    n82667, n82668, n82669, n82670, n82671, n82672, n82673, n82674, n82675,
    n82676, n82677, n82678, n82679, n82680, n82681, n82682, n82683, n82684,
    n82685, n82686, n82687, n82688, n82689, n82690, n82691, n82692, n82693,
    n82694, n82695, n82696, n82697, n82698, n82699, n82700, n82701, n82702,
    n82703, n82704, n82705, n82706, n82707, n82708, n82709, n82710, n82711,
    n82712, n82713, n82714, n82715, n82716, n82717, n82718, n82719, n82720,
    n82721, n82722, n82723, n82724, n82725, n82726, n82727, n82728, n82729,
    n82730, n82731, n82732, n82733, n82734, n82735, n82736, n82737, n82738,
    n82739, n82740, n82741, n82742, n82743, n82744, n82745, n82746, n82747,
    n82748, n82749, n82750, n82751, n82752, n82753, n82754, n82755, n82756,
    n82757, n82758, n82759, n82760, n82761, n82762, n82763, n82764, n82765,
    n82766, n82767, n82768, n82769, n82770, n82771, n82772, n82773, n82774,
    n82775, n82776, n82777, n82778, n82779, n82780, n82781, n82782, n82783,
    n82784, n82785, n82786, n82787, n82788, n82789, n82790, n82791, n82792,
    n82793, n82794, n82795, n82796, n82797, n82798, n82799, n82800, n82801,
    n82802, n82803, n82804, n82805, n82806, n82807, n82808, n82809, n82810,
    n82811, n82812, n82813, n82814, n82815, n82816, n82817, n82818, n82819,
    n82820, n82821, n82822, n82823, n82824, n82825, n82826, n82827, n82828,
    n82829, n82830, n82831, n82832, n82833, n82834, n82835, n82836, n82837,
    n82838, n82839, n82840, n82841, n82842, n82843, n82844, n82845, n82846,
    n82847, n82848, n82849, n82850, n82851, n82852, n82853, n82854, n82855,
    n82856, n82857, n82858, n82859, n82860, n82861, n82862, n82863, n82864,
    n82865, n82866, n82867, n82868, n82869, n82870, n82871, n82872, n82873,
    n82874, n82875, n82876, n82877, n82878, n82879, n82880, n82881, n82882,
    n82883, n82884, n82885, n82886, n82887, n82888, n82889, n82890, n82891,
    n82892, n82893, n82894, n82895, n82896, n82897, n82898, n82899, n82900,
    n82901, n82902, n82903, n82904, n82905, n82906, n82907, n82908, n82909,
    n82910, n82911, n82912, n82913, n82914, n82915, n82916, n82917, n82918,
    n82919, n82920, n82921, n82922, n82923, n82924, n82925, n82926, n82927,
    n82928, n82929, n82930, n82931, n82932, n82933, n82934, n82935, n82936,
    n82937, n82938, n82939, n82940, n82941, n82942, n82943, n82944, n82945,
    n82946, n82947, n82948, n82949, n82950, n82951, n82952, n82953, n82954,
    n82955, n82956, n82957, n82958, n82959, n82960, n82961, n82962, n82963,
    n82964, n82965, n82966, n82967, n82968, n82969, n82970, n82971, n82972,
    n82973, n82974, n82975, n82976, n82977, n82978, n82979, n82980, n82981,
    n82982, n82983, n82984, n82985, n82986, n82987, n82988, n82989, n82990,
    n82991, n82992, n82993, n82994, n82995, n82996, n82997, n82998, n82999,
    n83000, n83001, n83002, n83003, n83004, n83005, n83006, n83007, n83008,
    n83009, n83010, n83011, n83012, n83013, n83014, n83015, n83016, n83017,
    n83018, n83019, n83020, n83021, n83022, n83023, n83024, n83025, n83026,
    n83027, n83028, n83029, n83030, n83031, n83032, n83033, n83034, n83035,
    n83036, n83037, n83038, n83039, n83040, n83041, n83042, n83043, n83044,
    n83045, n83046, n83047, n83048, n83049, n83050, n83051, n83052, n83053,
    n83054, n83055, n83056, n83057, n83058, n83059, n83060, n83061, n83062,
    n83063, n83064, n83065, n83066, n83067, n83068, n83069, n83070, n83071,
    n83072, n83073, n83074, n83075, n83076, n83077, n83078, n83079, n83080,
    n83081, n83082, n83083, n83084, n83085, n83086, n83087, n83088, n83089,
    n83090, n83091, n83092, n83093, n83094, n83095, n83096, n83097, n83098,
    n83099, n83100, n83101, n83102, n83103, n83104, n83105, n83106, n83107,
    n83108, n83109, n83110, n83111, n83112, n83113, n83114, n83115, n83116,
    n83117, n83118, n83119, n83120, n83121, n83122, n83123, n83124, n83125,
    n83126, n83127, n83128, n83129, n83130, n83131, n83132, n83133, n83134,
    n83135, n83136, n83137, n83138, n83139, n83140, n83141, n83142, n83143,
    n83144, n83145, n83146, n83147, n83148, n83149, n83150, n83151, n83152,
    n83153, n83154, n83155, n83156, n83157, n83158, n83159, n83160, n83161,
    n83162, n83163, n83164, n83165, n83166, n83167, n83168, n83169, n83170,
    n83171, n83172, n83173, n83174, n83175, n83176, n83177, n83178, n83179,
    n83180, n83181, n83182, n83183, n83184, n83185, n83186, n83187, n83188,
    n83189, n83190, n83191, n83192, n83193, n83194, n83195, n83196, n83197,
    n83198, n83199, n83200, n83201, n83202, n83203, n83204, n83205, n83206,
    n83207, n83208, n83209, n83210, n83211, n83212, n83213, n83214, n83215,
    n83216, n83217, n83218, n83219, n83220, n83221, n83222, n83223, n83224,
    n83225, n83226, n83227, n83228, n83229, n83230, n83231, n83232, n83233,
    n83234, n83235, n83236, n83237, n83238, n83239, n83240, n83241, n83242,
    n83243, n83244, n83245, n83246, n83247, n83248, n83249, n83250, n83251,
    n83252, n83253, n83254, n83255, n83256, n83257, n83258, n83259, n83260,
    n83261, n83262, n83263, n83264, n83265, n83266, n83267, n83268, n83269,
    n83270, n83271, n83272, n83273, n83274, n83275, n83276, n83277, n83278,
    n83279, n83280, n83281, n83282, n83283, n83284, n83285, n83286, n83287,
    n83288, n83289, n83290, n83291, n83292, n83293, n83294, n83295, n83296,
    n83297, n83298, n83299, n83300, n83301, n83302, n83303, n83304, n83305,
    n83306, n83307, n83308, n83309, n83310, n83311, n83312, n83313, n83314,
    n83315, n83316, n83317, n83318, n83319, n83320, n83321, n83322, n83323,
    n83324, n83325, n83326, n83327, n83328, n83329, n83330, n83331, n83332,
    n83333, n83334, n83335, n83336, n83337, n83338, n83339, n83340, n83341,
    n83342, n83343, n83344, n83345, n83346, n83347, n83348, n83349, n83350,
    n83351, n83352, n83353, n83354, n83355, n83356, n83357, n83358, n83359,
    n83360, n83361, n83362, n83363, n83364, n83365, n83366, n83367, n83368,
    n83369, n83370, n83371, n83372, n83373, n83374, n83375, n83376, n83377,
    n83378, n83379, n83380, n83381, n83382, n83383, n83384, n83385, n83386,
    n83387, n83388, n83389, n83390, n83391, n83392, n83393, n83394, n83395,
    n83396, n83397, n83398, n83399, n83400, n83401, n83402, n83403, n83404,
    n83405, n83406, n83407, n83408, n83409, n83410, n83411, n83412, n83413,
    n83414, n83415, n83416, n83417, n83418, n83419, n83420, n83421, n83422,
    n83423, n83424, n83425, n83426, n83427, n83428, n83429, n83430, n83431,
    n83432, n83433, n83434, n83435, n83436, n83437, n83438, n83439, n83440,
    n83441, n83442, n83443, n83444, n83445, n83446, n83447, n83448, n83449,
    n83450, n83451, n83452, n83453, n83454, n83455, n83456, n83457, n83458,
    n83459, n83460, n83461, n83462, n83463, n83464, n83465, n83466, n83467,
    n83468, n83469, n83470, n83471, n83472, n83473, n83474, n83475, n83476,
    n83477, n83478, n83479, n83480, n83481, n83482, n83483, n83484, n83485,
    n83486, n83487, n83488, n83489, n83490, n83491, n83492, n83493, n83494,
    n83495, n83496, n83497, n83498, n83499, n83500, n83501, n83502, n83503,
    n83504, n83505, n83506, n83507, n83508, n83509, n83510, n83511, n83512,
    n83513, n83514, n83515, n83516, n83517, n83518, n83519, n83520, n83521,
    n83522, n83523, n83524, n83525, n83526, n83527, n83528, n83529, n83530,
    n83531, n83532, n83533, n83534, n83535, n83536, n83537, n83538, n83539,
    n83540, n83541, n83542, n83543, n83544, n83545, n83546, n83547, n83548,
    n83549, n83550, n83551, n83552, n83553, n83554, n83555, n83556, n83557,
    n83558, n83559, n83560, n83561, n83562, n83563, n83564, n83565, n83566,
    n83567, n83568, n83569, n83570, n83571, n83572, n83573, n83574, n83575,
    n83576, n83577, n83578, n83579, n83580, n83581, n83582, n83583, n83584,
    n83585, n83586, n83587, n83588, n83589, n83590, n83591, n83592, n83593,
    n83594, n83595, n83596, n83597, n83598, n83599, n83600, n83601, n83602,
    n83603, n83604, n83605, n83606, n83607, n83608, n83609, n83610, n83611,
    n83612, n83613, n83614, n83615, n83616, n83617, n83618, n83619, n83620,
    n83621, n83622, n83623, n83624, n83625, n83626, n83627, n83628, n83629,
    n83630, n83631, n83632, n83633, n83634, n83635, n83636, n83637, n83638,
    n83639, n83640, n83641, n83642, n83643, n83644, n83645, n83646, n83647,
    n83648, n83649, n83650, n83651, n83652, n83653, n83654, n83655, n83656,
    n83657, n83658, n83659, n83660, n83661, n83662, n83663, n83664, n83665,
    n83666, n83667, n83668, n83669, n83670, n83671, n83672, n83673, n83674,
    n83675, n83676, n83677, n83678, n83679, n83680, n83681, n83682, n83683,
    n83684, n83685, n83686, n83687, n83688, n83689, n83690, n83691, n83692,
    n83693, n83694, n83695, n83696, n83697, n83698, n83699, n83700, n83701,
    n83702, n83703, n83704, n83705, n83706, n83707, n83708, n83709, n83710,
    n83711, n83712, n83713, n83714, n83715, n83716, n83717, n83718, n83719,
    n83720, n83721, n83722, n83723, n83724, n83725, n83726, n83727, n83728,
    n83729, n83730, n83731, n83732, n83733, n83734, n83735, n83736, n83737,
    n83738, n83739, n83740, n83741, n83742, n83743, n83744, n83745, n83746,
    n83747, n83748, n83749, n83750, n83751, n83752, n83753, n83754, n83755,
    n83756, n83757, n83758, n83759, n83760, n83761, n83762, n83763, n83764,
    n83765, n83766, n83767, n83768, n83769, n83770, n83771, n83772, n83773,
    n83774, n83775, n83776, n83777, n83778, n83779, n83780, n83781, n83782,
    n83783, n83784, n83785, n83786, n83787, n83788, n83789, n83790, n83791,
    n83792, n83793, n83794, n83795, n83796, n83797, n83798, n83799, n83800,
    n83801, n83802, n83803, n83804, n83805, n83806, n83807, n83808, n83809,
    n83810, n83811, n83812, n83813, n83814, n83815, n83816, n83817, n83818,
    n83819, n83820, n83821, n83822, n83823, n83824, n83825, n83826, n83827,
    n83828, n83829, n83830, n83831, n83832, n83833, n83834, n83835, n83836,
    n83837, n83838, n83839, n83840, n83841, n83842, n83843, n83844, n83845,
    n83846, n83847, n83848, n83849, n83850, n83851, n83852, n83853, n83854,
    n83855, n83856, n83857, n83858, n83859, n83860, n83861, n83862, n83863,
    n83864, n83865, n83866, n83867, n83868, n83869, n83870, n83871, n83872,
    n83873, n83874, n83875, n83876, n83877, n83878, n83879, n83880, n83881,
    n83882, n83883, n83884, n83885, n83886, n83887, n83888, n83889, n83890,
    n83891, n83892, n83893, n83894, n83895, n83896, n83897, n83898, n83899,
    n83900, n83901, n83902, n83903, n83904, n83905, n83906, n83907, n83908,
    n83909, n83910, n83911, n83912, n83913, n83914, n83915, n83916, n83917,
    n83918, n83919, n83920, n83921, n83922, n83923, n83924, n83925, n83926,
    n83927, n83928, n83929, n83930, n83931, n83932, n83933, n83934, n83935,
    n83936, n83937, n83938, n83939, n83940, n83941, n83942, n83943, n83944,
    n83945, n83946, n83947, n83948, n83949, n83950, n83951, n83952, n83953,
    n83954, n83955, n83956, n83957, n83958, n83959, n83960, n83961, n83962,
    n83963, n83964, n83965, n83966, n83967, n83968, n83969, n83970, n83971,
    n83972, n83973, n83974, n83975, n83976, n83977, n83978, n83979, n83980,
    n83981, n83982, n83983, n83984, n83985, n83986, n83987, n83988, n83989,
    n83990, n83991, n83992, n83993, n83994, n83995, n83996, n83997, n83998,
    n83999, n84000, n84001, n84002, n84003, n84004, n84005, n84006, n84007,
    n84008, n84009, n84010, n84011, n84012, n84013, n84014, n84015, n84016,
    n84017, n84018, n84019, n84020, n84021, n84022, n84023, n84024, n84025,
    n84026, n84027, n84028, n84029, n84030, n84031, n84032, n84033, n84034,
    n84035, n84036, n84037, n84038, n84039, n84040, n84041, n84042, n84043,
    n84044, n84045, n84046, n84047, n84048, n84049, n84050, n84051, n84052,
    n84053, n84054, n84055, n84056, n84057, n84058, n84059, n84060, n84061,
    n84062, n84063, n84064, n84065, n84066, n84067, n84068, n84069, n84070,
    n84071, n84072, n84073, n84074, n84075, n84076, n84077, n84078, n84079,
    n84080, n84081, n84082, n84083, n84084, n84085, n84086, n84087, n84088,
    n84089, n84090, n84091, n84092, n84093, n84094, n84095, n84096, n84097,
    n84098, n84099, n84100, n84101, n84102, n84103, n84104, n84105, n84106,
    n84107, n84108, n84109, n84110, n84111, n84112, n84113, n84114, n84115,
    n84116, n84117, n84118, n84119, n84120, n84121, n84122, n84123, n84124,
    n84125, n84126, n84127, n84128, n84129, n84130, n84131, n84132, n84133,
    n84134, n84135, n84136, n84137, n84138, n84139, n84140, n84141, n84142,
    n84143, n84144, n84145, n84146, n84147, n84148, n84149, n84150, n84151,
    n84152, n84153, n84154, n84155, n84156, n84157, n84158, n84159, n84160,
    n84161, n84162, n84163, n84164, n84165, n84166, n84167, n84168, n84169,
    n84170, n84171, n84172, n84173, n84174, n84175, n84176, n84177, n84178,
    n84179, n84180, n84181, n84182, n84183, n84184, n84185, n84186, n84187,
    n84188, n84189, n84190, n84191, n84192, n84193, n84194, n84195, n84196,
    n84197, n84198, n84199, n84200, n84201, n84202, n84203, n84204, n84205,
    n84206, n84207, n84208, n84209, n84210, n84211, n84212, n84213, n84214,
    n84215, n84216, n84217, n84218, n84219, n84220, n84221, n84222, n84223,
    n84224, n84225, n84226, n84227, n84228, n84229, n84230, n84231, n84232,
    n84233, n84234, n84235, n84236, n84237, n84238, n84239, n84240, n84241,
    n84242, n84243, n84244, n84245, n84246, n84247, n84248, n84249, n84250,
    n84251, n84252, n84253, n84254, n84255, n84256, n84257, n84258, n84259,
    n84260, n84261, n84262, n84263, n84264, n84265, n84266, n84267, n84268,
    n84269, n84270, n84271, n84272, n84273, n84274, n84275, n84276, n84277,
    n84278, n84279, n84280, n84281, n84282, n84283, n84284, n84285, n84286,
    n84287, n84288, n84289, n84290, n84291, n84292, n84293, n84294, n84295,
    n84296, n84297, n84298, n84299, n84300, n84301, n84302, n84303, n84304,
    n84305, n84306, n84307, n84308, n84309, n84310, n84311, n84312, n84313,
    n84314, n84315, n84316, n84317, n84318, n84319, n84320, n84321, n84322,
    n84323, n84324, n84325, n84326, n84327, n84328, n84329, n84330, n84331,
    n84332, n84333, n84334, n84335, n84336, n84337, n84338, n84339, n84340,
    n84341, n84342, n84343, n84344, n84345, n84346, n84347, n84348, n84349,
    n84350, n84351, n84352, n84353, n84354, n84355, n84356, n84357, n84358,
    n84359, n84360, n84361, n84362, n84363, n84364, n84365, n84366, n84367,
    n84368, n84369, n84370, n84371, n84372, n84373, n84374, n84375, n84376,
    n84377, n84378, n84379, n84380, n84381, n84382, n84383, n84384, n84385,
    n84386, n84387, n84388, n84389, n84390, n84391, n84392, n84393, n84394,
    n84395, n84396, n84397, n84398, n84399, n84400, n84401, n84402, n84403,
    n84404, n84405, n84406, n84407, n84408, n84409, n84410, n84411, n84412,
    n84413, n84414, n84415, n84416, n84417, n84418, n84419, n84420, n84421,
    n84422, n84423, n84424, n84425, n84426, n84427, n84428, n84429, n84430,
    n84431, n84432, n84433, n84434, n84435, n84436, n84437, n84438, n84439,
    n84440, n84441, n84442, n84443, n84444, n84445, n84446, n84447, n84448,
    n84449, n84450, n84451, n84452, n84453, n84454, n84455, n84456, n84457,
    n84458, n84459, n84460, n84461, n84462, n84463, n84464, n84465, n84466,
    n84467, n84468, n84469, n84470, n84471, n84472, n84473, n84474, n84475,
    n84476, n84477, n84478, n84479, n84480, n84481, n84482, n84483, n84484,
    n84485, n84486, n84487, n84488, n84489, n84490, n84491, n84492, n84493,
    n84494, n84495, n84496, n84497, n84498, n84499, n84500, n84501, n84502,
    n84503, n84504, n84505, n84506, n84507, n84508, n84509, n84510, n84511,
    n84512, n84513, n84514, n84515, n84516, n84517, n84518, n84519, n84520,
    n84521, n84522, n84523, n84524, n84525, n84526, n84527, n84528, n84529,
    n84530, n84531, n84532, n84533, n84534, n84535, n84536, n84537, n84538,
    n84539, n84540, n84541, n84542, n84543, n84544, n84545, n84546, n84547,
    n84548, n84549, n84550, n84551, n84552, n84553, n84554, n84555, n84556,
    n84557, n84558, n84559, n84560, n84561, n84562, n84563, n84564, n84565,
    n84566, n84567, n84568, n84569, n84570, n84571, n84572, n84573, n84574,
    n84575, n84576, n84577, n84578, n84579, n84580, n84581, n84582, n84583,
    n84584, n84585, n84586, n84587, n84588, n84589, n84590, n84591, n84592,
    n84593, n84594, n84595, n84596, n84597, n84598, n84599, n84600, n84601,
    n84602, n84603, n84604, n84605, n84606, n84607, n84608, n84609, n84610,
    n84611, n84612, n84613, n84614, n84615, n84616, n84617, n84618, n84619,
    n84620, n84621, n84622, n84623, n84624, n84625, n84626, n84627, n84628,
    n84629, n84630, n84631, n84632, n84633, n84634, n84635, n84636, n84637,
    n84638, n84639, n84640, n84641, n84642, n84643, n84644, n84645, n84646,
    n84647, n84648, n84649, n84650, n84651, n84652, n84653, n84654, n84655,
    n84656, n84657, n84658, n84659, n84660, n84661, n84662, n84663, n84664,
    n84665, n84666, n84667, n84668, n84669, n84670, n84671, n84672, n84673,
    n84674, n84675, n84676, n84677, n84678, n84679, n84680, n84681, n84682,
    n84683, n84684, n84685, n84686, n84687, n84688, n84689, n84690, n84691,
    n84692, n84693, n84694, n84695, n84696, n84697, n84698, n84699, n84700,
    n84701, n84702, n84703, n84704, n84705, n84706, n84707, n84708, n84709,
    n84710, n84711, n84712, n84713, n84714, n84715, n84716, n84717, n84718,
    n84719, n84720, n84721, n84722, n84723, n84724, n84725, n84726, n84727,
    n84728, n84729, n84730, n84731, n84732, n84733, n84734, n84735, n84736,
    n84737, n84738, n84739, n84740, n84741, n84742, n84743, n84744, n84745,
    n84746, n84747, n84748, n84749, n84750, n84751, n84752, n84753, n84754,
    n84755, n84756, n84757, n84758, n84759, n84760, n84761, n84762, n84763,
    n84764, n84765, n84766, n84767, n84768, n84769, n84770, n84771, n84772,
    n84773, n84774, n84775, n84776, n84777, n84778, n84779, n84780, n84781,
    n84782, n84783, n84784, n84785, n84786, n84787, n84788, n84789, n84790,
    n84791, n84792, n84793, n84794, n84795, n84796, n84797, n84798, n84799,
    n84800, n84801, n84802, n84803, n84804, n84805, n84806, n84807, n84808,
    n84809, n84810, n84811, n84812, n84813, n84814, n84815, n84816, n84817,
    n84818, n84819, n84820, n84821, n84822, n84823, n84824, n84825, n84826,
    n84827, n84828, n84829, n84830, n84831, n84832, n84833, n84834, n84835,
    n84836, n84837, n84838, n84839, n84840, n84841, n84842, n84843, n84844,
    n84845, n84846, n84847, n84848, n84849, n84850, n84851, n84852, n84853,
    n84854, n84855, n84856, n84857, n84858, n84859;
  assign n32 = 1'b1;
  assign n33 = pi24 ? n32 : ~n32;
  assign n34 = pi23 ? n32 : n33;
  assign n35 = pi22 ? n34 : n32;
  assign n36 = pi21 ? n35 : n32;
  assign n37 = pi20 ? n36 : n32;
  assign n38 = pi19 ? n37 : n32;
  assign n39 = pi18 ? n32 : n38;
  assign n40 = pi17 ? n32 : n39;
  assign n41 = pi16 ? n32 : n40;
  assign n42 = pi15 ? n32 : n41;
  assign n43 = pi14 ? n42 : n32;
  assign n44 = pi13 ? n43 : n32;
  assign n45 = pi12 ? n32 : n44;
  assign n46 = pi11 ? n32 : n45;
  assign n47 = pi10 ? n32 : n46;
  assign n48 = pi09 ? n32 : n47;
  assign n49 = pi08 ? n48 : n32;
  assign n50 = pi23 ? n33 : ~n32;
  assign n51 = pi22 ? n32 : ~n50;
  assign n52 = pi21 ? n51 : n32;
  assign n53 = pi20 ? n52 : n32;
  assign n54 = pi19 ? n53 : n32;
  assign n55 = pi18 ? n32 : n54;
  assign n56 = pi17 ? n32 : n55;
  assign n57 = pi16 ? n32 : n56;
  assign n58 = pi15 ? n32 : n57;
  assign n59 = pi14 ? n58 : n32;
  assign n60 = pi13 ? n59 : n32;
  assign n61 = pi12 ? n32 : n60;
  assign n62 = pi11 ? n32 : n61;
  assign n63 = pi10 ? n32 : n62;
  assign n64 = pi09 ? n32 : n63;
  assign n65 = pi23 ? n33 : n32;
  assign n66 = pi22 ? n32 : n65;
  assign n67 = pi21 ? n32 : n66;
  assign n68 = pi20 ? n67 : n32;
  assign n69 = pi19 ? n68 : n32;
  assign n70 = pi18 ? n32 : n69;
  assign n71 = pi17 ? n32 : n70;
  assign n72 = pi16 ? n32 : n71;
  assign n73 = pi15 ? n32 : n72;
  assign n74 = pi14 ? n32 : n73;
  assign n75 = pi13 ? n74 : n32;
  assign n76 = pi12 ? n32 : n75;
  assign n77 = pi11 ? n32 : n76;
  assign n78 = pi10 ? n77 : n32;
  assign n79 = pi09 ? n32 : n78;
  assign n80 = pi08 ? n64 : n79;
  assign n81 = pi07 ? n49 : n80;
  assign n82 = pi06 ? n32 : n81;
  assign n83 = pi05 ? n32 : n82;
  assign n84 = pi23 ? n32 : ~n33;
  assign n85 = pi22 ? n84 : n32;
  assign n86 = pi21 ? n32 : n85;
  assign n87 = pi20 ? n86 : n32;
  assign n88 = pi19 ? n87 : n32;
  assign n89 = pi18 ? n32 : n88;
  assign n90 = pi17 ? n32 : n89;
  assign n91 = pi16 ? n32 : n90;
  assign n92 = pi15 ? n32 : n91;
  assign n93 = pi14 ? n32 : n92;
  assign n94 = pi13 ? n32 : n93;
  assign n95 = pi12 ? n94 : n32;
  assign n96 = pi11 ? n32 : n95;
  assign n97 = pi10 ? n32 : n96;
  assign n98 = pi09 ? n32 : n97;
  assign n99 = pi08 ? n32 : n98;
  assign n100 = pi22 ? n32 : n34;
  assign n101 = pi21 ? n32 : n100;
  assign n102 = pi20 ? n101 : n32;
  assign n103 = pi19 ? n102 : n32;
  assign n104 = pi18 ? n32 : n103;
  assign n105 = pi17 ? n32 : n104;
  assign n106 = pi16 ? n32 : n105;
  assign n107 = pi15 ? n106 : n32;
  assign n108 = pi14 ? n32 : n107;
  assign n109 = pi13 ? n108 : n32;
  assign n110 = pi12 ? n32 : n109;
  assign n111 = pi21 ? n32 : n51;
  assign n112 = pi20 ? n111 : n32;
  assign n113 = pi19 ? n112 : n32;
  assign n114 = pi18 ? n32 : n113;
  assign n115 = pi17 ? n32 : n114;
  assign n116 = pi16 ? n32 : n115;
  assign n117 = pi15 ? n32 : n116;
  assign n118 = pi14 ? n117 : n32;
  assign n119 = pi13 ? n32 : n118;
  assign n120 = pi12 ? n119 : n32;
  assign n121 = pi11 ? n110 : n120;
  assign n122 = pi10 ? n32 : n121;
  assign n123 = pi09 ? n32 : n122;
  assign n124 = pi22 ? n65 : n32;
  assign n125 = pi21 ? n124 : n32;
  assign n126 = pi20 ? n32 : n125;
  assign n127 = pi19 ? n32 : n126;
  assign n128 = pi18 ? n127 : n32;
  assign n129 = pi17 ? n32 : n128;
  assign n130 = pi16 ? n129 : n32;
  assign n131 = pi15 ? n130 : n32;
  assign n132 = pi14 ? n131 : n32;
  assign n133 = pi13 ? n32 : n132;
  assign n134 = pi12 ? n32 : n133;
  assign n135 = pi11 ? n32 : n134;
  assign n136 = pi10 ? n32 : n135;
  assign n137 = pi09 ? n32 : n136;
  assign n138 = pi08 ? n123 : n137;
  assign n139 = pi07 ? n99 : n138;
  assign n140 = pi22 ? n50 : ~n32;
  assign n141 = pi21 ? n140 : ~n32;
  assign n142 = pi20 ? n32 : ~n141;
  assign n143 = pi19 ? n142 : n32;
  assign n144 = pi18 ? n32 : n143;
  assign n145 = pi17 ? n32 : n144;
  assign n146 = pi16 ? n32 : n145;
  assign n147 = pi15 ? n146 : n32;
  assign n148 = pi14 ? n32 : n147;
  assign n149 = pi13 ? n148 : n32;
  assign n150 = pi12 ? n32 : n149;
  assign n151 = pi21 ? n32 : n35;
  assign n152 = pi20 ? n151 : n32;
  assign n153 = pi19 ? n152 : n32;
  assign n154 = pi18 ? n32 : n153;
  assign n155 = pi17 ? n32 : n154;
  assign n156 = pi16 ? n32 : n155;
  assign n157 = pi15 ? n32 : n156;
  assign n158 = pi14 ? n73 : n157;
  assign n159 = pi13 ? n32 : n158;
  assign n160 = pi21 ? n32 : ~n140;
  assign n161 = pi20 ? n160 : n32;
  assign n162 = pi19 ? n161 : n32;
  assign n163 = pi18 ? n32 : n162;
  assign n164 = pi17 ? n32 : n163;
  assign n165 = pi16 ? n32 : n164;
  assign n166 = pi15 ? n32 : n165;
  assign n167 = pi14 ? n32 : n166;
  assign n168 = pi13 ? n32 : n167;
  assign n169 = pi12 ? n159 : n168;
  assign n170 = pi11 ? n150 : n169;
  assign n171 = pi10 ? n32 : n170;
  assign n172 = pi09 ? n32 : n171;
  assign n173 = pi23 ? n32 : ~n32;
  assign n174 = pi22 ? n32 : ~n173;
  assign n175 = pi21 ? n32 : n174;
  assign n176 = pi20 ? n175 : n32;
  assign n177 = pi19 ? n176 : n32;
  assign n178 = pi18 ? n32 : n177;
  assign n179 = pi17 ? n32 : n178;
  assign n180 = pi16 ? n32 : n179;
  assign n181 = pi15 ? n32 : n180;
  assign n182 = pi14 ? n181 : n32;
  assign n183 = pi13 ? n32 : n182;
  assign n184 = pi12 ? n183 : n32;
  assign n185 = pi11 ? n32 : n184;
  assign n186 = pi10 ? n32 : n185;
  assign n187 = pi09 ? n32 : n186;
  assign n188 = pi08 ? n172 : n187;
  assign n189 = pi07 ? n188 : n32;
  assign n190 = pi06 ? n139 : n189;
  assign n191 = pi05 ? n32 : n190;
  assign n192 = pi04 ? n83 : n191;
  assign n193 = pi03 ? n32 : n192;
  assign n194 = pi15 ? n72 : n32;
  assign n195 = pi14 ? n32 : n194;
  assign n196 = pi13 ? n32 : n195;
  assign n197 = pi12 ? n32 : n196;
  assign n198 = pi11 ? n32 : n197;
  assign n199 = pi10 ? n32 : n198;
  assign n200 = pi09 ? n32 : n199;
  assign n201 = pi08 ? n32 : n200;
  assign n202 = pi07 ? n32 : n201;
  assign n203 = pi06 ? n32 : n202;
  assign n204 = pi08 ? n200 : n32;
  assign n205 = pi07 ? n204 : n32;
  assign n206 = pi22 ? n32 : ~n32;
  assign n207 = pi21 ? n206 : ~n32;
  assign n208 = pi20 ? n32 : n207;
  assign n209 = pi19 ? n32 : n208;
  assign n210 = pi18 ? n209 : n32;
  assign n211 = pi17 ? n32 : n210;
  assign n212 = pi16 ? n211 : n32;
  assign n213 = pi15 ? n32 : n212;
  assign n214 = pi14 ? n213 : n32;
  assign n215 = pi13 ? n32 : n214;
  assign n216 = pi12 ? n32 : n215;
  assign n217 = pi11 ? n32 : n216;
  assign n218 = pi10 ? n32 : n217;
  assign n219 = pi09 ? n218 : n32;
  assign n220 = pi21 ? n206 : ~n206;
  assign n221 = pi20 ? n32 : n220;
  assign n222 = pi19 ? n32 : n221;
  assign n223 = pi18 ? n222 : n32;
  assign n224 = pi17 ? n32 : n223;
  assign n225 = pi16 ? n224 : n32;
  assign n226 = pi15 ? n32 : n225;
  assign n227 = pi14 ? n213 : n226;
  assign n228 = pi13 ? n32 : n227;
  assign n229 = pi12 ? n32 : n228;
  assign n230 = pi11 ? n32 : n229;
  assign n231 = pi10 ? n32 : n230;
  assign n232 = pi09 ? n231 : n32;
  assign n233 = pi07 ? n219 : n232;
  assign n234 = pi06 ? n205 : n233;
  assign n235 = pi05 ? n203 : n234;
  assign n236 = pi20 ? n207 : ~n32;
  assign n237 = pi19 ? n236 : ~n32;
  assign n238 = pi18 ? n209 : ~n237;
  assign n239 = pi17 ? n32 : n238;
  assign n240 = pi16 ? n239 : n32;
  assign n241 = pi15 ? n32 : n240;
  assign n242 = pi22 ? n34 : ~n32;
  assign n243 = pi21 ? n242 : ~n32;
  assign n244 = pi20 ? n32 : n243;
  assign n245 = pi19 ? n32 : n244;
  assign n246 = pi21 ? n32 : ~n206;
  assign n247 = pi20 ? n246 : n32;
  assign n248 = pi19 ? n247 : n32;
  assign n249 = pi18 ? n245 : n248;
  assign n250 = pi17 ? n32 : n249;
  assign n251 = pi16 ? n250 : n32;
  assign n252 = pi15 ? n240 : n251;
  assign n253 = pi14 ? n241 : n252;
  assign n254 = pi13 ? n32 : n253;
  assign n255 = pi12 ? n32 : n254;
  assign n256 = pi11 ? n32 : n255;
  assign n257 = pi10 ? n32 : n256;
  assign n258 = pi15 ? n240 : n225;
  assign n259 = pi22 ? n173 : ~n32;
  assign n260 = pi21 ? n259 : ~n206;
  assign n261 = pi20 ? n32 : n260;
  assign n262 = pi19 ? n32 : n261;
  assign n263 = pi18 ? n262 : n32;
  assign n264 = pi17 ? n32 : n263;
  assign n265 = pi16 ? n264 : n32;
  assign n266 = pi21 ? n206 : n32;
  assign n267 = pi20 ? n32 : n266;
  assign n268 = pi19 ? n32 : n267;
  assign n269 = pi18 ? n268 : n32;
  assign n270 = pi17 ? n32 : n269;
  assign n271 = pi16 ? n270 : n32;
  assign n272 = pi15 ? n265 : n271;
  assign n273 = pi14 ? n258 : n272;
  assign n274 = pi21 ? n174 : n32;
  assign n275 = pi20 ? n32 : n274;
  assign n276 = pi19 ? n32 : n275;
  assign n277 = pi18 ? n276 : n32;
  assign n278 = pi17 ? n32 : n277;
  assign n279 = pi16 ? n278 : n32;
  assign n280 = pi15 ? n32 : n279;
  assign n281 = pi14 ? n280 : n32;
  assign n282 = pi13 ? n273 : n281;
  assign n283 = pi12 ? n282 : n32;
  assign n284 = pi11 ? n283 : n32;
  assign n285 = pi10 ? n284 : n32;
  assign n286 = pi09 ? n257 : n285;
  assign n287 = pi21 ? n206 : n259;
  assign n288 = pi20 ? n287 : ~n32;
  assign n289 = pi19 ? n288 : ~n32;
  assign n290 = pi18 ? n209 : ~n289;
  assign n291 = pi17 ? n32 : n290;
  assign n292 = pi16 ? n291 : n32;
  assign n293 = pi15 ? n292 : n225;
  assign n294 = pi14 ? n293 : n272;
  assign n295 = pi21 ? n140 : n173;
  assign n296 = pi20 ? n32 : n295;
  assign n297 = pi19 ? n32 : n296;
  assign n298 = pi18 ? n297 : n32;
  assign n299 = pi17 ? n32 : n298;
  assign n300 = pi16 ? n299 : n32;
  assign n301 = pi15 ? n32 : n300;
  assign n302 = pi14 ? n301 : n32;
  assign n303 = pi13 ? n294 : n302;
  assign n304 = pi12 ? n303 : n32;
  assign n305 = pi11 ? n304 : n32;
  assign n306 = pi10 ? n305 : n32;
  assign n307 = pi09 ? n257 : n306;
  assign n308 = pi08 ? n286 : n307;
  assign n309 = pi22 ? n173 : n32;
  assign n310 = pi21 ? n206 : n309;
  assign n311 = pi20 ? n32 : n310;
  assign n312 = pi19 ? n32 : n311;
  assign n313 = pi22 ? n173 : ~n173;
  assign n314 = pi21 ? n313 : ~n32;
  assign n315 = pi20 ? n314 : ~n32;
  assign n316 = pi19 ? n315 : ~n32;
  assign n317 = pi18 ? n312 : ~n316;
  assign n318 = pi17 ? n32 : n317;
  assign n319 = pi16 ? n318 : n32;
  assign n320 = pi15 ? n32 : n319;
  assign n321 = pi21 ? n32 : ~n32;
  assign n322 = pi20 ? n32 : n321;
  assign n323 = pi19 ? n322 : ~n32;
  assign n324 = pi18 ? n245 : ~n323;
  assign n325 = pi17 ? n32 : n324;
  assign n326 = pi16 ? n325 : n32;
  assign n327 = pi15 ? n326 : n279;
  assign n328 = pi14 ? n320 : n327;
  assign n329 = pi13 ? n32 : n328;
  assign n330 = pi12 ? n32 : n329;
  assign n331 = pi11 ? n32 : n330;
  assign n332 = pi10 ? n32 : n331;
  assign n333 = pi21 ? n174 : n309;
  assign n334 = pi20 ? n32 : n333;
  assign n335 = pi19 ? n32 : n334;
  assign n336 = pi18 ? n335 : n32;
  assign n337 = pi17 ? n32 : n336;
  assign n338 = pi16 ? n337 : n32;
  assign n339 = pi21 ? n259 : ~n32;
  assign n340 = pi20 ? n32 : n339;
  assign n341 = pi19 ? n32 : n340;
  assign n342 = pi21 ? n32 : n206;
  assign n343 = pi20 ? n342 : ~n32;
  assign n344 = pi19 ? n343 : ~n32;
  assign n345 = pi18 ? n341 : ~n344;
  assign n346 = pi17 ? n32 : n345;
  assign n347 = pi16 ? n346 : n32;
  assign n348 = pi15 ? n338 : n347;
  assign n349 = pi20 ? n321 : ~n32;
  assign n350 = pi19 ? n349 : ~n32;
  assign n351 = pi18 ? n262 : ~n350;
  assign n352 = pi17 ? n32 : n351;
  assign n353 = pi16 ? n352 : n32;
  assign n354 = pi21 ? n259 : ~n174;
  assign n355 = pi20 ? n32 : n354;
  assign n356 = pi19 ? n32 : n355;
  assign n357 = pi21 ? n309 : n32;
  assign n358 = pi20 ? n357 : n32;
  assign n359 = pi19 ? n358 : n32;
  assign n360 = pi18 ? n356 : n359;
  assign n361 = pi17 ? n32 : n360;
  assign n362 = pi16 ? n361 : n32;
  assign n363 = pi15 ? n353 : n362;
  assign n364 = pi14 ? n348 : n363;
  assign n365 = pi20 ? n32 : n141;
  assign n366 = pi19 ? n32 : n365;
  assign n367 = pi18 ? n366 : n32;
  assign n368 = pi17 ? n32 : n367;
  assign n369 = pi16 ? n368 : n32;
  assign n370 = pi15 ? n369 : n32;
  assign n371 = pi21 ? n259 : n309;
  assign n372 = pi20 ? n32 : n371;
  assign n373 = pi19 ? n32 : n372;
  assign n374 = pi18 ? n373 : n32;
  assign n375 = pi17 ? n32 : n374;
  assign n376 = pi16 ? n375 : n32;
  assign n377 = pi15 ? n32 : n376;
  assign n378 = pi14 ? n370 : n377;
  assign n379 = pi13 ? n364 : n378;
  assign n380 = pi12 ? n379 : n32;
  assign n381 = pi11 ? n380 : n32;
  assign n382 = pi21 ? n32 : n124;
  assign n383 = pi20 ? n32 : n382;
  assign n384 = pi19 ? n383 : n32;
  assign n385 = pi18 ? n32 : n384;
  assign n386 = pi17 ? n32 : n385;
  assign n387 = pi16 ? n32 : n386;
  assign n388 = pi15 ? n387 : n32;
  assign n389 = pi14 ? n32 : n388;
  assign n390 = pi13 ? n32 : n389;
  assign n391 = pi12 ? n32 : n390;
  assign n392 = pi11 ? n391 : n32;
  assign n393 = pi10 ? n381 : n392;
  assign n394 = pi09 ? n332 : n393;
  assign n395 = pi21 ? n259 : ~n173;
  assign n396 = pi20 ? n32 : ~n395;
  assign n397 = pi19 ? n396 : ~n32;
  assign n398 = pi18 ? n245 : ~n397;
  assign n399 = pi17 ? n32 : n398;
  assign n400 = pi16 ? n399 : n32;
  assign n401 = pi15 ? n32 : n400;
  assign n402 = pi21 ? n242 : ~n309;
  assign n403 = pi20 ? n32 : n402;
  assign n404 = pi19 ? n32 : n403;
  assign n405 = pi22 ? n32 : n173;
  assign n406 = pi21 ? n313 : n405;
  assign n407 = pi20 ? n406 : n357;
  assign n408 = pi19 ? n407 : n32;
  assign n409 = pi18 ? n404 : n408;
  assign n410 = pi17 ? n32 : n409;
  assign n411 = pi16 ? n410 : n32;
  assign n412 = pi15 ? n326 : n411;
  assign n413 = pi14 ? n401 : n412;
  assign n414 = pi13 ? n32 : n413;
  assign n415 = pi12 ? n32 : n414;
  assign n416 = pi11 ? n32 : n415;
  assign n417 = pi10 ? n32 : n416;
  assign n418 = pi19 ? n340 : ~n32;
  assign n419 = pi18 ? n341 : ~n418;
  assign n420 = pi17 ? n32 : n419;
  assign n421 = pi16 ? n420 : n32;
  assign n422 = pi20 ? n175 : ~n32;
  assign n423 = pi19 ? n422 : ~n32;
  assign n424 = pi18 ? n341 : ~n423;
  assign n425 = pi17 ? n32 : n424;
  assign n426 = pi16 ? n425 : n32;
  assign n427 = pi15 ? n421 : n426;
  assign n428 = pi21 ? n32 : n405;
  assign n429 = pi20 ? n428 : ~n32;
  assign n430 = pi19 ? n429 : ~n32;
  assign n431 = pi18 ? n341 : ~n430;
  assign n432 = pi17 ? n32 : n431;
  assign n433 = pi16 ? n432 : n32;
  assign n434 = pi18 ? n341 : ~n350;
  assign n435 = pi17 ? n32 : n434;
  assign n436 = pi16 ? n435 : n32;
  assign n437 = pi15 ? n433 : n436;
  assign n438 = pi14 ? n427 : n437;
  assign n439 = pi21 ? n313 : n32;
  assign n440 = pi20 ? n439 : n32;
  assign n441 = pi19 ? n440 : n32;
  assign n442 = pi18 ? n341 : n441;
  assign n443 = pi17 ? n32 : n442;
  assign n444 = pi16 ? n443 : n32;
  assign n445 = pi15 ? n444 : n369;
  assign n446 = pi14 ? n445 : n369;
  assign n447 = pi13 ? n438 : n446;
  assign n448 = pi21 ? n173 : n32;
  assign n449 = pi20 ? n32 : n448;
  assign n450 = pi19 ? n32 : n449;
  assign n451 = pi18 ? n450 : n32;
  assign n452 = pi17 ? n32 : n451;
  assign n453 = pi16 ? n452 : n32;
  assign n454 = pi22 ? n65 : ~n173;
  assign n455 = pi21 ? n454 : n32;
  assign n456 = pi20 ? n32 : n455;
  assign n457 = pi19 ? n32 : n456;
  assign n458 = pi18 ? n457 : n32;
  assign n459 = pi17 ? n32 : n458;
  assign n460 = pi16 ? n459 : n32;
  assign n461 = pi15 ? n453 : n460;
  assign n462 = pi20 ? n32 : n357;
  assign n463 = pi19 ? n32 : n462;
  assign n464 = pi18 ? n463 : n32;
  assign n465 = pi17 ? n32 : n464;
  assign n466 = pi16 ? n465 : n32;
  assign n467 = pi15 ? n460 : n466;
  assign n468 = pi14 ? n461 : n467;
  assign n469 = pi13 ? n468 : n32;
  assign n470 = pi12 ? n447 : n469;
  assign n471 = pi11 ? n470 : n32;
  assign n472 = pi20 ? n32 : n151;
  assign n473 = pi19 ? n472 : n32;
  assign n474 = pi18 ? n32 : n473;
  assign n475 = pi17 ? n32 : n474;
  assign n476 = pi16 ? n32 : n475;
  assign n477 = pi15 ? n476 : n32;
  assign n478 = pi14 ? n477 : n32;
  assign n479 = pi13 ? n478 : n32;
  assign n480 = pi12 ? n32 : n479;
  assign n481 = pi21 ? n85 : n32;
  assign n482 = pi20 ? n32 : n481;
  assign n483 = pi19 ? n482 : n32;
  assign n484 = pi18 ? n32 : n483;
  assign n485 = pi17 ? n32 : n484;
  assign n486 = pi16 ? n32 : n485;
  assign n487 = pi15 ? n32 : n486;
  assign n488 = pi14 ? n487 : n32;
  assign n489 = pi13 ? n32 : n488;
  assign n490 = pi12 ? n32 : n489;
  assign n491 = pi11 ? n480 : n490;
  assign n492 = pi10 ? n471 : n491;
  assign n493 = pi09 ? n417 : n492;
  assign n494 = pi08 ? n394 : n493;
  assign n495 = pi07 ? n308 : n494;
  assign n496 = pi19 ? n32 : n349;
  assign n497 = pi18 ? n245 : ~n496;
  assign n498 = pi17 ? n32 : n497;
  assign n499 = pi16 ? n498 : n32;
  assign n500 = pi15 ? n32 : n499;
  assign n501 = pi21 ? n174 : ~n32;
  assign n502 = pi20 ? n501 : ~n32;
  assign n503 = pi19 ? n32 : n502;
  assign n504 = pi18 ? n209 : ~n503;
  assign n505 = pi17 ? n32 : n504;
  assign n506 = pi16 ? n505 : n32;
  assign n507 = pi20 ? n32 : n342;
  assign n508 = pi19 ? n507 : ~n32;
  assign n509 = pi18 ? n245 : ~n508;
  assign n510 = pi17 ? n32 : n509;
  assign n511 = pi16 ? n510 : n32;
  assign n512 = pi15 ? n506 : n511;
  assign n513 = pi14 ? n500 : n512;
  assign n514 = pi13 ? n32 : n513;
  assign n515 = pi12 ? n32 : n514;
  assign n516 = pi11 ? n32 : n515;
  assign n517 = pi10 ? n32 : n516;
  assign n518 = pi21 ? n32 : n259;
  assign n519 = pi20 ? n32 : n518;
  assign n520 = pi19 ? n519 : ~n32;
  assign n521 = pi18 ? n341 : ~n520;
  assign n522 = pi17 ? n32 : n521;
  assign n523 = pi16 ? n522 : n32;
  assign n524 = pi18 ? n341 : ~n508;
  assign n525 = pi17 ? n32 : n524;
  assign n526 = pi16 ? n525 : n32;
  assign n527 = pi15 ? n523 : n526;
  assign n528 = pi18 ? n341 : ~n323;
  assign n529 = pi17 ? n32 : n528;
  assign n530 = pi16 ? n529 : n32;
  assign n531 = pi20 ? n32 : ~n32;
  assign n532 = pi19 ? n531 : ~n32;
  assign n533 = pi18 ? n366 : ~n532;
  assign n534 = pi17 ? n32 : n533;
  assign n535 = pi16 ? n534 : n32;
  assign n536 = pi15 ? n530 : n535;
  assign n537 = pi14 ? n527 : n536;
  assign n538 = pi18 ? n366 : ~n430;
  assign n539 = pi17 ? n32 : n538;
  assign n540 = pi16 ? n539 : n32;
  assign n541 = pi15 ? n535 : n540;
  assign n542 = pi18 ? n366 : ~n344;
  assign n543 = pi17 ? n32 : n542;
  assign n544 = pi16 ? n543 : n32;
  assign n545 = pi18 ? n366 : ~n350;
  assign n546 = pi17 ? n32 : n545;
  assign n547 = pi16 ? n546 : n32;
  assign n548 = pi15 ? n544 : n547;
  assign n549 = pi14 ? n541 : n548;
  assign n550 = pi13 ? n537 : n549;
  assign n551 = pi18 ? n341 : n32;
  assign n552 = pi17 ? n32 : n551;
  assign n553 = pi16 ? n552 : n32;
  assign n554 = pi18 ? n356 : n32;
  assign n555 = pi17 ? n32 : n554;
  assign n556 = pi16 ? n555 : n32;
  assign n557 = pi15 ? n553 : n556;
  assign n558 = pi21 ? n140 : ~n174;
  assign n559 = pi20 ? n32 : n558;
  assign n560 = pi19 ? n32 : n559;
  assign n561 = pi18 ? n560 : n32;
  assign n562 = pi17 ? n32 : n561;
  assign n563 = pi16 ? n562 : n32;
  assign n564 = pi21 ? n140 : n32;
  assign n565 = pi20 ? n32 : n564;
  assign n566 = pi19 ? n32 : n565;
  assign n567 = pi18 ? n566 : n32;
  assign n568 = pi17 ? n32 : n567;
  assign n569 = pi16 ? n568 : n32;
  assign n570 = pi15 ? n563 : n569;
  assign n571 = pi14 ? n557 : n570;
  assign n572 = pi20 ? n32 : n439;
  assign n573 = pi19 ? n32 : n572;
  assign n574 = pi18 ? n573 : n32;
  assign n575 = pi17 ? n32 : n574;
  assign n576 = pi16 ? n575 : n32;
  assign n577 = pi15 ? n569 : n576;
  assign n578 = pi15 ? n466 : n32;
  assign n579 = pi14 ? n577 : n578;
  assign n580 = pi13 ? n571 : n579;
  assign n581 = pi12 ? n550 : n580;
  assign n582 = pi11 ? n581 : n32;
  assign n583 = pi10 ? n582 : n32;
  assign n584 = pi09 ? n517 : n583;
  assign n585 = pi18 ? n209 : ~n496;
  assign n586 = pi17 ? n32 : n585;
  assign n587 = pi16 ? n586 : n32;
  assign n588 = pi15 ? n32 : n587;
  assign n589 = pi20 ? n518 : ~n32;
  assign n590 = pi19 ? n32 : n589;
  assign n591 = pi18 ? n245 : ~n590;
  assign n592 = pi17 ? n32 : n591;
  assign n593 = pi16 ? n592 : n32;
  assign n594 = pi20 ? n32 : n428;
  assign n595 = pi19 ? n594 : ~n32;
  assign n596 = pi18 ? n245 : ~n595;
  assign n597 = pi17 ? n32 : n596;
  assign n598 = pi16 ? n597 : n32;
  assign n599 = pi15 ? n593 : n598;
  assign n600 = pi14 ? n588 : n599;
  assign n601 = pi13 ? n32 : n600;
  assign n602 = pi12 ? n32 : n601;
  assign n603 = pi11 ? n32 : n602;
  assign n604 = pi10 ? n32 : n603;
  assign n605 = pi19 ? n208 : ~n32;
  assign n606 = pi18 ? n366 : ~n605;
  assign n607 = pi17 ? n32 : n606;
  assign n608 = pi16 ? n607 : n32;
  assign n609 = pi15 ? n530 : n608;
  assign n610 = pi14 ? n526 : n609;
  assign n611 = pi15 ? n347 : n436;
  assign n612 = pi14 ? n535 : n611;
  assign n613 = pi13 ? n610 : n612;
  assign n614 = pi18 ? n366 : ~n237;
  assign n615 = pi17 ? n32 : n614;
  assign n616 = pi16 ? n615 : n32;
  assign n617 = pi20 ? n339 : ~n32;
  assign n618 = pi19 ? n617 : ~n32;
  assign n619 = pi18 ? n366 : ~n618;
  assign n620 = pi17 ? n32 : n619;
  assign n621 = pi16 ? n620 : n32;
  assign n622 = pi15 ? n616 : n621;
  assign n623 = pi21 ? n259 : ~n259;
  assign n624 = pi20 ? n32 : n623;
  assign n625 = pi19 ? n32 : n624;
  assign n626 = pi18 ? n625 : n32;
  assign n627 = pi17 ? n32 : n626;
  assign n628 = pi16 ? n627 : n32;
  assign n629 = pi15 ? n621 : n628;
  assign n630 = pi14 ? n622 : n629;
  assign n631 = pi22 ? n50 : ~n173;
  assign n632 = pi21 ? n631 : n32;
  assign n633 = pi20 ? n32 : n632;
  assign n634 = pi19 ? n32 : n633;
  assign n635 = pi18 ? n634 : n32;
  assign n636 = pi17 ? n32 : n635;
  assign n637 = pi16 ? n636 : n32;
  assign n638 = pi15 ? n569 : n637;
  assign n639 = pi15 ? n637 : n32;
  assign n640 = pi14 ? n638 : n639;
  assign n641 = pi13 ? n630 : n640;
  assign n642 = pi12 ? n613 : n641;
  assign n643 = pi11 ? n642 : n32;
  assign n644 = pi20 ? n32 : n111;
  assign n645 = pi19 ? n644 : n32;
  assign n646 = pi18 ? n32 : n645;
  assign n647 = pi17 ? n32 : n646;
  assign n648 = pi16 ? n32 : n647;
  assign n649 = pi15 ? n648 : n32;
  assign n650 = pi14 ? n649 : n32;
  assign n651 = pi13 ? n650 : n32;
  assign n652 = pi12 ? n32 : n651;
  assign n653 = pi21 ? n100 : n32;
  assign n654 = pi20 ? n32 : n653;
  assign n655 = pi19 ? n654 : n32;
  assign n656 = pi18 ? n32 : n655;
  assign n657 = pi17 ? n32 : n656;
  assign n658 = pi16 ? n32 : n657;
  assign n659 = pi15 ? n32 : n658;
  assign n660 = pi14 ? n32 : n659;
  assign n661 = pi13 ? n660 : n32;
  assign n662 = pi20 ? n32 : n36;
  assign n663 = pi19 ? n662 : n32;
  assign n664 = pi18 ? n32 : n663;
  assign n665 = pi17 ? n32 : n664;
  assign n666 = pi16 ? n32 : n665;
  assign n667 = pi15 ? n32 : n666;
  assign n668 = pi19 ? n126 : n32;
  assign n669 = pi18 ? n32 : n668;
  assign n670 = pi17 ? n32 : n669;
  assign n671 = pi16 ? n32 : n670;
  assign n672 = pi15 ? n671 : n32;
  assign n673 = pi14 ? n667 : n672;
  assign n674 = pi13 ? n32 : n673;
  assign n675 = pi12 ? n661 : n674;
  assign n676 = pi11 ? n652 : n675;
  assign n677 = pi10 ? n643 : n676;
  assign n678 = pi09 ? n604 : n677;
  assign n679 = pi08 ? n584 : n678;
  assign n680 = pi18 ? n245 : ~n209;
  assign n681 = pi17 ? n32 : n680;
  assign n682 = pi16 ? n681 : n32;
  assign n683 = pi15 ? n32 : n682;
  assign n684 = pi19 ? n32 : n343;
  assign n685 = pi18 ? n245 : ~n684;
  assign n686 = pi17 ? n32 : n685;
  assign n687 = pi16 ? n686 : n32;
  assign n688 = pi15 ? n682 : n687;
  assign n689 = pi14 ? n683 : n688;
  assign n690 = pi13 ? n32 : n689;
  assign n691 = pi12 ? n32 : n690;
  assign n692 = pi11 ? n32 : n691;
  assign n693 = pi10 ? n32 : n692;
  assign n694 = pi18 ? n341 : ~n590;
  assign n695 = pi17 ? n32 : n694;
  assign n696 = pi16 ? n695 : n32;
  assign n697 = pi19 ? n32 : n236;
  assign n698 = pi18 ? n341 : ~n697;
  assign n699 = pi17 ? n32 : n698;
  assign n700 = pi16 ? n699 : n32;
  assign n701 = pi15 ? n696 : n700;
  assign n702 = pi19 ? n32 : ~n32;
  assign n703 = pi18 ? n341 : ~n702;
  assign n704 = pi17 ? n32 : n703;
  assign n705 = pi16 ? n704 : n32;
  assign n706 = pi18 ? n366 : ~n508;
  assign n707 = pi17 ? n32 : n706;
  assign n708 = pi16 ? n707 : n32;
  assign n709 = pi15 ? n705 : n708;
  assign n710 = pi14 ? n701 : n709;
  assign n711 = pi18 ? n341 : ~n605;
  assign n712 = pi17 ? n32 : n711;
  assign n713 = pi16 ? n712 : n32;
  assign n714 = pi15 ? n708 : n713;
  assign n715 = pi14 ? n714 : n608;
  assign n716 = pi13 ? n710 : n715;
  assign n717 = pi18 ? n341 : ~n237;
  assign n718 = pi17 ? n32 : n717;
  assign n719 = pi16 ? n718 : n32;
  assign n720 = pi15 ? n544 : n719;
  assign n721 = pi14 ? n535 : n720;
  assign n722 = pi18 ? n341 : ~n618;
  assign n723 = pi17 ? n32 : n722;
  assign n724 = pi16 ? n723 : n32;
  assign n725 = pi15 ? n724 : n621;
  assign n726 = pi21 ? n140 : ~n206;
  assign n727 = pi20 ? n32 : n726;
  assign n728 = pi19 ? n32 : n727;
  assign n729 = pi18 ? n728 : n32;
  assign n730 = pi17 ? n32 : n729;
  assign n731 = pi16 ? n730 : n32;
  assign n732 = pi15 ? n731 : n576;
  assign n733 = pi14 ? n725 : n732;
  assign n734 = pi13 ? n721 : n733;
  assign n735 = pi12 ? n716 : n734;
  assign n736 = pi11 ? n735 : n32;
  assign n737 = pi15 ? n32 : n476;
  assign n738 = pi14 ? n737 : n32;
  assign n739 = pi13 ? n32 : n738;
  assign n740 = pi12 ? n32 : n739;
  assign n741 = pi16 ? n129 : n485;
  assign n742 = pi15 ? n741 : n32;
  assign n743 = pi14 ? n32 : n742;
  assign n744 = pi13 ? n32 : n743;
  assign n745 = pi12 ? n32 : n744;
  assign n746 = pi11 ? n740 : n745;
  assign n747 = pi10 ? n736 : n746;
  assign n748 = pi09 ? n693 : n747;
  assign n749 = pi21 ? n405 : ~n32;
  assign n750 = pi20 ? n32 : n749;
  assign n751 = pi19 ? n32 : n750;
  assign n752 = pi18 ? n245 : ~n751;
  assign n753 = pi17 ? n32 : n752;
  assign n754 = pi16 ? n753 : n32;
  assign n755 = pi15 ? n32 : n754;
  assign n756 = pi18 ? n245 : ~n341;
  assign n757 = pi17 ? n32 : n756;
  assign n758 = pi16 ? n757 : n32;
  assign n759 = pi15 ? n682 : n758;
  assign n760 = pi14 ? n755 : n759;
  assign n761 = pi13 ? n32 : n760;
  assign n762 = pi12 ? n32 : n761;
  assign n763 = pi11 ? n32 : n762;
  assign n764 = pi10 ? n32 : n763;
  assign n765 = pi21 ? n405 : n259;
  assign n766 = pi20 ? n765 : ~n32;
  assign n767 = pi19 ? n32 : n766;
  assign n768 = pi18 ? n341 : ~n767;
  assign n769 = pi17 ? n32 : n768;
  assign n770 = pi16 ? n769 : n32;
  assign n771 = pi15 ? n696 : n770;
  assign n772 = pi19 ? n32 : ~n358;
  assign n773 = pi18 ? n341 : ~n772;
  assign n774 = pi17 ? n32 : n773;
  assign n775 = pi16 ? n774 : n32;
  assign n776 = pi19 ? n594 : n617;
  assign n777 = pi18 ? n366 : ~n776;
  assign n778 = pi17 ? n32 : n777;
  assign n779 = pi16 ? n778 : n32;
  assign n780 = pi15 ? n775 : n779;
  assign n781 = pi14 ? n771 : n780;
  assign n782 = pi18 ? n366 : ~n595;
  assign n783 = pi17 ? n32 : n782;
  assign n784 = pi16 ? n783 : n32;
  assign n785 = pi21 ? n206 : ~n309;
  assign n786 = pi20 ? n32 : n785;
  assign n787 = pi19 ? n786 : ~n32;
  assign n788 = pi18 ? n366 : ~n787;
  assign n789 = pi17 ? n32 : n788;
  assign n790 = pi16 ? n789 : n32;
  assign n791 = pi15 ? n784 : n790;
  assign n792 = pi20 ? n32 : n765;
  assign n793 = pi19 ? n792 : ~n32;
  assign n794 = pi18 ? n366 : ~n793;
  assign n795 = pi17 ? n32 : n794;
  assign n796 = pi16 ? n795 : n32;
  assign n797 = pi19 ? n750 : ~n32;
  assign n798 = pi18 ? n366 : ~n797;
  assign n799 = pi17 ? n32 : n798;
  assign n800 = pi16 ? n799 : n32;
  assign n801 = pi15 ? n796 : n800;
  assign n802 = pi14 ? n791 : n801;
  assign n803 = pi13 ? n781 : n802;
  assign n804 = pi20 ? n32 : ~n357;
  assign n805 = pi19 ? n804 : ~n32;
  assign n806 = pi18 ? n366 : ~n805;
  assign n807 = pi17 ? n32 : n806;
  assign n808 = pi16 ? n807 : n32;
  assign n809 = pi18 ? n341 : ~n532;
  assign n810 = pi17 ? n32 : n809;
  assign n811 = pi16 ? n810 : n32;
  assign n812 = pi15 ? n808 : n811;
  assign n813 = pi20 ? n749 : ~n32;
  assign n814 = pi19 ? n813 : ~n32;
  assign n815 = pi18 ? n366 : ~n814;
  assign n816 = pi17 ? n32 : n815;
  assign n817 = pi16 ? n816 : n32;
  assign n818 = pi15 ? n347 : n817;
  assign n819 = pi14 ? n812 : n818;
  assign n820 = pi21 ? n173 : ~n32;
  assign n821 = pi20 ? n820 : ~n32;
  assign n822 = pi19 ? n821 : ~n32;
  assign n823 = pi18 ? n366 : ~n822;
  assign n824 = pi17 ? n32 : n823;
  assign n825 = pi16 ? n824 : n32;
  assign n826 = pi19 ? n766 : ~n32;
  assign n827 = pi18 ? n366 : ~n826;
  assign n828 = pi17 ? n32 : n827;
  assign n829 = pi16 ? n828 : n32;
  assign n830 = pi15 ? n825 : n829;
  assign n831 = pi21 ? n259 : ~n405;
  assign n832 = pi20 ? n32 : n831;
  assign n833 = pi19 ? n32 : n832;
  assign n834 = pi18 ? n833 : n32;
  assign n835 = pi17 ? n32 : n834;
  assign n836 = pi16 ? n835 : n32;
  assign n837 = pi21 ? n140 : n309;
  assign n838 = pi20 ? n32 : n837;
  assign n839 = pi19 ? n32 : n838;
  assign n840 = pi18 ? n839 : n32;
  assign n841 = pi17 ? n32 : n840;
  assign n842 = pi16 ? n841 : n32;
  assign n843 = pi15 ? n836 : n842;
  assign n844 = pi14 ? n830 : n843;
  assign n845 = pi13 ? n819 : n844;
  assign n846 = pi12 ? n803 : n845;
  assign n847 = pi15 ? n453 : n130;
  assign n848 = pi14 ? n847 : n32;
  assign n849 = pi13 ? n848 : n32;
  assign n850 = pi12 ? n849 : n32;
  assign n851 = pi11 ? n846 : n850;
  assign n852 = pi10 ? n851 : n135;
  assign n853 = pi09 ? n764 : n852;
  assign n854 = pi08 ? n748 : n853;
  assign n855 = pi07 ? n679 : n854;
  assign n856 = pi06 ? n495 : n855;
  assign n857 = pi20 ? n32 : n175;
  assign n858 = pi19 ? n32 : n857;
  assign n859 = pi18 ? n245 : ~n858;
  assign n860 = pi17 ? n32 : n859;
  assign n861 = pi16 ? n860 : n32;
  assign n862 = pi15 ? n32 : n861;
  assign n863 = pi19 ? n32 : n507;
  assign n864 = pi18 ? n245 : ~n863;
  assign n865 = pi17 ? n32 : n864;
  assign n866 = pi16 ? n865 : n32;
  assign n867 = pi15 ? n866 : n754;
  assign n868 = pi14 ? n862 : n867;
  assign n869 = pi13 ? n32 : n868;
  assign n870 = pi12 ? n32 : n869;
  assign n871 = pi11 ? n32 : n870;
  assign n872 = pi10 ? n32 : n871;
  assign n873 = pi18 ? n341 : ~n209;
  assign n874 = pi17 ? n32 : n873;
  assign n875 = pi16 ? n874 : n32;
  assign n876 = pi18 ? n341 : ~n341;
  assign n877 = pi17 ? n32 : n876;
  assign n878 = pi16 ? n877 : n32;
  assign n879 = pi15 ? n875 : n878;
  assign n880 = pi19 ? n32 : n531;
  assign n881 = pi18 ? n341 : ~n880;
  assign n882 = pi17 ? n32 : n881;
  assign n883 = pi16 ? n882 : n32;
  assign n884 = pi18 ? n366 : ~n684;
  assign n885 = pi17 ? n32 : n884;
  assign n886 = pi16 ? n885 : n32;
  assign n887 = pi15 ? n883 : n886;
  assign n888 = pi14 ? n879 : n887;
  assign n889 = pi18 ? n341 : ~n496;
  assign n890 = pi17 ? n32 : n889;
  assign n891 = pi16 ? n890 : n32;
  assign n892 = pi18 ? n366 : ~n697;
  assign n893 = pi17 ? n32 : n892;
  assign n894 = pi16 ? n893 : n32;
  assign n895 = pi15 ? n891 : n894;
  assign n896 = pi18 ? n366 : ~n702;
  assign n897 = pi17 ? n32 : n896;
  assign n898 = pi16 ? n897 : n32;
  assign n899 = pi14 ? n895 : n898;
  assign n900 = pi13 ? n888 : n899;
  assign n901 = pi18 ? n366 : ~n323;
  assign n902 = pi17 ? n32 : n901;
  assign n903 = pi16 ? n902 : n32;
  assign n904 = pi15 ? n526 : n903;
  assign n905 = pi15 ? n903 : n608;
  assign n906 = pi14 ? n904 : n905;
  assign n907 = pi15 ? n608 : n544;
  assign n908 = pi15 ? n719 : n553;
  assign n909 = pi14 ? n907 : n908;
  assign n910 = pi13 ? n906 : n909;
  assign n911 = pi12 ? n900 : n910;
  assign n912 = pi15 ? n369 : n553;
  assign n913 = pi15 ? n369 : n731;
  assign n914 = pi14 ? n912 : n913;
  assign n915 = pi21 ? n259 : n32;
  assign n916 = pi20 ? n32 : n915;
  assign n917 = pi19 ? n32 : n916;
  assign n918 = pi18 ? n917 : n32;
  assign n919 = pi17 ? n32 : n918;
  assign n920 = pi16 ? n919 : n32;
  assign n921 = pi15 ? n920 : n569;
  assign n922 = pi14 ? n921 : n466;
  assign n923 = pi13 ? n914 : n922;
  assign n924 = pi14 ? n578 : n32;
  assign n925 = pi13 ? n924 : n32;
  assign n926 = pi12 ? n923 : n925;
  assign n927 = pi11 ? n911 : n926;
  assign n928 = pi10 ? n927 : n32;
  assign n929 = pi09 ? n872 : n928;
  assign n930 = pi18 ? n245 : ~n32;
  assign n931 = pi17 ? n32 : n930;
  assign n932 = pi18 ? n822 : ~n32;
  assign n933 = pi17 ? n932 : ~n32;
  assign n934 = pi16 ? n931 : ~n933;
  assign n935 = pi15 ? n32 : n934;
  assign n936 = pi19 ? n32 : n594;
  assign n937 = pi18 ? n245 : ~n936;
  assign n938 = pi17 ? n32 : n937;
  assign n939 = pi16 ? n938 : n32;
  assign n940 = pi19 ? n32 : n322;
  assign n941 = pi18 ? n245 : ~n940;
  assign n942 = pi17 ? n32 : n941;
  assign n943 = pi16 ? n942 : n32;
  assign n944 = pi15 ? n939 : n943;
  assign n945 = pi14 ? n935 : n944;
  assign n946 = pi13 ? n32 : n945;
  assign n947 = pi12 ? n32 : n946;
  assign n948 = pi11 ? n32 : n947;
  assign n949 = pi10 ? n32 : n948;
  assign n950 = pi18 ? n341 : ~n751;
  assign n951 = pi17 ? n32 : n950;
  assign n952 = pi16 ? n951 : n32;
  assign n953 = pi15 ? n952 : n878;
  assign n954 = pi18 ? n341 : ~n684;
  assign n955 = pi17 ? n32 : n954;
  assign n956 = pi16 ? n955 : n32;
  assign n957 = pi15 ? n883 : n956;
  assign n958 = pi14 ? n953 : n957;
  assign n959 = pi18 ? n366 : ~n496;
  assign n960 = pi17 ? n32 : n959;
  assign n961 = pi16 ? n960 : n32;
  assign n962 = pi19 ? n32 : n813;
  assign n963 = pi18 ? n366 : ~n962;
  assign n964 = pi17 ? n32 : n963;
  assign n965 = pi16 ? n964 : n32;
  assign n966 = pi15 ? n961 : n965;
  assign n967 = pi19 ? n32 : n821;
  assign n968 = pi18 ? n366 : ~n967;
  assign n969 = pi17 ? n32 : n968;
  assign n970 = pi16 ? n969 : n32;
  assign n971 = pi15 ? n970 : n898;
  assign n972 = pi14 ? n966 : n971;
  assign n973 = pi13 ? n958 : n972;
  assign n974 = pi21 ? n32 : n173;
  assign n975 = pi20 ? n32 : n974;
  assign n976 = pi19 ? n975 : ~n32;
  assign n977 = pi18 ? n366 : ~n976;
  assign n978 = pi17 ? n32 : n977;
  assign n979 = pi16 ? n978 : n32;
  assign n980 = pi15 ? n784 : n979;
  assign n981 = pi14 ? n980 : n903;
  assign n982 = pi15 ? n713 : n426;
  assign n983 = pi18 ? n341 : n359;
  assign n984 = pi17 ? n32 : n983;
  assign n985 = pi16 ? n984 : n32;
  assign n986 = pi15 ? n829 : n985;
  assign n987 = pi14 ? n982 : n986;
  assign n988 = pi13 ? n981 : n987;
  assign n989 = pi12 ? n973 : n988;
  assign n990 = pi15 ? n985 : n621;
  assign n991 = pi15 ? n369 : n563;
  assign n992 = pi14 ? n990 : n991;
  assign n993 = pi21 ? n140 : ~n173;
  assign n994 = pi20 ? n32 : n993;
  assign n995 = pi19 ? n32 : n994;
  assign n996 = pi18 ? n995 : n32;
  assign n997 = pi17 ? n32 : n996;
  assign n998 = pi16 ? n997 : n32;
  assign n999 = pi15 ? n300 : n998;
  assign n1000 = pi21 ? n631 : ~n259;
  assign n1001 = pi20 ? n32 : n1000;
  assign n1002 = pi19 ? n32 : n1001;
  assign n1003 = pi18 ? n1002 : n32;
  assign n1004 = pi17 ? n32 : n1003;
  assign n1005 = pi16 ? n1004 : n32;
  assign n1006 = pi15 ? n1005 : n466;
  assign n1007 = pi14 ? n999 : n1006;
  assign n1008 = pi13 ? n992 : n1007;
  assign n1009 = pi22 ? n50 : n32;
  assign n1010 = pi21 ? n1009 : n32;
  assign n1011 = pi20 ? n32 : n1010;
  assign n1012 = pi19 ? n32 : n1011;
  assign n1013 = pi18 ? n1012 : n32;
  assign n1014 = pi17 ? n32 : n1013;
  assign n1015 = pi16 ? n1014 : n32;
  assign n1016 = pi15 ? n1015 : n130;
  assign n1017 = pi14 ? n1016 : n32;
  assign n1018 = pi13 ? n1017 : n32;
  assign n1019 = pi12 ? n1008 : n1018;
  assign n1020 = pi11 ? n989 : n1019;
  assign n1021 = pi10 ? n1020 : n32;
  assign n1022 = pi09 ? n949 : n1021;
  assign n1023 = pi08 ? n929 : n1022;
  assign n1024 = pi18 ? n423 : ~n32;
  assign n1025 = pi17 ? n1024 : ~n32;
  assign n1026 = pi16 ? n931 : ~n1025;
  assign n1027 = pi15 ? n32 : n1026;
  assign n1028 = pi18 ? n237 : ~n32;
  assign n1029 = pi17 ? n1028 : ~n32;
  assign n1030 = pi16 ? n931 : ~n1029;
  assign n1031 = pi16 ? n931 : n32;
  assign n1032 = pi15 ? n1030 : n1031;
  assign n1033 = pi14 ? n1027 : n1032;
  assign n1034 = pi13 ? n32 : n1033;
  assign n1035 = pi12 ? n32 : n1034;
  assign n1036 = pi11 ? n32 : n1035;
  assign n1037 = pi10 ? n32 : n1036;
  assign n1038 = pi18 ? n341 : ~n863;
  assign n1039 = pi17 ? n32 : n1038;
  assign n1040 = pi16 ? n1039 : n32;
  assign n1041 = pi18 ? n341 : ~n936;
  assign n1042 = pi17 ? n32 : n1041;
  assign n1043 = pi16 ? n1042 : n32;
  assign n1044 = pi15 ? n1040 : n1043;
  assign n1045 = pi18 ? n341 : ~n940;
  assign n1046 = pi17 ? n32 : n1045;
  assign n1047 = pi16 ? n1046 : n32;
  assign n1048 = pi18 ? n366 : ~n209;
  assign n1049 = pi17 ? n32 : n1048;
  assign n1050 = pi16 ? n1049 : n32;
  assign n1051 = pi15 ? n1047 : n1050;
  assign n1052 = pi14 ? n1044 : n1051;
  assign n1053 = pi20 ? n32 : ~n274;
  assign n1054 = pi19 ? n32 : n1053;
  assign n1055 = pi18 ? n366 : ~n1054;
  assign n1056 = pi17 ? n32 : n1055;
  assign n1057 = pi16 ? n1056 : n32;
  assign n1058 = pi18 ? n366 : ~n880;
  assign n1059 = pi17 ? n32 : n1058;
  assign n1060 = pi16 ? n1059 : n32;
  assign n1061 = pi15 ? n1057 : n1060;
  assign n1062 = pi15 ? n886 : n891;
  assign n1063 = pi14 ? n1061 : n1062;
  assign n1064 = pi13 ? n1052 : n1063;
  assign n1065 = pi15 ? n961 : n970;
  assign n1066 = pi15 ? n961 : n705;
  assign n1067 = pi14 ? n1065 : n1066;
  assign n1068 = pi15 ? n979 : n903;
  assign n1069 = pi18 ? n366 : ~n418;
  assign n1070 = pi17 ? n32 : n1069;
  assign n1071 = pi16 ? n1070 : n32;
  assign n1072 = pi15 ? n903 : n1071;
  assign n1073 = pi14 ? n1068 : n1072;
  assign n1074 = pi13 ? n1067 : n1073;
  assign n1075 = pi12 ? n1064 : n1074;
  assign n1076 = pi21 ? n32 : ~n309;
  assign n1077 = pi20 ? n1076 : ~n32;
  assign n1078 = pi19 ? n1077 : ~n32;
  assign n1079 = pi18 ? n366 : ~n1078;
  assign n1080 = pi17 ? n32 : n1079;
  assign n1081 = pi16 ? n1080 : n32;
  assign n1082 = pi15 ? n544 : n1081;
  assign n1083 = pi18 ? n341 : ~n826;
  assign n1084 = pi17 ? n32 : n1083;
  assign n1085 = pi16 ? n1084 : n32;
  assign n1086 = pi14 ? n1082 : n1085;
  assign n1087 = pi15 ? n616 : n719;
  assign n1088 = pi14 ? n1087 : n622;
  assign n1089 = pi13 ? n1086 : n1088;
  assign n1090 = pi14 ? n913 : n731;
  assign n1091 = pi21 ? n313 : ~n259;
  assign n1092 = pi20 ? n32 : n1091;
  assign n1093 = pi19 ? n32 : n1092;
  assign n1094 = pi18 ? n1093 : n32;
  assign n1095 = pi17 ? n32 : n1094;
  assign n1096 = pi16 ? n1095 : n32;
  assign n1097 = pi15 ? n1096 : n920;
  assign n1098 = pi15 ? n569 : n466;
  assign n1099 = pi14 ? n1097 : n1098;
  assign n1100 = pi13 ? n1090 : n1099;
  assign n1101 = pi12 ? n1089 : n1100;
  assign n1102 = pi11 ? n1075 : n1101;
  assign n1103 = pi15 ? n279 : n32;
  assign n1104 = pi14 ? n1103 : n32;
  assign n1105 = pi20 ? n141 : ~n32;
  assign n1106 = pi19 ? n32 : ~n1105;
  assign n1107 = pi18 ? n32 : n1106;
  assign n1108 = pi17 ? n32 : n1107;
  assign n1109 = pi16 ? n32 : n1108;
  assign n1110 = pi15 ? n32 : n1109;
  assign n1111 = pi14 ? n32 : n1110;
  assign n1112 = pi13 ? n1104 : n1111;
  assign n1113 = pi12 ? n1112 : n32;
  assign n1114 = pi14 ? n32 : n131;
  assign n1115 = pi13 ? n1114 : n32;
  assign n1116 = pi12 ? n32 : n1115;
  assign n1117 = pi11 ? n1113 : n1116;
  assign n1118 = pi10 ? n1102 : n1117;
  assign n1119 = pi09 ? n1037 : n1118;
  assign n1120 = pi18 ? n418 : ~n32;
  assign n1121 = pi17 ? n1120 : ~n32;
  assign n1122 = pi16 ? n931 : ~n1121;
  assign n1123 = pi15 ? n32 : n1122;
  assign n1124 = pi18 ? n359 : n32;
  assign n1125 = pi17 ? n1124 : n32;
  assign n1126 = pi16 ? n931 : n1125;
  assign n1127 = pi15 ? n1030 : n1126;
  assign n1128 = pi14 ? n1123 : n1127;
  assign n1129 = pi13 ? n32 : n1128;
  assign n1130 = pi12 ? n32 : n1129;
  assign n1131 = pi11 ? n32 : n1130;
  assign n1132 = pi10 ? n32 : n1131;
  assign n1133 = pi16 ? n1042 : ~n933;
  assign n1134 = pi18 ? n341 : ~n32;
  assign n1135 = pi17 ? n32 : n1134;
  assign n1136 = pi16 ? n1135 : n32;
  assign n1137 = pi15 ? n1133 : n1136;
  assign n1138 = pi20 ? n32 : n501;
  assign n1139 = pi19 ? n32 : n1138;
  assign n1140 = pi18 ? n366 : ~n1139;
  assign n1141 = pi17 ? n32 : n1140;
  assign n1142 = pi16 ? n1141 : n32;
  assign n1143 = pi15 ? n1047 : n1142;
  assign n1144 = pi14 ? n1137 : n1143;
  assign n1145 = pi20 ? n32 : ~n439;
  assign n1146 = pi19 ? n32 : n1145;
  assign n1147 = pi18 ? n366 : ~n1146;
  assign n1148 = pi17 ? n32 : n1147;
  assign n1149 = pi16 ? n1148 : n32;
  assign n1150 = pi20 ? n32 : n820;
  assign n1151 = pi19 ? n32 : n1150;
  assign n1152 = pi18 ? n366 : ~n1151;
  assign n1153 = pi17 ? n32 : n1152;
  assign n1154 = pi16 ? n1153 : n32;
  assign n1155 = pi15 ? n1149 : n1154;
  assign n1156 = pi19 ? n32 : n1077;
  assign n1157 = pi18 ? n366 : ~n1156;
  assign n1158 = pi17 ? n32 : n1157;
  assign n1159 = pi16 ? n1158 : n32;
  assign n1160 = pi15 ? n956 : n1159;
  assign n1161 = pi14 ? n1155 : n1160;
  assign n1162 = pi13 ? n1144 : n1161;
  assign n1163 = pi15 ? n961 : n898;
  assign n1164 = pi14 ? n961 : n1163;
  assign n1165 = pi20 ? n32 : n1076;
  assign n1166 = pi19 ? n1165 : ~n32;
  assign n1167 = pi18 ? n366 : ~n1166;
  assign n1168 = pi17 ? n32 : n1167;
  assign n1169 = pi16 ? n1168 : n32;
  assign n1170 = pi15 ? n784 : n1169;
  assign n1171 = pi15 ? n903 : n713;
  assign n1172 = pi14 ? n1170 : n1171;
  assign n1173 = pi13 ? n1164 : n1172;
  assign n1174 = pi12 ? n1162 : n1173;
  assign n1175 = pi15 ? n347 : n433;
  assign n1176 = pi14 ? n1175 : n540;
  assign n1177 = pi18 ? n341 : ~n814;
  assign n1178 = pi17 ? n32 : n1177;
  assign n1179 = pi16 ? n1178 : n32;
  assign n1180 = pi15 ? n719 : n1179;
  assign n1181 = pi15 ? n1179 : n616;
  assign n1182 = pi14 ? n1180 : n1181;
  assign n1183 = pi13 ? n1176 : n1182;
  assign n1184 = pi18 ? n262 : ~n618;
  assign n1185 = pi17 ? n32 : n1184;
  assign n1186 = pi16 ? n1185 : n32;
  assign n1187 = pi15 ? n369 : n1186;
  assign n1188 = pi21 ? n140 : ~n405;
  assign n1189 = pi20 ? n32 : n1188;
  assign n1190 = pi19 ? n32 : n1189;
  assign n1191 = pi18 ? n1190 : ~n618;
  assign n1192 = pi17 ? n32 : n1191;
  assign n1193 = pi16 ? n1192 : n32;
  assign n1194 = pi14 ? n1187 : n1193;
  assign n1195 = pi15 ? n731 : n569;
  assign n1196 = pi15 ? n998 : n1005;
  assign n1197 = pi14 ? n1195 : n1196;
  assign n1198 = pi13 ? n1194 : n1197;
  assign n1199 = pi12 ? n1183 : n1198;
  assign n1200 = pi11 ? n1174 : n1199;
  assign n1201 = pi15 ? n466 : n130;
  assign n1202 = pi14 ? n1098 : n1201;
  assign n1203 = pi16 ? n465 : n1108;
  assign n1204 = pi15 ? n32 : n1203;
  assign n1205 = pi14 ? n32 : n1204;
  assign n1206 = pi13 ? n1202 : n1205;
  assign n1207 = pi12 ? n1206 : n32;
  assign n1208 = pi11 ? n1207 : n32;
  assign n1209 = pi10 ? n1200 : n1208;
  assign n1210 = pi09 ? n1132 : n1209;
  assign n1211 = pi08 ? n1119 : n1210;
  assign n1212 = pi07 ? n1023 : n1211;
  assign n1213 = pi18 ? n209 : ~n32;
  assign n1214 = pi17 ? n32 : n1213;
  assign n1215 = pi18 ? n323 : ~n32;
  assign n1216 = pi17 ? n1215 : ~n32;
  assign n1217 = pi16 ? n1214 : ~n1216;
  assign n1218 = pi15 ? n32 : n1217;
  assign n1219 = pi18 ? n532 : ~n32;
  assign n1220 = pi17 ? n1219 : ~n32;
  assign n1221 = pi16 ? n931 : ~n1220;
  assign n1222 = pi14 ? n1218 : n1221;
  assign n1223 = pi13 ? n32 : n1222;
  assign n1224 = pi12 ? n32 : n1223;
  assign n1225 = pi11 ? n32 : n1224;
  assign n1226 = pi10 ? n32 : n1225;
  assign n1227 = pi18 ? n344 : ~n32;
  assign n1228 = pi17 ? n1227 : ~n32;
  assign n1229 = pi16 ? n1135 : ~n1228;
  assign n1230 = pi16 ? n1135 : ~n1029;
  assign n1231 = pi15 ? n1229 : n1230;
  assign n1232 = pi18 ? n366 : ~n32;
  assign n1233 = pi17 ? n32 : n1232;
  assign n1234 = pi16 ? n1233 : ~n1029;
  assign n1235 = pi15 ? n1230 : n1234;
  assign n1236 = pi14 ? n1231 : n1235;
  assign n1237 = pi16 ? n1233 : n32;
  assign n1238 = pi18 ? n366 : ~n863;
  assign n1239 = pi17 ? n32 : n1238;
  assign n1240 = pi16 ? n1239 : n32;
  assign n1241 = pi15 ? n1237 : n1240;
  assign n1242 = pi18 ? n366 : ~n940;
  assign n1243 = pi17 ? n32 : n1242;
  assign n1244 = pi16 ? n1243 : n32;
  assign n1245 = pi15 ? n1244 : n1240;
  assign n1246 = pi14 ? n1241 : n1245;
  assign n1247 = pi13 ? n1236 : n1246;
  assign n1248 = pi20 ? n32 : ~n266;
  assign n1249 = pi19 ? n32 : n1248;
  assign n1250 = pi18 ? n366 : ~n1249;
  assign n1251 = pi17 ? n32 : n1250;
  assign n1252 = pi16 ? n1251 : n32;
  assign n1253 = pi15 ? n1252 : n1050;
  assign n1254 = pi15 ? n883 : n1060;
  assign n1255 = pi14 ? n1253 : n1254;
  assign n1256 = pi18 ? n209 : ~n508;
  assign n1257 = pi17 ? n32 : n1256;
  assign n1258 = pi16 ? n1257 : n32;
  assign n1259 = pi15 ? n891 : n1258;
  assign n1260 = pi14 ? n961 : n1259;
  assign n1261 = pi13 ? n1255 : n1260;
  assign n1262 = pi12 ? n1247 : n1261;
  assign n1263 = pi15 ? n705 : n1169;
  assign n1264 = pi14 ? n1263 : n905;
  assign n1265 = pi20 ? n974 : ~n32;
  assign n1266 = pi19 ? n1265 : ~n32;
  assign n1267 = pi18 ? n341 : ~n1266;
  assign n1268 = pi17 ? n32 : n1267;
  assign n1269 = pi16 ? n1268 : n32;
  assign n1270 = pi15 ? n608 : n1269;
  assign n1271 = pi14 ? n608 : n1270;
  assign n1272 = pi13 ? n1264 : n1271;
  assign n1273 = pi18 ? n341 : ~n1078;
  assign n1274 = pi17 ? n32 : n1273;
  assign n1275 = pi16 ? n1274 : n32;
  assign n1276 = pi15 ? n1275 : n1081;
  assign n1277 = pi15 ? n436 : n1179;
  assign n1278 = pi14 ? n1276 : n1277;
  assign n1279 = pi15 ? n817 : n616;
  assign n1280 = pi14 ? n1279 : n547;
  assign n1281 = pi13 ? n1278 : n1280;
  assign n1282 = pi12 ? n1272 : n1281;
  assign n1283 = pi11 ? n1262 : n1282;
  assign n1284 = pi14 ? n825 : n369;
  assign n1285 = pi18 ? n1190 : n32;
  assign n1286 = pi17 ? n32 : n1285;
  assign n1287 = pi16 ? n1286 : n32;
  assign n1288 = pi15 ? n369 : n1287;
  assign n1289 = pi15 ? n1287 : n265;
  assign n1290 = pi14 ? n1288 : n1289;
  assign n1291 = pi13 ? n1284 : n1290;
  assign n1292 = pi15 ? n731 : n628;
  assign n1293 = pi14 ? n731 : n1292;
  assign n1294 = pi15 ? n576 : n569;
  assign n1295 = pi14 ? n628 : n1294;
  assign n1296 = pi13 ? n1293 : n1295;
  assign n1297 = pi12 ? n1291 : n1296;
  assign n1298 = pi15 ? n842 : n466;
  assign n1299 = pi14 ? n1298 : n32;
  assign n1300 = pi15 ? n466 : n576;
  assign n1301 = pi15 ? n279 : n576;
  assign n1302 = pi14 ? n1300 : n1301;
  assign n1303 = pi13 ? n1299 : n1302;
  assign n1304 = pi15 ? n1096 : n466;
  assign n1305 = pi14 ? n1304 : n466;
  assign n1306 = pi15 ? n628 : n1287;
  assign n1307 = pi20 ? n32 : n395;
  assign n1308 = pi19 ? n32 : n1307;
  assign n1309 = pi18 ? n1308 : n32;
  assign n1310 = pi17 ? n32 : n1309;
  assign n1311 = pi16 ? n1310 : n32;
  assign n1312 = pi15 ? n1311 : n1287;
  assign n1313 = pi14 ? n1306 : n1312;
  assign n1314 = pi13 ? n1305 : n1313;
  assign n1315 = pi12 ? n1303 : n1314;
  assign n1316 = pi11 ? n1297 : n1315;
  assign n1317 = pi10 ? n1283 : n1316;
  assign n1318 = pi09 ? n1226 : n1317;
  assign n1319 = pi21 ? n32 : n242;
  assign n1320 = pi20 ? n32 : n1319;
  assign n1321 = pi19 ? n32 : n1320;
  assign n1322 = pi18 ? n1321 : ~n32;
  assign n1323 = pi17 ? n32 : n1322;
  assign n1324 = pi21 ? n32 : ~n174;
  assign n1325 = pi20 ? n32 : n1324;
  assign n1326 = pi19 ? n1325 : ~n32;
  assign n1327 = pi18 ? n1326 : ~n32;
  assign n1328 = pi17 ? n1327 : ~n32;
  assign n1329 = pi16 ? n1323 : ~n1328;
  assign n1330 = pi15 ? n32 : n1329;
  assign n1331 = pi21 ? n405 : n32;
  assign n1332 = pi20 ? n32 : ~n1331;
  assign n1333 = pi19 ? n1332 : ~n32;
  assign n1334 = pi18 ? n1333 : ~n32;
  assign n1335 = pi17 ? n1334 : ~n32;
  assign n1336 = pi16 ? n931 : ~n1335;
  assign n1337 = pi20 ? n32 : ~n448;
  assign n1338 = pi19 ? n1337 : ~n32;
  assign n1339 = pi18 ? n1338 : ~n32;
  assign n1340 = pi17 ? n1339 : ~n32;
  assign n1341 = pi16 ? n931 : ~n1340;
  assign n1342 = pi15 ? n1336 : n1341;
  assign n1343 = pi14 ? n1330 : n1342;
  assign n1344 = pi13 ? n32 : n1343;
  assign n1345 = pi12 ? n32 : n1344;
  assign n1346 = pi11 ? n32 : n1345;
  assign n1347 = pi10 ? n32 : n1346;
  assign n1348 = pi20 ? n428 : n339;
  assign n1349 = pi19 ? n1348 : ~n32;
  assign n1350 = pi18 ? n1349 : ~n32;
  assign n1351 = pi17 ? n1350 : ~n32;
  assign n1352 = pi16 ? n1135 : ~n1351;
  assign n1353 = pi19 ? n502 : ~n32;
  assign n1354 = pi18 ? n1353 : ~n32;
  assign n1355 = pi17 ? n1354 : ~n32;
  assign n1356 = pi16 ? n1135 : ~n1355;
  assign n1357 = pi15 ? n1352 : n1356;
  assign n1358 = pi18 ? n826 : ~n32;
  assign n1359 = pi17 ? n1358 : ~n32;
  assign n1360 = pi16 ? n1135 : ~n1359;
  assign n1361 = pi15 ? n1360 : n1234;
  assign n1362 = pi14 ? n1357 : n1361;
  assign n1363 = pi16 ? n1233 : n1125;
  assign n1364 = pi18 ? n366 : ~n936;
  assign n1365 = pi17 ? n32 : n1364;
  assign n1366 = pi16 ? n1365 : n32;
  assign n1367 = pi15 ? n1363 : n1366;
  assign n1368 = pi21 ? n32 : ~n173;
  assign n1369 = pi20 ? n32 : n1368;
  assign n1370 = pi19 ? n32 : n1369;
  assign n1371 = pi18 ? n366 : ~n1370;
  assign n1372 = pi17 ? n32 : n1371;
  assign n1373 = pi16 ? n1372 : n32;
  assign n1374 = pi15 ? n1373 : n1240;
  assign n1375 = pi14 ? n1367 : n1374;
  assign n1376 = pi13 ? n1362 : n1375;
  assign n1377 = pi21 ? n309 : n259;
  assign n1378 = pi20 ? n32 : n1377;
  assign n1379 = pi19 ? n32 : n1378;
  assign n1380 = pi18 ? n366 : ~n1379;
  assign n1381 = pi17 ? n32 : n1380;
  assign n1382 = pi16 ? n1381 : n32;
  assign n1383 = pi15 ? n1382 : n875;
  assign n1384 = pi14 ? n1383 : n1060;
  assign n1385 = pi21 ? n32 : ~n405;
  assign n1386 = pi20 ? n1385 : ~n32;
  assign n1387 = pi19 ? n32 : n1386;
  assign n1388 = pi18 ? n366 : ~n1387;
  assign n1389 = pi17 ? n32 : n1388;
  assign n1390 = pi16 ? n1389 : n32;
  assign n1391 = pi15 ? n1390 : n961;
  assign n1392 = pi22 ? n65 : ~n32;
  assign n1393 = pi21 ? n1392 : ~n32;
  assign n1394 = pi20 ? n32 : n1393;
  assign n1395 = pi19 ? n32 : n1394;
  assign n1396 = pi18 ? n1395 : ~n508;
  assign n1397 = pi17 ? n32 : n1396;
  assign n1398 = pi16 ? n1397 : n32;
  assign n1399 = pi15 ? n891 : n1398;
  assign n1400 = pi14 ? n1391 : n1399;
  assign n1401 = pi13 ? n1384 : n1400;
  assign n1402 = pi12 ? n1376 : n1401;
  assign n1403 = pi15 ? n898 : n784;
  assign n1404 = pi14 ? n1403 : n1171;
  assign n1405 = pi19 ? n1138 : ~n32;
  assign n1406 = pi18 ? n366 : ~n1405;
  assign n1407 = pi17 ? n32 : n1406;
  assign n1408 = pi16 ? n1407 : n32;
  assign n1409 = pi15 ? n1408 : n800;
  assign n1410 = pi15 ? n608 : n535;
  assign n1411 = pi14 ? n1409 : n1410;
  assign n1412 = pi13 ? n1404 : n1411;
  assign n1413 = pi14 ? n535 : n436;
  assign n1414 = pi18 ? n366 : ~n1353;
  assign n1415 = pi17 ? n32 : n1414;
  assign n1416 = pi16 ? n1415 : n32;
  assign n1417 = pi15 ? n436 : n1416;
  assign n1418 = pi14 ? n1417 : n547;
  assign n1419 = pi13 ? n1413 : n1418;
  assign n1420 = pi12 ? n1412 : n1419;
  assign n1421 = pi11 ? n1402 : n1420;
  assign n1422 = pi15 ? n436 : n817;
  assign n1423 = pi18 ? n366 : n359;
  assign n1424 = pi17 ? n32 : n1423;
  assign n1425 = pi16 ? n1424 : n32;
  assign n1426 = pi15 ? n1425 : n724;
  assign n1427 = pi14 ? n1422 : n1426;
  assign n1428 = pi15 ? n621 : n563;
  assign n1429 = pi14 ? n621 : n1428;
  assign n1430 = pi13 ? n1427 : n1429;
  assign n1431 = pi15 ? n1287 : n998;
  assign n1432 = pi14 ? n369 : n1431;
  assign n1433 = pi15 ? n842 : n731;
  assign n1434 = pi14 ? n1287 : n1433;
  assign n1435 = pi13 ? n1432 : n1434;
  assign n1436 = pi12 ? n1430 : n1435;
  assign n1437 = pi15 ? n731 : n1005;
  assign n1438 = pi14 ? n1437 : n1301;
  assign n1439 = pi21 ? n1392 : ~n259;
  assign n1440 = pi20 ? n32 : n1439;
  assign n1441 = pi19 ? n32 : n1440;
  assign n1442 = pi18 ? n1441 : n32;
  assign n1443 = pi17 ? n32 : n1442;
  assign n1444 = pi16 ? n1443 : n32;
  assign n1445 = pi21 ? n140 : ~n259;
  assign n1446 = pi20 ? n32 : n1445;
  assign n1447 = pi19 ? n32 : n1446;
  assign n1448 = pi18 ? n1447 : n32;
  assign n1449 = pi17 ? n32 : n1448;
  assign n1450 = pi16 ? n1449 : n32;
  assign n1451 = pi15 ? n1444 : n1450;
  assign n1452 = pi14 ? n1005 : n1451;
  assign n1453 = pi13 ? n1438 : n1452;
  assign n1454 = pi15 ? n731 : n453;
  assign n1455 = pi14 ? n1454 : n453;
  assign n1456 = pi15 ? n1287 : n369;
  assign n1457 = pi14 ? n1456 : n369;
  assign n1458 = pi13 ? n1455 : n1457;
  assign n1459 = pi12 ? n1453 : n1458;
  assign n1460 = pi11 ? n1436 : n1459;
  assign n1461 = pi10 ? n1421 : n1460;
  assign n1462 = pi09 ? n1347 : n1461;
  assign n1463 = pi08 ? n1318 : n1462;
  assign n1464 = pi20 ? n32 : n246;
  assign n1465 = pi19 ? n1464 : n236;
  assign n1466 = pi18 ? n1465 : ~n32;
  assign n1467 = pi17 ? n1466 : ~n32;
  assign n1468 = pi16 ? n1323 : ~n1467;
  assign n1469 = pi15 ? n32 : n1468;
  assign n1470 = pi18 ? n940 : ~n32;
  assign n1471 = pi17 ? n32 : n1470;
  assign n1472 = pi18 ? n697 : ~n32;
  assign n1473 = pi17 ? n1472 : ~n32;
  assign n1474 = pi16 ? n1471 : ~n1473;
  assign n1475 = pi21 ? n100 : ~n32;
  assign n1476 = pi20 ? n32 : n1475;
  assign n1477 = pi19 ? n32 : n1476;
  assign n1478 = pi18 ? n1477 : ~n32;
  assign n1479 = pi17 ? n32 : n1478;
  assign n1480 = pi18 ? n702 : ~n32;
  assign n1481 = pi17 ? n1480 : ~n32;
  assign n1482 = pi16 ? n1479 : ~n1481;
  assign n1483 = pi15 ? n1474 : n1482;
  assign n1484 = pi14 ? n1469 : n1483;
  assign n1485 = pi13 ? n32 : n1484;
  assign n1486 = pi12 ? n32 : n1485;
  assign n1487 = pi11 ? n32 : n1486;
  assign n1488 = pi10 ? n32 : n1487;
  assign n1489 = pi16 ? n931 : ~n1481;
  assign n1490 = pi20 ? n342 : n321;
  assign n1491 = pi19 ? n1490 : ~n32;
  assign n1492 = pi18 ? n1491 : ~n32;
  assign n1493 = pi17 ? n1492 : ~n32;
  assign n1494 = pi16 ? n1135 : ~n1493;
  assign n1495 = pi15 ? n1489 : n1494;
  assign n1496 = pi16 ? n1135 : ~n1216;
  assign n1497 = pi16 ? n1233 : ~n1220;
  assign n1498 = pi15 ? n1496 : n1497;
  assign n1499 = pi14 ? n1495 : n1498;
  assign n1500 = pi18 ? n350 : ~n32;
  assign n1501 = pi17 ? n1500 : ~n32;
  assign n1502 = pi16 ? n1233 : ~n1501;
  assign n1503 = pi16 ? n1233 : ~n1228;
  assign n1504 = pi15 ? n1502 : n1503;
  assign n1505 = pi15 ? n1234 : n1363;
  assign n1506 = pi14 ? n1504 : n1505;
  assign n1507 = pi13 ? n1499 : n1506;
  assign n1508 = pi20 ? n32 : ~n220;
  assign n1509 = pi19 ? n32 : n1508;
  assign n1510 = pi18 ? n366 : ~n1509;
  assign n1511 = pi17 ? n32 : n1510;
  assign n1512 = pi16 ? n1511 : n32;
  assign n1513 = pi15 ? n1244 : n1512;
  assign n1514 = pi14 ? n1237 : n1513;
  assign n1515 = pi15 ? n1050 : n956;
  assign n1516 = pi14 ? n1515 : n1163;
  assign n1517 = pi13 ? n1514 : n1516;
  assign n1518 = pi12 ? n1507 : n1517;
  assign n1519 = pi15 ? n700 : n961;
  assign n1520 = pi14 ? n1163 : n1519;
  assign n1521 = pi15 ? n898 : n708;
  assign n1522 = pi15 ? n898 : n979;
  assign n1523 = pi14 ? n1521 : n1522;
  assign n1524 = pi13 ? n1520 : n1523;
  assign n1525 = pi14 ? n903 : n800;
  assign n1526 = pi19 ? n32 : n53;
  assign n1527 = pi18 ? n32 : n1526;
  assign n1528 = pi17 ? n32 : n1527;
  assign n1529 = pi16 ? n607 : n1528;
  assign n1530 = pi15 ? n1529 : n426;
  assign n1531 = pi15 ? n713 : n808;
  assign n1532 = pi14 ? n1530 : n1531;
  assign n1533 = pi13 ? n1525 : n1532;
  assign n1534 = pi12 ? n1524 : n1533;
  assign n1535 = pi11 ? n1518 : n1534;
  assign n1536 = pi15 ? n544 : n347;
  assign n1537 = pi15 ? n347 : n544;
  assign n1538 = pi14 ? n1536 : n1537;
  assign n1539 = pi18 ? n366 : ~n1266;
  assign n1540 = pi17 ? n32 : n1539;
  assign n1541 = pi19 ? n32 : ~n617;
  assign n1542 = pi18 ? n32 : n1541;
  assign n1543 = pi17 ? n32 : n1542;
  assign n1544 = pi16 ? n1540 : n1543;
  assign n1545 = pi15 ? n1269 : n1544;
  assign n1546 = pi14 ? n544 : n1545;
  assign n1547 = pi13 ? n1538 : n1546;
  assign n1548 = pi19 ? n589 : ~n32;
  assign n1549 = pi18 ? n366 : ~n1548;
  assign n1550 = pi17 ? n32 : n1549;
  assign n1551 = pi16 ? n1550 : n32;
  assign n1552 = pi15 ? n1551 : n544;
  assign n1553 = pi15 ? n1081 : n547;
  assign n1554 = pi14 ? n1552 : n1553;
  assign n1555 = pi15 ? n1551 : n829;
  assign n1556 = pi14 ? n1555 : n817;
  assign n1557 = pi13 ? n1554 : n1556;
  assign n1558 = pi12 ? n1547 : n1557;
  assign n1559 = pi15 ? n547 : n369;
  assign n1560 = pi15 ? n369 : n616;
  assign n1561 = pi14 ? n1559 : n1560;
  assign n1562 = pi14 ? n616 : n547;
  assign n1563 = pi13 ? n1561 : n1562;
  assign n1564 = pi15 ? n547 : n817;
  assign n1565 = pi14 ? n1564 : n817;
  assign n1566 = pi16 ? n1540 : n32;
  assign n1567 = pi15 ? n1551 : n1566;
  assign n1568 = pi14 ? n1567 : n1566;
  assign n1569 = pi13 ? n1565 : n1568;
  assign n1570 = pi12 ? n1563 : n1569;
  assign n1571 = pi11 ? n1558 : n1570;
  assign n1572 = pi10 ? n1535 : n1571;
  assign n1573 = pi09 ? n1488 : n1572;
  assign n1574 = pi20 ? n32 : n101;
  assign n1575 = pi19 ? n32 : n1574;
  assign n1576 = pi18 ? n1575 : ~n32;
  assign n1577 = pi17 ? n32 : n1576;
  assign n1578 = pi16 ? n1577 : ~n1467;
  assign n1579 = pi15 ? n32 : n1578;
  assign n1580 = pi18 ? n863 : ~n32;
  assign n1581 = pi17 ? n32 : n1580;
  assign n1582 = pi18 ? n503 : ~n32;
  assign n1583 = pi17 ? n1582 : ~n32;
  assign n1584 = pi16 ? n1581 : ~n1583;
  assign n1585 = pi16 ? n1323 : ~n1481;
  assign n1586 = pi15 ? n1584 : n1585;
  assign n1587 = pi14 ? n1579 : n1586;
  assign n1588 = pi13 ? n32 : n1587;
  assign n1589 = pi12 ? n32 : n1588;
  assign n1590 = pi11 ? n32 : n1589;
  assign n1591 = pi10 ? n32 : n1590;
  assign n1592 = pi19 ? n32 : n519;
  assign n1593 = pi18 ? n1592 : ~n32;
  assign n1594 = pi17 ? n32 : n1593;
  assign n1595 = pi16 ? n1594 : ~n1481;
  assign n1596 = pi15 ? n1595 : n1494;
  assign n1597 = pi16 ? n1233 : ~n1340;
  assign n1598 = pi15 ? n1496 : n1597;
  assign n1599 = pi14 ? n1596 : n1598;
  assign n1600 = pi20 ? n321 : n339;
  assign n1601 = pi19 ? n1600 : ~n32;
  assign n1602 = pi18 ? n1601 : ~n32;
  assign n1603 = pi17 ? n1602 : ~n32;
  assign n1604 = pi16 ? n1233 : ~n1603;
  assign n1605 = pi18 ? n430 : ~n32;
  assign n1606 = pi17 ? n1605 : ~n32;
  assign n1607 = pi16 ? n1233 : ~n1606;
  assign n1608 = pi15 ? n1604 : n1607;
  assign n1609 = pi14 ? n1608 : n1234;
  assign n1610 = pi13 ? n1599 : n1609;
  assign n1611 = pi21 ? n309 : n206;
  assign n1612 = pi20 ? n32 : n1611;
  assign n1613 = pi19 ? n32 : n1612;
  assign n1614 = pi18 ? n366 : ~n1613;
  assign n1615 = pi17 ? n32 : n1614;
  assign n1616 = pi16 ? n1615 : n32;
  assign n1617 = pi15 ? n1244 : n1616;
  assign n1618 = pi14 ? n1237 : n1617;
  assign n1619 = pi15 ? n875 : n886;
  assign n1620 = pi14 ? n1619 : n1066;
  assign n1621 = pi13 ? n1618 : n1620;
  assign n1622 = pi12 ? n1610 : n1621;
  assign n1623 = pi15 ? n894 : n961;
  assign n1624 = pi14 ? n1163 : n1623;
  assign n1625 = pi15 ? n898 : n526;
  assign n1626 = pi14 ? n1625 : n898;
  assign n1627 = pi13 ? n1624 : n1626;
  assign n1628 = pi14 ? n530 : n796;
  assign n1629 = pi21 ? n66 : n32;
  assign n1630 = pi20 ? n1629 : n32;
  assign n1631 = pi19 ? n32 : n1630;
  assign n1632 = pi18 ? n32 : n1631;
  assign n1633 = pi17 ? n32 : n1632;
  assign n1634 = pi16 ? n607 : n1633;
  assign n1635 = pi15 ? n1634 : n608;
  assign n1636 = pi14 ? n1635 : n800;
  assign n1637 = pi13 ? n1628 : n1636;
  assign n1638 = pi12 ? n1627 : n1637;
  assign n1639 = pi11 ? n1622 : n1638;
  assign n1640 = pi18 ? n366 : ~n423;
  assign n1641 = pi17 ? n32 : n1640;
  assign n1642 = pi16 ? n1641 : n32;
  assign n1643 = pi15 ? n544 : n1642;
  assign n1644 = pi15 ? n1642 : n540;
  assign n1645 = pi14 ? n1643 : n1644;
  assign n1646 = pi15 ? n540 : n535;
  assign n1647 = pi14 ? n540 : n1646;
  assign n1648 = pi13 ? n1645 : n1647;
  assign n1649 = pi15 ? n1642 : n347;
  assign n1650 = pi15 ? n540 : n1566;
  assign n1651 = pi14 ? n1649 : n1650;
  assign n1652 = pi15 ? n1566 : n1551;
  assign n1653 = pi14 ? n1652 : n1081;
  assign n1654 = pi13 ? n1651 : n1653;
  assign n1655 = pi12 ? n1648 : n1654;
  assign n1656 = pi15 ? n547 : n621;
  assign n1657 = pi15 ? n825 : n817;
  assign n1658 = pi14 ? n1656 : n1657;
  assign n1659 = pi15 ? n817 : n829;
  assign n1660 = pi14 ? n1659 : n1551;
  assign n1661 = pi13 ? n1658 : n1660;
  assign n1662 = pi15 ? n1551 : n547;
  assign n1663 = pi14 ? n1662 : n436;
  assign n1664 = pi15 ? n1566 : n535;
  assign n1665 = pi14 ? n1664 : n535;
  assign n1666 = pi13 ? n1663 : n1665;
  assign n1667 = pi12 ? n1661 : n1666;
  assign n1668 = pi11 ? n1655 : n1667;
  assign n1669 = pi10 ? n1639 : n1668;
  assign n1670 = pi09 ? n1591 : n1669;
  assign n1671 = pi08 ? n1573 : n1670;
  assign n1672 = pi07 ? n1463 : n1671;
  assign n1673 = pi06 ? n1212 : n1672;
  assign n1674 = pi05 ? n856 : n1673;
  assign n1675 = pi04 ? n235 : n1674;
  assign n1676 = pi19 ? n1105 : ~n32;
  assign n1677 = pi18 ? n32 : n1676;
  assign n1678 = pi17 ? n32 : n1677;
  assign n1679 = pi17 ? n1470 : ~n32;
  assign n1680 = pi16 ? n1678 : ~n1679;
  assign n1681 = pi15 ? n32 : n1680;
  assign n1682 = pi18 ? n32 : ~n32;
  assign n1683 = pi17 ? n32 : n1682;
  assign n1684 = pi16 ? n1683 : ~n1679;
  assign n1685 = pi21 ? n206 : ~n259;
  assign n1686 = pi20 ? n1685 : ~n32;
  assign n1687 = pi19 ? n857 : n1686;
  assign n1688 = pi18 ? n1687 : ~n32;
  assign n1689 = pi17 ? n1688 : ~n32;
  assign n1690 = pi16 ? n1323 : ~n1689;
  assign n1691 = pi15 ? n1684 : n1690;
  assign n1692 = pi14 ? n1681 : n1691;
  assign n1693 = pi13 ? n32 : n1692;
  assign n1694 = pi12 ? n32 : n1693;
  assign n1695 = pi11 ? n32 : n1694;
  assign n1696 = pi10 ? n32 : n1695;
  assign n1697 = pi18 ? n880 : ~n32;
  assign n1698 = pi17 ? n1697 : ~n32;
  assign n1699 = pi16 ? n1594 : ~n1698;
  assign n1700 = pi18 ? n590 : ~n32;
  assign n1701 = pi17 ? n1700 : ~n32;
  assign n1702 = pi16 ? n1479 : ~n1701;
  assign n1703 = pi15 ? n1699 : n1702;
  assign n1704 = pi18 ? n751 : ~n32;
  assign n1705 = pi17 ? n32 : n1704;
  assign n1706 = pi18 ? n684 : ~n32;
  assign n1707 = pi17 ? n1706 : ~n32;
  assign n1708 = pi16 ? n1705 : ~n1707;
  assign n1709 = pi16 ? n1135 : ~n1481;
  assign n1710 = pi15 ? n1708 : n1709;
  assign n1711 = pi14 ? n1703 : n1710;
  assign n1712 = pi19 ? n322 : n236;
  assign n1713 = pi18 ? n1712 : ~n32;
  assign n1714 = pi17 ? n1713 : ~n32;
  assign n1715 = pi16 ? n1233 : ~n1714;
  assign n1716 = pi16 ? n1233 : ~n1481;
  assign n1717 = pi15 ? n1715 : n1716;
  assign n1718 = pi18 ? n508 : ~n32;
  assign n1719 = pi17 ? n1718 : ~n32;
  assign n1720 = pi16 ? n1233 : ~n1719;
  assign n1721 = pi14 ? n1717 : n1720;
  assign n1722 = pi13 ? n1711 : n1721;
  assign n1723 = pi16 ? n1233 : ~n1216;
  assign n1724 = pi16 ? n1233 : ~n1121;
  assign n1725 = pi15 ? n1723 : n1724;
  assign n1726 = pi18 ? n1548 : ~n32;
  assign n1727 = pi17 ? n1726 : ~n32;
  assign n1728 = pi16 ? n1233 : ~n1727;
  assign n1729 = pi15 ? n1503 : n1728;
  assign n1730 = pi14 ? n1725 : n1729;
  assign n1731 = pi15 ? n1234 : n1244;
  assign n1732 = pi18 ? n366 : ~n268;
  assign n1733 = pi17 ? n32 : n1732;
  assign n1734 = pi16 ? n1733 : n32;
  assign n1735 = pi15 ? n875 : n1734;
  assign n1736 = pi14 ? n1731 : n1735;
  assign n1737 = pi13 ? n1730 : n1736;
  assign n1738 = pi12 ? n1722 : n1737;
  assign n1739 = pi14 ? n1513 : n1245;
  assign n1740 = pi20 ? n342 : n207;
  assign n1741 = pi19 ? n32 : n1740;
  assign n1742 = pi18 ? n366 : ~n1741;
  assign n1743 = pi17 ? n32 : n1742;
  assign n1744 = pi16 ? n1743 : n32;
  assign n1745 = pi15 ? n1252 : n1744;
  assign n1746 = pi15 ? n1050 : n886;
  assign n1747 = pi14 ? n1745 : n1746;
  assign n1748 = pi13 ? n1739 : n1747;
  assign n1749 = pi15 ? n886 : n1744;
  assign n1750 = pi19 ? n32 : n617;
  assign n1751 = pi18 ? n366 : ~n1750;
  assign n1752 = pi17 ? n32 : n1751;
  assign n1753 = pi16 ? n1752 : n32;
  assign n1754 = pi15 ? n961 : n1753;
  assign n1755 = pi14 ? n1749 : n1754;
  assign n1756 = pi16 ? n893 : n1633;
  assign n1757 = pi20 ? n266 : n32;
  assign n1758 = pi19 ? n32 : ~n1757;
  assign n1759 = pi18 ? n366 : ~n1758;
  assign n1760 = pi17 ? n32 : n1759;
  assign n1761 = pi16 ? n1760 : n32;
  assign n1762 = pi15 ? n1756 : n1761;
  assign n1763 = pi14 ? n1762 : n1623;
  assign n1764 = pi13 ? n1755 : n1763;
  assign n1765 = pi12 ? n1748 : n1764;
  assign n1766 = pi11 ? n1738 : n1765;
  assign n1767 = pi18 ? n366 : ~n520;
  assign n1768 = pi17 ? n32 : n1767;
  assign n1769 = pi16 ? n1768 : n32;
  assign n1770 = pi15 ? n1769 : n979;
  assign n1771 = pi15 ? n784 : n530;
  assign n1772 = pi14 ? n1770 : n1771;
  assign n1773 = pi18 ? n341 : ~n1405;
  assign n1774 = pi17 ? n32 : n1773;
  assign n1775 = pi16 ? n1774 : n32;
  assign n1776 = pi15 ? n1775 : n523;
  assign n1777 = pi15 ? n1769 : n608;
  assign n1778 = pi14 ? n1776 : n1777;
  assign n1779 = pi13 ? n1772 : n1778;
  assign n1780 = pi15 ? n903 : n1769;
  assign n1781 = pi15 ? n1769 : n708;
  assign n1782 = pi14 ? n1780 : n1781;
  assign n1783 = pi13 ? n1782 : n903;
  assign n1784 = pi12 ? n1779 : n1783;
  assign n1785 = pi20 ? n32 : n67;
  assign n1786 = pi19 ? n1785 : n32;
  assign n1787 = pi18 ? n32 : n1786;
  assign n1788 = pi17 ? n32 : n1787;
  assign n1789 = pi16 ? n810 : n1788;
  assign n1790 = pi15 ? n800 : n1789;
  assign n1791 = pi14 ? n1790 : n713;
  assign n1792 = pi13 ? n1791 : n608;
  assign n1793 = pi15 ? n608 : n800;
  assign n1794 = pi14 ? n1793 : n800;
  assign n1795 = pi16 ? n707 : n657;
  assign n1796 = pi15 ? n1795 : n898;
  assign n1797 = pi18 ? n366 : ~n772;
  assign n1798 = pi17 ? n32 : n1797;
  assign n1799 = pi16 ? n1798 : n32;
  assign n1800 = pi15 ? n898 : n1799;
  assign n1801 = pi14 ? n1796 : n1800;
  assign n1802 = pi13 ? n1794 : n1801;
  assign n1803 = pi12 ? n1792 : n1802;
  assign n1804 = pi11 ? n1784 : n1803;
  assign n1805 = pi10 ? n1766 : n1804;
  assign n1806 = pi09 ? n1696 : n1805;
  assign n1807 = pi18 ? n32 : n350;
  assign n1808 = pi17 ? n32 : n1807;
  assign n1809 = pi17 ? n1593 : ~n32;
  assign n1810 = pi16 ? n1808 : ~n1809;
  assign n1811 = pi15 ? n32 : n1810;
  assign n1812 = pi20 ? n1475 : ~n32;
  assign n1813 = pi19 ? n1812 : ~n32;
  assign n1814 = pi18 ? n32 : n1813;
  assign n1815 = pi17 ? n32 : n1814;
  assign n1816 = pi16 ? n1815 : ~n1679;
  assign n1817 = pi21 ? n32 : ~n259;
  assign n1818 = pi20 ? n32 : n1817;
  assign n1819 = pi19 ? n32 : n1818;
  assign n1820 = pi18 ? n32 : ~n1819;
  assign n1821 = pi17 ? n32 : n1820;
  assign n1822 = pi20 ? n1331 : n1377;
  assign n1823 = pi19 ? n1822 : n1686;
  assign n1824 = pi18 ? n1823 : ~n32;
  assign n1825 = pi17 ? n1824 : ~n32;
  assign n1826 = pi16 ? n1821 : ~n1825;
  assign n1827 = pi15 ? n1816 : n1826;
  assign n1828 = pi14 ? n1811 : n1827;
  assign n1829 = pi13 ? n32 : n1828;
  assign n1830 = pi12 ? n32 : n1829;
  assign n1831 = pi11 ? n32 : n1830;
  assign n1832 = pi10 ? n32 : n1831;
  assign n1833 = pi18 ? n936 : ~n32;
  assign n1834 = pi17 ? n32 : n1833;
  assign n1835 = pi16 ? n1834 : ~n1698;
  assign n1836 = pi16 ? n1323 : ~n1707;
  assign n1837 = pi15 ? n1835 : n1836;
  assign n1838 = pi16 ? n1594 : ~n1707;
  assign n1839 = pi21 ? n32 : n140;
  assign n1840 = pi20 ? n32 : n1839;
  assign n1841 = pi19 ? n32 : n1840;
  assign n1842 = pi18 ? n1841 : ~n32;
  assign n1843 = pi17 ? n32 : n1842;
  assign n1844 = pi20 ? n1331 : n32;
  assign n1845 = pi19 ? n32 : ~n1844;
  assign n1846 = pi18 ? n1845 : ~n32;
  assign n1847 = pi17 ? n1846 : ~n32;
  assign n1848 = pi16 ? n1843 : ~n1847;
  assign n1849 = pi15 ? n1838 : n1848;
  assign n1850 = pi14 ? n1837 : n1849;
  assign n1851 = pi13 ? n1850 : n1721;
  assign n1852 = pi16 ? n1233 : ~n1351;
  assign n1853 = pi15 ? n1852 : n1728;
  assign n1854 = pi14 ? n1725 : n1853;
  assign n1855 = pi18 ? n341 : ~n268;
  assign n1856 = pi17 ? n32 : n1855;
  assign n1857 = pi16 ? n1856 : n32;
  assign n1858 = pi15 ? n1050 : n1857;
  assign n1859 = pi14 ? n1731 : n1858;
  assign n1860 = pi13 ? n1854 : n1859;
  assign n1861 = pi12 ? n1851 : n1860;
  assign n1862 = pi19 ? n32 : n1165;
  assign n1863 = pi18 ? n366 : ~n1862;
  assign n1864 = pi17 ? n32 : n1863;
  assign n1865 = pi16 ? n1864 : n32;
  assign n1866 = pi15 ? n1865 : n1240;
  assign n1867 = pi14 ? n1617 : n1866;
  assign n1868 = pi20 ? n428 : n749;
  assign n1869 = pi19 ? n32 : n1868;
  assign n1870 = pi18 ? n366 : ~n1869;
  assign n1871 = pi17 ? n32 : n1870;
  assign n1872 = pi16 ? n1871 : n32;
  assign n1873 = pi15 ? n1252 : n1872;
  assign n1874 = pi18 ? n366 : ~n1592;
  assign n1875 = pi17 ? n32 : n1874;
  assign n1876 = pi16 ? n1875 : n32;
  assign n1877 = pi15 ? n1876 : n886;
  assign n1878 = pi14 ? n1873 : n1877;
  assign n1879 = pi13 ? n1867 : n1878;
  assign n1880 = pi18 ? n366 : ~n590;
  assign n1881 = pi17 ? n32 : n1880;
  assign n1882 = pi16 ? n1881 : n32;
  assign n1883 = pi15 ? n1882 : n894;
  assign n1884 = pi14 ? n1749 : n1883;
  assign n1885 = pi20 ? n915 : n32;
  assign n1886 = pi19 ? n32 : ~n1885;
  assign n1887 = pi18 ? n366 : ~n1886;
  assign n1888 = pi17 ? n32 : n1887;
  assign n1889 = pi16 ? n1888 : n32;
  assign n1890 = pi15 ? n894 : n1889;
  assign n1891 = pi14 ? n1890 : n961;
  assign n1892 = pi13 ? n1884 : n1891;
  assign n1893 = pi12 ? n1879 : n1892;
  assign n1894 = pi11 ? n1861 : n1893;
  assign n1895 = pi15 ? n784 : n898;
  assign n1896 = pi15 ? n1799 : n1769;
  assign n1897 = pi14 ? n1895 : n1896;
  assign n1898 = pi19 ? n975 : n617;
  assign n1899 = pi18 ? n366 : ~n1898;
  assign n1900 = pi17 ? n32 : n1899;
  assign n1901 = pi16 ? n1900 : n32;
  assign n1902 = pi15 ? n979 : n1901;
  assign n1903 = pi15 ? n1753 : n713;
  assign n1904 = pi14 ? n1902 : n1903;
  assign n1905 = pi13 ? n1897 : n1904;
  assign n1906 = pi18 ? n341 : ~n1166;
  assign n1907 = pi17 ? n32 : n1906;
  assign n1908 = pi16 ? n1907 : n32;
  assign n1909 = pi15 ? n1908 : n708;
  assign n1910 = pi14 ? n1909 : n708;
  assign n1911 = pi14 ? n979 : n1169;
  assign n1912 = pi13 ? n1910 : n1911;
  assign n1913 = pi12 ? n1905 : n1912;
  assign n1914 = pi19 ? n1150 : ~n32;
  assign n1915 = pi18 ? n366 : ~n1914;
  assign n1916 = pi17 ? n32 : n1915;
  assign n1917 = pi16 ? n1916 : n32;
  assign n1918 = pi15 ? n1169 : n1917;
  assign n1919 = pi14 ? n1918 : n800;
  assign n1920 = pi13 ? n1919 : n796;
  assign n1921 = pi15 ? n796 : n1769;
  assign n1922 = pi14 ? n1921 : n1769;
  assign n1923 = pi16 ? n783 : n657;
  assign n1924 = pi15 ? n1923 : n1753;
  assign n1925 = pi15 ? n1753 : n894;
  assign n1926 = pi14 ? n1924 : n1925;
  assign n1927 = pi13 ? n1922 : n1926;
  assign n1928 = pi12 ? n1920 : n1927;
  assign n1929 = pi11 ? n1913 : n1928;
  assign n1930 = pi10 ? n1894 : n1929;
  assign n1931 = pi09 ? n1832 : n1930;
  assign n1932 = pi08 ? n1806 : n1931;
  assign n1933 = pi18 ? n32 : n344;
  assign n1934 = pi17 ? n32 : n1933;
  assign n1935 = pi17 ? n1682 : ~n32;
  assign n1936 = pi16 ? n1934 : ~n1935;
  assign n1937 = pi15 ? n32 : n1936;
  assign n1938 = pi16 ? n1815 : ~n1935;
  assign n1939 = pi22 ? n32 : n50;
  assign n1940 = pi21 ? n1939 : ~n32;
  assign n1941 = pi20 ? n1940 : ~n32;
  assign n1942 = pi19 ? n1941 : ~n32;
  assign n1943 = pi18 ? n32 : n1942;
  assign n1944 = pi17 ? n32 : n1943;
  assign n1945 = pi17 ? n1833 : ~n32;
  assign n1946 = pi16 ? n1944 : ~n1945;
  assign n1947 = pi15 ? n1938 : n1946;
  assign n1948 = pi14 ? n1937 : n1947;
  assign n1949 = pi13 ? n32 : n1948;
  assign n1950 = pi12 ? n32 : n1949;
  assign n1951 = pi11 ? n32 : n1950;
  assign n1952 = pi10 ? n32 : n1951;
  assign n1953 = pi17 ? n1580 : ~n32;
  assign n1954 = pi16 ? n1683 : ~n1953;
  assign n1955 = pi16 ? n1577 : ~n1953;
  assign n1956 = pi15 ? n1954 : n1955;
  assign n1957 = pi19 ? n32 : n792;
  assign n1958 = pi18 ? n1957 : ~n32;
  assign n1959 = pi17 ? n1958 : ~n32;
  assign n1960 = pi16 ? n1594 : ~n1959;
  assign n1961 = pi17 ? n1213 : ~n32;
  assign n1962 = pi16 ? n1471 : ~n1961;
  assign n1963 = pi15 ? n1960 : n1962;
  assign n1964 = pi14 ? n1956 : n1963;
  assign n1965 = pi19 ? n32 : n429;
  assign n1966 = pi18 ? n1965 : ~n32;
  assign n1967 = pi17 ? n1966 : ~n32;
  assign n1968 = pi16 ? n1705 : ~n1967;
  assign n1969 = pi20 ? n32 : n1940;
  assign n1970 = pi19 ? n32 : n1969;
  assign n1971 = pi18 ? n1970 : ~n32;
  assign n1972 = pi17 ? n32 : n1971;
  assign n1973 = pi16 ? n1972 : ~n1967;
  assign n1974 = pi15 ? n1968 : n1973;
  assign n1975 = pi18 ? n1156 : ~n32;
  assign n1976 = pi17 ? n1975 : ~n32;
  assign n1977 = pi16 ? n1135 : ~n1976;
  assign n1978 = pi18 ? n496 : ~n32;
  assign n1979 = pi17 ? n1978 : ~n32;
  assign n1980 = pi16 ? n1233 : ~n1979;
  assign n1981 = pi15 ? n1977 : n1980;
  assign n1982 = pi14 ? n1974 : n1981;
  assign n1983 = pi13 ? n1964 : n1982;
  assign n1984 = pi18 ? n1750 : ~n32;
  assign n1985 = pi17 ? n1984 : ~n32;
  assign n1986 = pi16 ? n1233 : ~n1985;
  assign n1987 = pi16 ? n1233 : ~n1473;
  assign n1988 = pi15 ? n1986 : n1987;
  assign n1989 = pi18 ? n595 : ~n32;
  assign n1990 = pi17 ? n1989 : ~n32;
  assign n1991 = pi16 ? n1233 : ~n1990;
  assign n1992 = pi15 ? n1987 : n1991;
  assign n1993 = pi14 ? n1988 : n1992;
  assign n1994 = pi18 ? n1166 : ~n32;
  assign n1995 = pi17 ? n1994 : ~n32;
  assign n1996 = pi16 ? n1233 : ~n1995;
  assign n1997 = pi18 ? n1405 : ~n32;
  assign n1998 = pi17 ? n1997 : ~n32;
  assign n1999 = pi16 ? n1233 : ~n1998;
  assign n2000 = pi15 ? n1996 : n1999;
  assign n2001 = pi15 ? n1497 : n1503;
  assign n2002 = pi14 ? n2000 : n2001;
  assign n2003 = pi13 ? n1993 : n2002;
  assign n2004 = pi12 ? n1983 : n2003;
  assign n2005 = pi18 ? n814 : ~n32;
  assign n2006 = pi17 ? n2005 : ~n32;
  assign n2007 = pi16 ? n1233 : ~n2006;
  assign n2008 = pi18 ? n618 : ~n32;
  assign n2009 = pi17 ? n2008 : ~n32;
  assign n2010 = pi16 ? n1233 : ~n2009;
  assign n2011 = pi15 ? n2007 : n2010;
  assign n2012 = pi14 ? n1503 : n2011;
  assign n2013 = pi15 ? n1363 : n1234;
  assign n2014 = pi16 ? n1365 : ~n2009;
  assign n2015 = pi15 ? n2014 : n1616;
  assign n2016 = pi14 ? n2013 : n2015;
  assign n2017 = pi13 ? n2012 : n2016;
  assign n2018 = pi15 ? n1240 : n1237;
  assign n2019 = pi21 ? n173 : ~n259;
  assign n2020 = pi20 ? n32 : ~n2019;
  assign n2021 = pi19 ? n32 : n2020;
  assign n2022 = pi18 ? n366 : ~n2021;
  assign n2023 = pi17 ? n32 : n2022;
  assign n2024 = pi16 ? n2023 : n32;
  assign n2025 = pi20 ? n428 : n207;
  assign n2026 = pi19 ? n32 : n2025;
  assign n2027 = pi18 ? n366 : ~n2026;
  assign n2028 = pi17 ? n32 : n2027;
  assign n2029 = pi16 ? n2028 : n32;
  assign n2030 = pi15 ? n2024 : n2029;
  assign n2031 = pi14 ? n2018 : n2030;
  assign n2032 = pi15 ? n1050 : n1244;
  assign n2033 = pi20 ? n175 : ~n266;
  assign n2034 = pi19 ? n32 : n2033;
  assign n2035 = pi18 ? n366 : ~n2034;
  assign n2036 = pi17 ? n32 : n2035;
  assign n2037 = pi16 ? n2036 : n32;
  assign n2038 = pi15 ? n2037 : n886;
  assign n2039 = pi14 ? n2032 : n2038;
  assign n2040 = pi13 ? n2031 : n2039;
  assign n2041 = pi12 ? n2017 : n2040;
  assign n2042 = pi11 ? n2004 : n2041;
  assign n2043 = pi19 ? n32 : n422;
  assign n2044 = pi18 ? n366 : ~n2043;
  assign n2045 = pi17 ? n32 : n2044;
  assign n2046 = pi16 ? n2045 : n32;
  assign n2047 = pi15 ? n2046 : n1050;
  assign n2048 = pi15 ? n891 : n961;
  assign n2049 = pi14 ? n2047 : n2048;
  assign n2050 = pi15 ? n1159 : n1050;
  assign n2051 = pi18 ? n366 : ~n767;
  assign n2052 = pi17 ? n32 : n2051;
  assign n2053 = pi19 ? n32 : n37;
  assign n2054 = pi18 ? n32 : n2053;
  assign n2055 = pi17 ? n32 : n2054;
  assign n2056 = pi16 ? n2052 : n2055;
  assign n2057 = pi16 ? n2052 : n32;
  assign n2058 = pi15 ? n2056 : n2057;
  assign n2059 = pi14 ? n2050 : n2058;
  assign n2060 = pi13 ? n2049 : n2059;
  assign n2061 = pi18 ? n341 : ~n503;
  assign n2062 = pi17 ? n32 : n2061;
  assign n2063 = pi16 ? n2062 : n32;
  assign n2064 = pi15 ? n2063 : n891;
  assign n2065 = pi14 ? n1882 : n2064;
  assign n2066 = pi15 ? n961 : n886;
  assign n2067 = pi16 ? n893 : n1108;
  assign n2068 = pi15 ? n961 : n2067;
  assign n2069 = pi14 ? n2066 : n2068;
  assign n2070 = pi13 ? n2065 : n2069;
  assign n2071 = pi12 ? n2060 : n2070;
  assign n2072 = pi19 ? n1574 : n32;
  assign n2073 = pi18 ? n32 : n2072;
  assign n2074 = pi17 ? n32 : n2073;
  assign n2075 = pi16 ? n960 : n2074;
  assign n2076 = pi22 ? n32 : n84;
  assign n2077 = pi21 ? n32 : n2076;
  assign n2078 = pi20 ? n32 : n2077;
  assign n2079 = pi19 ? n2078 : n32;
  assign n2080 = pi18 ? n32 : n2079;
  assign n2081 = pi17 ? n32 : n2080;
  assign n2082 = pi16 ? n704 : n2081;
  assign n2083 = pi15 ? n2075 : n2082;
  assign n2084 = pi15 ? n705 : n894;
  assign n2085 = pi14 ? n2083 : n2084;
  assign n2086 = pi15 ? n894 : n898;
  assign n2087 = pi15 ? n961 : n1882;
  assign n2088 = pi14 ? n2086 : n2087;
  assign n2089 = pi13 ? n2085 : n2088;
  assign n2090 = pi16 ? n960 : n475;
  assign n2091 = pi15 ? n961 : n2090;
  assign n2092 = pi20 ? n32 : n86;
  assign n2093 = pi19 ? n2092 : n32;
  assign n2094 = pi18 ? n32 : n2093;
  assign n2095 = pi17 ? n32 : n2094;
  assign n2096 = pi16 ? n890 : n2095;
  assign n2097 = pi16 ? n885 : n386;
  assign n2098 = pi15 ? n2096 : n2097;
  assign n2099 = pi14 ? n2091 : n2098;
  assign n2100 = pi18 ? n366 : ~n1965;
  assign n2101 = pi17 ? n32 : n2100;
  assign n2102 = pi21 ? n100 : ~n140;
  assign n2103 = pi20 ? n32 : n2102;
  assign n2104 = pi19 ? n2103 : n32;
  assign n2105 = pi18 ? n32 : n2104;
  assign n2106 = pi17 ? n32 : n2105;
  assign n2107 = pi16 ? n2101 : n2106;
  assign n2108 = pi19 ? n32 : n804;
  assign n2109 = pi18 ? n366 : ~n2108;
  assign n2110 = pi17 ? n32 : n2109;
  assign n2111 = pi16 ? n2110 : n32;
  assign n2112 = pi15 ? n2107 : n2111;
  assign n2113 = pi14 ? n2112 : n2111;
  assign n2114 = pi13 ? n2099 : n2113;
  assign n2115 = pi12 ? n2089 : n2114;
  assign n2116 = pi11 ? n2071 : n2115;
  assign n2117 = pi10 ? n2042 : n2116;
  assign n2118 = pi09 ? n1952 : n2117;
  assign n2119 = pi18 ? n32 : n605;
  assign n2120 = pi17 ? n32 : n2119;
  assign n2121 = pi16 ? n2120 : ~n1935;
  assign n2122 = pi15 ? n32 : n2121;
  assign n2123 = pi18 ? n32 : n618;
  assign n2124 = pi17 ? n2123 : ~n32;
  assign n2125 = pi16 ? n1934 : ~n2124;
  assign n2126 = pi16 ? n1808 : ~n1935;
  assign n2127 = pi15 ? n2125 : n2126;
  assign n2128 = pi14 ? n2122 : n2127;
  assign n2129 = pi13 ? n32 : n2128;
  assign n2130 = pi12 ? n32 : n2129;
  assign n2131 = pi11 ? n32 : n2130;
  assign n2132 = pi10 ? n32 : n2131;
  assign n2133 = pi18 ? n858 : ~n32;
  assign n2134 = pi17 ? n2133 : ~n32;
  assign n2135 = pi16 ? n1815 : ~n2134;
  assign n2136 = pi18 ? n32 : n814;
  assign n2137 = pi17 ? n32 : n2136;
  assign n2138 = pi16 ? n2137 : ~n1945;
  assign n2139 = pi15 ? n2135 : n2138;
  assign n2140 = pi21 ? n32 : n1939;
  assign n2141 = pi20 ? n32 : n2140;
  assign n2142 = pi19 ? n32 : n2141;
  assign n2143 = pi18 ? n2142 : ~n32;
  assign n2144 = pi17 ? n32 : n2143;
  assign n2145 = pi16 ? n2144 : ~n1961;
  assign n2146 = pi15 ? n1955 : n2145;
  assign n2147 = pi14 ? n2139 : n2146;
  assign n2148 = pi17 ? n1134 : ~n32;
  assign n2149 = pi16 ? n1594 : ~n2148;
  assign n2150 = pi18 ? n2108 : ~n32;
  assign n2151 = pi17 ? n2150 : ~n32;
  assign n2152 = pi16 ? n1843 : ~n2151;
  assign n2153 = pi15 ? n2149 : n2152;
  assign n2154 = pi16 ? n1843 : ~n1967;
  assign n2155 = pi16 ? n1233 : ~n1701;
  assign n2156 = pi15 ? n2154 : n2155;
  assign n2157 = pi14 ? n2153 : n2156;
  assign n2158 = pi13 ? n2147 : n2157;
  assign n2159 = pi18 ? n962 : ~n32;
  assign n2160 = pi17 ? n2159 : ~n32;
  assign n2161 = pi16 ? n1233 : ~n2160;
  assign n2162 = pi15 ? n2161 : n1991;
  assign n2163 = pi14 ? n1987 : n2162;
  assign n2164 = pi15 ? n1996 : n1723;
  assign n2165 = pi18 ? n805 : ~n32;
  assign n2166 = pi17 ? n2165 : ~n32;
  assign n2167 = pi16 ? n1233 : ~n2166;
  assign n2168 = pi20 ? n175 : n207;
  assign n2169 = pi19 ? n2168 : ~n32;
  assign n2170 = pi18 ? n2169 : ~n32;
  assign n2171 = pi17 ? n2170 : ~n32;
  assign n2172 = pi16 ? n1233 : ~n2171;
  assign n2173 = pi15 ? n2167 : n2172;
  assign n2174 = pi14 ? n2164 : n2173;
  assign n2175 = pi13 ? n2163 : n2174;
  assign n2176 = pi12 ? n2158 : n2175;
  assign n2177 = pi18 ? n1078 : ~n32;
  assign n2178 = pi17 ? n2177 : ~n32;
  assign n2179 = pi16 ? n1233 : ~n2178;
  assign n2180 = pi21 ? n174 : ~n309;
  assign n2181 = pi20 ? n2180 : ~n32;
  assign n2182 = pi19 ? n2181 : ~n32;
  assign n2183 = pi18 ? n2182 : ~n32;
  assign n2184 = pi17 ? n2183 : ~n32;
  assign n2185 = pi16 ? n1233 : ~n2184;
  assign n2186 = pi15 ? n2179 : n2185;
  assign n2187 = pi14 ? n1852 : n2186;
  assign n2188 = pi16 ? n1233 : ~n1359;
  assign n2189 = pi15 ? n2188 : n2007;
  assign n2190 = pi18 ? n366 : ~n858;
  assign n2191 = pi17 ? n32 : n2190;
  assign n2192 = pi16 ? n2191 : n1125;
  assign n2193 = pi15 ? n1234 : n2192;
  assign n2194 = pi14 ? n2189 : n2193;
  assign n2195 = pi13 ? n2187 : n2194;
  assign n2196 = pi15 ? n2010 : n1237;
  assign n2197 = pi19 ? n32 : n975;
  assign n2198 = pi18 ? n366 : ~n2197;
  assign n2199 = pi17 ? n32 : n2198;
  assign n2200 = pi16 ? n2199 : n32;
  assign n2201 = pi20 ? n32 : n2180;
  assign n2202 = pi19 ? n32 : n2201;
  assign n2203 = pi18 ? n366 : ~n2202;
  assign n2204 = pi17 ? n32 : n2203;
  assign n2205 = pi16 ? n2204 : n32;
  assign n2206 = pi15 ? n2200 : n2205;
  assign n2207 = pi14 ? n2196 : n2206;
  assign n2208 = pi15 ? n2205 : n1373;
  assign n2209 = pi19 ? n32 : n1348;
  assign n2210 = pi18 ? n366 : ~n2209;
  assign n2211 = pi17 ? n32 : n2210;
  assign n2212 = pi16 ? n2211 : n32;
  assign n2213 = pi15 ? n1382 : n2212;
  assign n2214 = pi14 ? n2208 : n2213;
  assign n2215 = pi13 ? n2207 : n2214;
  assign n2216 = pi12 ? n2195 : n2215;
  assign n2217 = pi11 ? n2176 : n2216;
  assign n2218 = pi15 ? n1154 : n1876;
  assign n2219 = pi15 ? n1159 : n2212;
  assign n2220 = pi14 ? n2218 : n2219;
  assign n2221 = pi20 ? n428 : n820;
  assign n2222 = pi19 ? n32 : n2221;
  assign n2223 = pi18 ? n366 : ~n2222;
  assign n2224 = pi17 ? n32 : n2223;
  assign n2225 = pi16 ? n2224 : n32;
  assign n2226 = pi18 ? n366 : ~n751;
  assign n2227 = pi17 ? n32 : n2226;
  assign n2228 = pi16 ? n2227 : n32;
  assign n2229 = pi15 ? n2225 : n2228;
  assign n2230 = pi15 ? n1882 : n2046;
  assign n2231 = pi14 ? n2229 : n2230;
  assign n2232 = pi13 ? n2220 : n2231;
  assign n2233 = pi19 ? n32 : n1265;
  assign n2234 = pi18 ? n366 : ~n2233;
  assign n2235 = pi17 ? n32 : n2234;
  assign n2236 = pi16 ? n2235 : n32;
  assign n2237 = pi14 ? n2046 : n2236;
  assign n2238 = pi15 ? n2236 : n2212;
  assign n2239 = pi18 ? n341 : ~n1156;
  assign n2240 = pi17 ? n32 : n2239;
  assign n2241 = pi16 ? n2240 : n32;
  assign n2242 = pi19 ? n32 : n2181;
  assign n2243 = pi18 ? n366 : ~n2242;
  assign n2244 = pi17 ? n32 : n2243;
  assign n2245 = pi16 ? n2244 : n32;
  assign n2246 = pi15 ? n2241 : n2245;
  assign n2247 = pi14 ? n2238 : n2246;
  assign n2248 = pi13 ? n2237 : n2247;
  assign n2249 = pi12 ? n2232 : n2248;
  assign n2250 = pi20 ? n448 : n32;
  assign n2251 = pi19 ? n32 : ~n2250;
  assign n2252 = pi18 ? n366 : ~n2251;
  assign n2253 = pi17 ? n32 : n2252;
  assign n2254 = pi16 ? n2253 : n32;
  assign n2255 = pi15 ? n961 : n2254;
  assign n2256 = pi21 ? n173 : n309;
  assign n2257 = pi20 ? n2256 : n32;
  assign n2258 = pi19 ? n32 : ~n2257;
  assign n2259 = pi18 ? n366 : ~n2258;
  assign n2260 = pi17 ? n32 : n2259;
  assign n2261 = pi16 ? n2260 : n32;
  assign n2262 = pi15 ? n2261 : n2245;
  assign n2263 = pi14 ? n2255 : n2262;
  assign n2264 = pi15 ? n2245 : n898;
  assign n2265 = pi20 ? n1368 : ~n32;
  assign n2266 = pi19 ? n32 : n2265;
  assign n2267 = pi18 ? n366 : ~n2266;
  assign n2268 = pi17 ? n32 : n2267;
  assign n2269 = pi16 ? n2268 : n32;
  assign n2270 = pi15 ? n2269 : n2046;
  assign n2271 = pi14 ? n2264 : n2270;
  assign n2272 = pi13 ? n2263 : n2271;
  assign n2273 = pi15 ? n2269 : n2236;
  assign n2274 = pi16 ? n2101 : n32;
  assign n2275 = pi15 ? n2236 : n2274;
  assign n2276 = pi14 ? n2273 : n2275;
  assign n2277 = pi20 ? n32 : n160;
  assign n2278 = pi19 ? n2277 : n32;
  assign n2279 = pi18 ? n32 : n2278;
  assign n2280 = pi17 ? n32 : n2279;
  assign n2281 = pi16 ? n2110 : n2280;
  assign n2282 = pi15 ? n2281 : n1050;
  assign n2283 = pi14 ? n2282 : n1050;
  assign n2284 = pi13 ? n2276 : n2283;
  assign n2285 = pi12 ? n2272 : n2284;
  assign n2286 = pi11 ? n2249 : n2285;
  assign n2287 = pi10 ? n2217 : n2286;
  assign n2288 = pi09 ? n2132 : n2287;
  assign n2289 = pi08 ? n2118 : n2288;
  assign n2290 = pi07 ? n1932 : n2289;
  assign n2291 = pi19 ? n1476 : ~n32;
  assign n2292 = pi18 ? n32 : n2291;
  assign n2293 = pi17 ? n32 : n2292;
  assign n2294 = pi17 ? n2119 : ~n32;
  assign n2295 = pi16 ? n2293 : ~n2294;
  assign n2296 = pi15 ? n32 : n2295;
  assign n2297 = pi20 ? n101 : ~n32;
  assign n2298 = pi19 ? n2297 : ~n32;
  assign n2299 = pi18 ? n32 : n2298;
  assign n2300 = pi17 ? n32 : n2299;
  assign n2301 = pi17 ? n1933 : ~n32;
  assign n2302 = pi16 ? n2300 : ~n2301;
  assign n2303 = pi20 ? n2140 : ~n32;
  assign n2304 = pi19 ? n2303 : ~n32;
  assign n2305 = pi18 ? n32 : n2304;
  assign n2306 = pi17 ? n32 : n2305;
  assign n2307 = pi16 ? n2306 : ~n2301;
  assign n2308 = pi15 ? n2302 : n2307;
  assign n2309 = pi14 ? n2296 : n2308;
  assign n2310 = pi13 ? n32 : n2309;
  assign n2311 = pi12 ? n32 : n2310;
  assign n2312 = pi11 ? n32 : n2311;
  assign n2313 = pi10 ? n32 : n2312;
  assign n2314 = pi18 ? n32 : n1353;
  assign n2315 = pi17 ? n2314 : ~n32;
  assign n2316 = pi16 ? n1934 : ~n2315;
  assign n2317 = pi20 ? n1319 : ~n32;
  assign n2318 = pi19 ? n2317 : ~n32;
  assign n2319 = pi18 ? n32 : n2318;
  assign n2320 = pi17 ? n32 : n2319;
  assign n2321 = pi17 ? n1807 : ~n32;
  assign n2322 = pi16 ? n2320 : ~n2321;
  assign n2323 = pi15 ? n2316 : n2322;
  assign n2324 = pi16 ? n2137 : ~n2124;
  assign n2325 = pi18 ? n32 : n237;
  assign n2326 = pi17 ? n32 : n2325;
  assign n2327 = pi16 ? n2326 : ~n2134;
  assign n2328 = pi15 ? n2324 : n2327;
  assign n2329 = pi14 ? n2323 : n2328;
  assign n2330 = pi16 ? n1834 : ~n1945;
  assign n2331 = pi15 ? n1955 : n2330;
  assign n2332 = pi18 ? n1862 : ~n32;
  assign n2333 = pi17 ? n2332 : ~n32;
  assign n2334 = pi16 ? n1843 : ~n2333;
  assign n2335 = pi16 ? n1471 : ~n1679;
  assign n2336 = pi15 ? n2334 : n2335;
  assign n2337 = pi14 ? n2331 : n2336;
  assign n2338 = pi13 ? n2329 : n2337;
  assign n2339 = pi16 ? n1705 : ~n2148;
  assign n2340 = pi16 ? n1972 : ~n2151;
  assign n2341 = pi15 ? n2339 : n2340;
  assign n2342 = pi16 ? n1135 : ~n1707;
  assign n2343 = pi15 ? n2342 : n2155;
  assign n2344 = pi14 ? n2341 : n2343;
  assign n2345 = pi18 ? n776 : ~n32;
  assign n2346 = pi17 ? n2345 : ~n32;
  assign n2347 = pi16 ? n1233 : ~n2346;
  assign n2348 = pi15 ? n2347 : n1991;
  assign n2349 = pi14 ? n1987 : n2348;
  assign n2350 = pi13 ? n2344 : n2349;
  assign n2351 = pi12 ? n2338 : n2350;
  assign n2352 = pi15 ? n1996 : n1720;
  assign n2353 = pi14 ? n2352 : n1720;
  assign n2354 = pi15 ? n1723 : n1999;
  assign n2355 = pi18 ? n605 : ~n32;
  assign n2356 = pi17 ? n2355 : ~n32;
  assign n2357 = pi16 ? n1233 : ~n2356;
  assign n2358 = pi21 ? n309 : ~n32;
  assign n2359 = pi20 ? n32 : n2358;
  assign n2360 = pi19 ? n2359 : ~n32;
  assign n2361 = pi18 ? n2360 : ~n32;
  assign n2362 = pi17 ? n2361 : ~n32;
  assign n2363 = pi16 ? n1233 : ~n2362;
  assign n2364 = pi15 ? n2357 : n2363;
  assign n2365 = pi14 ? n2354 : n2364;
  assign n2366 = pi13 ? n2353 : n2365;
  assign n2367 = pi15 ? n1497 : n1607;
  assign n2368 = pi14 ? n2367 : n1503;
  assign n2369 = pi15 ? n1503 : n1502;
  assign n2370 = pi15 ? n1502 : n1234;
  assign n2371 = pi14 ? n2369 : n2370;
  assign n2372 = pi13 ? n2368 : n2371;
  assign n2373 = pi12 ? n2366 : n2372;
  assign n2374 = pi11 ? n2351 : n2373;
  assign n2375 = pi15 ? n2014 : n1237;
  assign n2376 = pi14 ? n1234 : n2375;
  assign n2377 = pi14 ? n1234 : n2018;
  assign n2378 = pi13 ? n2376 : n2377;
  assign n2379 = pi15 ? n1876 : n1240;
  assign n2380 = pi14 ? n1237 : n2379;
  assign n2381 = pi15 ? n1240 : n1366;
  assign n2382 = pi14 ? n2381 : n1245;
  assign n2383 = pi13 ? n2380 : n2382;
  assign n2384 = pi12 ? n2378 : n2383;
  assign n2385 = pi21 ? n405 : n206;
  assign n2386 = pi20 ? n32 : n2385;
  assign n2387 = pi19 ? n32 : n2386;
  assign n2388 = pi18 ? n366 : ~n2387;
  assign n2389 = pi17 ? n32 : n2388;
  assign n2390 = pi16 ? n2389 : n32;
  assign n2391 = pi15 ? n2390 : n2228;
  assign n2392 = pi14 ? n2391 : n2228;
  assign n2393 = pi18 ? n366 : ~n1957;
  assign n2394 = pi17 ? n32 : n2393;
  assign n2395 = pi16 ? n2394 : n32;
  assign n2396 = pi15 ? n1244 : n2395;
  assign n2397 = pi14 ? n2396 : n1876;
  assign n2398 = pi13 ? n2392 : n2397;
  assign n2399 = pi15 ? n1244 : n1876;
  assign n2400 = pi14 ? n1876 : n2399;
  assign n2401 = pi15 ? n1366 : n1234;
  assign n2402 = pi14 ? n2401 : n1234;
  assign n2403 = pi13 ? n2400 : n2402;
  assign n2404 = pi12 ? n2398 : n2403;
  assign n2405 = pi11 ? n2384 : n2404;
  assign n2406 = pi10 ? n2374 : n2405;
  assign n2407 = pi09 ? n2313 : n2406;
  assign n2408 = pi18 ? n32 : n797;
  assign n2409 = pi17 ? n32 : n2408;
  assign n2410 = pi18 ? n32 : n430;
  assign n2411 = pi17 ? n2410 : ~n32;
  assign n2412 = pi16 ? n2409 : ~n2411;
  assign n2413 = pi19 ? n1969 : ~n32;
  assign n2414 = pi18 ? n32 : n2413;
  assign n2415 = pi17 ? n32 : n2414;
  assign n2416 = pi16 ? n2415 : ~n2301;
  assign n2417 = pi15 ? n2412 : n2416;
  assign n2418 = pi14 ? n2296 : n2417;
  assign n2419 = pi13 ? n32 : n2418;
  assign n2420 = pi12 ? n32 : n2419;
  assign n2421 = pi11 ? n32 : n2420;
  assign n2422 = pi10 ? n32 : n2421;
  assign n2423 = pi16 ? n2120 : ~n2301;
  assign n2424 = pi19 ? n244 : ~n32;
  assign n2425 = pi18 ? n32 : n2424;
  assign n2426 = pi17 ? n32 : n2425;
  assign n2427 = pi16 ? n2426 : ~n2321;
  assign n2428 = pi15 ? n2423 : n2427;
  assign n2429 = pi16 ? n2320 : ~n2315;
  assign n2430 = pi16 ? n1815 : ~n2124;
  assign n2431 = pi15 ? n2429 : n2430;
  assign n2432 = pi14 ? n2428 : n2431;
  assign n2433 = pi18 ? n936 : n618;
  assign n2434 = pi17 ? n2433 : ~n32;
  assign n2435 = pi16 ? n2137 : ~n2434;
  assign n2436 = pi16 ? n1944 : ~n1935;
  assign n2437 = pi15 ? n2435 : n2436;
  assign n2438 = pi16 ? n1834 : ~n1953;
  assign n2439 = pi16 ? n2144 : ~n1679;
  assign n2440 = pi15 ? n2438 : n2439;
  assign n2441 = pi14 ? n2437 : n2440;
  assign n2442 = pi13 ? n2432 : n2441;
  assign n2443 = pi16 ? n1594 : ~n1961;
  assign n2444 = pi16 ? n1843 : ~n1961;
  assign n2445 = pi15 ? n2443 : n2444;
  assign n2446 = pi18 ? n2209 : ~n32;
  assign n2447 = pi17 ? n2446 : ~n32;
  assign n2448 = pi16 ? n1843 : ~n2447;
  assign n2449 = pi18 ? n2233 : ~n32;
  assign n2450 = pi17 ? n2449 : ~n32;
  assign n2451 = pi16 ? n1233 : ~n2450;
  assign n2452 = pi15 ? n2448 : n2451;
  assign n2453 = pi14 ? n2445 : n2452;
  assign n2454 = pi15 ? n1987 : n2161;
  assign n2455 = pi15 ? n1987 : n1716;
  assign n2456 = pi14 ? n2454 : n2455;
  assign n2457 = pi13 ? n2453 : n2456;
  assign n2458 = pi12 ? n2442 : n2457;
  assign n2459 = pi15 ? n1991 : n1720;
  assign n2460 = pi14 ? n1991 : n2459;
  assign n2461 = pi18 ? n520 : ~n32;
  assign n2462 = pi17 ? n2461 : ~n32;
  assign n2463 = pi16 ? n1233 : ~n2462;
  assign n2464 = pi15 ? n1723 : n2463;
  assign n2465 = pi18 ? n797 : ~n32;
  assign n2466 = pi17 ? n2465 : ~n32;
  assign n2467 = pi16 ? n1233 : ~n2466;
  assign n2468 = pi15 ? n2467 : n1723;
  assign n2469 = pi14 ? n2464 : n2468;
  assign n2470 = pi13 ? n2460 : n2469;
  assign n2471 = pi14 ? n2167 : n1607;
  assign n2472 = pi19 ? n2265 : ~n32;
  assign n2473 = pi18 ? n2472 : ~n32;
  assign n2474 = pi17 ? n2473 : ~n32;
  assign n2475 = pi16 ? n1233 : ~n2474;
  assign n2476 = pi15 ? n1852 : n2475;
  assign n2477 = pi15 ? n2179 : n2007;
  assign n2478 = pi14 ? n2476 : n2477;
  assign n2479 = pi13 ? n2471 : n2478;
  assign n2480 = pi12 ? n2470 : n2479;
  assign n2481 = pi11 ? n2458 : n2480;
  assign n2482 = pi14 ? n2007 : n1505;
  assign n2483 = pi16 ? n1233 : ~n1355;
  assign n2484 = pi15 ? n2014 : n2010;
  assign n2485 = pi14 ? n2483 : n2484;
  assign n2486 = pi13 ? n2482 : n2485;
  assign n2487 = pi16 ? n1233 : ~n933;
  assign n2488 = pi15 ? n2010 : n2487;
  assign n2489 = pi16 ? n2191 : n32;
  assign n2490 = pi14 ? n2488 : n2489;
  assign n2491 = pi15 ? n2489 : n1363;
  assign n2492 = pi15 ? n2200 : n1366;
  assign n2493 = pi14 ? n2491 : n2492;
  assign n2494 = pi13 ? n2490 : n2493;
  assign n2495 = pi12 ? n2486 : n2494;
  assign n2496 = pi15 ? n1240 : n1865;
  assign n2497 = pi14 ? n2496 : n1865;
  assign n2498 = pi15 ? n1865 : n2489;
  assign n2499 = pi14 ? n2498 : n2489;
  assign n2500 = pi13 ? n2497 : n2499;
  assign n2501 = pi15 ? n1373 : n2489;
  assign n2502 = pi14 ? n2489 : n2501;
  assign n2503 = pi15 ? n1363 : n2483;
  assign n2504 = pi15 ? n2483 : n1234;
  assign n2505 = pi14 ? n2503 : n2504;
  assign n2506 = pi13 ? n2502 : n2505;
  assign n2507 = pi12 ? n2500 : n2506;
  assign n2508 = pi11 ? n2495 : n2507;
  assign n2509 = pi10 ? n2481 : n2508;
  assign n2510 = pi09 ? n2422 : n2509;
  assign n2511 = pi08 ? n2407 : n2510;
  assign n2512 = pi18 ? n32 : n508;
  assign n2513 = pi17 ? n32 : n2512;
  assign n2514 = pi17 ? n2512 : ~n32;
  assign n2515 = pi16 ? n2513 : ~n2514;
  assign n2516 = pi15 ? n32 : n2515;
  assign n2517 = pi18 ? n32 : n520;
  assign n2518 = pi17 ? n32 : n2517;
  assign n2519 = pi18 ? n32 : n323;
  assign n2520 = pi17 ? n2519 : ~n32;
  assign n2521 = pi16 ? n2518 : ~n2520;
  assign n2522 = pi14 ? n2516 : n2521;
  assign n2523 = pi13 ? n32 : n2522;
  assign n2524 = pi12 ? n32 : n2523;
  assign n2525 = pi11 ? n32 : n2524;
  assign n2526 = pi10 ? n32 : n2525;
  assign n2527 = pi16 ? n2293 : ~n2520;
  assign n2528 = pi16 ? n2409 : ~n2294;
  assign n2529 = pi15 ? n2527 : n2528;
  assign n2530 = pi17 ? n32 : n2410;
  assign n2531 = pi18 ? n32 : n532;
  assign n2532 = pi17 ? n2531 : ~n32;
  assign n2533 = pi16 ? n2530 : ~n2532;
  assign n2534 = pi16 ? n1934 : ~n2411;
  assign n2535 = pi15 ? n2533 : n2534;
  assign n2536 = pi14 ? n2529 : n2535;
  assign n2537 = pi18 ? n32 : n1548;
  assign n2538 = pi17 ? n2537 : ~n32;
  assign n2539 = pi16 ? n2320 : ~n2538;
  assign n2540 = pi17 ? n32 : n2537;
  assign n2541 = pi16 ? n2540 : ~n2321;
  assign n2542 = pi15 ? n2539 : n2541;
  assign n2543 = pi16 ? n1944 : ~n2315;
  assign n2544 = pi17 ? n2325 : ~n32;
  assign n2545 = pi16 ? n2326 : ~n2544;
  assign n2546 = pi15 ? n2543 : n2545;
  assign n2547 = pi14 ? n2542 : n2546;
  assign n2548 = pi13 ? n2536 : n2547;
  assign n2549 = pi16 ? n1577 : ~n2124;
  assign n2550 = pi16 ? n1834 : ~n1935;
  assign n2551 = pi15 ? n2549 : n2550;
  assign n2552 = pi16 ? n1843 : ~n1953;
  assign n2553 = pi15 ? n2552 : n2335;
  assign n2554 = pi14 ? n2551 : n2553;
  assign n2555 = pi18 ? n2043 : ~n32;
  assign n2556 = pi17 ? n2555 : ~n32;
  assign n2557 = pi16 ? n1705 : ~n2556;
  assign n2558 = pi16 ? n1972 : ~n1698;
  assign n2559 = pi15 ? n2557 : n2558;
  assign n2560 = pi18 ? n2026 : ~n32;
  assign n2561 = pi17 ? n2560 : ~n32;
  assign n2562 = pi16 ? n1135 : ~n2561;
  assign n2563 = pi15 ? n2562 : n2451;
  assign n2564 = pi14 ? n2559 : n2563;
  assign n2565 = pi13 ? n2554 : n2564;
  assign n2566 = pi12 ? n2548 : n2565;
  assign n2567 = pi18 ? n772 : ~n32;
  assign n2568 = pi17 ? n2567 : ~n32;
  assign n2569 = pi16 ? n1233 : ~n2568;
  assign n2570 = pi15 ? n2569 : n1716;
  assign n2571 = pi14 ? n1988 : n2570;
  assign n2572 = pi13 ? n1980 : n2571;
  assign n2573 = pi18 ? n976 : ~n32;
  assign n2574 = pi17 ? n2573 : ~n32;
  assign n2575 = pi16 ? n1233 : ~n2574;
  assign n2576 = pi15 ? n2575 : n1991;
  assign n2577 = pi14 ? n2576 : n1720;
  assign n2578 = pi15 ? n1723 : n1716;
  assign n2579 = pi15 ? n2463 : n2357;
  assign n2580 = pi14 ? n2578 : n2579;
  assign n2581 = pi13 ? n2577 : n2580;
  assign n2582 = pi12 ? n2572 : n2581;
  assign n2583 = pi11 ? n2566 : n2582;
  assign n2584 = pi15 ? n2357 : n1999;
  assign n2585 = pi15 ? n2357 : n1724;
  assign n2586 = pi14 ? n2584 : n2585;
  assign n2587 = pi15 ? n2467 : n1497;
  assign n2588 = pi14 ? n2587 : n1497;
  assign n2589 = pi13 ? n2586 : n2588;
  assign n2590 = pi14 ? n1497 : n1607;
  assign n2591 = pi15 ? n1607 : n1852;
  assign n2592 = pi15 ? n2179 : n1503;
  assign n2593 = pi14 ? n2591 : n2592;
  assign n2594 = pi13 ? n2590 : n2593;
  assign n2595 = pi12 ? n2589 : n2594;
  assign n2596 = pi13 ? n1502 : n1503;
  assign n2597 = pi18 ? n1266 : ~n32;
  assign n2598 = pi17 ? n2597 : ~n32;
  assign n2599 = pi16 ? n1233 : ~n2598;
  assign n2600 = pi15 ? n1503 : n2599;
  assign n2601 = pi15 ? n2599 : n1497;
  assign n2602 = pi14 ? n2600 : n2601;
  assign n2603 = pi15 ? n1497 : n2363;
  assign n2604 = pi18 ? n1914 : ~n32;
  assign n2605 = pi17 ? n2604 : ~n32;
  assign n2606 = pi16 ? n1233 : ~n2605;
  assign n2607 = pi15 ? n2363 : n2606;
  assign n2608 = pi14 ? n2603 : n2607;
  assign n2609 = pi13 ? n2602 : n2608;
  assign n2610 = pi12 ? n2596 : n2609;
  assign n2611 = pi11 ? n2595 : n2610;
  assign n2612 = pi10 ? n2583 : n2611;
  assign n2613 = pi09 ? n2526 : n2612;
  assign n2614 = pi20 ? n243 : ~n32;
  assign n2615 = pi19 ? n32 : n2614;
  assign n2616 = pi18 ? n32 : n2615;
  assign n2617 = pi17 ? n32 : n2616;
  assign n2618 = pi18 ? n32 : n595;
  assign n2619 = pi17 ? n2618 : ~n32;
  assign n2620 = pi16 ? n2617 : ~n2619;
  assign n2621 = pi15 ? n32 : n2620;
  assign n2622 = pi19 ? n32 : n1105;
  assign n2623 = pi18 ? n32 : n2622;
  assign n2624 = pi17 ? n32 : n2623;
  assign n2625 = pi17 ? n2517 : ~n32;
  assign n2626 = pi16 ? n2624 : ~n2625;
  assign n2627 = pi19 ? n2141 : ~n32;
  assign n2628 = pi18 ? n32 : n2627;
  assign n2629 = pi17 ? n32 : n2628;
  assign n2630 = pi16 ? n2629 : ~n2520;
  assign n2631 = pi15 ? n2626 : n2630;
  assign n2632 = pi14 ? n2621 : n2631;
  assign n2633 = pi13 ? n32 : n2632;
  assign n2634 = pi12 ? n32 : n2633;
  assign n2635 = pi11 ? n32 : n2634;
  assign n2636 = pi10 ? n32 : n2635;
  assign n2637 = pi18 ? n32 : n1166;
  assign n2638 = pi17 ? n2637 : ~n32;
  assign n2639 = pi16 ? n2513 : ~n2638;
  assign n2640 = pi18 ? n32 : n793;
  assign n2641 = pi17 ? n2640 : ~n32;
  assign n2642 = pi16 ? n2409 : ~n2641;
  assign n2643 = pi15 ? n2639 : n2642;
  assign n2644 = pi18 ? n32 : n805;
  assign n2645 = pi17 ? n2644 : ~n32;
  assign n2646 = pi16 ? n2415 : ~n2645;
  assign n2647 = pi16 ? n2120 : ~n2411;
  assign n2648 = pi15 ? n2646 : n2647;
  assign n2649 = pi14 ? n2643 : n2648;
  assign n2650 = pi18 ? n32 : n1266;
  assign n2651 = pi17 ? n2650 : ~n32;
  assign n2652 = pi16 ? n2426 : ~n2651;
  assign n2653 = pi18 ? n32 : n418;
  assign n2654 = pi17 ? n32 : n2653;
  assign n2655 = pi16 ? n2654 : ~n2321;
  assign n2656 = pi15 ? n2652 : n2655;
  assign n2657 = pi17 ? n2136 : ~n32;
  assign n2658 = pi16 ? n1815 : ~n2657;
  assign n2659 = pi15 ? n2541 : n2658;
  assign n2660 = pi14 ? n2656 : n2659;
  assign n2661 = pi13 ? n2649 : n2660;
  assign n2662 = pi19 ? n2250 : n32;
  assign n2663 = pi18 ? n32 : ~n2662;
  assign n2664 = pi17 ? n2663 : ~n32;
  assign n2665 = pi16 ? n1944 : ~n2664;
  assign n2666 = pi15 ? n2324 : n2665;
  assign n2667 = pi16 ? n1834 : ~n2434;
  assign n2668 = pi15 ? n2667 : n2439;
  assign n2669 = pi14 ? n2666 : n2668;
  assign n2670 = pi18 ? n1151 : ~n32;
  assign n2671 = pi17 ? n2670 : ~n32;
  assign n2672 = pi16 ? n1843 : ~n2671;
  assign n2673 = pi15 ? n1699 : n2672;
  assign n2674 = pi16 ? n1233 : ~n1698;
  assign n2675 = pi15 ? n2444 : n2674;
  assign n2676 = pi14 ? n2673 : n2675;
  assign n2677 = pi13 ? n2669 : n2676;
  assign n2678 = pi12 ? n2661 : n2677;
  assign n2679 = pi16 ? n1233 : ~n1583;
  assign n2680 = pi15 ? n1987 : n2679;
  assign n2681 = pi15 ? n2161 : n1986;
  assign n2682 = pi14 ? n2680 : n2681;
  assign n2683 = pi13 ? n2155 : n2682;
  assign n2684 = pi19 ? n857 : ~n32;
  assign n2685 = pi18 ? n2684 : ~n32;
  assign n2686 = pi17 ? n2685 : ~n32;
  assign n2687 = pi16 ? n1233 : ~n2686;
  assign n2688 = pi15 ? n2687 : n1991;
  assign n2689 = pi14 ? n1716 : n2688;
  assign n2690 = pi15 ? n2575 : n1716;
  assign n2691 = pi15 ? n1720 : n1999;
  assign n2692 = pi14 ? n2690 : n2691;
  assign n2693 = pi13 ? n2689 : n2692;
  assign n2694 = pi12 ? n2683 : n2693;
  assign n2695 = pi11 ? n2678 : n2694;
  assign n2696 = pi15 ? n1999 : n2463;
  assign n2697 = pi14 ? n2696 : n2467;
  assign n2698 = pi15 ? n1723 : n1597;
  assign n2699 = pi14 ? n2698 : n2357;
  assign n2700 = pi13 ? n2697 : n2699;
  assign n2701 = pi14 ? n2585 : n1724;
  assign n2702 = pi15 ? n1724 : n2357;
  assign n2703 = pi14 ? n2702 : n1497;
  assign n2704 = pi13 ? n2701 : n2703;
  assign n2705 = pi12 ? n2700 : n2704;
  assign n2706 = pi15 ? n1728 : n2599;
  assign n2707 = pi14 ? n2706 : n2599;
  assign n2708 = pi14 ? n2591 : n1852;
  assign n2709 = pi13 ? n2707 : n2708;
  assign n2710 = pi15 ? n1852 : n1497;
  assign n2711 = pi15 ? n1497 : n2606;
  assign n2712 = pi14 ? n2710 : n2711;
  assign n2713 = pi15 ? n2606 : n1723;
  assign n2714 = pi15 ? n1723 : n2467;
  assign n2715 = pi14 ? n2713 : n2714;
  assign n2716 = pi13 ? n2712 : n2715;
  assign n2717 = pi12 ? n2709 : n2716;
  assign n2718 = pi11 ? n2705 : n2717;
  assign n2719 = pi10 ? n2695 : n2718;
  assign n2720 = pi09 ? n2636 : n2719;
  assign n2721 = pi08 ? n2613 : n2720;
  assign n2722 = pi07 ? n2511 : n2721;
  assign n2723 = pi06 ? n2290 : n2722;
  assign n2724 = pi18 ? n32 : n962;
  assign n2725 = pi17 ? n32 : n2724;
  assign n2726 = pi18 ? n32 : n880;
  assign n2727 = pi17 ? n2726 : ~n32;
  assign n2728 = pi16 ? n2725 : ~n2727;
  assign n2729 = pi15 ? n32 : n2728;
  assign n2730 = pi19 ? n32 : n1941;
  assign n2731 = pi18 ? n32 : n2730;
  assign n2732 = pi17 ? n32 : n2731;
  assign n2733 = pi18 ? n32 : n684;
  assign n2734 = pi17 ? n2733 : ~n32;
  assign n2735 = pi16 ? n2732 : ~n2734;
  assign n2736 = pi18 ? n32 : n697;
  assign n2737 = pi17 ? n2736 : ~n32;
  assign n2738 = pi16 ? n2732 : ~n2737;
  assign n2739 = pi15 ? n2735 : n2738;
  assign n2740 = pi14 ? n2729 : n2739;
  assign n2741 = pi13 ? n32 : n2740;
  assign n2742 = pi12 ? n32 : n2741;
  assign n2743 = pi11 ? n32 : n2742;
  assign n2744 = pi10 ? n32 : n2743;
  assign n2745 = pi17 ? n32 : n2736;
  assign n2746 = pi16 ? n2745 : ~n2737;
  assign n2747 = pi19 ? n1320 : ~n32;
  assign n2748 = pi18 ? n32 : n2747;
  assign n2749 = pi17 ? n32 : n2748;
  assign n2750 = pi18 ? n32 : n702;
  assign n2751 = pi17 ? n2750 : ~n32;
  assign n2752 = pi16 ? n2749 : ~n2751;
  assign n2753 = pi15 ? n2746 : n2752;
  assign n2754 = pi19 ? n1840 : ~n32;
  assign n2755 = pi18 ? n32 : n2754;
  assign n2756 = pi17 ? n32 : n2755;
  assign n2757 = pi16 ? n2756 : ~n2514;
  assign n2758 = pi14 ? n2753 : n2757;
  assign n2759 = pi16 ? n2409 : ~n2514;
  assign n2760 = pi16 ? n2415 : ~n2520;
  assign n2761 = pi15 ? n2759 : n2760;
  assign n2762 = pi16 ? n2306 : ~n2294;
  assign n2763 = pi16 ? n1934 : ~n2294;
  assign n2764 = pi15 ? n2762 : n2763;
  assign n2765 = pi14 ? n2761 : n2764;
  assign n2766 = pi13 ? n2758 : n2765;
  assign n2767 = pi16 ? n2320 : ~n2651;
  assign n2768 = pi16 ? n2540 : ~n2301;
  assign n2769 = pi15 ? n2767 : n2768;
  assign n2770 = pi16 ? n1944 : ~n2321;
  assign n2771 = pi15 ? n2770 : n2545;
  assign n2772 = pi14 ? n2769 : n2771;
  assign n2773 = pi15 ? n1955 : n2550;
  assign n2774 = pi16 ? n1843 : ~n1935;
  assign n2775 = pi16 ? n1471 : ~n1953;
  assign n2776 = pi15 ? n2774 : n2775;
  assign n2777 = pi14 ? n2773 : n2776;
  assign n2778 = pi13 ? n2772 : n2777;
  assign n2779 = pi12 ? n2766 : n2778;
  assign n2780 = pi16 ? n1705 : ~n1679;
  assign n2781 = pi16 ? n1705 : ~n2333;
  assign n2782 = pi15 ? n2780 : n2781;
  assign n2783 = pi16 ? n931 : ~n1679;
  assign n2784 = pi16 ? n1135 : ~n1961;
  assign n2785 = pi15 ? n2783 : n2784;
  assign n2786 = pi14 ? n2782 : n2785;
  assign n2787 = pi16 ? n1233 : ~n1967;
  assign n2788 = pi15 ? n2787 : n2674;
  assign n2789 = pi16 ? n1233 : ~n2151;
  assign n2790 = pi16 ? n1233 : ~n2556;
  assign n2791 = pi15 ? n2789 : n2790;
  assign n2792 = pi14 ? n2788 : n2791;
  assign n2793 = pi13 ? n2786 : n2792;
  assign n2794 = pi16 ? n1233 : ~n1976;
  assign n2795 = pi15 ? n2155 : n2794;
  assign n2796 = pi14 ? n2155 : n2795;
  assign n2797 = pi14 ? n1980 : n2454;
  assign n2798 = pi13 ? n2796 : n2797;
  assign n2799 = pi12 ? n2793 : n2798;
  assign n2800 = pi11 ? n2779 : n2799;
  assign n2801 = pi15 ? n2569 : n1986;
  assign n2802 = pi14 ? n1988 : n2801;
  assign n2803 = pi15 ? n1986 : n2347;
  assign n2804 = pi15 ? n1991 : n1716;
  assign n2805 = pi14 ? n2803 : n2804;
  assign n2806 = pi13 ? n2802 : n2805;
  assign n2807 = pi15 ? n1716 : n2687;
  assign n2808 = pi15 ? n1720 : n1991;
  assign n2809 = pi14 ? n2807 : n2808;
  assign n2810 = pi15 ? n1991 : n2575;
  assign n2811 = pi15 ? n2463 : n1723;
  assign n2812 = pi14 ? n2810 : n2811;
  assign n2813 = pi13 ? n2809 : n2812;
  assign n2814 = pi12 ? n2806 : n2813;
  assign n2815 = pi13 ? n1723 : n1996;
  assign n2816 = pi19 ? n519 : ~n358;
  assign n2817 = pi18 ? n2816 : ~n32;
  assign n2818 = pi17 ? n2817 : ~n32;
  assign n2819 = pi16 ? n1233 : ~n2818;
  assign n2820 = pi15 ? n1996 : n2819;
  assign n2821 = pi15 ? n2463 : n1716;
  assign n2822 = pi14 ? n2820 : n2821;
  assign n2823 = pi15 ? n1716 : n1987;
  assign n2824 = pi14 ? n2823 : n1987;
  assign n2825 = pi13 ? n2822 : n2824;
  assign n2826 = pi12 ? n2815 : n2825;
  assign n2827 = pi11 ? n2814 : n2826;
  assign n2828 = pi10 ? n2800 : n2827;
  assign n2829 = pi09 ? n2744 : n2828;
  assign n2830 = pi19 ? n32 : n2303;
  assign n2831 = pi18 ? n32 : n2830;
  assign n2832 = pi17 ? n32 : n2831;
  assign n2833 = pi16 ? n2832 : ~n2727;
  assign n2834 = pi15 ? n32 : n2833;
  assign n2835 = pi19 ? n32 : n2317;
  assign n2836 = pi18 ? n32 : n2835;
  assign n2837 = pi17 ? n32 : n2836;
  assign n2838 = pi16 ? n2837 : ~n2734;
  assign n2839 = pi18 ? n32 : n590;
  assign n2840 = pi17 ? n32 : n2839;
  assign n2841 = pi16 ? n2840 : ~n2737;
  assign n2842 = pi15 ? n2838 : n2841;
  assign n2843 = pi14 ? n2834 : n2842;
  assign n2844 = pi13 ? n32 : n2843;
  assign n2845 = pi12 ? n32 : n2844;
  assign n2846 = pi11 ? n32 : n2845;
  assign n2847 = pi10 ? n32 : n2846;
  assign n2848 = pi20 ? n1839 : ~n32;
  assign n2849 = pi19 ? n32 : n2848;
  assign n2850 = pi18 ? n32 : n2849;
  assign n2851 = pi17 ? n32 : n2850;
  assign n2852 = pi18 ? n32 : n503;
  assign n2853 = pi17 ? n2852 : ~n32;
  assign n2854 = pi16 ? n2851 : ~n2853;
  assign n2855 = pi18 ? n32 : n1750;
  assign n2856 = pi17 ? n32 : n2855;
  assign n2857 = pi17 ? n2855 : ~n32;
  assign n2858 = pi16 ? n2856 : ~n2857;
  assign n2859 = pi15 ? n2854 : n2858;
  assign n2860 = pi17 ? n32 : n2750;
  assign n2861 = pi18 ? n32 : n2684;
  assign n2862 = pi17 ? n2861 : ~n32;
  assign n2863 = pi16 ? n2860 : ~n2862;
  assign n2864 = pi15 ? n2863 : n2515;
  assign n2865 = pi14 ? n2859 : n2864;
  assign n2866 = pi16 ? n2749 : ~n2619;
  assign n2867 = pi15 ? n2866 : n2760;
  assign n2868 = pi18 ? n32 : n1405;
  assign n2869 = pi17 ? n2868 : ~n32;
  assign n2870 = pi16 ? n2415 : ~n2869;
  assign n2871 = pi16 ? n2120 : ~n2294;
  assign n2872 = pi15 ? n2870 : n2871;
  assign n2873 = pi14 ? n2867 : n2872;
  assign n2874 = pi13 ? n2865 : n2873;
  assign n2875 = pi17 ? n2653 : ~n32;
  assign n2876 = pi16 ? n2426 : ~n2875;
  assign n2877 = pi16 ? n2654 : ~n2301;
  assign n2878 = pi15 ? n2876 : n2877;
  assign n2879 = pi16 ? n2540 : ~n2651;
  assign n2880 = pi18 ? n32 : n826;
  assign n2881 = pi17 ? n2880 : ~n32;
  assign n2882 = pi16 ? n1815 : ~n2881;
  assign n2883 = pi15 ? n2879 : n2882;
  assign n2884 = pi14 ? n2878 : n2883;
  assign n2885 = pi18 ? n858 : ~n359;
  assign n2886 = pi17 ? n2885 : ~n32;
  assign n2887 = pi16 ? n2137 : ~n2886;
  assign n2888 = pi16 ? n1944 : ~n2124;
  assign n2889 = pi15 ? n2887 : n2888;
  assign n2890 = pi16 ? n1834 : ~n2124;
  assign n2891 = pi16 ? n2144 : ~n1953;
  assign n2892 = pi15 ? n2890 : n2891;
  assign n2893 = pi14 ? n2889 : n2892;
  assign n2894 = pi13 ? n2884 : n2893;
  assign n2895 = pi12 ? n2874 : n2894;
  assign n2896 = pi16 ? n1594 : ~n2333;
  assign n2897 = pi16 ? n1594 : ~n1953;
  assign n2898 = pi15 ? n2896 : n2897;
  assign n2899 = pi18 ? n2197 : ~n32;
  assign n2900 = pi17 ? n2899 : ~n32;
  assign n2901 = pi16 ? n1594 : ~n2900;
  assign n2902 = pi16 ? n1843 : ~n1959;
  assign n2903 = pi15 ? n2901 : n2902;
  assign n2904 = pi14 ? n2898 : n2903;
  assign n2905 = pi16 ? n1479 : ~n1698;
  assign n2906 = pi19 ? n32 : n1337;
  assign n2907 = pi18 ? n2906 : ~n32;
  assign n2908 = pi17 ? n2907 : ~n32;
  assign n2909 = pi16 ? n1479 : ~n2908;
  assign n2910 = pi15 ? n2905 : n2909;
  assign n2911 = pi16 ? n1214 : ~n1961;
  assign n2912 = pi16 ? n931 : ~n2148;
  assign n2913 = pi15 ? n2911 : n2912;
  assign n2914 = pi14 ? n2910 : n2913;
  assign n2915 = pi13 ? n2904 : n2914;
  assign n2916 = pi16 ? n1233 : ~n1707;
  assign n2917 = pi15 ? n2155 : n2451;
  assign n2918 = pi18 ? n767 : ~n32;
  assign n2919 = pi17 ? n2918 : ~n32;
  assign n2920 = pi16 ? n1233 : ~n2919;
  assign n2921 = pi15 ? n2920 : n1980;
  assign n2922 = pi14 ? n2917 : n2921;
  assign n2923 = pi13 ? n2916 : n2922;
  assign n2924 = pi12 ? n2915 : n2923;
  assign n2925 = pi11 ? n2895 : n2924;
  assign n2926 = pi18 ? n967 : ~n32;
  assign n2927 = pi17 ? n2926 : ~n32;
  assign n2928 = pi16 ? n1233 : ~n2927;
  assign n2929 = pi15 ? n2161 : n2928;
  assign n2930 = pi14 ? n2680 : n2929;
  assign n2931 = pi14 ? n1987 : n2569;
  assign n2932 = pi13 ? n2930 : n2931;
  assign n2933 = pi15 ? n1716 : n1986;
  assign n2934 = pi14 ? n2933 : n2347;
  assign n2935 = pi15 ? n2347 : n1716;
  assign n2936 = pi15 ? n2687 : n2463;
  assign n2937 = pi14 ? n2935 : n2936;
  assign n2938 = pi13 ? n2934 : n2937;
  assign n2939 = pi12 ? n2932 : n2938;
  assign n2940 = pi13 ? n2463 : n1991;
  assign n2941 = pi15 ? n1991 : n2161;
  assign n2942 = pi15 ? n1991 : n1986;
  assign n2943 = pi14 ? n2941 : n2942;
  assign n2944 = pi15 ? n1986 : n2161;
  assign n2945 = pi14 ? n2944 : n2161;
  assign n2946 = pi13 ? n2943 : n2945;
  assign n2947 = pi12 ? n2940 : n2946;
  assign n2948 = pi11 ? n2939 : n2947;
  assign n2949 = pi10 ? n2925 : n2948;
  assign n2950 = pi09 ? n2847 : n2949;
  assign n2951 = pi08 ? n2829 : n2950;
  assign n2952 = pi18 ? n32 : n341;
  assign n2953 = pi17 ? n32 : n2952;
  assign n2954 = pi18 ? n32 : n863;
  assign n2955 = pi17 ? n2954 : ~n32;
  assign n2956 = pi16 ? n2953 : ~n2955;
  assign n2957 = pi15 ? n32 : n2956;
  assign n2958 = pi17 ? n32 : n2726;
  assign n2959 = pi18 ? n32 : n209;
  assign n2960 = pi17 ? n2959 : ~n32;
  assign n2961 = pi16 ? n2958 : ~n2960;
  assign n2962 = pi19 ? n32 : n2297;
  assign n2963 = pi18 ? n32 : n2962;
  assign n2964 = pi17 ? n32 : n2963;
  assign n2965 = pi16 ? n2964 : ~n2734;
  assign n2966 = pi15 ? n2961 : n2965;
  assign n2967 = pi14 ? n2957 : n2966;
  assign n2968 = pi13 ? n32 : n2967;
  assign n2969 = pi12 ? n32 : n2968;
  assign n2970 = pi11 ? n32 : n2969;
  assign n2971 = pi10 ? n32 : n2970;
  assign n2972 = pi16 ? n2732 : ~n2727;
  assign n2973 = pi15 ? n2965 : n2972;
  assign n2974 = pi14 ? n2973 : n2746;
  assign n2975 = pi16 ? n2617 : ~n2734;
  assign n2976 = pi16 ? n2518 : ~n2751;
  assign n2977 = pi15 ? n2975 : n2976;
  assign n2978 = pi16 ? n2756 : ~n2751;
  assign n2979 = pi14 ? n2977 : n2978;
  assign n2980 = pi13 ? n2974 : n2979;
  assign n2981 = pi16 ? n2409 : ~n2737;
  assign n2982 = pi16 ? n2415 : ~n2625;
  assign n2983 = pi15 ? n2981 : n2982;
  assign n2984 = pi16 ? n2306 : ~n2520;
  assign n2985 = pi16 ? n1934 : ~n2532;
  assign n2986 = pi15 ? n2984 : n2985;
  assign n2987 = pi14 ? n2983 : n2986;
  assign n2988 = pi16 ? n2320 : ~n2301;
  assign n2989 = pi15 ? n2988 : n2768;
  assign n2990 = pi16 ? n1944 : ~n2301;
  assign n2991 = pi16 ? n2326 : ~n2301;
  assign n2992 = pi15 ? n2990 : n2991;
  assign n2993 = pi14 ? n2989 : n2992;
  assign n2994 = pi13 ? n2987 : n2993;
  assign n2995 = pi12 ? n2980 : n2994;
  assign n2996 = pi16 ? n1577 : ~n2321;
  assign n2997 = pi16 ? n1577 : ~n2544;
  assign n2998 = pi15 ? n2997 : n2550;
  assign n2999 = pi14 ? n2996 : n2998;
  assign n3000 = pi16 ? n1323 : ~n2434;
  assign n3001 = pi16 ? n1323 : ~n1935;
  assign n3002 = pi15 ? n3000 : n3001;
  assign n3003 = pi16 ? n1594 : ~n1935;
  assign n3004 = pi15 ? n3001 : n3003;
  assign n3005 = pi14 ? n3002 : n3004;
  assign n3006 = pi13 ? n2999 : n3005;
  assign n3007 = pi16 ? n1471 : ~n1809;
  assign n3008 = pi16 ? n1471 : ~n2900;
  assign n3009 = pi15 ? n3007 : n3008;
  assign n3010 = pi16 ? n1972 : ~n1809;
  assign n3011 = pi16 ? n1214 : ~n1679;
  assign n3012 = pi15 ? n3010 : n3011;
  assign n3013 = pi14 ? n3009 : n3012;
  assign n3014 = pi16 ? n931 : ~n1961;
  assign n3015 = pi16 ? n931 : ~n1953;
  assign n3016 = pi15 ? n3014 : n3015;
  assign n3017 = pi16 ? n1233 : ~n2671;
  assign n3018 = pi15 ? n2784 : n3017;
  assign n3019 = pi14 ? n3016 : n3018;
  assign n3020 = pi13 ? n3013 : n3019;
  assign n3021 = pi12 ? n3006 : n3020;
  assign n3022 = pi11 ? n2995 : n3021;
  assign n3023 = pi16 ? n1233 : ~n2148;
  assign n3024 = pi16 ? n1233 : ~n2447;
  assign n3025 = pi15 ? n3023 : n3024;
  assign n3026 = pi14 ? n3025 : n2787;
  assign n3027 = pi13 ? n2674 : n3026;
  assign n3028 = pi15 ? n2916 : n2155;
  assign n3029 = pi15 ? n2155 : n1987;
  assign n3030 = pi14 ? n3028 : n3029;
  assign n3031 = pi13 ? n2916 : n3030;
  assign n3032 = pi12 ? n3027 : n3031;
  assign n3033 = pi15 ? n2679 : n1980;
  assign n3034 = pi14 ? n2679 : n3033;
  assign n3035 = pi13 ? n3034 : n2794;
  assign n3036 = pi15 ? n1980 : n2790;
  assign n3037 = pi14 ? n2916 : n3036;
  assign n3038 = pi16 ? n1233 : ~n1961;
  assign n3039 = pi15 ? n2790 : n3038;
  assign n3040 = pi14 ? n3039 : n3038;
  assign n3041 = pi13 ? n3037 : n3040;
  assign n3042 = pi12 ? n3035 : n3041;
  assign n3043 = pi11 ? n3032 : n3042;
  assign n3044 = pi10 ? n3022 : n3043;
  assign n3045 = pi09 ? n2971 : n3044;
  assign n3046 = pi18 ? n32 : n1477;
  assign n3047 = pi17 ? n32 : n3046;
  assign n3048 = pi16 ? n3047 : ~n2955;
  assign n3049 = pi15 ? n32 : n3048;
  assign n3050 = pi18 ? n32 : n245;
  assign n3051 = pi17 ? n32 : n3050;
  assign n3052 = pi16 ? n3051 : ~n2960;
  assign n3053 = pi16 ? n3051 : ~n2734;
  assign n3054 = pi15 ? n3052 : n3053;
  assign n3055 = pi14 ? n3049 : n3054;
  assign n3056 = pi13 ? n32 : n3055;
  assign n3057 = pi12 ? n32 : n3056;
  assign n3058 = pi11 ? n32 : n3057;
  assign n3059 = pi10 ? n32 : n3058;
  assign n3060 = pi16 ? n2953 : ~n2734;
  assign n3061 = pi17 ? n32 : n2733;
  assign n3062 = pi17 ? n2952 : ~n32;
  assign n3063 = pi16 ? n3061 : ~n3062;
  assign n3064 = pi15 ? n3060 : n3063;
  assign n3065 = pi15 ? n2841 : n2854;
  assign n3066 = pi14 ? n3064 : n3065;
  assign n3067 = pi18 ? n32 : n496;
  assign n3068 = pi17 ? n32 : n3067;
  assign n3069 = pi16 ? n3068 : ~n2734;
  assign n3070 = pi18 ? n32 : n772;
  assign n3071 = pi17 ? n3070 : ~n32;
  assign n3072 = pi16 ? n2624 : ~n3071;
  assign n3073 = pi15 ? n3069 : n3072;
  assign n3074 = pi16 ? n2860 : ~n2751;
  assign n3075 = pi16 ? n2513 : ~n2751;
  assign n3076 = pi15 ? n3074 : n3075;
  assign n3077 = pi14 ? n3073 : n3076;
  assign n3078 = pi13 ? n3066 : n3077;
  assign n3079 = pi16 ? n2749 : ~n2737;
  assign n3080 = pi16 ? n2415 : ~n2862;
  assign n3081 = pi15 ? n3079 : n3080;
  assign n3082 = pi16 ? n2120 : ~n2875;
  assign n3083 = pi15 ? n2982 : n3082;
  assign n3084 = pi14 ? n3081 : n3083;
  assign n3085 = pi16 ? n2426 : ~n2301;
  assign n3086 = pi15 ? n3085 : n2877;
  assign n3087 = pi16 ? n2540 : ~n2411;
  assign n3088 = pi16 ? n1815 : ~n2411;
  assign n3089 = pi15 ? n3087 : n3088;
  assign n3090 = pi14 ? n3086 : n3089;
  assign n3091 = pi13 ? n3084 : n3090;
  assign n3092 = pi12 ? n3078 : n3091;
  assign n3093 = pi18 ? n32 : n1078;
  assign n3094 = pi17 ? n3093 : ~n32;
  assign n3095 = pi16 ? n2137 : ~n3094;
  assign n3096 = pi16 ? n2137 : ~n2544;
  assign n3097 = pi15 ? n3096 : n2888;
  assign n3098 = pi14 ? n3095 : n3097;
  assign n3099 = pi16 ? n1683 : ~n2544;
  assign n3100 = pi18 ? n32 : ~n359;
  assign n3101 = pi17 ? n3100 : ~n32;
  assign n3102 = pi16 ? n1683 : ~n3101;
  assign n3103 = pi15 ? n3099 : n3102;
  assign n3104 = pi16 ? n1577 : ~n1935;
  assign n3105 = pi15 ? n3102 : n3104;
  assign n3106 = pi14 ? n3103 : n3105;
  assign n3107 = pi13 ? n3098 : n3106;
  assign n3108 = pi16 ? n1581 : ~n2900;
  assign n3109 = pi16 ? n1581 : ~n1945;
  assign n3110 = pi15 ? n3108 : n3109;
  assign n3111 = pi16 ? n1581 : ~n2134;
  assign n3112 = pi18 ? n1370 : ~n32;
  assign n3113 = pi17 ? n3112 : ~n32;
  assign n3114 = pi16 ? n1323 : ~n3113;
  assign n3115 = pi15 ? n3111 : n3114;
  assign n3116 = pi14 ? n3110 : n3115;
  assign n3117 = pi15 ? n1960 : n2897;
  assign n3118 = pi17 ? n1704 : ~n32;
  assign n3119 = pi16 ? n1479 : ~n3118;
  assign n3120 = pi16 ? n1705 : ~n3118;
  assign n3121 = pi15 ? n3119 : n3120;
  assign n3122 = pi14 ? n3117 : n3121;
  assign n3123 = pi13 ? n3116 : n3122;
  assign n3124 = pi12 ? n3107 : n3123;
  assign n3125 = pi11 ? n3092 : n3124;
  assign n3126 = pi15 ? n2558 : n2340;
  assign n3127 = pi14 ? n3126 : n2913;
  assign n3128 = pi16 ? n1135 : ~n2148;
  assign n3129 = pi14 ? n3128 : n2674;
  assign n3130 = pi13 ? n3127 : n3129;
  assign n3131 = pi15 ? n2790 : n2674;
  assign n3132 = pi14 ? n3131 : n2787;
  assign n3133 = pi15 ? n2916 : n1980;
  assign n3134 = pi14 ? n2787 : n3133;
  assign n3135 = pi13 ? n3132 : n3134;
  assign n3136 = pi12 ? n3130 : n3135;
  assign n3137 = pi15 ? n1980 : n2155;
  assign n3138 = pi14 ? n3137 : n2155;
  assign n3139 = pi15 ? n2916 : n2787;
  assign n3140 = pi14 ? n3139 : n2787;
  assign n3141 = pi13 ? n3138 : n3140;
  assign n3142 = pi15 ? n2787 : n3024;
  assign n3143 = pi15 ? n2451 : n3023;
  assign n3144 = pi14 ? n3142 : n3143;
  assign n3145 = pi16 ? n1233 : ~n3118;
  assign n3146 = pi15 ? n3023 : n3145;
  assign n3147 = pi14 ? n3146 : n3145;
  assign n3148 = pi13 ? n3144 : n3147;
  assign n3149 = pi12 ? n3141 : n3148;
  assign n3150 = pi11 ? n3136 : n3149;
  assign n3151 = pi10 ? n3125 : n3150;
  assign n3152 = pi09 ? n3059 : n3151;
  assign n3153 = pi08 ? n3045 : n3152;
  assign n3154 = pi07 ? n2951 : n3153;
  assign n3155 = pi18 ? n32 : n2142;
  assign n3156 = pi17 ? n32 : n3155;
  assign n3157 = pi17 ? n32 : n1227;
  assign n3158 = pi16 ? n3156 : ~n3157;
  assign n3159 = pi15 ? n32 : n3158;
  assign n3160 = pi18 ? n32 : n1841;
  assign n3161 = pi17 ? n32 : n3160;
  assign n3162 = pi17 ? n32 : n1500;
  assign n3163 = pi16 ? n3161 : ~n3162;
  assign n3164 = pi18 ? n32 : n940;
  assign n3165 = pi17 ? n32 : n3164;
  assign n3166 = pi17 ? n32 : ~n32;
  assign n3167 = pi16 ? n3165 : ~n3166;
  assign n3168 = pi15 ? n3163 : n3167;
  assign n3169 = pi14 ? n3159 : n3168;
  assign n3170 = pi13 ? n32 : n3169;
  assign n3171 = pi12 ? n32 : n3170;
  assign n3172 = pi11 ? n32 : n3171;
  assign n3173 = pi10 ? n32 : n3172;
  assign n3174 = pi16 ? n2953 : ~n3166;
  assign n3175 = pi18 ? n32 : n366;
  assign n3176 = pi17 ? n32 : n3175;
  assign n3177 = pi17 ? n32 : n1028;
  assign n3178 = pi16 ? n3176 : ~n3177;
  assign n3179 = pi15 ? n3174 : n3178;
  assign n3180 = pi17 ? n3164 : ~n32;
  assign n3181 = pi16 ? n2964 : ~n3180;
  assign n3182 = pi18 ? n32 : n1965;
  assign n3183 = pi17 ? n32 : n3182;
  assign n3184 = pi16 ? n3183 : ~n2960;
  assign n3185 = pi15 ? n3181 : n3184;
  assign n3186 = pi14 ? n3179 : n3185;
  assign n3187 = pi16 ? n3183 : ~n3166;
  assign n3188 = pi16 ? n2745 : ~n3180;
  assign n3189 = pi15 ? n3187 : n3188;
  assign n3190 = pi16 ? n2745 : ~n2734;
  assign n3191 = pi14 ? n3189 : n3190;
  assign n3192 = pi13 ? n3186 : n3191;
  assign n3193 = pi16 ? n2617 : ~n2727;
  assign n3194 = pi17 ? n3067 : ~n32;
  assign n3195 = pi16 ? n2518 : ~n3194;
  assign n3196 = pi15 ? n3193 : n3195;
  assign n3197 = pi16 ? n2756 : ~n2737;
  assign n3198 = pi15 ? n3197 : n2978;
  assign n3199 = pi14 ? n3196 : n3198;
  assign n3200 = pi19 ? n594 : n236;
  assign n3201 = pi18 ? n32 : n3200;
  assign n3202 = pi17 ? n3201 : ~n32;
  assign n3203 = pi16 ? n2409 : ~n3202;
  assign n3204 = pi16 ? n2415 : ~n2751;
  assign n3205 = pi15 ? n3203 : n3204;
  assign n3206 = pi16 ? n2306 : ~n2514;
  assign n3207 = pi16 ? n1934 : ~n2514;
  assign n3208 = pi15 ? n3206 : n3207;
  assign n3209 = pi14 ? n3205 : n3208;
  assign n3210 = pi13 ? n3199 : n3209;
  assign n3211 = pi12 ? n3192 : n3210;
  assign n3212 = pi16 ? n2320 : ~n2875;
  assign n3213 = pi16 ? n2320 : ~n2294;
  assign n3214 = pi15 ? n3212 : n3213;
  assign n3215 = pi16 ? n1808 : ~n2645;
  assign n3216 = pi15 ? n3213 : n3215;
  assign n3217 = pi14 ? n3214 : n3216;
  assign n3218 = pi16 ? n1815 : ~n2532;
  assign n3219 = pi16 ? n1815 : ~n2301;
  assign n3220 = pi16 ? n2137 : ~n2301;
  assign n3221 = pi15 ? n3219 : n3220;
  assign n3222 = pi14 ? n3218 : n3221;
  assign n3223 = pi13 ? n3217 : n3222;
  assign n3224 = pi16 ? n1678 : ~n2301;
  assign n3225 = pi15 ? n3224 : n3099;
  assign n3226 = pi14 ? n3224 : n3225;
  assign n3227 = pi16 ? n1834 : ~n2321;
  assign n3228 = pi16 ? n1834 : ~n2315;
  assign n3229 = pi16 ? n2144 : ~n2544;
  assign n3230 = pi15 ? n3228 : n3229;
  assign n3231 = pi14 ? n3227 : n3230;
  assign n3232 = pi13 ? n3226 : n3231;
  assign n3233 = pi12 ? n3223 : n3232;
  assign n3234 = pi11 ? n3211 : n3233;
  assign n3235 = pi16 ? n1581 : ~n2434;
  assign n3236 = pi16 ? n1581 : ~n2124;
  assign n3237 = pi15 ? n3235 : n3236;
  assign n3238 = pi16 ? n1471 : ~n3101;
  assign n3239 = pi15 ? n2774 : n3238;
  assign n3240 = pi14 ? n3237 : n3239;
  assign n3241 = pi16 ? n1479 : ~n1935;
  assign n3242 = pi19 ? n32 : n161;
  assign n3243 = pi18 ? n32 : n3242;
  assign n3244 = pi17 ? n1580 : ~n3243;
  assign n3245 = pi16 ? n1479 : ~n3244;
  assign n3246 = pi15 ? n3241 : n3245;
  assign n3247 = pi16 ? n1705 : ~n2434;
  assign n3248 = pi14 ? n3246 : n3247;
  assign n3249 = pi13 ? n3240 : n3248;
  assign n3250 = pi16 ? n1972 : ~n1953;
  assign n3251 = pi16 ? n1214 : ~n2134;
  assign n3252 = pi14 ? n3250 : n3251;
  assign n3253 = pi16 ? n1233 : ~n1953;
  assign n3254 = pi16 ? n1233 : ~n1679;
  assign n3255 = pi17 ? n1213 : ~n2054;
  assign n3256 = pi16 ? n1233 : ~n3255;
  assign n3257 = pi15 ? n3254 : n3256;
  assign n3258 = pi14 ? n3253 : n3257;
  assign n3259 = pi13 ? n3252 : n3258;
  assign n3260 = pi12 ? n3249 : n3259;
  assign n3261 = pi14 ? n3038 : n3254;
  assign n3262 = pi14 ? n3254 : n3253;
  assign n3263 = pi13 ? n3261 : n3262;
  assign n3264 = pi17 ? n1580 : ~n1787;
  assign n3265 = pi16 ? n1233 : ~n3264;
  assign n3266 = pi15 ? n3253 : n3265;
  assign n3267 = pi16 ? n1135 : ~n1935;
  assign n3268 = pi15 ? n3253 : n3267;
  assign n3269 = pi14 ? n3266 : n3268;
  assign n3270 = pi16 ? n1135 : ~n2544;
  assign n3271 = pi15 ? n3267 : n3270;
  assign n3272 = pi16 ? n1972 : ~n2544;
  assign n3273 = pi15 ? n3270 : n3272;
  assign n3274 = pi14 ? n3271 : n3273;
  assign n3275 = pi13 ? n3269 : n3274;
  assign n3276 = pi12 ? n3263 : n3275;
  assign n3277 = pi11 ? n3260 : n3276;
  assign n3278 = pi10 ? n3234 : n3277;
  assign n3279 = pi09 ? n3173 : n3278;
  assign n3280 = pi16 ? n32 : ~n3157;
  assign n3281 = pi15 ? n32 : n3280;
  assign n3282 = pi18 ? n32 : n936;
  assign n3283 = pi17 ? n32 : n3282;
  assign n3284 = pi16 ? n3283 : ~n3162;
  assign n3285 = pi15 ? n3284 : n3167;
  assign n3286 = pi14 ? n3281 : n3285;
  assign n3287 = pi13 ? n32 : n3286;
  assign n3288 = pi12 ? n32 : n3287;
  assign n3289 = pi11 ? n32 : n3288;
  assign n3290 = pi10 ? n32 : n3289;
  assign n3291 = pi16 ? n3047 : ~n3166;
  assign n3292 = pi18 ? n32 : n751;
  assign n3293 = pi17 ? n32 : n3292;
  assign n3294 = pi16 ? n3293 : ~n3177;
  assign n3295 = pi15 ? n3291 : n3294;
  assign n3296 = pi18 ? n32 : n1370;
  assign n3297 = pi17 ? n3296 : ~n32;
  assign n3298 = pi16 ? n2953 : ~n3297;
  assign n3299 = pi16 ? n2953 : ~n2960;
  assign n3300 = pi15 ? n3298 : n3299;
  assign n3301 = pi14 ? n3295 : n3300;
  assign n3302 = pi16 ? n3176 : ~n3166;
  assign n3303 = pi16 ? n2837 : ~n3180;
  assign n3304 = pi15 ? n3302 : n3303;
  assign n3305 = pi16 ? n2840 : ~n2734;
  assign n3306 = pi16 ? n2851 : ~n2734;
  assign n3307 = pi15 ? n3305 : n3306;
  assign n3308 = pi14 ? n3304 : n3307;
  assign n3309 = pi13 ? n3301 : n3308;
  assign n3310 = pi16 ? n3068 : ~n2727;
  assign n3311 = pi16 ? n2624 : ~n3194;
  assign n3312 = pi15 ? n3310 : n3311;
  assign n3313 = pi16 ? n2860 : ~n2737;
  assign n3314 = pi16 ? n2513 : ~n2857;
  assign n3315 = pi15 ? n3313 : n3314;
  assign n3316 = pi14 ? n3312 : n3315;
  assign n3317 = pi15 ? n3079 : n3204;
  assign n3318 = pi16 ? n2415 : ~n2619;
  assign n3319 = pi16 ? n2120 : ~n2514;
  assign n3320 = pi15 ? n3318 : n3319;
  assign n3321 = pi14 ? n3317 : n3320;
  assign n3322 = pi13 ? n3316 : n3321;
  assign n3323 = pi12 ? n3309 : n3322;
  assign n3324 = pi16 ? n2426 : ~n2869;
  assign n3325 = pi19 ? n2201 : ~n32;
  assign n3326 = pi18 ? n32 : n3325;
  assign n3327 = pi17 ? n3326 : ~n32;
  assign n3328 = pi16 ? n2426 : ~n3327;
  assign n3329 = pi15 ? n3324 : n3328;
  assign n3330 = pi16 ? n2530 : ~n2869;
  assign n3331 = pi15 ? n3330 : n2762;
  assign n3332 = pi14 ? n3329 : n3331;
  assign n3333 = pi18 ? n32 : n423;
  assign n3334 = pi17 ? n3333 : ~n32;
  assign n3335 = pi16 ? n1934 : ~n3334;
  assign n3336 = pi19 ? n2848 : ~n32;
  assign n3337 = pi18 ? n32 : n3336;
  assign n3338 = pi17 ? n32 : n3337;
  assign n3339 = pi16 ? n3338 : ~n3334;
  assign n3340 = pi15 ? n3335 : n3339;
  assign n3341 = pi14 ? n2985 : n3340;
  assign n3342 = pi13 ? n3332 : n3341;
  assign n3343 = pi16 ? n1808 : ~n2411;
  assign n3344 = pi16 ? n1808 : ~n2301;
  assign n3345 = pi18 ? n32 : n2182;
  assign n3346 = pi17 ? n3345 : ~n32;
  assign n3347 = pi16 ? n1815 : ~n3346;
  assign n3348 = pi15 ? n3344 : n3347;
  assign n3349 = pi14 ? n3343 : n3348;
  assign n3350 = pi19 ? n2614 : ~n32;
  assign n3351 = pi18 ? n32 : n3350;
  assign n3352 = pi17 ? n32 : n3351;
  assign n3353 = pi16 ? n3352 : ~n3094;
  assign n3354 = pi16 ? n3352 : ~n2321;
  assign n3355 = pi15 ? n3353 : n3354;
  assign n3356 = pi17 ? n32 : n2123;
  assign n3357 = pi16 ? n3356 : ~n2544;
  assign n3358 = pi15 ? n3354 : n3357;
  assign n3359 = pi14 ? n3355 : n3358;
  assign n3360 = pi13 ? n3349 : n3359;
  assign n3361 = pi12 ? n3342 : n3360;
  assign n3362 = pi11 ? n3323 : n3361;
  assign n3363 = pi16 ? n1683 : ~n2315;
  assign n3364 = pi15 ? n3099 : n3363;
  assign n3365 = pi15 ? n3102 : n2997;
  assign n3366 = pi14 ? n3364 : n3365;
  assign n3367 = pi18 ? n936 : n822;
  assign n3368 = pi17 ? n3367 : ~n3243;
  assign n3369 = pi16 ? n1834 : ~n3368;
  assign n3370 = pi15 ? n2550 : n3369;
  assign n3371 = pi16 ? n1323 : ~n2124;
  assign n3372 = pi14 ? n3370 : n3371;
  assign n3373 = pi13 ? n3366 : n3372;
  assign n3374 = pi16 ? n1594 : ~n2134;
  assign n3375 = pi15 ? n2897 : n3374;
  assign n3376 = pi14 ? n3375 : n2774;
  assign n3377 = pi16 ? n1471 : ~n1945;
  assign n3378 = pi15 ? n2775 : n3377;
  assign n3379 = pi16 ? n1479 : ~n1679;
  assign n3380 = pi18 ? n1139 : ~n32;
  assign n3381 = pi17 ? n3380 : ~n32;
  assign n3382 = pi16 ? n1479 : ~n3381;
  assign n3383 = pi15 ? n3379 : n3382;
  assign n3384 = pi14 ? n3378 : n3383;
  assign n3385 = pi13 ? n3376 : n3384;
  assign n3386 = pi12 ? n3373 : n3385;
  assign n3387 = pi16 ? n931 : ~n3381;
  assign n3388 = pi18 ? n2202 : ~n32;
  assign n3389 = pi17 ? n3388 : ~n32;
  assign n3390 = pi16 ? n1135 : ~n3389;
  assign n3391 = pi15 ? n3387 : n3390;
  assign n3392 = pi16 ? n1135 : ~n2333;
  assign n3393 = pi14 ? n3391 : n3392;
  assign n3394 = pi16 ? n931 : ~n2333;
  assign n3395 = pi16 ? n931 : ~n3113;
  assign n3396 = pi15 ? n3394 : n3395;
  assign n3397 = pi16 ? n1705 : ~n2134;
  assign n3398 = pi17 ? n2133 : ~n2073;
  assign n3399 = pi16 ? n1705 : ~n3398;
  assign n3400 = pi15 ? n3397 : n3399;
  assign n3401 = pi14 ? n3396 : n3400;
  assign n3402 = pi13 ? n3393 : n3401;
  assign n3403 = pi16 ? n1705 : ~n2886;
  assign n3404 = pi15 ? n3397 : n3403;
  assign n3405 = pi16 ? n1972 : ~n1945;
  assign n3406 = pi17 ? n3100 : ~n646;
  assign n3407 = pi16 ? n1479 : ~n3406;
  assign n3408 = pi15 ? n3405 : n3407;
  assign n3409 = pi14 ? n3404 : n3408;
  assign n3410 = pi16 ? n1479 : ~n3101;
  assign n3411 = pi16 ? n1594 : ~n2544;
  assign n3412 = pi15 ? n3410 : n3411;
  assign n3413 = pi16 ? n1594 : ~n2315;
  assign n3414 = pi16 ? n1594 : ~n2321;
  assign n3415 = pi15 ? n3413 : n3414;
  assign n3416 = pi14 ? n3412 : n3415;
  assign n3417 = pi13 ? n3409 : n3416;
  assign n3418 = pi12 ? n3402 : n3417;
  assign n3419 = pi11 ? n3386 : n3418;
  assign n3420 = pi10 ? n3362 : n3419;
  assign n3421 = pi09 ? n3290 : n3420;
  assign n3422 = pi08 ? n3279 : n3421;
  assign n3423 = pi17 ? n2005 : ~n1718;
  assign n3424 = pi16 ? n32 : n3423;
  assign n3425 = pi15 ? n32 : n3424;
  assign n3426 = pi17 ? n1028 : ~n1718;
  assign n3427 = pi16 ? n32 : n3426;
  assign n3428 = pi17 ? n32 : n2355;
  assign n3429 = pi16 ? n3283 : ~n3428;
  assign n3430 = pi15 ? n3427 : n3429;
  assign n3431 = pi14 ? n3425 : n3430;
  assign n3432 = pi13 ? n32 : n3431;
  assign n3433 = pi12 ? n32 : n3432;
  assign n3434 = pi11 ? n32 : n3433;
  assign n3435 = pi10 ? n32 : n3434;
  assign n3436 = pi17 ? n32 : n1219;
  assign n3437 = pi16 ? n3156 : ~n3436;
  assign n3438 = pi17 ? n32 : n2954;
  assign n3439 = pi16 ? n3438 : ~n3428;
  assign n3440 = pi15 ? n3437 : n3439;
  assign n3441 = pi16 ? n3165 : ~n3162;
  assign n3442 = pi15 ? n3441 : n3291;
  assign n3443 = pi14 ? n3440 : n3442;
  assign n3444 = pi16 ? n2958 : ~n3162;
  assign n3445 = pi15 ? n3178 : n3444;
  assign n3446 = pi16 ? n2964 : ~n3166;
  assign n3447 = pi18 ? n32 : n1139;
  assign n3448 = pi17 ? n3447 : ~n32;
  assign n3449 = pi16 ? n3183 : ~n3448;
  assign n3450 = pi15 ? n3446 : n3449;
  assign n3451 = pi14 ? n3445 : n3450;
  assign n3452 = pi13 ? n3443 : n3451;
  assign n3453 = pi16 ? n3183 : ~n2727;
  assign n3454 = pi15 ? n3453 : n3188;
  assign n3455 = pi14 ? n3454 : n3190;
  assign n3456 = pi16 ? n2518 : ~n2737;
  assign n3457 = pi15 ? n2975 : n3456;
  assign n3458 = pi14 ? n3457 : n3197;
  assign n3459 = pi13 ? n3455 : n3458;
  assign n3460 = pi12 ? n3452 : n3459;
  assign n3461 = pi16 ? n2409 : ~n3194;
  assign n3462 = pi15 ? n3461 : n2981;
  assign n3463 = pi16 ? n2409 : ~n2751;
  assign n3464 = pi15 ? n3463 : n3204;
  assign n3465 = pi14 ? n3462 : n3464;
  assign n3466 = pi16 ? n2120 : ~n2751;
  assign n3467 = pi16 ? n2120 : ~n2737;
  assign n3468 = pi15 ? n3466 : n3467;
  assign n3469 = pi16 ? n2300 : ~n2514;
  assign n3470 = pi16 ? n2530 : ~n2514;
  assign n3471 = pi15 ? n3469 : n3470;
  assign n3472 = pi14 ? n3468 : n3471;
  assign n3473 = pi13 ? n3465 : n3472;
  assign n3474 = pi15 ? n2762 : n2984;
  assign n3475 = pi17 ? n2408 : ~n32;
  assign n3476 = pi16 ? n2540 : ~n3475;
  assign n3477 = pi15 ? n3206 : n3476;
  assign n3478 = pi14 ? n3474 : n3477;
  assign n3479 = pi16 ? n2540 : ~n2294;
  assign n3480 = pi16 ? n2540 : ~n2645;
  assign n3481 = pi16 ? n3338 : ~n2532;
  assign n3482 = pi15 ? n3480 : n3481;
  assign n3483 = pi14 ? n3479 : n3482;
  assign n3484 = pi13 ? n3478 : n3483;
  assign n3485 = pi12 ? n3473 : n3484;
  assign n3486 = pi11 ? n3460 : n3485;
  assign n3487 = pi16 ? n1944 : ~n2294;
  assign n3488 = pi16 ? n1944 : ~n2875;
  assign n3489 = pi15 ? n3487 : n3488;
  assign n3490 = pi16 ? n1944 : ~n2532;
  assign n3491 = pi16 ? n2326 : ~n3334;
  assign n3492 = pi15 ? n3490 : n3491;
  assign n3493 = pi14 ? n3489 : n3492;
  assign n3494 = pi16 ? n3356 : ~n2532;
  assign n3495 = pi20 ? n1817 : n32;
  assign n3496 = pi19 ? n32 : n3495;
  assign n3497 = pi18 ? n32 : n3496;
  assign n3498 = pi17 ? n2531 : ~n3497;
  assign n3499 = pi16 ? n3356 : ~n3498;
  assign n3500 = pi15 ? n3494 : n3499;
  assign n3501 = pi14 ? n3500 : n3494;
  assign n3502 = pi13 ? n3493 : n3501;
  assign n3503 = pi16 ? n1678 : ~n2651;
  assign n3504 = pi16 ? n1834 : ~n2301;
  assign n3505 = pi14 ? n3503 : n3504;
  assign n3506 = pi16 ? n2144 : ~n3094;
  assign n3507 = pi20 ? n2385 : ~n32;
  assign n3508 = pi19 ? n3507 : ~n32;
  assign n3509 = pi18 ? n32 : n3508;
  assign n3510 = pi17 ? n3509 : ~n32;
  assign n3511 = pi16 ? n1581 : ~n3510;
  assign n3512 = pi17 ? n3509 : ~n1527;
  assign n3513 = pi16 ? n1581 : ~n3512;
  assign n3514 = pi15 ? n3511 : n3513;
  assign n3515 = pi14 ? n3506 : n3514;
  assign n3516 = pi13 ? n3505 : n3515;
  assign n3517 = pi12 ? n3502 : n3516;
  assign n3518 = pi16 ? n1323 : ~n3510;
  assign n3519 = pi16 ? n1479 : ~n2881;
  assign n3520 = pi15 ? n3518 : n3519;
  assign n3521 = pi16 ? n1479 : ~n2538;
  assign n3522 = pi14 ? n3520 : n3521;
  assign n3523 = pi21 ? n32 : n309;
  assign n3524 = pi20 ? n3523 : ~n32;
  assign n3525 = pi19 ? n3524 : ~n32;
  assign n3526 = pi18 ? n32 : n3525;
  assign n3527 = pi17 ? n3526 : ~n32;
  assign n3528 = pi16 ? n1323 : ~n3527;
  assign n3529 = pi16 ? n1323 : ~n2651;
  assign n3530 = pi15 ? n3528 : n3529;
  assign n3531 = pi16 ? n1323 : ~n2411;
  assign n3532 = pi17 ? n2410 : ~n2073;
  assign n3533 = pi16 ? n1323 : ~n3532;
  assign n3534 = pi15 ? n3531 : n3533;
  assign n3535 = pi14 ? n3530 : n3534;
  assign n3536 = pi13 ? n3522 : n3535;
  assign n3537 = pi17 ? n2410 : ~n2080;
  assign n3538 = pi16 ? n1323 : ~n3537;
  assign n3539 = pi15 ? n3531 : n3538;
  assign n3540 = pi16 ? n1594 : ~n2301;
  assign n3541 = pi16 ? n1577 : ~n2875;
  assign n3542 = pi15 ? n3540 : n3541;
  assign n3543 = pi14 ? n3539 : n3542;
  assign n3544 = pi16 ? n1577 : ~n3475;
  assign n3545 = pi16 ? n1577 : ~n2294;
  assign n3546 = pi15 ? n3544 : n3545;
  assign n3547 = pi14 ? n3541 : n3546;
  assign n3548 = pi13 ? n3543 : n3547;
  assign n3549 = pi12 ? n3536 : n3548;
  assign n3550 = pi11 ? n3517 : n3549;
  assign n3551 = pi10 ? n3486 : n3550;
  assign n3552 = pi09 ? n3435 : n3551;
  assign n3553 = pi18 ? n2318 : ~n32;
  assign n3554 = pi17 ? n3553 : ~n1718;
  assign n3555 = pi16 ? n32 : n3554;
  assign n3556 = pi15 ? n32 : n3555;
  assign n3557 = pi18 ? n1676 : ~n32;
  assign n3558 = pi18 ? n3325 : ~n32;
  assign n3559 = pi17 ? n3557 : ~n3558;
  assign n3560 = pi16 ? n32 : n3559;
  assign n3561 = pi15 ? n3427 : n3560;
  assign n3562 = pi14 ? n3556 : n3561;
  assign n3563 = pi13 ? n32 : n3562;
  assign n3564 = pi12 ? n32 : n3563;
  assign n3565 = pi11 ? n32 : n3564;
  assign n3566 = pi10 ? n32 : n3565;
  assign n3567 = pi17 ? n32 : n1339;
  assign n3568 = pi16 ? n32 : ~n3567;
  assign n3569 = pi18 ? n32 : n1575;
  assign n3570 = pi17 ? n32 : n3569;
  assign n3571 = pi18 ? n793 : ~n32;
  assign n3572 = pi17 ? n32 : n3571;
  assign n3573 = pi16 ? n3570 : ~n3572;
  assign n3574 = pi15 ? n3568 : n3573;
  assign n3575 = pi20 ? n1368 : ~n448;
  assign n3576 = pi19 ? n3575 : ~n32;
  assign n3577 = pi18 ? n3576 : ~n32;
  assign n3578 = pi17 ? n32 : n3577;
  assign n3579 = pi16 ? n3156 : ~n3578;
  assign n3580 = pi18 ? n2662 : n32;
  assign n3581 = pi17 ? n32 : ~n3580;
  assign n3582 = pi16 ? n3047 : ~n3581;
  assign n3583 = pi15 ? n3579 : n3582;
  assign n3584 = pi14 ? n3574 : n3583;
  assign n3585 = pi17 ? n32 : n2005;
  assign n3586 = pi16 ? n3293 : ~n3585;
  assign n3587 = pi18 ? n32 : n1970;
  assign n3588 = pi17 ? n32 : n3587;
  assign n3589 = pi16 ? n3588 : ~n3162;
  assign n3590 = pi15 ? n3586 : n3589;
  assign n3591 = pi16 ? n2953 : ~n3448;
  assign n3592 = pi15 ? n3174 : n3591;
  assign n3593 = pi14 ? n3590 : n3592;
  assign n3594 = pi13 ? n3584 : n3593;
  assign n3595 = pi16 ? n3176 : ~n3062;
  assign n3596 = pi16 ? n2837 : ~n3297;
  assign n3597 = pi15 ? n3595 : n3596;
  assign n3598 = pi14 ? n3597 : n3307;
  assign n3599 = pi16 ? n2624 : ~n2737;
  assign n3600 = pi15 ? n3069 : n3599;
  assign n3601 = pi16 ? n2860 : ~n2853;
  assign n3602 = pi17 ? n2724 : ~n32;
  assign n3603 = pi16 ? n2513 : ~n3602;
  assign n3604 = pi15 ? n3601 : n3603;
  assign n3605 = pi14 ? n3600 : n3604;
  assign n3606 = pi13 ? n3598 : n3605;
  assign n3607 = pi12 ? n3594 : n3606;
  assign n3608 = pi16 ? n2749 : ~n3194;
  assign n3609 = pi15 ? n3608 : n3079;
  assign n3610 = pi16 ? n2518 : ~n3071;
  assign n3611 = pi15 ? n2976 : n3610;
  assign n3612 = pi14 ? n3609 : n3611;
  assign n3613 = pi16 ? n2293 : ~n2857;
  assign n3614 = pi16 ? n2293 : ~n2737;
  assign n3615 = pi15 ? n3613 : n3614;
  assign n3616 = pi16 ? n2293 : ~n2862;
  assign n3617 = pi15 ? n3616 : n2759;
  assign n3618 = pi14 ? n3615 : n3617;
  assign n3619 = pi13 ? n3612 : n3618;
  assign n3620 = pi16 ? n2415 : ~n2641;
  assign n3621 = pi18 ? n32 : n976;
  assign n3622 = pi17 ? n3621 : ~n32;
  assign n3623 = pi16 ? n2415 : ~n3622;
  assign n3624 = pi15 ? n3620 : n3623;
  assign n3625 = pi17 ? n32 : n2531;
  assign n3626 = pi16 ? n3625 : ~n2514;
  assign n3627 = pi16 ? n2300 : ~n2638;
  assign n3628 = pi15 ? n3626 : n3627;
  assign n3629 = pi14 ? n3624 : n3628;
  assign n3630 = pi16 ? n2300 : ~n2294;
  assign n3631 = pi16 ? n1934 : ~n2875;
  assign n3632 = pi15 ? n3630 : n3631;
  assign n3633 = pi14 ? n3630 : n3632;
  assign n3634 = pi13 ? n3629 : n3633;
  assign n3635 = pi12 ? n3619 : n3634;
  assign n3636 = pi11 ? n3607 : n3635;
  assign n3637 = pi16 ? n1934 : ~n3475;
  assign n3638 = pi16 ? n2320 : ~n2532;
  assign n3639 = pi15 ? n2985 : n3638;
  assign n3640 = pi14 ? n3637 : n3639;
  assign n3641 = pi16 ? n1815 : ~n2875;
  assign n3642 = pi15 ? n3218 : n3641;
  assign n3643 = pi15 ? n3641 : n3218;
  assign n3644 = pi14 ? n3642 : n3643;
  assign n3645 = pi13 ? n3640 : n3644;
  assign n3646 = pi16 ? n1944 : ~n2411;
  assign n3647 = pi15 ? n3646 : n3490;
  assign n3648 = pi16 ? n1944 : ~n3334;
  assign n3649 = pi14 ? n3647 : n3648;
  assign n3650 = pi16 ? n2326 : ~n2411;
  assign n3651 = pi15 ? n3224 : n3650;
  assign n3652 = pi17 ? n1933 : ~n1632;
  assign n3653 = pi16 ? n1678 : ~n3652;
  assign n3654 = pi15 ? n3653 : n3224;
  assign n3655 = pi14 ? n3651 : n3654;
  assign n3656 = pi13 ? n3649 : n3655;
  assign n3657 = pi12 ? n3645 : n3656;
  assign n3658 = pi16 ? n1683 : ~n2301;
  assign n3659 = pi16 ? n1577 : ~n2301;
  assign n3660 = pi15 ? n3658 : n3659;
  assign n3661 = pi14 ? n3660 : n3659;
  assign n3662 = pi16 ? n1683 : ~n2532;
  assign n3663 = pi16 ? n3352 : ~n2532;
  assign n3664 = pi17 ? n2531 : ~n1107;
  assign n3665 = pi16 ? n3352 : ~n3664;
  assign n3666 = pi15 ? n3663 : n3665;
  assign n3667 = pi14 ? n3662 : n3666;
  assign n3668 = pi13 ? n3661 : n3667;
  assign n3669 = pi16 ? n3352 : ~n2645;
  assign n3670 = pi15 ? n3663 : n3669;
  assign n3671 = pi16 ? n3356 : ~n3334;
  assign n3672 = pi17 ? n2119 : ~n1787;
  assign n3673 = pi16 ? n2326 : ~n3672;
  assign n3674 = pi15 ? n3671 : n3673;
  assign n3675 = pi14 ? n3670 : n3674;
  assign n3676 = pi16 ? n2326 : ~n2294;
  assign n3677 = pi16 ? n1815 : ~n2294;
  assign n3678 = pi15 ? n3676 : n3677;
  assign n3679 = pi16 ? n2137 : ~n2520;
  assign n3680 = pi16 ? n2137 : ~n2869;
  assign n3681 = pi15 ? n3679 : n3680;
  assign n3682 = pi14 ? n3678 : n3681;
  assign n3683 = pi13 ? n3675 : n3682;
  assign n3684 = pi12 ? n3668 : n3683;
  assign n3685 = pi11 ? n3657 : n3684;
  assign n3686 = pi10 ? n3636 : n3685;
  assign n3687 = pi09 ? n3566 : n3686;
  assign n3688 = pi08 ? n3552 : n3687;
  assign n3689 = pi07 ? n3422 : n3688;
  assign n3690 = pi06 ? n3154 : n3689;
  assign n3691 = pi05 ? n2723 : n3690;
  assign n3692 = pi20 ? n220 : n32;
  assign n3693 = pi19 ? n975 : n3692;
  assign n3694 = pi18 ? n532 : ~n3693;
  assign n3695 = pi21 ? n309 : ~n405;
  assign n3696 = pi20 ? n3695 : ~n820;
  assign n3697 = pi19 ? n3696 : n32;
  assign n3698 = pi18 ? n3697 : n32;
  assign n3699 = pi17 ? n3694 : n3698;
  assign n3700 = pi16 ? n32 : n3699;
  assign n3701 = pi15 ? n32 : n3700;
  assign n3702 = pi17 ? n1726 : ~n1718;
  assign n3703 = pi16 ? n32 : n3702;
  assign n3704 = pi18 ? n1813 : ~n32;
  assign n3705 = pi17 ? n3704 : ~n1480;
  assign n3706 = pi16 ? n32 : n3705;
  assign n3707 = pi15 ? n3703 : n3706;
  assign n3708 = pi14 ? n3701 : n3707;
  assign n3709 = pi13 ? n32 : n3708;
  assign n3710 = pi12 ? n32 : n3709;
  assign n3711 = pi11 ? n32 : n3710;
  assign n3712 = pi10 ? n32 : n3711;
  assign n3713 = pi17 ? n2005 : ~n1472;
  assign n3714 = pi16 ? n32 : n3713;
  assign n3715 = pi18 ? n1942 : ~n32;
  assign n3716 = pi17 ? n3715 : ~n1700;
  assign n3717 = pi16 ? n32 : n3716;
  assign n3718 = pi15 ? n3714 : n3717;
  assign n3719 = pi18 ? n3350 : ~n32;
  assign n3720 = pi17 ? n3719 : ~n1480;
  assign n3721 = pi16 ? n32 : n3720;
  assign n3722 = pi17 ? n32 : n2345;
  assign n3723 = pi16 ? n3156 : ~n3722;
  assign n3724 = pi15 ? n3721 : n3723;
  assign n3725 = pi14 ? n3718 : n3724;
  assign n3726 = pi17 ? n32 : n1215;
  assign n3727 = pi16 ? n3438 : ~n3726;
  assign n3728 = pi18 ? n32 : n1321;
  assign n3729 = pi17 ? n32 : n3728;
  assign n3730 = pi17 ? n32 : n2685;
  assign n3731 = pi16 ? n3729 : ~n3730;
  assign n3732 = pi15 ? n3727 : n3731;
  assign n3733 = pi16 ? n3165 : ~n3726;
  assign n3734 = pi17 ? n32 : n2465;
  assign n3735 = pi16 ? n3047 : ~n3734;
  assign n3736 = pi15 ? n3733 : n3735;
  assign n3737 = pi14 ? n3732 : n3736;
  assign n3738 = pi13 ? n3725 : n3737;
  assign n3739 = pi16 ? n3176 : ~n3436;
  assign n3740 = pi17 ? n32 : n1997;
  assign n3741 = pi16 ? n2958 : ~n3740;
  assign n3742 = pi15 ? n3739 : n3741;
  assign n3743 = pi15 ? n3446 : n3453;
  assign n3744 = pi14 ? n3742 : n3743;
  assign n3745 = pi16 ? n2745 : ~n3166;
  assign n3746 = pi15 ? n3453 : n3745;
  assign n3747 = pi15 ? n3745 : n3190;
  assign n3748 = pi14 ? n3746 : n3747;
  assign n3749 = pi13 ? n3744 : n3748;
  assign n3750 = pi12 ? n3738 : n3749;
  assign n3751 = pi18 ? n32 : n2233;
  assign n3752 = pi17 ? n3751 : ~n32;
  assign n3753 = pi16 ? n2856 : ~n3752;
  assign n3754 = pi15 ? n2975 : n3753;
  assign n3755 = pi17 ? n3182 : ~n32;
  assign n3756 = pi16 ? n2624 : ~n3755;
  assign n3757 = pi16 ? n2629 : ~n2960;
  assign n3758 = pi15 ? n3756 : n3757;
  assign n3759 = pi14 ? n3754 : n3758;
  assign n3760 = pi16 ? n2513 : ~n3166;
  assign n3761 = pi16 ? n2513 : ~n2955;
  assign n3762 = pi15 ? n3760 : n3761;
  assign n3763 = pi18 ? n32 : n767;
  assign n3764 = pi17 ? n3763 : ~n32;
  assign n3765 = pi16 ? n2749 : ~n3764;
  assign n3766 = pi15 ? n3608 : n3765;
  assign n3767 = pi14 ? n3762 : n3766;
  assign n3768 = pi13 ? n3759 : n3767;
  assign n3769 = pi17 ? n32 : n2519;
  assign n3770 = pi16 ? n3769 : ~n2734;
  assign n3771 = pi16 ? n3769 : ~n3194;
  assign n3772 = pi16 ? n2293 : ~n3194;
  assign n3773 = pi15 ? n3771 : n3772;
  assign n3774 = pi14 ? n3770 : n3773;
  assign n3775 = pi20 ? n1331 : ~n32;
  assign n3776 = pi19 ? n32 : n3775;
  assign n3777 = pi18 ? n32 : n3776;
  assign n3778 = pi17 ? n3777 : ~n32;
  assign n3779 = pi16 ? n2293 : ~n3778;
  assign n3780 = pi19 ? n32 : n3507;
  assign n3781 = pi18 ? n32 : n3780;
  assign n3782 = pi17 ? n3781 : ~n32;
  assign n3783 = pi16 ? n2293 : ~n3782;
  assign n3784 = pi15 ? n3779 : n3783;
  assign n3785 = pi16 ? n2654 : ~n2737;
  assign n3786 = pi19 ? n365 : ~n32;
  assign n3787 = pi18 ? n32 : n3786;
  assign n3788 = pi17 ? n32 : n3787;
  assign n3789 = pi16 ? n3788 : ~n2737;
  assign n3790 = pi15 ? n3785 : n3789;
  assign n3791 = pi14 ? n3784 : n3790;
  assign n3792 = pi13 ? n3774 : n3791;
  assign n3793 = pi12 ? n3768 : n3792;
  assign n3794 = pi11 ? n3750 : n3793;
  assign n3795 = pi16 ? n3788 : ~n3202;
  assign n3796 = pi15 ? n3789 : n3795;
  assign n3797 = pi19 ? n594 : n821;
  assign n3798 = pi18 ? n32 : n3797;
  assign n3799 = pi17 ? n3798 : ~n32;
  assign n3800 = pi16 ? n3788 : ~n3799;
  assign n3801 = pi16 ? n2530 : ~n2619;
  assign n3802 = pi15 ? n3800 : n3801;
  assign n3803 = pi14 ? n3796 : n3802;
  assign n3804 = pi16 ? n2530 : ~n2751;
  assign n3805 = pi15 ? n3470 : n3804;
  assign n3806 = pi15 ? n3804 : n3470;
  assign n3807 = pi14 ? n3805 : n3806;
  assign n3808 = pi13 ? n3803 : n3807;
  assign n3809 = pi16 ? n2540 : ~n2514;
  assign n3810 = pi16 ? n2540 : ~n2751;
  assign n3811 = pi15 ? n3809 : n3810;
  assign n3812 = pi18 ? n32 : n776;
  assign n3813 = pi17 ? n3812 : ~n32;
  assign n3814 = pi16 ? n2540 : ~n3813;
  assign n3815 = pi15 ? n3814 : n3809;
  assign n3816 = pi14 ? n3811 : n3815;
  assign n3817 = pi16 ? n1808 : ~n2520;
  assign n3818 = pi16 ? n1808 : ~n2625;
  assign n3819 = pi15 ? n3817 : n3818;
  assign n3820 = pi14 ? n3819 : n3817;
  assign n3821 = pi13 ? n3816 : n3820;
  assign n3822 = pi12 ? n3808 : n3821;
  assign n3823 = pi16 ? n2326 : ~n2520;
  assign n3824 = pi16 ? n2326 : ~n2514;
  assign n3825 = pi14 ? n3823 : n3824;
  assign n3826 = pi16 ? n1815 : ~n2514;
  assign n3827 = pi16 ? n1808 : ~n2751;
  assign n3828 = pi14 ? n3826 : n3827;
  assign n3829 = pi13 ? n3825 : n3828;
  assign n3830 = pi16 ? n1815 : ~n3202;
  assign n3831 = pi16 ? n2320 : ~n2737;
  assign n3832 = pi15 ? n3830 : n3831;
  assign n3833 = pi14 ? n3827 : n3832;
  assign n3834 = pi16 ? n1934 : ~n2737;
  assign n3835 = pi15 ? n3831 : n3834;
  assign n3836 = pi16 ? n2320 : ~n3194;
  assign n3837 = pi14 ? n3835 : n3836;
  assign n3838 = pi13 ? n3833 : n3837;
  assign n3839 = pi12 ? n3829 : n3838;
  assign n3840 = pi11 ? n3822 : n3839;
  assign n3841 = pi10 ? n3794 : n3840;
  assign n3842 = pi09 ? n3712 : n3841;
  assign n3843 = pi21 ? n405 : n309;
  assign n3844 = pi20 ? n3843 : n32;
  assign n3845 = pi19 ? n32 : n3844;
  assign n3846 = pi18 ? n2298 : ~n3845;
  assign n3847 = pi21 ? n405 : n173;
  assign n3848 = pi20 ? n274 : n3847;
  assign n3849 = pi20 ? n173 : n339;
  assign n3850 = pi19 ? n3848 : n3849;
  assign n3851 = pi18 ? n3850 : ~n32;
  assign n3852 = pi17 ? n3846 : ~n3851;
  assign n3853 = pi16 ? n32 : n3852;
  assign n3854 = pi15 ? n32 : n3853;
  assign n3855 = pi18 ? n2304 : ~n32;
  assign n3856 = pi20 ? n173 : n820;
  assign n3857 = pi19 ? n594 : n3856;
  assign n3858 = pi18 ? n3857 : ~n32;
  assign n3859 = pi17 ? n3855 : ~n3858;
  assign n3860 = pi16 ? n32 : n3859;
  assign n3861 = pi20 ? n173 : n357;
  assign n3862 = pi19 ? n32 : ~n3861;
  assign n3863 = pi18 ? n3862 : ~n32;
  assign n3864 = pi17 ? n1227 : ~n3863;
  assign n3865 = pi16 ? n32 : n3864;
  assign n3866 = pi15 ? n3860 : n3865;
  assign n3867 = pi14 ? n3854 : n3866;
  assign n3868 = pi13 ? n32 : n3867;
  assign n3869 = pi12 ? n32 : n3868;
  assign n3870 = pi11 ? n32 : n3869;
  assign n3871 = pi10 ? n32 : n3870;
  assign n3872 = pi17 ? n3553 : ~n1472;
  assign n3873 = pi16 ? n32 : n3872;
  assign n3874 = pi17 ? n1726 : ~n1700;
  assign n3875 = pi16 ? n32 : n3874;
  assign n3876 = pi15 ? n3873 : n3875;
  assign n3877 = pi17 ? n3719 : ~n2567;
  assign n3878 = pi16 ? n32 : n3877;
  assign n3879 = pi17 ? n32 : n1582;
  assign n3880 = pi16 ? n32 : ~n3879;
  assign n3881 = pi15 ? n3878 : n3880;
  assign n3882 = pi14 ? n3876 : n3881;
  assign n3883 = pi19 ? n975 : n821;
  assign n3884 = pi18 ? n3883 : ~n32;
  assign n3885 = pi17 ? n32 : n3884;
  assign n3886 = pi16 ? n3570 : ~n3885;
  assign n3887 = pi17 ? n32 : n2926;
  assign n3888 = pi16 ? n3283 : ~n3887;
  assign n3889 = pi15 ? n3886 : n3888;
  assign n3890 = pi19 ? n1369 : ~n32;
  assign n3891 = pi18 ? n3890 : ~n32;
  assign n3892 = pi17 ? n32 : n3891;
  assign n3893 = pi16 ? n3156 : ~n3892;
  assign n3894 = pi15 ? n3893 : n3735;
  assign n3895 = pi14 ? n3889 : n3894;
  assign n3896 = pi13 ? n3882 : n3895;
  assign n3897 = pi21 ? n173 : n259;
  assign n3898 = pi20 ? n32 : n3897;
  assign n3899 = pi19 ? n3898 : ~n32;
  assign n3900 = pi18 ? n3899 : ~n32;
  assign n3901 = pi17 ? n32 : n3900;
  assign n3902 = pi16 ? n3293 : ~n3901;
  assign n3903 = pi16 ? n3588 : ~n3740;
  assign n3904 = pi15 ? n3902 : n3903;
  assign n3905 = pi19 ? n3861 : n32;
  assign n3906 = pi18 ? n3905 : n32;
  assign n3907 = pi17 ? n32 : ~n3906;
  assign n3908 = pi16 ? n2953 : ~n3907;
  assign n3909 = pi16 ? n2953 : ~n3062;
  assign n3910 = pi15 ? n3908 : n3909;
  assign n3911 = pi14 ? n3904 : n3910;
  assign n3912 = pi20 ? n32 : n173;
  assign n3913 = pi19 ? n32 : n3912;
  assign n3914 = pi18 ? n32 : n3913;
  assign n3915 = pi20 ? n3897 : ~n32;
  assign n3916 = pi19 ? n3915 : ~n32;
  assign n3917 = pi18 ? n3916 : ~n32;
  assign n3918 = pi17 ? n3914 : n3917;
  assign n3919 = pi16 ? n3176 : ~n3918;
  assign n3920 = pi16 ? n2837 : ~n3581;
  assign n3921 = pi15 ? n3919 : n3920;
  assign n3922 = pi16 ? n2840 : ~n3166;
  assign n3923 = pi20 ? n428 : n173;
  assign n3924 = pi19 ? n32 : n3923;
  assign n3925 = pi18 ? n32 : n3924;
  assign n3926 = pi17 ? n3925 : n2008;
  assign n3927 = pi16 ? n2851 : ~n3926;
  assign n3928 = pi15 ? n3922 : n3927;
  assign n3929 = pi14 ? n3921 : n3928;
  assign n3930 = pi13 ? n3911 : n3929;
  assign n3931 = pi12 ? n3896 : n3930;
  assign n3932 = pi16 ? n3068 : ~n3926;
  assign n3933 = pi20 ? n32 : ~n173;
  assign n3934 = pi19 ? n32 : n3933;
  assign n3935 = pi18 ? n32 : n3934;
  assign n3936 = pi17 ? n3935 : ~n32;
  assign n3937 = pi16 ? n2732 : ~n3936;
  assign n3938 = pi15 ? n3932 : n3937;
  assign n3939 = pi16 ? n2732 : ~n2960;
  assign n3940 = pi15 ? n3937 : n3939;
  assign n3941 = pi14 ? n3938 : n3940;
  assign n3942 = pi16 ? n2617 : ~n2955;
  assign n3943 = pi15 ? n3745 : n3942;
  assign n3944 = pi17 ? n2839 : ~n32;
  assign n3945 = pi16 ? n2856 : ~n3944;
  assign n3946 = pi17 ? n32 : n2618;
  assign n3947 = pi16 ? n3946 : ~n2734;
  assign n3948 = pi15 ? n3945 : n3947;
  assign n3949 = pi14 ? n3943 : n3948;
  assign n3950 = pi13 ? n3941 : n3949;
  assign n3951 = pi16 ? n2629 : ~n2734;
  assign n3952 = pi16 ? n2513 : ~n3194;
  assign n3953 = pi14 ? n3951 : n3952;
  assign n3954 = pi16 ? n2518 : ~n2727;
  assign n3955 = pi16 ? n2518 : ~n2734;
  assign n3956 = pi15 ? n3954 : n3955;
  assign n3957 = pi15 ? n3456 : n3197;
  assign n3958 = pi14 ? n3956 : n3957;
  assign n3959 = pi13 ? n3953 : n3958;
  assign n3960 = pi12 ? n3950 : n3959;
  assign n3961 = pi11 ? n3931 : n3960;
  assign n3962 = pi19 ? n594 : n813;
  assign n3963 = pi18 ? n32 : n3962;
  assign n3964 = pi17 ? n3963 : ~n32;
  assign n3965 = pi16 ? n2756 : ~n3964;
  assign n3966 = pi15 ? n3197 : n3965;
  assign n3967 = pi18 ? n32 : n967;
  assign n3968 = pi17 ? n3967 : ~n32;
  assign n3969 = pi16 ? n2120 : ~n3968;
  assign n3970 = pi18 ? n32 : n2251;
  assign n3971 = pi17 ? n3970 : ~n32;
  assign n3972 = pi16 ? n2426 : ~n3971;
  assign n3973 = pi15 ? n3969 : n3972;
  assign n3974 = pi14 ? n3966 : n3973;
  assign n3975 = pi19 ? n857 : ~n358;
  assign n3976 = pi18 ? n32 : n3975;
  assign n3977 = pi17 ? n3976 : ~n32;
  assign n3978 = pi16 ? n2426 : ~n3977;
  assign n3979 = pi16 ? n2426 : ~n2751;
  assign n3980 = pi15 ? n3978 : n3979;
  assign n3981 = pi16 ? n3788 : ~n2619;
  assign n3982 = pi15 ? n3979 : n3981;
  assign n3983 = pi14 ? n3980 : n3982;
  assign n3984 = pi13 ? n3974 : n3983;
  assign n3985 = pi16 ? n3788 : ~n2857;
  assign n3986 = pi15 ? n3981 : n3985;
  assign n3987 = pi16 ? n3788 : ~n2514;
  assign n3988 = pi15 ? n3985 : n3987;
  assign n3989 = pi14 ? n3986 : n3988;
  assign n3990 = pi16 ? n2306 : ~n2638;
  assign n3991 = pi16 ? n2306 : ~n2862;
  assign n3992 = pi15 ? n3990 : n3991;
  assign n3993 = pi16 ? n2306 : ~n2625;
  assign n3994 = pi14 ? n3992 : n3993;
  assign n3995 = pi13 ? n3989 : n3994;
  assign n3996 = pi12 ? n3984 : n3995;
  assign n3997 = pi16 ? n2320 : ~n2625;
  assign n3998 = pi16 ? n2320 : ~n2619;
  assign n3999 = pi14 ? n3997 : n3998;
  assign n4000 = pi16 ? n1934 : ~n2619;
  assign n4001 = pi16 ? n2300 : ~n2857;
  assign n4002 = pi14 ? n4000 : n4001;
  assign n4003 = pi13 ? n3999 : n4002;
  assign n4004 = pi16 ? n2530 : ~n2737;
  assign n4005 = pi16 ? n3625 : ~n3602;
  assign n4006 = pi15 ? n4004 : n4005;
  assign n4007 = pi14 ? n4001 : n4006;
  assign n4008 = pi16 ? n2426 : ~n3602;
  assign n4009 = pi15 ? n4005 : n4008;
  assign n4010 = pi16 ? n3625 : ~n3944;
  assign n4011 = pi16 ? n2654 : ~n3752;
  assign n4012 = pi15 ? n4010 : n4011;
  assign n4013 = pi14 ? n4009 : n4012;
  assign n4014 = pi13 ? n4007 : n4013;
  assign n4015 = pi12 ? n4003 : n4014;
  assign n4016 = pi11 ? n3996 : n4015;
  assign n4017 = pi10 ? n3961 : n4016;
  assign n4018 = pi09 ? n3871 : n4017;
  assign n4019 = pi08 ? n3842 : n4018;
  assign n4020 = pi17 ? n2355 : ~n1580;
  assign n4021 = pi16 ? n32 : n4020;
  assign n4022 = pi15 ? n32 : n4021;
  assign n4023 = pi18 ? n2424 : ~n32;
  assign n4024 = pi17 ? n4023 : ~n2136;
  assign n4025 = pi16 ? n32 : n4024;
  assign n4026 = pi17 ? n1120 : ~n2325;
  assign n4027 = pi16 ? n32 : n4026;
  assign n4028 = pi15 ? n4025 : n4027;
  assign n4029 = pi14 ? n4022 : n4028;
  assign n4030 = pi13 ? n32 : n4029;
  assign n4031 = pi12 ? n32 : n4030;
  assign n4032 = pi11 ? n32 : n4031;
  assign n4033 = pi10 ? n32 : n4032;
  assign n4034 = pi18 ? n3786 : ~n32;
  assign n4035 = pi17 ? n4034 : ~n1470;
  assign n4036 = pi16 ? n32 : n4035;
  assign n4037 = pi18 ? n2298 : ~n32;
  assign n4038 = pi17 ? n4037 : ~n1580;
  assign n4039 = pi16 ? n32 : n4038;
  assign n4040 = pi15 ? n4036 : n4039;
  assign n4041 = pi18 ? n3336 : ~n32;
  assign n4042 = pi17 ? n4041 : ~n1213;
  assign n4043 = pi16 ? n32 : n4042;
  assign n4044 = pi17 ? n2005 : ~n1470;
  assign n4045 = pi16 ? n32 : n4044;
  assign n4046 = pi15 ? n4043 : n4045;
  assign n4047 = pi14 ? n4040 : n4046;
  assign n4048 = pi17 ? n3715 : ~n1470;
  assign n4049 = pi16 ? n32 : n4048;
  assign n4050 = pi17 ? n1028 : ~n1978;
  assign n4051 = pi16 ? n32 : n4050;
  assign n4052 = pi15 ? n4049 : n4051;
  assign n4053 = pi17 ? n3719 : ~n1697;
  assign n4054 = pi16 ? n32 : n4053;
  assign n4055 = pi17 ? n32 : n1472;
  assign n4056 = pi16 ? n3156 : ~n4055;
  assign n4057 = pi15 ? n4054 : n4056;
  assign n4058 = pi14 ? n4052 : n4057;
  assign n4059 = pi13 ? n4047 : n4058;
  assign n4060 = pi17 ? n32 : n1978;
  assign n4061 = pi16 ? n3438 : ~n4060;
  assign n4062 = pi16 ? n3729 : ~n4060;
  assign n4063 = pi15 ? n4061 : n4062;
  assign n4064 = pi17 ? n32 : n1480;
  assign n4065 = pi16 ? n3165 : ~n4064;
  assign n4066 = pi17 ? n32 : n1718;
  assign n4067 = pi16 ? n3047 : ~n4066;
  assign n4068 = pi15 ? n4065 : n4067;
  assign n4069 = pi14 ? n4063 : n4068;
  assign n4070 = pi16 ? n3176 : ~n3726;
  assign n4071 = pi16 ? n2958 : ~n4066;
  assign n4072 = pi15 ? n4070 : n4071;
  assign n4073 = pi16 ? n2964 : ~n3726;
  assign n4074 = pi16 ? n3183 : ~n3428;
  assign n4075 = pi15 ? n4073 : n4074;
  assign n4076 = pi14 ? n4072 : n4075;
  assign n4077 = pi13 ? n4069 : n4076;
  assign n4078 = pi12 ? n4059 : n4077;
  assign n4079 = pi16 ? n3183 : ~n3436;
  assign n4080 = pi16 ? n3061 : ~n3428;
  assign n4081 = pi15 ? n4079 : n4080;
  assign n4082 = pi16 ? n3061 : ~n3726;
  assign n4083 = pi16 ? n2837 : ~n3726;
  assign n4084 = pi15 ? n4082 : n4083;
  assign n4085 = pi14 ? n4081 : n4084;
  assign n4086 = pi16 ? n2840 : ~n3436;
  assign n4087 = pi16 ? n2851 : ~n3157;
  assign n4088 = pi15 ? n4086 : n4087;
  assign n4089 = pi16 ? n2725 : ~n3162;
  assign n4090 = pi16 ? n2725 : ~n3157;
  assign n4091 = pi15 ? n4089 : n4090;
  assign n4092 = pi14 ? n4088 : n4091;
  assign n4093 = pi13 ? n4085 : n4092;
  assign n4094 = pi16 ? n2732 : ~n3157;
  assign n4095 = pi16 ? n2745 : ~n3162;
  assign n4096 = pi15 ? n4094 : n4095;
  assign n4097 = pi16 ? n2617 : ~n3162;
  assign n4098 = pi19 ? n1574 : ~n32;
  assign n4099 = pi18 ? n32 : n4098;
  assign n4100 = pi17 ? n32 : n4099;
  assign n4101 = pi16 ? n4100 : ~n3177;
  assign n4102 = pi15 ? n4097 : n4101;
  assign n4103 = pi14 ? n4096 : n4102;
  assign n4104 = pi16 ? n3946 : ~n3166;
  assign n4105 = pi16 ? n3946 : ~n3180;
  assign n4106 = pi15 ? n4104 : n4105;
  assign n4107 = pi14 ? n4101 : n4106;
  assign n4108 = pi13 ? n4103 : n4107;
  assign n4109 = pi12 ? n4093 : n4108;
  assign n4110 = pi11 ? n4078 : n4109;
  assign n4111 = pi18 ? n32 : n1592;
  assign n4112 = pi17 ? n4111 : ~n32;
  assign n4113 = pi16 ? n2513 : ~n4112;
  assign n4114 = pi15 ? n4113 : n3760;
  assign n4115 = pi16 ? n2749 : ~n3180;
  assign n4116 = pi15 ? n3760 : n4115;
  assign n4117 = pi14 ? n4114 : n4116;
  assign n4118 = pi18 ? n32 : n2202;
  assign n4119 = pi17 ? n4118 : ~n32;
  assign n4120 = pi16 ? n2749 : ~n4119;
  assign n4121 = pi16 ? n2749 : ~n2960;
  assign n4122 = pi15 ? n4120 : n4121;
  assign n4123 = pi16 ? n2409 : ~n2960;
  assign n4124 = pi14 ? n4122 : n4123;
  assign n4125 = pi13 ? n4117 : n4124;
  assign n4126 = pi20 ? n32 : n206;
  assign n4127 = pi19 ? n32 : n4126;
  assign n4128 = pi18 ? n32 : n4127;
  assign n4129 = pi17 ? n4128 : ~n32;
  assign n4130 = pi16 ? n2409 : ~n4129;
  assign n4131 = pi16 ? n2409 : ~n4112;
  assign n4132 = pi15 ? n4130 : n4131;
  assign n4133 = pi16 ? n2409 : ~n2727;
  assign n4134 = pi16 ? n2120 : ~n2727;
  assign n4135 = pi15 ? n4133 : n4134;
  assign n4136 = pi14 ? n4132 : n4135;
  assign n4137 = pi16 ? n2120 : ~n2734;
  assign n4138 = pi15 ? n4134 : n4137;
  assign n4139 = pi14 ? n4138 : n4137;
  assign n4140 = pi13 ? n4136 : n4139;
  assign n4141 = pi12 ? n4125 : n4140;
  assign n4142 = pi16 ? n3625 : ~n2734;
  assign n4143 = pi16 ? n3625 : ~n2727;
  assign n4144 = pi15 ? n4142 : n4143;
  assign n4145 = pi14 ? n4144 : n4143;
  assign n4146 = pi16 ? n2426 : ~n2727;
  assign n4147 = pi16 ? n2120 : ~n2960;
  assign n4148 = pi16 ? n2426 : ~n2960;
  assign n4149 = pi15 ? n4147 : n4148;
  assign n4150 = pi14 ? n4146 : n4149;
  assign n4151 = pi13 ? n4145 : n4150;
  assign n4152 = pi16 ? n2293 : ~n3180;
  assign n4153 = pi15 ? n4148 : n4152;
  assign n4154 = pi14 ? n4147 : n4153;
  assign n4155 = pi16 ? n3769 : ~n3180;
  assign n4156 = pi15 ? n4152 : n4155;
  assign n4157 = pi16 ? n2293 : ~n2955;
  assign n4158 = pi14 ? n4156 : n4157;
  assign n4159 = pi13 ? n4154 : n4158;
  assign n4160 = pi12 ? n4151 : n4159;
  assign n4161 = pi11 ? n4141 : n4160;
  assign n4162 = pi10 ? n4110 : n4161;
  assign n4163 = pi09 ? n4033 : n4162;
  assign n4164 = pi17 ? n2461 : ~n2885;
  assign n4165 = pi16 ? n32 : n4164;
  assign n4166 = pi15 ? n32 : n4165;
  assign n4167 = pi18 ? n2754 : ~n32;
  assign n4168 = pi17 ? n4167 : ~n2136;
  assign n4169 = pi16 ? n32 : n4168;
  assign n4170 = pi17 ? n1215 : ~n2136;
  assign n4171 = pi16 ? n32 : n4170;
  assign n4172 = pi15 ? n4169 : n4171;
  assign n4173 = pi14 ? n4166 : n4172;
  assign n4174 = pi13 ? n32 : n4173;
  assign n4175 = pi12 ? n32 : n4174;
  assign n4176 = pi11 ? n32 : n4175;
  assign n4177 = pi10 ? n32 : n4176;
  assign n4178 = pi17 ? n2355 : ~n1470;
  assign n4179 = pi16 ? n32 : n4178;
  assign n4180 = pi15 ? n4179 : n4039;
  assign n4181 = pi17 ? n1605 : ~n1704;
  assign n4182 = pi16 ? n32 : n4181;
  assign n4183 = pi17 ? n1227 : ~n1470;
  assign n4184 = pi16 ? n32 : n4183;
  assign n4185 = pi15 ? n4182 : n4184;
  assign n4186 = pi14 ? n4180 : n4185;
  assign n4187 = pi17 ? n3553 : ~n1470;
  assign n4188 = pi16 ? n32 : n4187;
  assign n4189 = pi17 ? n1726 : ~n1978;
  assign n4190 = pi16 ? n32 : n4189;
  assign n4191 = pi15 ? n4188 : n4190;
  assign n4192 = pi17 ? n4041 : ~n1134;
  assign n4193 = pi16 ? n32 : n4192;
  assign n4194 = pi17 ? n3719 : ~n1582;
  assign n4195 = pi16 ? n32 : n4194;
  assign n4196 = pi15 ? n4193 : n4195;
  assign n4197 = pi14 ? n4191 : n4196;
  assign n4198 = pi13 ? n4186 : n4197;
  assign n4199 = pi17 ? n32 : n1975;
  assign n4200 = pi16 ? n32 : ~n4199;
  assign n4201 = pi17 ? n32 : n1700;
  assign n4202 = pi16 ? n3570 : ~n4201;
  assign n4203 = pi15 ? n4200 : n4202;
  assign n4204 = pi16 ? n3283 : ~n4064;
  assign n4205 = pi16 ? n3156 : ~n3730;
  assign n4206 = pi15 ? n4204 : n4205;
  assign n4207 = pi14 ? n4203 : n4206;
  assign n4208 = pi16 ? n3047 : ~n3726;
  assign n4209 = pi16 ? n3293 : ~n4066;
  assign n4210 = pi15 ? n4208 : n4209;
  assign n4211 = pi16 ? n3588 : ~n3726;
  assign n4212 = pi16 ? n2953 : ~n3428;
  assign n4213 = pi15 ? n4211 : n4212;
  assign n4214 = pi14 ? n4210 : n4213;
  assign n4215 = pi13 ? n4207 : n4214;
  assign n4216 = pi12 ? n4198 : n4215;
  assign n4217 = pi17 ? n32 : n2604;
  assign n4218 = pi16 ? n2953 : ~n4217;
  assign n4219 = pi16 ? n3176 : ~n3734;
  assign n4220 = pi15 ? n4218 : n4219;
  assign n4221 = pi17 ? n32 : n2461;
  assign n4222 = pi16 ? n3176 : ~n4221;
  assign n4223 = pi16 ? n2958 : ~n4221;
  assign n4224 = pi15 ? n4222 : n4223;
  assign n4225 = pi14 ? n4220 : n4224;
  assign n4226 = pi17 ? n32 : n2165;
  assign n4227 = pi16 ? n2964 : ~n4226;
  assign n4228 = pi16 ? n2964 : ~n3157;
  assign n4229 = pi15 ? n4227 : n4228;
  assign n4230 = pi17 ? n32 : n1726;
  assign n4231 = pi16 ? n2832 : ~n4230;
  assign n4232 = pi17 ? n32 : n1605;
  assign n4233 = pi16 ? n2832 : ~n4232;
  assign n4234 = pi15 ? n4231 : n4233;
  assign n4235 = pi14 ? n4229 : n4234;
  assign n4236 = pi13 ? n4225 : n4235;
  assign n4237 = pi17 ? n32 : n1350;
  assign n4238 = pi16 ? n3061 : ~n4237;
  assign n4239 = pi17 ? n32 : n2473;
  assign n4240 = pi16 ? n2837 : ~n4239;
  assign n4241 = pi15 ? n4238 : n4240;
  assign n4242 = pi17 ? n32 : n2177;
  assign n4243 = pi16 ? n2840 : ~n4242;
  assign n4244 = pi19 ? n32 : n1812;
  assign n4245 = pi18 ? n32 : n4244;
  assign n4246 = pi17 ? n32 : n4245;
  assign n4247 = pi16 ? n4246 : ~n3585;
  assign n4248 = pi15 ? n4243 : n4247;
  assign n4249 = pi14 ? n4241 : n4248;
  assign n4250 = pi16 ? n4246 : ~n3177;
  assign n4251 = pi15 ? n4250 : n4247;
  assign n4252 = pi17 ? n32 : n932;
  assign n4253 = pi16 ? n2725 : ~n4252;
  assign n4254 = pi17 ? n3296 : ~n1124;
  assign n4255 = pi16 ? n2732 : ~n4254;
  assign n4256 = pi15 ? n4253 : n4255;
  assign n4257 = pi14 ? n4251 : n4256;
  assign n4258 = pi13 ? n4249 : n4257;
  assign n4259 = pi12 ? n4236 : n4258;
  assign n4260 = pi11 ? n4216 : n4259;
  assign n4261 = pi18 ? n32 : n858;
  assign n4262 = pi17 ? n4261 : ~n32;
  assign n4263 = pi16 ? n2624 : ~n4262;
  assign n4264 = pi16 ? n2624 : ~n3166;
  assign n4265 = pi15 ? n4263 : n4264;
  assign n4266 = pi17 ? n32 : ~n1124;
  assign n4267 = pi16 ? n2624 : ~n4266;
  assign n4268 = pi18 ? n32 : n2197;
  assign n4269 = pi17 ? n4268 : n2008;
  assign n4270 = pi16 ? n2860 : ~n4269;
  assign n4271 = pi15 ? n4267 : n4270;
  assign n4272 = pi14 ? n4265 : n4271;
  assign n4273 = pi17 ? n3282 : n2008;
  assign n4274 = pi16 ? n2860 : ~n4273;
  assign n4275 = pi16 ? n3946 : ~n4119;
  assign n4276 = pi15 ? n4274 : n4275;
  assign n4277 = pi14 ? n4276 : n4275;
  assign n4278 = pi13 ? n4272 : n4277;
  assign n4279 = pi21 ? n174 : n206;
  assign n4280 = pi20 ? n32 : n4279;
  assign n4281 = pi19 ? n32 : n4280;
  assign n4282 = pi18 ? n32 : n4281;
  assign n4283 = pi17 ? n4282 : ~n32;
  assign n4284 = pi16 ? n3946 : ~n4283;
  assign n4285 = pi16 ? n3946 : ~n4262;
  assign n4286 = pi15 ? n4284 : n4285;
  assign n4287 = pi19 ? n32 : n3898;
  assign n4288 = pi18 ? n32 : n4287;
  assign n4289 = pi17 ? n4288 : ~n32;
  assign n4290 = pi16 ? n3946 : ~n4289;
  assign n4291 = pi16 ? n2756 : ~n4289;
  assign n4292 = pi15 ? n4290 : n4291;
  assign n4293 = pi14 ? n4286 : n4292;
  assign n4294 = pi18 ? n32 : n2043;
  assign n4295 = pi17 ? n4294 : ~n32;
  assign n4296 = pi16 ? n2756 : ~n4295;
  assign n4297 = pi15 ? n4291 : n4296;
  assign n4298 = pi14 ? n4297 : n4296;
  assign n4299 = pi13 ? n4293 : n4298;
  assign n4300 = pi12 ? n4278 : n4299;
  assign n4301 = pi16 ? n2293 : ~n4295;
  assign n4302 = pi18 ? n32 : n2108;
  assign n4303 = pi17 ? n4302 : ~n32;
  assign n4304 = pi16 ? n2293 : ~n4303;
  assign n4305 = pi15 ? n4301 : n4304;
  assign n4306 = pi14 ? n4305 : n4304;
  assign n4307 = pi16 ? n3769 : ~n4303;
  assign n4308 = pi18 ? n32 : n2906;
  assign n4309 = pi17 ? n4308 : ~n32;
  assign n4310 = pi16 ? n3769 : ~n4309;
  assign n4311 = pi15 ? n4307 : n4310;
  assign n4312 = pi16 ? n2749 : ~n3448;
  assign n4313 = pi16 ? n3769 : ~n3448;
  assign n4314 = pi15 ? n4312 : n4313;
  assign n4315 = pi14 ? n4311 : n4314;
  assign n4316 = pi13 ? n4306 : n4315;
  assign n4317 = pi17 ? n3292 : ~n32;
  assign n4318 = pi16 ? n2518 : ~n4317;
  assign n4319 = pi18 ? n32 : n1862;
  assign n4320 = pi17 ? n4319 : ~n32;
  assign n4321 = pi16 ? n2513 : ~n4320;
  assign n4322 = pi15 ? n4318 : n4321;
  assign n4323 = pi14 ? n4312 : n4322;
  assign n4324 = pi16 ? n4100 : ~n4320;
  assign n4325 = pi15 ? n4321 : n4324;
  assign n4326 = pi16 ? n2513 : ~n4262;
  assign n4327 = pi17 ? n4261 : ~n1124;
  assign n4328 = pi16 ? n4100 : ~n4327;
  assign n4329 = pi15 ? n4326 : n4328;
  assign n4330 = pi14 ? n4325 : n4329;
  assign n4331 = pi13 ? n4323 : n4330;
  assign n4332 = pi12 ? n4316 : n4331;
  assign n4333 = pi11 ? n4300 : n4332;
  assign n4334 = pi10 ? n4260 : n4333;
  assign n4335 = pi09 ? n4177 : n4334;
  assign n4336 = pi08 ? n4163 : n4335;
  assign n4337 = pi07 ? n4019 : n4336;
  assign n4338 = pi17 ? n1480 : ~n1682;
  assign n4339 = pi16 ? n32 : n4338;
  assign n4340 = pi15 ? n32 : n4339;
  assign n4341 = pi18 ? n4098 : ~n32;
  assign n4342 = pi20 ? n321 : n32;
  assign n4343 = pi19 ? n4342 : n32;
  assign n4344 = pi18 ? n32 : ~n4343;
  assign n4345 = pi17 ? n4341 : ~n4344;
  assign n4346 = pi16 ? n32 : n4345;
  assign n4347 = pi17 ? n1989 : ~n4344;
  assign n4348 = pi16 ? n32 : n4347;
  assign n4349 = pi15 ? n4346 : n4348;
  assign n4350 = pi14 ? n4340 : n4349;
  assign n4351 = pi13 ? n32 : n4350;
  assign n4352 = pi12 ? n32 : n4351;
  assign n4353 = pi11 ? n32 : n4352;
  assign n4354 = pi10 ? n32 : n4353;
  assign n4355 = pi17 ? n2461 : ~n1682;
  assign n4356 = pi16 ? n32 : n4355;
  assign n4357 = pi17 ? n2355 : ~n1682;
  assign n4358 = pi16 ? n32 : n4357;
  assign n4359 = pi15 ? n4356 : n4358;
  assign n4360 = pi17 ? n4023 : ~n1807;
  assign n4361 = pi16 ? n32 : n4360;
  assign n4362 = pi17 ? n1120 : ~n1807;
  assign n4363 = pi16 ? n32 : n4362;
  assign n4364 = pi15 ? n4361 : n4363;
  assign n4365 = pi14 ? n4359 : n4364;
  assign n4366 = pi17 ? n4034 : ~n2325;
  assign n4367 = pi16 ? n32 : n4366;
  assign n4368 = pi17 ? n1219 : ~n1470;
  assign n4369 = pi16 ? n32 : n4368;
  assign n4370 = pi15 ? n4367 : n4369;
  assign n4371 = pi17 ? n1605 : ~n2123;
  assign n4372 = pi16 ? n32 : n4371;
  assign n4373 = pi17 ? n4041 : ~n1580;
  assign n4374 = pi16 ? n32 : n4373;
  assign n4375 = pi15 ? n4372 : n4374;
  assign n4376 = pi14 ? n4370 : n4375;
  assign n4377 = pi13 ? n4365 : n4376;
  assign n4378 = pi17 ? n2005 : ~n2325;
  assign n4379 = pi16 ? n32 : n4378;
  assign n4380 = pi19 ? n32 : n1464;
  assign n4381 = pi18 ? n4380 : ~n32;
  assign n4382 = pi17 ? n3715 : ~n4381;
  assign n4383 = pi16 ? n32 : n4382;
  assign n4384 = pi15 ? n4379 : n4383;
  assign n4385 = pi17 ? n1028 : ~n1697;
  assign n4386 = pi16 ? n32 : n4385;
  assign n4387 = pi17 ? n3719 : ~n1213;
  assign n4388 = pi16 ? n32 : n4387;
  assign n4389 = pi15 ? n4386 : n4388;
  assign n4390 = pi14 ? n4384 : n4389;
  assign n4391 = pi20 ? n321 : n207;
  assign n4392 = pi19 ? n32 : n4391;
  assign n4393 = pi18 ? n4392 : ~n32;
  assign n4394 = pi17 ? n32 : n4393;
  assign n4395 = pi16 ? n3156 : ~n4394;
  assign n4396 = pi18 ? n1741 : ~n32;
  assign n4397 = pi17 ? n32 : n4396;
  assign n4398 = pi16 ? n3438 : ~n4397;
  assign n4399 = pi15 ? n4395 : n4398;
  assign n4400 = pi16 ? n3729 : ~n4397;
  assign n4401 = pi16 ? n3165 : ~n4060;
  assign n4402 = pi15 ? n4400 : n4401;
  assign n4403 = pi14 ? n4399 : n4402;
  assign n4404 = pi13 ? n4390 : n4403;
  assign n4405 = pi12 ? n4377 : n4404;
  assign n4406 = pi20 ? n206 : ~n32;
  assign n4407 = pi19 ? n32 : n4406;
  assign n4408 = pi18 ? n4407 : ~n32;
  assign n4409 = pi17 ? n32 : n4408;
  assign n4410 = pi16 ? n3047 : ~n4409;
  assign n4411 = pi16 ? n3047 : ~n4064;
  assign n4412 = pi15 ? n4410 : n4411;
  assign n4413 = pi16 ? n3047 : ~n4055;
  assign n4414 = pi16 ? n3293 : ~n4055;
  assign n4415 = pi15 ? n4413 : n4414;
  assign n4416 = pi14 ? n4412 : n4415;
  assign n4417 = pi16 ? n3051 : ~n4055;
  assign n4418 = pi16 ? n3051 : ~n4066;
  assign n4419 = pi15 ? n4417 : n4418;
  assign n4420 = pi16 ? n2953 : ~n4066;
  assign n4421 = pi16 ? n2953 : ~n4064;
  assign n4422 = pi15 ? n4420 : n4421;
  assign n4423 = pi14 ? n4419 : n4422;
  assign n4424 = pi13 ? n4416 : n4423;
  assign n4425 = pi16 ? n3176 : ~n4064;
  assign n4426 = pi16 ? n2958 : ~n4064;
  assign n4427 = pi15 ? n4425 : n4426;
  assign n4428 = pi19 ? n1464 : ~n32;
  assign n4429 = pi18 ? n4428 : ~n32;
  assign n4430 = pi17 ? n32 : n4429;
  assign n4431 = pi16 ? n2958 : ~n4430;
  assign n4432 = pi16 ? n3183 : ~n4430;
  assign n4433 = pi15 ? n4431 : n4432;
  assign n4434 = pi14 ? n4427 : n4433;
  assign n4435 = pi16 ? n3183 : ~n3726;
  assign n4436 = pi16 ? n2832 : ~n3726;
  assign n4437 = pi15 ? n4436 : n4080;
  assign n4438 = pi14 ? n4435 : n4437;
  assign n4439 = pi13 ? n4434 : n4438;
  assign n4440 = pi12 ? n4424 : n4439;
  assign n4441 = pi11 ? n4405 : n4440;
  assign n4442 = pi16 ? n2851 : ~n3436;
  assign n4443 = pi16 ? n2851 : ~n3726;
  assign n4444 = pi15 ? n4442 : n4443;
  assign n4445 = pi16 ? n3068 : ~n3428;
  assign n4446 = pi15 ? n4443 : n4445;
  assign n4447 = pi14 ? n4444 : n4446;
  assign n4448 = pi17 ? n32 : n1120;
  assign n4449 = pi16 ? n4246 : ~n4448;
  assign n4450 = pi16 ? n2617 : ~n3157;
  assign n4451 = pi15 ? n4449 : n4450;
  assign n4452 = pi16 ? n2617 : ~n3436;
  assign n4453 = pi14 ? n4451 : n4452;
  assign n4454 = pi13 ? n4447 : n4453;
  assign n4455 = pi16 ? n2617 : ~n3428;
  assign n4456 = pi15 ? n4455 : n4452;
  assign n4457 = pi16 ? n2624 : ~n3162;
  assign n4458 = pi16 ? n2624 : ~n3157;
  assign n4459 = pi15 ? n4457 : n4458;
  assign n4460 = pi14 ? n4456 : n4459;
  assign n4461 = pi15 ? n4458 : n4457;
  assign n4462 = pi14 ? n4461 : n4457;
  assign n4463 = pi13 ? n4460 : n4462;
  assign n4464 = pi12 ? n4454 : n4463;
  assign n4465 = pi16 ? n2513 : ~n3157;
  assign n4466 = pi16 ? n2513 : ~n3162;
  assign n4467 = pi15 ? n4465 : n4466;
  assign n4468 = pi15 ? n4466 : n4465;
  assign n4469 = pi14 ? n4467 : n4468;
  assign n4470 = pi16 ? n2860 : ~n3157;
  assign n4471 = pi16 ? n2860 : ~n3436;
  assign n4472 = pi15 ? n4470 : n4471;
  assign n4473 = pi14 ? n4472 : n4470;
  assign n4474 = pi13 ? n4469 : n4473;
  assign n4475 = pi20 ? n3523 : ~n448;
  assign n4476 = pi20 ? n339 : ~n274;
  assign n4477 = pi19 ? n4475 : n4476;
  assign n4478 = pi18 ? n4477 : ~n32;
  assign n4479 = pi17 ? n32 : n4478;
  assign n4480 = pi16 ? n4100 : ~n4479;
  assign n4481 = pi16 ? n2745 : ~n3436;
  assign n4482 = pi15 ? n4480 : n4481;
  assign n4483 = pi14 ? n4470 : n4482;
  assign n4484 = pi16 ? n2745 : ~n3428;
  assign n4485 = pi14 ? n4481 : n4484;
  assign n4486 = pi13 ? n4483 : n4485;
  assign n4487 = pi12 ? n4474 : n4486;
  assign n4488 = pi11 ? n4464 : n4487;
  assign n4489 = pi10 ? n4441 : n4488;
  assign n4490 = pi09 ? n4354 : n4489;
  assign n4491 = pi20 ? n428 : n32;
  assign n4492 = pi19 ? n4491 : n32;
  assign n4493 = pi18 ? n32 : ~n4492;
  assign n4494 = pi17 ? n2159 : ~n4493;
  assign n4495 = pi16 ? n32 : n4494;
  assign n4496 = pi15 ? n32 : n4495;
  assign n4497 = pi18 ? n2730 : ~n32;
  assign n4498 = pi17 ? n4497 : ~n4344;
  assign n4499 = pi16 ? n32 : n4498;
  assign n4500 = pi17 ? n1472 : ~n4344;
  assign n4501 = pi16 ? n32 : n4500;
  assign n4502 = pi15 ? n4499 : n4501;
  assign n4503 = pi14 ? n4496 : n4502;
  assign n4504 = pi13 ? n32 : n4503;
  assign n4505 = pi12 ? n32 : n4504;
  assign n4506 = pi11 ? n32 : n4505;
  assign n4507 = pi10 ? n32 : n4506;
  assign n4508 = pi15 ? n4339 : n4356;
  assign n4509 = pi17 ? n4167 : ~n1807;
  assign n4510 = pi16 ? n32 : n4509;
  assign n4511 = pi17 ? n1215 : ~n2537;
  assign n4512 = pi16 ? n32 : n4511;
  assign n4513 = pi15 ? n4510 : n4512;
  assign n4514 = pi14 ? n4508 : n4513;
  assign n4515 = pi18 ? n2291 : ~n32;
  assign n4516 = pi17 ? n4515 : ~n2314;
  assign n4517 = pi16 ? n32 : n4516;
  assign n4518 = pi20 ? n32 : n1385;
  assign n4519 = pi19 ? n32 : n4518;
  assign n4520 = pi18 ? n4519 : ~n32;
  assign n4521 = pi17 ? n4023 : ~n4520;
  assign n4522 = pi16 ? n32 : n4521;
  assign n4523 = pi15 ? n4517 : n4522;
  assign n4524 = pi17 ? n1605 : ~n1833;
  assign n4525 = pi16 ? n32 : n4524;
  assign n4526 = pi15 ? n4372 : n4525;
  assign n4527 = pi14 ? n4523 : n4526;
  assign n4528 = pi13 ? n4514 : n4527;
  assign n4529 = pi17 ? n1227 : ~n2325;
  assign n4530 = pi16 ? n32 : n4529;
  assign n4531 = pi18 ? n1819 : ~n32;
  assign n4532 = pi17 ? n3553 : ~n4531;
  assign n4533 = pi16 ? n32 : n4532;
  assign n4534 = pi15 ? n4530 : n4533;
  assign n4535 = pi17 ? n1726 : ~n1697;
  assign n4536 = pi16 ? n32 : n4535;
  assign n4537 = pi17 ? n4041 : ~n1704;
  assign n4538 = pi16 ? n32 : n4537;
  assign n4539 = pi15 ? n4536 : n4538;
  assign n4540 = pi14 ? n4534 : n4539;
  assign n4541 = pi20 ? n1368 : n207;
  assign n4542 = pi19 ? n32 : n4541;
  assign n4543 = pi18 ? n4542 : ~n32;
  assign n4544 = pi17 ? n3719 : ~n4543;
  assign n4545 = pi16 ? n32 : n4544;
  assign n4546 = pi19 ? n32 : n2168;
  assign n4547 = pi18 ? n4546 : ~n32;
  assign n4548 = pi17 ? n32 : n4547;
  assign n4549 = pi16 ? n32 : ~n4548;
  assign n4550 = pi15 ? n4545 : n4549;
  assign n4551 = pi17 ? n32 : n2560;
  assign n4552 = pi16 ? n3570 : ~n4551;
  assign n4553 = pi16 ? n3283 : ~n4201;
  assign n4554 = pi15 ? n4552 : n4553;
  assign n4555 = pi14 ? n4550 : n4554;
  assign n4556 = pi13 ? n4540 : n4555;
  assign n4557 = pi12 ? n4528 : n4556;
  assign n4558 = pi20 ? n4279 : ~n32;
  assign n4559 = pi19 ? n32 : n4558;
  assign n4560 = pi18 ? n4559 : ~n32;
  assign n4561 = pi17 ? n32 : n4560;
  assign n4562 = pi16 ? n3156 : ~n4561;
  assign n4563 = pi17 ? n32 : n2567;
  assign n4564 = pi16 ? n3156 : ~n4563;
  assign n4565 = pi15 ? n4562 : n4564;
  assign n4566 = pi16 ? n3156 : ~n3879;
  assign n4567 = pi17 ? n32 : n2159;
  assign n4568 = pi16 ? n3438 : ~n4567;
  assign n4569 = pi15 ? n4566 : n4568;
  assign n4570 = pi14 ? n4565 : n4569;
  assign n4571 = pi16 ? n3161 : ~n4055;
  assign n4572 = pi16 ? n3165 : ~n3730;
  assign n4573 = pi15 ? n4571 : n4572;
  assign n4574 = pi16 ? n3165 : ~n4066;
  assign n4575 = pi15 ? n4574 : n4065;
  assign n4576 = pi14 ? n4573 : n4575;
  assign n4577 = pi13 ? n4570 : n4576;
  assign n4578 = pi17 ? n32 : n2959;
  assign n4579 = pi16 ? n4578 : ~n4064;
  assign n4580 = pi15 ? n4411 : n4579;
  assign n4581 = pi19 ? n1818 : ~n32;
  assign n4582 = pi18 ? n4581 : ~n32;
  assign n4583 = pi17 ? n32 : n4582;
  assign n4584 = pi16 ? n4578 : ~n4583;
  assign n4585 = pi16 ? n3051 : ~n4583;
  assign n4586 = pi15 ? n4584 : n4585;
  assign n4587 = pi14 ? n4580 : n4586;
  assign n4588 = pi17 ? n32 : n1994;
  assign n4589 = pi16 ? n3051 : ~n4588;
  assign n4590 = pi16 ? n2953 : ~n4588;
  assign n4591 = pi16 ? n2953 : ~n3734;
  assign n4592 = pi15 ? n4590 : n4591;
  assign n4593 = pi14 ? n4589 : n4592;
  assign n4594 = pi13 ? n4587 : n4593;
  assign n4595 = pi12 ? n4577 : n4594;
  assign n4596 = pi11 ? n4557 : n4595;
  assign n4597 = pi16 ? n2958 : ~n4217;
  assign n4598 = pi16 ? n2958 : ~n3726;
  assign n4599 = pi15 ? n4597 : n4598;
  assign n4600 = pi16 ? n2964 : ~n3740;
  assign n4601 = pi15 ? n4223 : n4600;
  assign n4602 = pi14 ? n4599 : n4601;
  assign n4603 = pi16 ? n3183 : ~n3740;
  assign n4604 = pi16 ? n2840 : ~n4237;
  assign n4605 = pi15 ? n4603 : n4604;
  assign n4606 = pi16 ? n2837 : ~n4448;
  assign n4607 = pi14 ? n4605 : n4606;
  assign n4608 = pi13 ? n4602 : n4607;
  assign n4609 = pi16 ? n2837 : ~n3428;
  assign n4610 = pi16 ? n2840 : ~n4217;
  assign n4611 = pi15 ? n4609 : n4610;
  assign n4612 = pi16 ? n2725 : ~n4239;
  assign n4613 = pi17 ? n32 : n1024;
  assign n4614 = pi16 ? n2725 : ~n4613;
  assign n4615 = pi15 ? n4612 : n4614;
  assign n4616 = pi14 ? n4611 : n4615;
  assign n4617 = pi16 ? n2725 : ~n4242;
  assign n4618 = pi15 ? n4614 : n4617;
  assign n4619 = pi16 ? n2725 : ~n4230;
  assign n4620 = pi16 ? n2745 : ~n4230;
  assign n4621 = pi15 ? n4619 : n4620;
  assign n4622 = pi14 ? n4618 : n4621;
  assign n4623 = pi13 ? n4616 : n4622;
  assign n4624 = pi12 ? n4608 : n4623;
  assign n4625 = pi16 ? n2745 : ~n4232;
  assign n4626 = pi15 ? n4625 : n4620;
  assign n4627 = pi15 ? n4620 : n4625;
  assign n4628 = pi14 ? n4626 : n4627;
  assign n4629 = pi16 ? n2732 : ~n4232;
  assign n4630 = pi16 ? n3068 : ~n4448;
  assign n4631 = pi15 ? n4629 : n4630;
  assign n4632 = pi16 ? n3068 : ~n4232;
  assign n4633 = pi14 ? n4631 : n4632;
  assign n4634 = pi13 ? n4628 : n4633;
  assign n4635 = pi19 ? n975 : n4476;
  assign n4636 = pi18 ? n4635 : ~n32;
  assign n4637 = pi17 ? n32 : n4636;
  assign n4638 = pi16 ? n4246 : ~n4637;
  assign n4639 = pi16 ? n2851 : ~n4448;
  assign n4640 = pi15 ? n4638 : n4639;
  assign n4641 = pi14 ? n4632 : n4640;
  assign n4642 = pi16 ? n3061 : ~n4448;
  assign n4643 = pi15 ? n4642 : n4639;
  assign n4644 = pi16 ? n2837 : ~n3572;
  assign n4645 = pi15 ? n4080 : n4644;
  assign n4646 = pi14 ? n4643 : n4645;
  assign n4647 = pi13 ? n4641 : n4646;
  assign n4648 = pi12 ? n4634 : n4647;
  assign n4649 = pi11 ? n4624 : n4648;
  assign n4650 = pi10 ? n4596 : n4649;
  assign n4651 = pi09 ? n4507 : n4650;
  assign n4652 = pi08 ? n4490 : n4651;
  assign n4653 = pi17 ? n1706 : ~n1682;
  assign n4654 = pi16 ? n32 : n4653;
  assign n4655 = pi15 ? n32 : n4654;
  assign n4656 = pi18 ? n2835 : ~n32;
  assign n4657 = pi17 ? n4656 : ~n4344;
  assign n4658 = pi16 ? n32 : n4657;
  assign n4659 = pi18 ? n4244 : ~n32;
  assign n4660 = pi17 ? n4659 : ~n4344;
  assign n4661 = pi16 ? n32 : n4660;
  assign n4662 = pi15 ? n4658 : n4661;
  assign n4663 = pi14 ? n4655 : n4662;
  assign n4664 = pi13 ? n32 : n4663;
  assign n4665 = pi12 ? n32 : n4664;
  assign n4666 = pi11 ? n32 : n4665;
  assign n4667 = pi10 ? n32 : n4666;
  assign n4668 = pi17 ? n2159 : ~n1682;
  assign n4669 = pi16 ? n32 : n4668;
  assign n4670 = pi20 ? n342 : n32;
  assign n4671 = pi19 ? n4670 : n32;
  assign n4672 = pi18 ? n32 : ~n4671;
  assign n4673 = pi17 ? n1480 : ~n4672;
  assign n4674 = pi16 ? n32 : n4673;
  assign n4675 = pi15 ? n4669 : n4674;
  assign n4676 = pi17 ? n4341 : ~n2119;
  assign n4677 = pi16 ? n32 : n4676;
  assign n4678 = pi17 ? n1989 : ~n2119;
  assign n4679 = pi16 ? n32 : n4678;
  assign n4680 = pi15 ? n4677 : n4679;
  assign n4681 = pi14 ? n4675 : n4680;
  assign n4682 = pi18 ? n2627 : ~n32;
  assign n4683 = pi17 ? n4682 : ~n1933;
  assign n4684 = pi16 ? n32 : n4683;
  assign n4685 = pi18 ? n4380 : n237;
  assign n4686 = pi17 ? n4167 : ~n4685;
  assign n4687 = pi16 ? n32 : n4686;
  assign n4688 = pi15 ? n4684 : n4687;
  assign n4689 = pi19 ? n3692 : n32;
  assign n4690 = pi18 ? n32 : ~n4689;
  assign n4691 = pi17 ? n4023 : ~n4690;
  assign n4692 = pi16 ? n32 : n4691;
  assign n4693 = pi15 ? n4692 : n4361;
  assign n4694 = pi14 ? n4688 : n4693;
  assign n4695 = pi13 ? n4681 : n4694;
  assign n4696 = pi17 ? n1120 : ~n1933;
  assign n4697 = pi16 ? n32 : n4696;
  assign n4698 = pi17 ? n4034 : ~n4685;
  assign n4699 = pi16 ? n32 : n4698;
  assign n4700 = pi15 ? n4697 : n4699;
  assign n4701 = pi17 ? n1605 : ~n2325;
  assign n4702 = pi16 ? n32 : n4701;
  assign n4703 = pi15 ? n4369 : n4702;
  assign n4704 = pi14 ? n4700 : n4703;
  assign n4705 = pi17 ? n4041 : ~n1682;
  assign n4706 = pi16 ? n32 : n4705;
  assign n4707 = pi17 ? n2005 : ~n1580;
  assign n4708 = pi16 ? n32 : n4707;
  assign n4709 = pi15 ? n4706 : n4708;
  assign n4710 = pi17 ? n3715 : ~n1580;
  assign n4711 = pi16 ? n32 : n4710;
  assign n4712 = pi17 ? n1028 : ~n1706;
  assign n4713 = pi16 ? n32 : n4712;
  assign n4714 = pi15 ? n4711 : n4713;
  assign n4715 = pi14 ? n4709 : n4714;
  assign n4716 = pi13 ? n4704 : n4715;
  assign n4717 = pi12 ? n4695 : n4716;
  assign n4718 = pi17 ? n3719 : ~n1580;
  assign n4719 = pi16 ? n32 : n4718;
  assign n4720 = pi15 ? n4719 : n4054;
  assign n4721 = pi20 ? n32 : ~n246;
  assign n4722 = pi19 ? n32 : n4721;
  assign n4723 = pi18 ? n4722 : ~n32;
  assign n4724 = pi17 ? n3557 : ~n4723;
  assign n4725 = pi16 ? n32 : n4724;
  assign n4726 = pi16 ? n32 : ~n1471;
  assign n4727 = pi15 ? n4725 : n4726;
  assign n4728 = pi14 ? n4720 : n4727;
  assign n4729 = pi17 ? n32 : n1697;
  assign n4730 = pi16 ? n3570 : ~n4729;
  assign n4731 = pi16 ? n3283 : ~n1214;
  assign n4732 = pi15 ? n4730 : n4731;
  assign n4733 = pi17 ? n32 : n1706;
  assign n4734 = pi16 ? n3283 : ~n4733;
  assign n4735 = pi16 ? n3283 : ~n4729;
  assign n4736 = pi15 ? n4734 : n4735;
  assign n4737 = pi14 ? n4732 : n4736;
  assign n4738 = pi13 ? n4728 : n4737;
  assign n4739 = pi16 ? n3156 : ~n4729;
  assign n4740 = pi17 ? n32 : n4111;
  assign n4741 = pi16 ? n4740 : ~n4733;
  assign n4742 = pi15 ? n4739 : n4741;
  assign n4743 = pi16 ? n3161 : ~n4733;
  assign n4744 = pi16 ? n3161 : ~n4060;
  assign n4745 = pi15 ? n4743 : n4744;
  assign n4746 = pi14 ? n4742 : n4745;
  assign n4747 = pi14 ? n4744 : n4414;
  assign n4748 = pi13 ? n4746 : n4747;
  assign n4749 = pi12 ? n4738 : n4748;
  assign n4750 = pi11 ? n4717 : n4749;
  assign n4751 = pi16 ? n3588 : ~n4055;
  assign n4752 = pi16 ? n3588 : ~n4060;
  assign n4753 = pi15 ? n4751 : n4752;
  assign n4754 = pi16 ? n4578 : ~n4060;
  assign n4755 = pi15 ? n4752 : n4754;
  assign n4756 = pi14 ? n4753 : n4755;
  assign n4757 = pi15 ? n4579 : n4421;
  assign n4758 = pi16 ? n2953 : ~n4055;
  assign n4759 = pi14 ? n4757 : n4758;
  assign n4760 = pi13 ? n4756 : n4759;
  assign n4761 = pi16 ? n3176 : ~n4055;
  assign n4762 = pi15 ? n4758 : n4761;
  assign n4763 = pi16 ? n2832 : ~n4064;
  assign n4764 = pi16 ? n2832 : ~n4055;
  assign n4765 = pi15 ? n4763 : n4764;
  assign n4766 = pi14 ? n4762 : n4765;
  assign n4767 = pi16 ? n3183 : ~n4064;
  assign n4768 = pi15 ? n4764 : n4767;
  assign n4769 = pi16 ? n2832 : ~n4066;
  assign n4770 = pi16 ? n2851 : ~n4066;
  assign n4771 = pi15 ? n4769 : n4770;
  assign n4772 = pi14 ? n4768 : n4771;
  assign n4773 = pi13 ? n4766 : n4772;
  assign n4774 = pi12 ? n4760 : n4773;
  assign n4775 = pi16 ? n2851 : ~n4064;
  assign n4776 = pi15 ? n4775 : n4770;
  assign n4777 = pi16 ? n3061 : ~n4064;
  assign n4778 = pi15 ? n4770 : n4777;
  assign n4779 = pi14 ? n4776 : n4778;
  assign n4780 = pi15 ? n4777 : n4764;
  assign n4781 = pi14 ? n4780 : n4763;
  assign n4782 = pi13 ? n4779 : n4781;
  assign n4783 = pi15 ? n4777 : n4763;
  assign n4784 = pi16 ? n2958 : ~n4055;
  assign n4785 = pi14 ? n4783 : n4784;
  assign n4786 = pi18 ? n697 : ~n2079;
  assign n4787 = pi17 ? n32 : n4786;
  assign n4788 = pi16 ? n2958 : ~n4787;
  assign n4789 = pi15 ? n4761 : n4788;
  assign n4790 = pi16 ? n2958 : ~n4060;
  assign n4791 = pi15 ? n4784 : n4790;
  assign n4792 = pi14 ? n4789 : n4791;
  assign n4793 = pi13 ? n4785 : n4792;
  assign n4794 = pi12 ? n4782 : n4793;
  assign n4795 = pi11 ? n4774 : n4794;
  assign n4796 = pi10 ? n4750 : n4795;
  assign n4797 = pi09 ? n4667 : n4796;
  assign n4798 = pi18 ? n2962 : ~n32;
  assign n4799 = pi17 ? n4798 : ~n1682;
  assign n4800 = pi16 ? n32 : n4799;
  assign n4801 = pi15 ? n32 : n4800;
  assign n4802 = pi17 ? n1966 : ~n4344;
  assign n4803 = pi16 ? n32 : n4802;
  assign n4804 = pi18 ? n2830 : ~n32;
  assign n4805 = pi17 ? n4804 : ~n4344;
  assign n4806 = pi16 ? n32 : n4805;
  assign n4807 = pi15 ? n4803 : n4806;
  assign n4808 = pi14 ? n4801 : n4807;
  assign n4809 = pi13 ? n32 : n4808;
  assign n4810 = pi12 ? n32 : n4809;
  assign n4811 = pi11 ? n32 : n4810;
  assign n4812 = pi10 ? n32 : n4811;
  assign n4813 = pi17 ? n2159 : ~n4672;
  assign n4814 = pi16 ? n32 : n4813;
  assign n4815 = pi15 ? n4654 : n4814;
  assign n4816 = pi17 ? n4497 : ~n2119;
  assign n4817 = pi16 ? n32 : n4816;
  assign n4818 = pi17 ? n1472 : ~n2119;
  assign n4819 = pi16 ? n32 : n4818;
  assign n4820 = pi15 ? n4817 : n4819;
  assign n4821 = pi14 ? n4815 : n4820;
  assign n4822 = pi18 ? n2615 : ~n32;
  assign n4823 = pi17 ? n4822 : ~n1933;
  assign n4824 = pi16 ? n32 : n4823;
  assign n4825 = pi17 ? n4341 : ~n4685;
  assign n4826 = pi16 ? n32 : n4825;
  assign n4827 = pi15 ? n4824 : n4826;
  assign n4828 = pi17 ? n4167 : ~n4690;
  assign n4829 = pi16 ? n32 : n4828;
  assign n4830 = pi17 ? n4167 : ~n2537;
  assign n4831 = pi16 ? n32 : n4830;
  assign n4832 = pi15 ? n4829 : n4831;
  assign n4833 = pi14 ? n4827 : n4832;
  assign n4834 = pi13 ? n4821 : n4833;
  assign n4835 = pi17 ? n1215 : ~n1933;
  assign n4836 = pi16 ? n32 : n4835;
  assign n4837 = pi17 ? n4515 : ~n4685;
  assign n4838 = pi16 ? n32 : n4837;
  assign n4839 = pi15 ? n4836 : n4838;
  assign n4840 = pi17 ? n4023 : ~n1470;
  assign n4841 = pi16 ? n32 : n4840;
  assign n4842 = pi17 ? n1605 : ~n2136;
  assign n4843 = pi16 ? n32 : n4842;
  assign n4844 = pi15 ? n4841 : n4843;
  assign n4845 = pi14 ? n4839 : n4844;
  assign n4846 = pi17 ? n1605 : ~n1682;
  assign n4847 = pi16 ? n32 : n4846;
  assign n4848 = pi17 ? n1227 : ~n1580;
  assign n4849 = pi16 ? n32 : n4848;
  assign n4850 = pi15 ? n4847 : n4849;
  assign n4851 = pi17 ? n3553 : ~n1580;
  assign n4852 = pi16 ? n32 : n4851;
  assign n4853 = pi17 ? n1726 : ~n1706;
  assign n4854 = pi16 ? n32 : n4853;
  assign n4855 = pi15 ? n4852 : n4854;
  assign n4856 = pi14 ? n4850 : n4855;
  assign n4857 = pi13 ? n4845 : n4856;
  assign n4858 = pi12 ? n4834 : n4857;
  assign n4859 = pi17 ? n4041 : ~n2433;
  assign n4860 = pi16 ? n32 : n4859;
  assign n4861 = pi20 ? n32 : ~n1368;
  assign n4862 = pi19 ? n32 : n4861;
  assign n4863 = pi18 ? n4862 : ~n32;
  assign n4864 = pi17 ? n4041 : ~n4863;
  assign n4865 = pi16 ? n32 : n4864;
  assign n4866 = pi15 ? n4860 : n4865;
  assign n4867 = pi20 ? n32 : ~n1385;
  assign n4868 = pi19 ? n32 : n4867;
  assign n4869 = pi18 ? n4868 : ~n32;
  assign n4870 = pi17 ? n3704 : ~n4869;
  assign n4871 = pi16 ? n32 : n4870;
  assign n4872 = pi17 ? n2005 : ~n2332;
  assign n4873 = pi16 ? n32 : n4872;
  assign n4874 = pi15 ? n4871 : n4873;
  assign n4875 = pi14 ? n4866 : n4874;
  assign n4876 = pi17 ? n3715 : ~n1697;
  assign n4877 = pi16 ? n32 : n4876;
  assign n4878 = pi17 ? n1028 : ~n1704;
  assign n4879 = pi16 ? n32 : n4878;
  assign n4880 = pi15 ? n4877 : n4879;
  assign n4881 = pi17 ? n1028 : ~n2446;
  assign n4882 = pi16 ? n32 : n4881;
  assign n4883 = pi17 ? n2008 : ~n1134;
  assign n4884 = pi16 ? n32 : n4883;
  assign n4885 = pi15 ? n4882 : n4884;
  assign n4886 = pi14 ? n4880 : n4885;
  assign n4887 = pi13 ? n4875 : n4886;
  assign n4888 = pi17 ? n3557 : ~n2150;
  assign n4889 = pi16 ? n32 : n4888;
  assign n4890 = pi17 ? n32 : n2555;
  assign n4891 = pi16 ? n32 : ~n4890;
  assign n4892 = pi15 ? n4889 : n4891;
  assign n4893 = pi16 ? n3570 : ~n4733;
  assign n4894 = pi16 ? n3570 : ~n4060;
  assign n4895 = pi15 ? n4893 : n4894;
  assign n4896 = pi14 ? n4892 : n4895;
  assign n4897 = pi16 ? n3438 : ~n3879;
  assign n4898 = pi16 ? n3729 : ~n3879;
  assign n4899 = pi15 ? n4897 : n4898;
  assign n4900 = pi14 ? n4202 : n4899;
  assign n4901 = pi13 ? n4896 : n4900;
  assign n4902 = pi12 ? n4887 : n4901;
  assign n4903 = pi11 ? n4858 : n4902;
  assign n4904 = pi16 ? n3729 : ~n4055;
  assign n4905 = pi18 ? n1387 : ~n32;
  assign n4906 = pi17 ? n32 : n4905;
  assign n4907 = pi16 ? n3729 : ~n4906;
  assign n4908 = pi15 ? n4904 : n4907;
  assign n4909 = pi15 ? n4062 : n4401;
  assign n4910 = pi14 ? n4908 : n4909;
  assign n4911 = pi16 ? n3165 : ~n4563;
  assign n4912 = pi16 ? n3047 : ~n4563;
  assign n4913 = pi15 ? n4911 : n4912;
  assign n4914 = pi16 ? n3047 : ~n3879;
  assign n4915 = pi14 ? n4913 : n4914;
  assign n4916 = pi13 ? n4910 : n4915;
  assign n4917 = pi18 ? n2242 : ~n32;
  assign n4918 = pi17 ? n32 : n4917;
  assign n4919 = pi16 ? n3047 : ~n4918;
  assign n4920 = pi15 ? n4919 : n4413;
  assign n4921 = pi17 ? n32 : n1984;
  assign n4922 = pi16 ? n2953 : ~n4921;
  assign n4923 = pi15 ? n4922 : n4751;
  assign n4924 = pi14 ? n4920 : n4923;
  assign n4925 = pi16 ? n3588 : ~n4921;
  assign n4926 = pi15 ? n4751 : n4925;
  assign n4927 = pi16 ? n4578 : ~n3730;
  assign n4928 = pi16 ? n2832 : ~n3730;
  assign n4929 = pi15 ? n4927 : n4928;
  assign n4930 = pi14 ? n4926 : n4929;
  assign n4931 = pi13 ? n4924 : n4930;
  assign n4932 = pi12 ? n4916 : n4931;
  assign n4933 = pi16 ? n2958 : ~n3730;
  assign n4934 = pi15 ? n4426 : n4933;
  assign n4935 = pi18 ? n3975 : ~n32;
  assign n4936 = pi17 ? n32 : n4935;
  assign n4937 = pi16 ? n2958 : ~n4936;
  assign n4938 = pi16 ? n3176 : ~n4563;
  assign n4939 = pi15 ? n4937 : n4938;
  assign n4940 = pi14 ? n4934 : n4939;
  assign n4941 = pi15 ? n4938 : n4761;
  assign n4942 = pi16 ? n4578 : ~n4563;
  assign n4943 = pi15 ? n4938 : n4942;
  assign n4944 = pi14 ? n4941 : n4943;
  assign n4945 = pi13 ? n4940 : n4944;
  assign n4946 = pi16 ? n3588 : ~n3879;
  assign n4947 = pi15 ? n4946 : n4751;
  assign n4948 = pi14 ? n4942 : n4947;
  assign n4949 = pi18 ? n503 : ~n2079;
  assign n4950 = pi17 ? n32 : n4949;
  assign n4951 = pi16 ? n3165 : ~n4950;
  assign n4952 = pi15 ? n4946 : n4951;
  assign n4953 = pi16 ? n3047 : ~n4199;
  assign n4954 = pi15 ? n4914 : n4953;
  assign n4955 = pi14 ? n4952 : n4954;
  assign n4956 = pi13 ? n4948 : n4955;
  assign n4957 = pi12 ? n4945 : n4956;
  assign n4958 = pi11 ? n4932 : n4957;
  assign n4959 = pi10 ? n4903 : n4958;
  assign n4960 = pi09 ? n4812 : n4959;
  assign n4961 = pi08 ? n4797 : n4960;
  assign n4962 = pi07 ? n4652 : n4961;
  assign n4963 = pi06 ? n4337 : n4962;
  assign n4964 = pi20 ? n321 : ~n321;
  assign n4965 = pi19 ? n4964 : n322;
  assign n4966 = pi18 ? n4965 : ~n32;
  assign n4967 = pi17 ? n1971 : ~n4966;
  assign n4968 = pi16 ? n32 : n4967;
  assign n4969 = pi15 ? n32 : n4968;
  assign n4970 = pi19 ? n4670 : n208;
  assign n4971 = pi18 ? n4970 : ~n32;
  assign n4972 = pi17 ? n930 : ~n4971;
  assign n4973 = pi16 ? n32 : n4972;
  assign n4974 = pi17 ? n1134 : ~n1697;
  assign n4975 = pi16 ? n32 : n4974;
  assign n4976 = pi15 ? n4973 : n4975;
  assign n4977 = pi14 ? n4969 : n4976;
  assign n4978 = pi13 ? n32 : n4977;
  assign n4979 = pi12 ? n32 : n4978;
  assign n4980 = pi11 ? n32 : n4979;
  assign n4981 = pi10 ? n32 : n4980;
  assign n4982 = pi20 ? n32 : ~n342;
  assign n4983 = pi19 ? n4982 : n32;
  assign n4984 = pi18 ? n863 : ~n4983;
  assign n4985 = pi17 ? n1706 : ~n4984;
  assign n4986 = pi16 ? n32 : n4985;
  assign n4987 = pi18 ? n940 : ~n4983;
  assign n4988 = pi17 ? n1706 : ~n4987;
  assign n4989 = pi16 ? n32 : n4988;
  assign n4990 = pi15 ? n4986 : n4989;
  assign n4991 = pi17 ? n4656 : ~n1697;
  assign n4992 = pi16 ? n32 : n4991;
  assign n4993 = pi19 ? n4342 : n531;
  assign n4994 = pi18 ? n4993 : ~n32;
  assign n4995 = pi17 ? n1700 : ~n4994;
  assign n4996 = pi16 ? n32 : n4995;
  assign n4997 = pi15 ? n4992 : n4996;
  assign n4998 = pi14 ? n4990 : n4997;
  assign n4999 = pi17 ? n2159 : ~n1697;
  assign n5000 = pi16 ? n32 : n4999;
  assign n5001 = pi17 ? n4497 : ~n1470;
  assign n5002 = pi16 ? n32 : n5001;
  assign n5003 = pi15 ? n5000 : n5002;
  assign n5004 = pi20 ? n321 : ~n207;
  assign n5005 = pi19 ? n5004 : n32;
  assign n5006 = pi18 ? n32 : ~n5005;
  assign n5007 = pi17 ? n4341 : ~n5006;
  assign n5008 = pi16 ? n32 : n5007;
  assign n5009 = pi19 ? n4964 : n32;
  assign n5010 = pi18 ? n32 : ~n5009;
  assign n5011 = pi17 ? n4341 : ~n5010;
  assign n5012 = pi16 ? n32 : n5011;
  assign n5013 = pi15 ? n5008 : n5012;
  assign n5014 = pi14 ? n5003 : n5013;
  assign n5015 = pi13 ? n4998 : n5014;
  assign n5016 = pi17 ? n4682 : ~n2531;
  assign n5017 = pi16 ? n32 : n5016;
  assign n5018 = pi15 ? n4679 : n5017;
  assign n5019 = pi17 ? n4023 : ~n1933;
  assign n5020 = pi16 ? n32 : n5019;
  assign n5021 = pi15 ? n4510 : n5020;
  assign n5022 = pi14 ? n5018 : n5021;
  assign n5023 = pi17 ? n4023 : ~n2531;
  assign n5024 = pi16 ? n32 : n5023;
  assign n5025 = pi17 ? n1120 : ~n2531;
  assign n5026 = pi16 ? n32 : n5025;
  assign n5027 = pi15 ? n5024 : n5026;
  assign n5028 = pi17 ? n4034 : ~n1933;
  assign n5029 = pi16 ? n32 : n5028;
  assign n5030 = pi17 ? n1219 : ~n1807;
  assign n5031 = pi16 ? n32 : n5030;
  assign n5032 = pi15 ? n5029 : n5031;
  assign n5033 = pi14 ? n5027 : n5032;
  assign n5034 = pi13 ? n5022 : n5033;
  assign n5035 = pi12 ? n5015 : n5034;
  assign n5036 = pi17 ? n1605 : ~n1807;
  assign n5037 = pi16 ? n32 : n5036;
  assign n5038 = pi17 ? n3855 : ~n1933;
  assign n5039 = pi16 ? n32 : n5038;
  assign n5040 = pi17 ? n1227 : ~n1807;
  assign n5041 = pi16 ? n32 : n5040;
  assign n5042 = pi15 ? n5039 : n5041;
  assign n5043 = pi14 ? n5037 : n5042;
  assign n5044 = pi17 ? n3553 : ~n1682;
  assign n5045 = pi16 ? n32 : n5044;
  assign n5046 = pi17 ? n1726 : ~n2325;
  assign n5047 = pi16 ? n32 : n5046;
  assign n5048 = pi15 ? n5045 : n5047;
  assign n5049 = pi17 ? n1500 : ~n1807;
  assign n5050 = pi16 ? n32 : n5049;
  assign n5051 = pi15 ? n5047 : n5050;
  assign n5052 = pi14 ? n5048 : n5051;
  assign n5053 = pi13 ? n5043 : n5052;
  assign n5054 = pi17 ? n3704 : ~n2325;
  assign n5055 = pi16 ? n32 : n5054;
  assign n5056 = pi17 ? n2005 : ~n1682;
  assign n5057 = pi16 ? n32 : n5056;
  assign n5058 = pi15 ? n5055 : n5057;
  assign n5059 = pi17 ? n3715 : ~n2325;
  assign n5060 = pi16 ? n32 : n5059;
  assign n5061 = pi15 ? n5060 : n4049;
  assign n5062 = pi14 ? n5058 : n5061;
  assign n5063 = pi17 ? n3719 : ~n1682;
  assign n5064 = pi16 ? n32 : n5063;
  assign n5065 = pi15 ? n4719 : n5064;
  assign n5066 = pi17 ? n2008 : ~n1580;
  assign n5067 = pi16 ? n32 : n5066;
  assign n5068 = pi17 ? n3557 : ~n1580;
  assign n5069 = pi16 ? n32 : n5068;
  assign n5070 = pi15 ? n5067 : n5069;
  assign n5071 = pi14 ? n5065 : n5070;
  assign n5072 = pi13 ? n5062 : n5071;
  assign n5073 = pi12 ? n5053 : n5072;
  assign n5074 = pi11 ? n5035 : n5073;
  assign n5075 = pi17 ? n3557 : ~n1213;
  assign n5076 = pi16 ? n32 : n5075;
  assign n5077 = pi18 ? n940 : n237;
  assign n5078 = pi17 ? n3557 : ~n5077;
  assign n5079 = pi16 ? n32 : n5078;
  assign n5080 = pi15 ? n5079 : n4731;
  assign n5081 = pi14 ? n5076 : n5080;
  assign n5082 = pi16 ? n3156 : ~n1581;
  assign n5083 = pi16 ? n3156 : ~n1471;
  assign n5084 = pi15 ? n5082 : n5083;
  assign n5085 = pi14 ? n5084 : n5083;
  assign n5086 = pi13 ? n5081 : n5085;
  assign n5087 = pi16 ? n3729 : ~n1471;
  assign n5088 = pi17 ? n32 : n1958;
  assign n5089 = pi16 ? n3729 : ~n5088;
  assign n5090 = pi15 ? n5087 : n5089;
  assign n5091 = pi16 ? n4740 : ~n1214;
  assign n5092 = pi14 ? n5090 : n5091;
  assign n5093 = pi16 ? n4740 : ~n4729;
  assign n5094 = pi16 ? n3588 : ~n1214;
  assign n5095 = pi15 ? n5091 : n5094;
  assign n5096 = pi14 ? n5093 : n5095;
  assign n5097 = pi13 ? n5092 : n5096;
  assign n5098 = pi12 ? n5086 : n5097;
  assign n5099 = pi16 ? n3588 : ~n4729;
  assign n5100 = pi15 ? n5094 : n5099;
  assign n5101 = pi16 ? n3165 : ~n1214;
  assign n5102 = pi16 ? n3165 : ~n4729;
  assign n5103 = pi15 ? n5101 : n5102;
  assign n5104 = pi14 ? n5100 : n5103;
  assign n5105 = pi16 ? n3165 : ~n1471;
  assign n5106 = pi15 ? n5105 : n5101;
  assign n5107 = pi16 ? n3161 : ~n1214;
  assign n5108 = pi15 ? n5101 : n5107;
  assign n5109 = pi14 ? n5106 : n5108;
  assign n5110 = pi13 ? n5104 : n5109;
  assign n5111 = pi16 ? n3161 : ~n1471;
  assign n5112 = pi18 ? n940 : ~n1106;
  assign n5113 = pi17 ? n32 : n5112;
  assign n5114 = pi16 ? n3438 : ~n5113;
  assign n5115 = pi16 ? n3438 : ~n4729;
  assign n5116 = pi15 ? n5114 : n5115;
  assign n5117 = pi14 ? n5111 : n5116;
  assign n5118 = pi16 ? n3438 : ~n1471;
  assign n5119 = pi18 ? n940 : ~n2079;
  assign n5120 = pi17 ? n32 : n5119;
  assign n5121 = pi16 ? n3156 : ~n5120;
  assign n5122 = pi15 ? n5118 : n5121;
  assign n5123 = pi16 ? n3438 : ~n1581;
  assign n5124 = pi16 ? n3438 : ~n1683;
  assign n5125 = pi15 ? n5123 : n5124;
  assign n5126 = pi14 ? n5122 : n5125;
  assign n5127 = pi13 ? n5117 : n5126;
  assign n5128 = pi12 ? n5110 : n5127;
  assign n5129 = pi11 ? n5098 : n5128;
  assign n5130 = pi10 ? n5074 : n5129;
  assign n5131 = pi09 ? n4981 : n5130;
  assign n5132 = pi17 ? n1593 : ~n4966;
  assign n5133 = pi16 ? n32 : n5132;
  assign n5134 = pi15 ? n32 : n5133;
  assign n5135 = pi17 ? n1470 : ~n4971;
  assign n5136 = pi16 ? n32 : n5135;
  assign n5137 = pi17 ? n1470 : ~n1697;
  assign n5138 = pi16 ? n32 : n5137;
  assign n5139 = pi15 ? n5136 : n5138;
  assign n5140 = pi14 ? n5134 : n5139;
  assign n5141 = pi13 ? n32 : n5140;
  assign n5142 = pi12 ? n32 : n5141;
  assign n5143 = pi11 ? n32 : n5142;
  assign n5144 = pi10 ? n32 : n5143;
  assign n5145 = pi17 ? n1134 : ~n4984;
  assign n5146 = pi16 ? n32 : n5145;
  assign n5147 = pi17 ? n1134 : ~n4987;
  assign n5148 = pi16 ? n32 : n5147;
  assign n5149 = pi15 ? n5146 : n5148;
  assign n5150 = pi17 ? n1966 : ~n1697;
  assign n5151 = pi16 ? n32 : n5150;
  assign n5152 = pi17 ? n4804 : ~n4994;
  assign n5153 = pi16 ? n32 : n5152;
  assign n5154 = pi15 ? n5151 : n5153;
  assign n5155 = pi14 ? n5149 : n5154;
  assign n5156 = pi17 ? n1706 : ~n1697;
  assign n5157 = pi16 ? n32 : n5156;
  assign n5158 = pi19 ? n275 : n32;
  assign n5159 = pi18 ? n940 : ~n5158;
  assign n5160 = pi17 ? n4656 : ~n5159;
  assign n5161 = pi16 ? n32 : n5160;
  assign n5162 = pi15 ? n5157 : n5161;
  assign n5163 = pi20 ? n321 : ~n749;
  assign n5164 = pi19 ? n5163 : n32;
  assign n5165 = pi18 ? n32 : ~n5164;
  assign n5166 = pi17 ? n4497 : ~n5165;
  assign n5167 = pi16 ? n32 : n5166;
  assign n5168 = pi17 ? n4497 : ~n5010;
  assign n5169 = pi16 ? n32 : n5168;
  assign n5170 = pi15 ? n5167 : n5169;
  assign n5171 = pi14 ? n5162 : n5170;
  assign n5172 = pi13 ? n5155 : n5171;
  assign n5173 = pi17 ? n4822 : ~n2531;
  assign n5174 = pi16 ? n32 : n5173;
  assign n5175 = pi15 ? n4819 : n5174;
  assign n5176 = pi17 ? n4341 : ~n1807;
  assign n5177 = pi16 ? n32 : n5176;
  assign n5178 = pi17 ? n4167 : ~n1933;
  assign n5179 = pi16 ? n32 : n5178;
  assign n5180 = pi15 ? n5177 : n5179;
  assign n5181 = pi14 ? n5175 : n5180;
  assign n5182 = pi17 ? n4167 : ~n2531;
  assign n5183 = pi16 ? n32 : n5182;
  assign n5184 = pi17 ? n1215 : ~n2531;
  assign n5185 = pi16 ? n32 : n5184;
  assign n5186 = pi15 ? n5183 : n5185;
  assign n5187 = pi17 ? n4515 : ~n1933;
  assign n5188 = pi16 ? n32 : n5187;
  assign n5189 = pi15 ? n5188 : n4361;
  assign n5190 = pi14 ? n5186 : n5189;
  assign n5191 = pi13 ? n5181 : n5190;
  assign n5192 = pi12 ? n5172 : n5191;
  assign n5193 = pi17 ? n4023 : ~n2537;
  assign n5194 = pi16 ? n32 : n5193;
  assign n5195 = pi15 ? n5194 : n4361;
  assign n5196 = pi15 ? n5020 : n4363;
  assign n5197 = pi14 ? n5195 : n5196;
  assign n5198 = pi17 ? n4034 : ~n3100;
  assign n5199 = pi16 ? n32 : n5198;
  assign n5200 = pi17 ? n4037 : ~n2314;
  assign n5201 = pi16 ? n32 : n5200;
  assign n5202 = pi15 ? n5199 : n5201;
  assign n5203 = pi17 ? n4037 : ~n2325;
  assign n5204 = pi16 ? n32 : n5203;
  assign n5205 = pi19 ? n349 : ~n482;
  assign n5206 = pi18 ? n32 : n5205;
  assign n5207 = pi17 ? n1605 : ~n5206;
  assign n5208 = pi16 ? n32 : n5207;
  assign n5209 = pi15 ? n5204 : n5208;
  assign n5210 = pi14 ? n5202 : n5209;
  assign n5211 = pi13 ? n5197 : n5210;
  assign n5212 = pi17 ? n3855 : ~n2136;
  assign n5213 = pi16 ? n32 : n5212;
  assign n5214 = pi17 ? n1227 : ~n3100;
  assign n5215 = pi16 ? n32 : n5214;
  assign n5216 = pi15 ? n5213 : n5215;
  assign n5217 = pi17 ? n3553 : ~n2325;
  assign n5218 = pi16 ? n32 : n5217;
  assign n5219 = pi17 ? n3553 : ~n3112;
  assign n5220 = pi16 ? n32 : n5219;
  assign n5221 = pi15 ? n5218 : n5220;
  assign n5222 = pi14 ? n5216 : n5221;
  assign n5223 = pi17 ? n4041 : ~n2133;
  assign n5224 = pi16 ? n32 : n5223;
  assign n5225 = pi17 ? n4041 : ~n3100;
  assign n5226 = pi16 ? n32 : n5225;
  assign n5227 = pi15 ? n5224 : n5226;
  assign n5228 = pi17 ? n1500 : ~n1833;
  assign n5229 = pi16 ? n32 : n5228;
  assign n5230 = pi17 ? n3704 : ~n1833;
  assign n5231 = pi16 ? n32 : n5230;
  assign n5232 = pi15 ? n5229 : n5231;
  assign n5233 = pi14 ? n5227 : n5232;
  assign n5234 = pi13 ? n5222 : n5233;
  assign n5235 = pi12 ? n5211 : n5234;
  assign n5236 = pi11 ? n5192 : n5235;
  assign n5237 = pi17 ? n3704 : ~n3380;
  assign n5238 = pi16 ? n32 : n5237;
  assign n5239 = pi17 ? n3715 : ~n3380;
  assign n5240 = pi16 ? n32 : n5239;
  assign n5241 = pi15 ? n5238 : n5240;
  assign n5242 = pi18 ? n1862 : n237;
  assign n5243 = pi17 ? n3715 : ~n5242;
  assign n5244 = pi16 ? n32 : n5243;
  assign n5245 = pi17 ? n1028 : ~n3388;
  assign n5246 = pi16 ? n32 : n5245;
  assign n5247 = pi15 ? n5244 : n5246;
  assign n5248 = pi14 ? n5241 : n5247;
  assign n5249 = pi17 ? n3719 : ~n1470;
  assign n5250 = pi16 ? n32 : n5249;
  assign n5251 = pi15 ? n4719 : n5250;
  assign n5252 = pi17 ? n3719 : ~n1593;
  assign n5253 = pi16 ? n32 : n5252;
  assign n5254 = pi15 ? n5250 : n5253;
  assign n5255 = pi14 ? n5251 : n5254;
  assign n5256 = pi13 ? n5248 : n5255;
  assign n5257 = pi17 ? n3557 : ~n1593;
  assign n5258 = pi16 ? n32 : n5257;
  assign n5259 = pi17 ? n32 : n2899;
  assign n5260 = pi16 ? n3283 : ~n5259;
  assign n5261 = pi15 ? n5258 : n5260;
  assign n5262 = pi17 ? n32 : n3380;
  assign n5263 = pi16 ? n32 : ~n5262;
  assign n5264 = pi16 ? n3283 : ~n5262;
  assign n5265 = pi15 ? n5263 : n5264;
  assign n5266 = pi14 ? n5261 : n5265;
  assign n5267 = pi19 ? n32 : n87;
  assign n5268 = pi18 ? n2906 : ~n5267;
  assign n5269 = pi17 ? n32 : n5268;
  assign n5270 = pi16 ? n32 : ~n5269;
  assign n5271 = pi17 ? n32 : n2907;
  assign n5272 = pi16 ? n3283 : ~n5271;
  assign n5273 = pi15 ? n5270 : n5272;
  assign n5274 = pi16 ? n3283 : ~n1705;
  assign n5275 = pi16 ? n3729 : ~n1705;
  assign n5276 = pi15 ? n5274 : n5275;
  assign n5277 = pi14 ? n5273 : n5276;
  assign n5278 = pi13 ? n5266 : n5277;
  assign n5279 = pi12 ? n5256 : n5278;
  assign n5280 = pi16 ? n3438 : ~n1705;
  assign n5281 = pi17 ? n32 : n2670;
  assign n5282 = pi16 ? n3438 : ~n5281;
  assign n5283 = pi15 ? n5280 : n5282;
  assign n5284 = pi16 ? n3156 : ~n5088;
  assign n5285 = pi16 ? n3156 : ~n5281;
  assign n5286 = pi15 ? n5284 : n5285;
  assign n5287 = pi14 ? n5283 : n5286;
  assign n5288 = pi16 ? n3156 : ~n1594;
  assign n5289 = pi18 ? n1957 : ~n1526;
  assign n5290 = pi17 ? n32 : n5289;
  assign n5291 = pi16 ? n3570 : ~n5290;
  assign n5292 = pi15 ? n5288 : n5291;
  assign n5293 = pi16 ? n3570 : ~n5088;
  assign n5294 = pi15 ? n5284 : n5293;
  assign n5295 = pi14 ? n5292 : n5294;
  assign n5296 = pi13 ? n5287 : n5295;
  assign n5297 = pi16 ? n32 : ~n1594;
  assign n5298 = pi17 ? n3557 : ~n2899;
  assign n5299 = pi16 ? n32 : n5298;
  assign n5300 = pi17 ? n3557 : ~n2907;
  assign n5301 = pi16 ? n32 : n5300;
  assign n5302 = pi15 ? n5299 : n5301;
  assign n5303 = pi14 ? n5297 : n5302;
  assign n5304 = pi18 ? n2197 : ~n2079;
  assign n5305 = pi17 ? n3719 : ~n5304;
  assign n5306 = pi16 ? n32 : n5305;
  assign n5307 = pi15 ? n5299 : n5306;
  assign n5308 = pi17 ? n1028 : ~n1833;
  assign n5309 = pi16 ? n32 : n5308;
  assign n5310 = pi17 ? n1028 : ~n2123;
  assign n5311 = pi16 ? n32 : n5310;
  assign n5312 = pi15 ? n5309 : n5311;
  assign n5313 = pi14 ? n5307 : n5312;
  assign n5314 = pi13 ? n5303 : n5313;
  assign n5315 = pi12 ? n5296 : n5314;
  assign n5316 = pi11 ? n5279 : n5315;
  assign n5317 = pi10 ? n5236 : n5316;
  assign n5318 = pi09 ? n5144 : n5317;
  assign n5319 = pi08 ? n5131 : n5318;
  assign n5320 = pi17 ? n1833 : ~n4966;
  assign n5321 = pi16 ? n32 : n5320;
  assign n5322 = pi15 ? n32 : n5321;
  assign n5323 = pi19 ? n4491 : n208;
  assign n5324 = pi18 ? n5323 : ~n32;
  assign n5325 = pi17 ? n2143 : ~n5324;
  assign n5326 = pi16 ? n32 : n5325;
  assign n5327 = pi17 ? n1322 : ~n1697;
  assign n5328 = pi16 ? n32 : n5327;
  assign n5329 = pi15 ? n5326 : n5328;
  assign n5330 = pi14 ? n5322 : n5329;
  assign n5331 = pi13 ? n32 : n5330;
  assign n5332 = pi12 ? n32 : n5331;
  assign n5333 = pi11 ? n32 : n5332;
  assign n5334 = pi10 ? n32 : n5333;
  assign n5335 = pi19 ? n531 : n32;
  assign n5336 = pi18 ? n863 : ~n5335;
  assign n5337 = pi17 ? n1971 : ~n5336;
  assign n5338 = pi16 ? n32 : n5337;
  assign n5339 = pi17 ? n1971 : ~n4987;
  assign n5340 = pi16 ? n32 : n5339;
  assign n5341 = pi15 ? n5338 : n5340;
  assign n5342 = pi17 ? n1213 : ~n1697;
  assign n5343 = pi16 ? n32 : n5342;
  assign n5344 = pi17 ? n1134 : ~n4994;
  assign n5345 = pi16 ? n32 : n5344;
  assign n5346 = pi15 ? n5343 : n5345;
  assign n5347 = pi14 ? n5341 : n5346;
  assign n5348 = pi17 ? n1232 : ~n1697;
  assign n5349 = pi16 ? n32 : n5348;
  assign n5350 = pi20 ? n32 : n1685;
  assign n5351 = pi19 ? n5350 : n32;
  assign n5352 = pi18 ? n940 : ~n5351;
  assign n5353 = pi17 ? n4656 : ~n5352;
  assign n5354 = pi16 ? n32 : n5353;
  assign n5355 = pi15 ? n5349 : n5354;
  assign n5356 = pi20 ? n321 : ~n342;
  assign n5357 = pi19 ? n5356 : n32;
  assign n5358 = pi18 ? n32 : ~n5357;
  assign n5359 = pi17 ? n4656 : ~n5358;
  assign n5360 = pi16 ? n32 : n5359;
  assign n5361 = pi17 ? n4656 : ~n5010;
  assign n5362 = pi16 ? n32 : n5361;
  assign n5363 = pi15 ? n5360 : n5362;
  assign n5364 = pi14 ? n5355 : n5363;
  assign n5365 = pi13 ? n5347 : n5364;
  assign n5366 = pi17 ? n1700 : ~n2119;
  assign n5367 = pi16 ? n32 : n5366;
  assign n5368 = pi17 ? n2159 : ~n2531;
  assign n5369 = pi16 ? n32 : n5368;
  assign n5370 = pi15 ? n5367 : n5369;
  assign n5371 = pi20 ? n321 : ~n266;
  assign n5372 = pi19 ? n5371 : ~n32;
  assign n5373 = pi18 ? n32 : n5372;
  assign n5374 = pi17 ? n4497 : ~n5373;
  assign n5375 = pi16 ? n32 : n5374;
  assign n5376 = pi17 ? n4341 : ~n2519;
  assign n5377 = pi16 ? n32 : n5376;
  assign n5378 = pi15 ? n5375 : n5377;
  assign n5379 = pi14 ? n5370 : n5378;
  assign n5380 = pi15 ? n4684 : n4510;
  assign n5381 = pi14 ? n4680 : n5380;
  assign n5382 = pi13 ? n5379 : n5381;
  assign n5383 = pi12 ? n5365 : n5382;
  assign n5384 = pi17 ? n4167 : ~n2119;
  assign n5385 = pi16 ? n32 : n5384;
  assign n5386 = pi15 ? n5183 : n5385;
  assign n5387 = pi15 ? n5385 : n5185;
  assign n5388 = pi14 ? n5386 : n5387;
  assign n5389 = pi17 ? n2355 : ~n1933;
  assign n5390 = pi16 ? n32 : n5389;
  assign n5391 = pi13 ? n5388 : n5390;
  assign n5392 = pi15 ? n5024 : n4363;
  assign n5393 = pi17 ? n1219 : ~n1933;
  assign n5394 = pi16 ? n32 : n5393;
  assign n5395 = pi15 ? n5394 : n5031;
  assign n5396 = pi14 ? n5392 : n5395;
  assign n5397 = pi17 ? n4037 : ~n1807;
  assign n5398 = pi16 ? n32 : n5397;
  assign n5399 = pi17 ? n4037 : ~n1933;
  assign n5400 = pi16 ? n32 : n5399;
  assign n5401 = pi15 ? n5398 : n5400;
  assign n5402 = pi15 ? n5037 : n5039;
  assign n5403 = pi14 ? n5401 : n5402;
  assign n5404 = pi13 ? n5396 : n5403;
  assign n5405 = pi12 ? n5391 : n5404;
  assign n5406 = pi11 ? n5383 : n5405;
  assign n5407 = pi17 ? n3855 : ~n1807;
  assign n5408 = pi16 ? n32 : n5407;
  assign n5409 = pi17 ? n3553 : ~n1807;
  assign n5410 = pi16 ? n32 : n5409;
  assign n5411 = pi15 ? n5408 : n5410;
  assign n5412 = pi17 ? n1726 : ~n1807;
  assign n5413 = pi16 ? n32 : n5412;
  assign n5414 = pi15 ? n5410 : n5413;
  assign n5415 = pi14 ? n5411 : n5414;
  assign n5416 = pi17 ? n4041 : ~n1807;
  assign n5417 = pi16 ? n32 : n5416;
  assign n5418 = pi17 ? n3704 : ~n1807;
  assign n5419 = pi16 ? n32 : n5418;
  assign n5420 = pi14 ? n5417 : n5419;
  assign n5421 = pi13 ? n5415 : n5420;
  assign n5422 = pi17 ? n1028 : ~n1933;
  assign n5423 = pi16 ? n32 : n5422;
  assign n5424 = pi15 ? n5419 : n5423;
  assign n5425 = pi17 ? n1028 : ~n2325;
  assign n5426 = pi16 ? n32 : n5425;
  assign n5427 = pi15 ? n4379 : n5426;
  assign n5428 = pi14 ? n5424 : n5427;
  assign n5429 = pi18 ? n32 : ~n5267;
  assign n5430 = pi17 ? n2005 : ~n5429;
  assign n5431 = pi16 ? n32 : n5430;
  assign n5432 = pi17 ? n1028 : ~n2133;
  assign n5433 = pi16 ? n32 : n5432;
  assign n5434 = pi15 ? n5431 : n5433;
  assign n5435 = pi20 ? n246 : n207;
  assign n5436 = pi19 ? n5435 : ~n32;
  assign n5437 = pi18 ? n32 : n5436;
  assign n5438 = pi17 ? n3557 : ~n5437;
  assign n5439 = pi16 ? n32 : n5438;
  assign n5440 = pi17 ? n3557 : ~n1682;
  assign n5441 = pi16 ? n32 : n5440;
  assign n5442 = pi15 ? n5439 : n5441;
  assign n5443 = pi14 ? n5434 : n5442;
  assign n5444 = pi13 ? n5428 : n5443;
  assign n5445 = pi12 ? n5421 : n5444;
  assign n5446 = pi20 ? n653 : n32;
  assign n5447 = pi19 ? n236 : ~n5446;
  assign n5448 = pi18 ? n32 : n5447;
  assign n5449 = pi17 ? n3557 : ~n5448;
  assign n5450 = pi16 ? n32 : n5449;
  assign n5451 = pi15 ? n5441 : n5450;
  assign n5452 = pi17 ? n3719 : ~n2325;
  assign n5453 = pi16 ? n32 : n5452;
  assign n5454 = pi15 ? n5453 : n5060;
  assign n5455 = pi14 ? n5451 : n5454;
  assign n5456 = pi17 ? n3715 : ~n1807;
  assign n5457 = pi16 ? n32 : n5456;
  assign n5458 = pi14 ? n5060 : n5457;
  assign n5459 = pi13 ? n5455 : n5458;
  assign n5460 = pi15 ? n5419 : n5417;
  assign n5461 = pi14 ? n5457 : n5460;
  assign n5462 = pi17 ? n4041 : ~n3093;
  assign n5463 = pi16 ? n32 : n5462;
  assign n5464 = pi15 ? n5419 : n5463;
  assign n5465 = pi17 ? n4041 : ~n1933;
  assign n5466 = pi16 ? n32 : n5465;
  assign n5467 = pi17 ? n1500 : ~n3333;
  assign n5468 = pi16 ? n32 : n5467;
  assign n5469 = pi15 ? n5466 : n5468;
  assign n5470 = pi14 ? n5464 : n5469;
  assign n5471 = pi13 ? n5461 : n5470;
  assign n5472 = pi12 ? n5459 : n5471;
  assign n5473 = pi11 ? n5445 : n5472;
  assign n5474 = pi10 ? n5406 : n5473;
  assign n5475 = pi09 ? n5334 : n5474;
  assign n5476 = pi17 ? n1943 : ~n4966;
  assign n5477 = pi16 ? n32 : n5476;
  assign n5478 = pi15 ? n32 : n5477;
  assign n5479 = pi17 ? n2325 : ~n5324;
  assign n5480 = pi16 ? n32 : n5479;
  assign n5481 = pi17 ? n1682 : ~n1697;
  assign n5482 = pi16 ? n32 : n5481;
  assign n5483 = pi15 ? n5480 : n5482;
  assign n5484 = pi14 ? n5478 : n5483;
  assign n5485 = pi13 ? n32 : n5484;
  assign n5486 = pi12 ? n32 : n5485;
  assign n5487 = pi11 ? n32 : n5486;
  assign n5488 = pi10 ? n32 : n5487;
  assign n5489 = pi17 ? n1322 : ~n5336;
  assign n5490 = pi16 ? n32 : n5489;
  assign n5491 = pi17 ? n1322 : ~n4987;
  assign n5492 = pi16 ? n32 : n5491;
  assign n5493 = pi15 ? n5490 : n5492;
  assign n5494 = pi17 ? n1842 : ~n1697;
  assign n5495 = pi16 ? n32 : n5494;
  assign n5496 = pi17 ? n1478 : ~n4994;
  assign n5497 = pi16 ? n32 : n5496;
  assign n5498 = pi15 ? n5495 : n5497;
  assign n5499 = pi14 ? n5493 : n5498;
  assign n5500 = pi17 ? n1478 : ~n1697;
  assign n5501 = pi16 ? n32 : n5500;
  assign n5502 = pi19 ? n221 : n32;
  assign n5503 = pi18 ? n940 : ~n5502;
  assign n5504 = pi17 ? n1232 : ~n5503;
  assign n5505 = pi16 ? n32 : n5504;
  assign n5506 = pi15 ? n5501 : n5505;
  assign n5507 = pi17 ? n1232 : ~n5358;
  assign n5508 = pi16 ? n32 : n5507;
  assign n5509 = pi17 ? n1966 : ~n5010;
  assign n5510 = pi16 ? n32 : n5509;
  assign n5511 = pi15 ? n5508 : n5510;
  assign n5512 = pi14 ? n5506 : n5511;
  assign n5513 = pi13 ? n5499 : n5512;
  assign n5514 = pi17 ? n4804 : ~n2119;
  assign n5515 = pi16 ? n32 : n5514;
  assign n5516 = pi17 ? n1706 : ~n2531;
  assign n5517 = pi16 ? n32 : n5516;
  assign n5518 = pi15 ? n5515 : n5517;
  assign n5519 = pi17 ? n4656 : ~n5373;
  assign n5520 = pi16 ? n32 : n5519;
  assign n5521 = pi17 ? n4497 : ~n2519;
  assign n5522 = pi16 ? n32 : n5521;
  assign n5523 = pi15 ? n5520 : n5522;
  assign n5524 = pi14 ? n5518 : n5523;
  assign n5525 = pi15 ? n4824 : n5177;
  assign n5526 = pi14 ? n4820 : n5525;
  assign n5527 = pi13 ? n5524 : n5526;
  assign n5528 = pi12 ? n5513 : n5527;
  assign n5529 = pi17 ? n4341 : ~n2653;
  assign n5530 = pi16 ? n32 : n5529;
  assign n5531 = pi15 ? n5530 : n4677;
  assign n5532 = pi17 ? n1989 : ~n2531;
  assign n5533 = pi16 ? n32 : n5532;
  assign n5534 = pi15 ? n4677 : n5533;
  assign n5535 = pi14 ? n5531 : n5534;
  assign n5536 = pi17 ? n2461 : ~n1933;
  assign n5537 = pi16 ? n32 : n5536;
  assign n5538 = pi13 ? n5535 : n5537;
  assign n5539 = pi17 ? n4167 : ~n2653;
  assign n5540 = pi16 ? n32 : n5539;
  assign n5541 = pi18 ? n2413 : ~n32;
  assign n5542 = pi17 ? n5541 : ~n3093;
  assign n5543 = pi16 ? n32 : n5542;
  assign n5544 = pi15 ? n5540 : n5543;
  assign n5545 = pi17 ? n5541 : ~n1933;
  assign n5546 = pi16 ? n32 : n5545;
  assign n5547 = pi17 ? n5541 : ~n1807;
  assign n5548 = pi16 ? n32 : n5547;
  assign n5549 = pi15 ? n5546 : n5548;
  assign n5550 = pi14 ? n5544 : n5549;
  assign n5551 = pi17 ? n5541 : ~n3333;
  assign n5552 = pi16 ? n32 : n5551;
  assign n5553 = pi15 ? n5543 : n5552;
  assign n5554 = pi17 ? n2355 : ~n2537;
  assign n5555 = pi16 ? n32 : n5554;
  assign n5556 = pi15 ? n5555 : n4697;
  assign n5557 = pi14 ? n5553 : n5556;
  assign n5558 = pi13 ? n5550 : n5557;
  assign n5559 = pi12 ? n5538 : n5558;
  assign n5560 = pi11 ? n5528 : n5559;
  assign n5561 = pi17 ? n1120 : ~n2537;
  assign n5562 = pi16 ? n32 : n5561;
  assign n5563 = pi17 ? n4034 : ~n2650;
  assign n5564 = pi16 ? n32 : n5563;
  assign n5565 = pi15 ? n5562 : n5564;
  assign n5566 = pi19 ? n1265 : ~n102;
  assign n5567 = pi18 ? n32 : n5566;
  assign n5568 = pi17 ? n4034 : ~n5567;
  assign n5569 = pi16 ? n32 : n5568;
  assign n5570 = pi15 ? n5569 : n5031;
  assign n5571 = pi14 ? n5565 : n5570;
  assign n5572 = pi19 ? n349 : ~n102;
  assign n5573 = pi18 ? n32 : n5572;
  assign n5574 = pi17 ? n4037 : ~n5573;
  assign n5575 = pi16 ? n32 : n5574;
  assign n5576 = pi15 ? n5575 : n5398;
  assign n5577 = pi14 ? n5576 : n5408;
  assign n5578 = pi13 ? n5571 : n5577;
  assign n5579 = pi17 ? n1726 : ~n1933;
  assign n5580 = pi16 ? n32 : n5579;
  assign n5581 = pi15 ? n5408 : n5580;
  assign n5582 = pi17 ? n1227 : ~n2136;
  assign n5583 = pi16 ? n32 : n5582;
  assign n5584 = pi17 ? n1726 : ~n2136;
  assign n5585 = pi16 ? n32 : n5584;
  assign n5586 = pi15 ? n5583 : n5585;
  assign n5587 = pi14 ? n5581 : n5586;
  assign n5588 = pi19 ? n358 : n87;
  assign n5589 = pi18 ? n32 : ~n5588;
  assign n5590 = pi17 ? n1726 : ~n5589;
  assign n5591 = pi16 ? n32 : n5590;
  assign n5592 = pi17 ? n1726 : ~n2885;
  assign n5593 = pi16 ? n32 : n5592;
  assign n5594 = pi15 ? n5591 : n5593;
  assign n5595 = pi17 ? n3715 : ~n5437;
  assign n5596 = pi16 ? n32 : n5595;
  assign n5597 = pi20 ? n382 : n32;
  assign n5598 = pi19 ? n358 : n5597;
  assign n5599 = pi18 ? n32 : ~n5598;
  assign n5600 = pi17 ? n3704 : ~n5599;
  assign n5601 = pi16 ? n32 : n5600;
  assign n5602 = pi15 ? n5596 : n5601;
  assign n5603 = pi14 ? n5594 : n5602;
  assign n5604 = pi13 ? n5587 : n5603;
  assign n5605 = pi12 ? n5578 : n5604;
  assign n5606 = pi17 ? n3704 : ~n3100;
  assign n5607 = pi16 ? n32 : n5606;
  assign n5608 = pi17 ? n3704 : ~n2314;
  assign n5609 = pi16 ? n32 : n5608;
  assign n5610 = pi15 ? n5607 : n5609;
  assign n5611 = pi17 ? n4041 : ~n2314;
  assign n5612 = pi16 ? n32 : n5611;
  assign n5613 = pi14 ? n5610 : n5612;
  assign n5614 = pi20 ? n274 : n32;
  assign n5615 = pi19 ? n502 : ~n5614;
  assign n5616 = pi18 ? n32 : n5615;
  assign n5617 = pi17 ? n4041 : ~n5616;
  assign n5618 = pi16 ? n32 : n5617;
  assign n5619 = pi15 ? n5618 : n5612;
  assign n5620 = pi17 ? n3553 : ~n3093;
  assign n5621 = pi16 ? n32 : n5620;
  assign n5622 = pi15 ? n5417 : n5621;
  assign n5623 = pi14 ? n5619 : n5622;
  assign n5624 = pi13 ? n5613 : n5623;
  assign n5625 = pi15 ? n5410 : n5621;
  assign n5626 = pi20 ? n481 : n32;
  assign n5627 = pi19 ? n349 : ~n5626;
  assign n5628 = pi18 ? n32 : n5627;
  assign n5629 = pi17 ? n3855 : ~n5628;
  assign n5630 = pi16 ? n32 : n5629;
  assign n5631 = pi17 ? n3855 : ~n2537;
  assign n5632 = pi16 ? n32 : n5631;
  assign n5633 = pi15 ? n5630 : n5632;
  assign n5634 = pi14 ? n5625 : n5633;
  assign n5635 = pi20 ? n125 : n32;
  assign n5636 = pi19 ? n589 : ~n5635;
  assign n5637 = pi18 ? n32 : n5636;
  assign n5638 = pi17 ? n3855 : ~n5637;
  assign n5639 = pi16 ? n32 : n5638;
  assign n5640 = pi15 ? n5639 : n5400;
  assign n5641 = pi17 ? n1605 : ~n2531;
  assign n5642 = pi16 ? n32 : n5641;
  assign n5643 = pi15 ? n5400 : n5642;
  assign n5644 = pi14 ? n5640 : n5643;
  assign n5645 = pi13 ? n5634 : n5644;
  assign n5646 = pi12 ? n5624 : n5645;
  assign n5647 = pi11 ? n5605 : n5646;
  assign n5648 = pi10 ? n5560 : n5647;
  assign n5649 = pi09 ? n5488 : n5648;
  assign n5650 = pi08 ? n5475 : n5649;
  assign n5651 = pi07 ? n5319 : n5650;
  assign n5652 = pi17 ? n3337 : ~n1593;
  assign n5653 = pi16 ? n32 : n5652;
  assign n5654 = pi15 ? n32 : n5653;
  assign n5655 = pi17 ? n1814 : ~n3380;
  assign n5656 = pi16 ? n32 : n5655;
  assign n5657 = pi19 ? n32 : n1757;
  assign n5658 = pi18 ? n5657 : n605;
  assign n5659 = pi17 ? n1814 : ~n5658;
  assign n5660 = pi16 ? n32 : n5659;
  assign n5661 = pi15 ? n5656 : n5660;
  assign n5662 = pi14 ? n5654 : n5661;
  assign n5663 = pi13 ? n32 : n5662;
  assign n5664 = pi12 ? n32 : n5663;
  assign n5665 = pi11 ? n32 : n5664;
  assign n5666 = pi10 ? n32 : n5665;
  assign n5667 = pi19 ? n507 : ~n236;
  assign n5668 = pi18 ? n5667 : ~n32;
  assign n5669 = pi17 ? n1682 : ~n5668;
  assign n5670 = pi16 ? n32 : n5669;
  assign n5671 = pi18 ? n507 : ~n32;
  assign n5672 = pi17 ? n1576 : ~n5671;
  assign n5673 = pi16 ? n32 : n5672;
  assign n5674 = pi15 ? n5670 : n5673;
  assign n5675 = pi20 ? n342 : n266;
  assign n5676 = pi19 ? n5675 : n208;
  assign n5677 = pi18 ? n5676 : ~n32;
  assign n5678 = pi17 ? n2143 : ~n5677;
  assign n5679 = pi16 ? n32 : n5678;
  assign n5680 = pi19 ? n4670 : n531;
  assign n5681 = pi18 ? n5680 : ~n32;
  assign n5682 = pi17 ? n1580 : ~n5681;
  assign n5683 = pi16 ? n32 : n5682;
  assign n5684 = pi15 ? n5679 : n5683;
  assign n5685 = pi14 ? n5674 : n5684;
  assign n5686 = pi17 ? n1593 : ~n1580;
  assign n5687 = pi16 ? n32 : n5686;
  assign n5688 = pi20 ? n266 : n321;
  assign n5689 = pi19 ? n5688 : ~n236;
  assign n5690 = pi18 ? n863 : ~n5689;
  assign n5691 = pi17 ? n1213 : ~n5690;
  assign n5692 = pi16 ? n32 : n5691;
  assign n5693 = pi15 ? n5687 : n5692;
  assign n5694 = pi20 ? n32 : ~n321;
  assign n5695 = pi19 ? n5694 : n208;
  assign n5696 = pi18 ? n5695 : ~n32;
  assign n5697 = pi17 ? n1213 : ~n5696;
  assign n5698 = pi16 ? n32 : n5697;
  assign n5699 = pi18 ? n209 : ~n5657;
  assign n5700 = pi19 ? n4964 : n343;
  assign n5701 = pi18 ? n5700 : ~n32;
  assign n5702 = pi17 ? n5699 : ~n5701;
  assign n5703 = pi16 ? n32 : n5702;
  assign n5704 = pi15 ? n5698 : n5703;
  assign n5705 = pi14 ? n5693 : n5704;
  assign n5706 = pi13 ? n5685 : n5705;
  assign n5707 = pi20 ? n207 : n32;
  assign n5708 = pi19 ? n5707 : n4406;
  assign n5709 = pi18 ? n5708 : ~n32;
  assign n5710 = pi17 ? n1134 : ~n5709;
  assign n5711 = pi16 ? n32 : n5710;
  assign n5712 = pi15 ? n5711 : n5349;
  assign n5713 = pi17 ? n4656 : ~n4984;
  assign n5714 = pi16 ? n32 : n5713;
  assign n5715 = pi19 ? n208 : n32;
  assign n5716 = pi18 ? n32 : ~n5715;
  assign n5717 = pi17 ? n4656 : ~n5716;
  assign n5718 = pi16 ? n32 : n5717;
  assign n5719 = pi15 ? n5714 : n5718;
  assign n5720 = pi14 ? n5712 : n5719;
  assign n5721 = pi19 ? n247 : n343;
  assign n5722 = pi18 ? n5721 : ~n32;
  assign n5723 = pi17 ? n4656 : ~n5722;
  assign n5724 = pi16 ? n32 : n5723;
  assign n5725 = pi19 ? n531 : ~n236;
  assign n5726 = pi18 ? n5725 : n32;
  assign n5727 = pi17 ? n1700 : n5726;
  assign n5728 = pi16 ? n32 : n5727;
  assign n5729 = pi15 ? n5724 : n5728;
  assign n5730 = pi20 ? n32 : ~n518;
  assign n5731 = pi19 ? n5730 : n32;
  assign n5732 = pi18 ? n863 : ~n5731;
  assign n5733 = pi17 ? n4497 : ~n5732;
  assign n5734 = pi16 ? n32 : n5733;
  assign n5735 = pi15 ? n5000 : n5734;
  assign n5736 = pi14 ? n5729 : n5735;
  assign n5737 = pi13 ? n5720 : n5736;
  assign n5738 = pi12 ? n5706 : n5737;
  assign n5739 = pi17 ? n4497 : ~n5358;
  assign n5740 = pi16 ? n32 : n5739;
  assign n5741 = pi20 ? n342 : ~n342;
  assign n5742 = pi19 ? n5741 : n32;
  assign n5743 = pi18 ? n940 : ~n5742;
  assign n5744 = pi17 ? n4497 : ~n5743;
  assign n5745 = pi16 ? n32 : n5744;
  assign n5746 = pi15 ? n5740 : n5745;
  assign n5747 = pi19 ? n349 : ~n349;
  assign n5748 = pi20 ? n342 : ~n207;
  assign n5749 = pi19 ? n5748 : n32;
  assign n5750 = pi18 ? n5747 : n5749;
  assign n5751 = pi17 ? n4497 : n5750;
  assign n5752 = pi16 ? n32 : n5751;
  assign n5753 = pi18 ? n5747 : n4671;
  assign n5754 = pi17 ? n1472 : n5753;
  assign n5755 = pi16 ? n32 : n5754;
  assign n5756 = pi15 ? n5752 : n5755;
  assign n5757 = pi14 ? n5746 : n5756;
  assign n5758 = pi18 ? n940 : ~n5009;
  assign n5759 = pi17 ? n1480 : ~n5758;
  assign n5760 = pi16 ? n32 : n5759;
  assign n5761 = pi17 ? n1480 : ~n5358;
  assign n5762 = pi16 ? n32 : n5761;
  assign n5763 = pi14 ? n5760 : n5762;
  assign n5764 = pi13 ? n5757 : n5763;
  assign n5765 = pi18 ? n2747 : ~n32;
  assign n5766 = pi18 ? n940 : n323;
  assign n5767 = pi17 ? n5765 : ~n5766;
  assign n5768 = pi16 ? n32 : n5767;
  assign n5769 = pi15 ? n5008 : n5768;
  assign n5770 = pi17 ? n5765 : ~n2531;
  assign n5771 = pi16 ? n32 : n5770;
  assign n5772 = pi17 ? n5765 : ~n2519;
  assign n5773 = pi16 ? n32 : n5772;
  assign n5774 = pi15 ? n5771 : n5773;
  assign n5775 = pi14 ? n5769 : n5774;
  assign n5776 = pi17 ? n5765 : ~n2119;
  assign n5777 = pi16 ? n32 : n5776;
  assign n5778 = pi19 ? n4126 : ~n32;
  assign n5779 = pi18 ? n32 : n5778;
  assign n5780 = pi17 ? n5765 : ~n5779;
  assign n5781 = pi16 ? n32 : n5780;
  assign n5782 = pi15 ? n5777 : n5781;
  assign n5783 = pi17 ? n4515 : ~n2531;
  assign n5784 = pi16 ? n32 : n5783;
  assign n5785 = pi17 ? n4515 : ~n2119;
  assign n5786 = pi16 ? n32 : n5785;
  assign n5787 = pi15 ? n5784 : n5786;
  assign n5788 = pi14 ? n5782 : n5787;
  assign n5789 = pi13 ? n5775 : n5788;
  assign n5790 = pi12 ? n5764 : n5789;
  assign n5791 = pi11 ? n5738 : n5790;
  assign n5792 = pi17 ? n2465 : ~n2531;
  assign n5793 = pi16 ? n32 : n5792;
  assign n5794 = pi15 ? n5786 : n5793;
  assign n5795 = pi14 ? n5786 : n5794;
  assign n5796 = pi17 ? n2355 : ~n2119;
  assign n5797 = pi16 ? n32 : n5796;
  assign n5798 = pi17 ? n4023 : ~n2119;
  assign n5799 = pi16 ? n32 : n5798;
  assign n5800 = pi14 ? n5797 : n5799;
  assign n5801 = pi13 ? n5795 : n5800;
  assign n5802 = pi17 ? n4023 : ~n2519;
  assign n5803 = pi16 ? n32 : n5802;
  assign n5804 = pi17 ? n1219 : ~n2519;
  assign n5805 = pi16 ? n32 : n5804;
  assign n5806 = pi15 ? n5803 : n5805;
  assign n5807 = pi17 ? n1120 : ~n2519;
  assign n5808 = pi16 ? n32 : n5807;
  assign n5809 = pi15 ? n5808 : n5805;
  assign n5810 = pi14 ? n5806 : n5809;
  assign n5811 = pi17 ? n1227 : ~n2519;
  assign n5812 = pi16 ? n32 : n5811;
  assign n5813 = pi17 ? n3855 : ~n2512;
  assign n5814 = pi16 ? n32 : n5813;
  assign n5815 = pi15 ? n5812 : n5814;
  assign n5816 = pi14 ? n5805 : n5815;
  assign n5817 = pi13 ? n5810 : n5816;
  assign n5818 = pi12 ? n5801 : n5817;
  assign n5819 = pi17 ? n4037 : ~n2512;
  assign n5820 = pi16 ? n32 : n5819;
  assign n5821 = pi14 ? n5814 : n5820;
  assign n5822 = pi17 ? n4034 : ~n2512;
  assign n5823 = pi16 ? n32 : n5822;
  assign n5824 = pi15 ? n5820 : n5823;
  assign n5825 = pi14 ? n5820 : n5824;
  assign n5826 = pi13 ? n5821 : n5825;
  assign n5827 = pi17 ? n4034 : ~n2750;
  assign n5828 = pi16 ? n32 : n5827;
  assign n5829 = pi19 ? n176 : ~n32;
  assign n5830 = pi18 ? n32 : n5829;
  assign n5831 = pi17 ? n4034 : ~n5830;
  assign n5832 = pi16 ? n32 : n5831;
  assign n5833 = pi15 ? n5828 : n5832;
  assign n5834 = pi17 ? n4023 : ~n2750;
  assign n5835 = pi16 ? n32 : n5834;
  assign n5836 = pi14 ? n5833 : n5835;
  assign n5837 = pi17 ? n5541 : ~n2623;
  assign n5838 = pi16 ? n32 : n5837;
  assign n5839 = pi15 ? n5835 : n5838;
  assign n5840 = pi17 ? n5541 : ~n2512;
  assign n5841 = pi16 ? n32 : n5840;
  assign n5842 = pi17 ? n2355 : ~n2512;
  assign n5843 = pi16 ? n32 : n5842;
  assign n5844 = pi15 ? n5841 : n5843;
  assign n5845 = pi14 ? n5839 : n5844;
  assign n5846 = pi13 ? n5836 : n5845;
  assign n5847 = pi12 ? n5826 : n5846;
  assign n5848 = pi11 ? n5818 : n5847;
  assign n5849 = pi10 ? n5791 : n5848;
  assign n5850 = pi09 ? n5666 : n5849;
  assign n5851 = pi17 ? n2305 : ~n1580;
  assign n5852 = pi16 ? n32 : n5851;
  assign n5853 = pi15 ? n32 : n5852;
  assign n5854 = pi21 ? n174 : ~n206;
  assign n5855 = pi20 ? n5854 : n32;
  assign n5856 = pi19 ? n5855 : n32;
  assign n5857 = pi18 ? n940 : ~n5856;
  assign n5858 = pi17 ? n1933 : ~n5857;
  assign n5859 = pi16 ? n32 : n5858;
  assign n5860 = pi15 ? n5859 : n5660;
  assign n5861 = pi14 ? n5853 : n5860;
  assign n5862 = pi13 ? n32 : n5861;
  assign n5863 = pi12 ? n32 : n5862;
  assign n5864 = pi11 ? n32 : n5863;
  assign n5865 = pi10 ? n32 : n5864;
  assign n5866 = pi17 ? n1814 : ~n5668;
  assign n5867 = pi16 ? n32 : n5866;
  assign n5868 = pi17 ? n2136 : ~n5671;
  assign n5869 = pi16 ? n32 : n5868;
  assign n5870 = pi15 ? n5867 : n5869;
  assign n5871 = pi17 ? n2325 : ~n5677;
  assign n5872 = pi16 ? n32 : n5871;
  assign n5873 = pi19 ? n176 : n340;
  assign n5874 = pi18 ? n5873 : ~n32;
  assign n5875 = pi17 ? n3351 : ~n5874;
  assign n5876 = pi16 ? n32 : n5875;
  assign n5877 = pi15 ? n5872 : n5876;
  assign n5878 = pi14 ? n5870 : n5877;
  assign n5879 = pi17 ? n1576 : ~n1580;
  assign n5880 = pi16 ? n32 : n5879;
  assign n5881 = pi18 ? n858 : ~n5689;
  assign n5882 = pi17 ? n1593 : ~n5881;
  assign n5883 = pi16 ? n32 : n5882;
  assign n5884 = pi15 ? n5880 : n5883;
  assign n5885 = pi17 ? n1593 : ~n5696;
  assign n5886 = pi16 ? n32 : n5885;
  assign n5887 = pi18 ? n1841 : ~n5657;
  assign n5888 = pi17 ? n5887 : ~n5701;
  assign n5889 = pi16 ? n32 : n5888;
  assign n5890 = pi15 ? n5886 : n5889;
  assign n5891 = pi14 ? n5884 : n5890;
  assign n5892 = pi13 ? n5878 : n5891;
  assign n5893 = pi17 ? n1478 : ~n5709;
  assign n5894 = pi16 ? n32 : n5893;
  assign n5895 = pi15 ? n5894 : n5501;
  assign n5896 = pi17 ? n1232 : ~n4984;
  assign n5897 = pi16 ? n32 : n5896;
  assign n5898 = pi17 ? n1232 : ~n5716;
  assign n5899 = pi16 ? n32 : n5898;
  assign n5900 = pi15 ? n5897 : n5899;
  assign n5901 = pi14 ? n5895 : n5900;
  assign n5902 = pi17 ? n1966 : ~n5722;
  assign n5903 = pi16 ? n32 : n5902;
  assign n5904 = pi17 ? n4804 : n5726;
  assign n5905 = pi16 ? n32 : n5904;
  assign n5906 = pi15 ? n5903 : n5905;
  assign n5907 = pi17 ? n4656 : ~n5732;
  assign n5908 = pi16 ? n32 : n5907;
  assign n5909 = pi15 ? n5157 : n5908;
  assign n5910 = pi14 ? n5906 : n5909;
  assign n5911 = pi13 ? n5901 : n5910;
  assign n5912 = pi12 ? n5892 : n5911;
  assign n5913 = pi17 ? n4656 : ~n5743;
  assign n5914 = pi16 ? n32 : n5913;
  assign n5915 = pi15 ? n5360 : n5914;
  assign n5916 = pi17 ? n4656 : n5750;
  assign n5917 = pi16 ? n32 : n5916;
  assign n5918 = pi17 ? n4659 : n5753;
  assign n5919 = pi16 ? n32 : n5918;
  assign n5920 = pi15 ? n5917 : n5919;
  assign n5921 = pi14 ? n5915 : n5920;
  assign n5922 = pi17 ? n2159 : ~n5758;
  assign n5923 = pi16 ? n32 : n5922;
  assign n5924 = pi17 ? n2159 : ~n5358;
  assign n5925 = pi16 ? n32 : n5924;
  assign n5926 = pi14 ? n5923 : n5925;
  assign n5927 = pi13 ? n5921 : n5926;
  assign n5928 = pi17 ? n4497 : ~n5006;
  assign n5929 = pi16 ? n32 : n5928;
  assign n5930 = pi18 ? n2622 : ~n32;
  assign n5931 = pi17 ? n5930 : ~n5766;
  assign n5932 = pi16 ? n32 : n5931;
  assign n5933 = pi15 ? n5929 : n5932;
  assign n5934 = pi17 ? n5930 : ~n2644;
  assign n5935 = pi16 ? n32 : n5934;
  assign n5936 = pi17 ? n5930 : ~n2519;
  assign n5937 = pi16 ? n32 : n5936;
  assign n5938 = pi15 ? n5935 : n5937;
  assign n5939 = pi14 ? n5933 : n5938;
  assign n5940 = pi17 ? n5930 : ~n2119;
  assign n5941 = pi16 ? n32 : n5940;
  assign n5942 = pi17 ? n5930 : ~n5779;
  assign n5943 = pi16 ? n32 : n5942;
  assign n5944 = pi15 ? n5941 : n5943;
  assign n5945 = pi18 ? n32 : n1914;
  assign n5946 = pi17 ? n4682 : ~n5945;
  assign n5947 = pi16 ? n32 : n5946;
  assign n5948 = pi17 ? n4682 : ~n2119;
  assign n5949 = pi16 ? n32 : n5948;
  assign n5950 = pi15 ? n5947 : n5949;
  assign n5951 = pi14 ? n5944 : n5950;
  assign n5952 = pi13 ? n5939 : n5951;
  assign n5953 = pi12 ? n5927 : n5952;
  assign n5954 = pi11 ? n5912 : n5953;
  assign n5955 = pi17 ? n4682 : ~n2408;
  assign n5956 = pi16 ? n32 : n5955;
  assign n5957 = pi15 ? n5956 : n5183;
  assign n5958 = pi14 ? n5956 : n5957;
  assign n5959 = pi13 ? n5958 : n5385;
  assign n5960 = pi17 ? n4167 : ~n2519;
  assign n5961 = pi16 ? n32 : n5960;
  assign n5962 = pi17 ? n2465 : ~n2519;
  assign n5963 = pi16 ? n32 : n5962;
  assign n5964 = pi15 ? n5961 : n5963;
  assign n5965 = pi17 ? n4515 : ~n2519;
  assign n5966 = pi16 ? n32 : n5965;
  assign n5967 = pi15 ? n5966 : n5963;
  assign n5968 = pi14 ? n5964 : n5967;
  assign n5969 = pi17 ? n1120 : ~n2512;
  assign n5970 = pi16 ? n32 : n5969;
  assign n5971 = pi15 ? n5808 : n5970;
  assign n5972 = pi14 ? n5963 : n5971;
  assign n5973 = pi13 ? n5968 : n5972;
  assign n5974 = pi12 ? n5959 : n5973;
  assign n5975 = pi17 ? n4023 : ~n2512;
  assign n5976 = pi16 ? n32 : n5975;
  assign n5977 = pi19 ? n507 : ~n5635;
  assign n5978 = pi18 ? n32 : n5977;
  assign n5979 = pi17 ? n4023 : ~n5978;
  assign n5980 = pi16 ? n32 : n5979;
  assign n5981 = pi15 ? n5976 : n5980;
  assign n5982 = pi14 ? n5981 : n5841;
  assign n5983 = pi19 ? n507 : ~n358;
  assign n5984 = pi18 ? n32 : n5983;
  assign n5985 = pi17 ? n5541 : ~n5984;
  assign n5986 = pi16 ? n32 : n5985;
  assign n5987 = pi15 ? n5841 : n5986;
  assign n5988 = pi17 ? n2465 : ~n2512;
  assign n5989 = pi16 ? n32 : n5988;
  assign n5990 = pi15 ? n5841 : n5989;
  assign n5991 = pi14 ? n5987 : n5990;
  assign n5992 = pi13 ? n5982 : n5991;
  assign n5993 = pi17 ? n4515 : ~n2750;
  assign n5994 = pi16 ? n32 : n5993;
  assign n5995 = pi17 ? n4515 : ~n5830;
  assign n5996 = pi16 ? n32 : n5995;
  assign n5997 = pi15 ? n5994 : n5996;
  assign n5998 = pi17 ? n4167 : ~n2750;
  assign n5999 = pi16 ? n32 : n5998;
  assign n6000 = pi14 ? n5997 : n5999;
  assign n6001 = pi17 ? n4167 : ~n2623;
  assign n6002 = pi16 ? n32 : n6001;
  assign n6003 = pi17 ? n2461 : ~n2623;
  assign n6004 = pi16 ? n32 : n6003;
  assign n6005 = pi15 ? n6002 : n6004;
  assign n6006 = pi17 ? n5765 : ~n2512;
  assign n6007 = pi16 ? n32 : n6006;
  assign n6008 = pi17 ? n2461 : ~n2512;
  assign n6009 = pi16 ? n32 : n6008;
  assign n6010 = pi15 ? n6007 : n6009;
  assign n6011 = pi14 ? n6005 : n6010;
  assign n6012 = pi13 ? n6000 : n6011;
  assign n6013 = pi12 ? n5992 : n6012;
  assign n6014 = pi11 ? n5974 : n6013;
  assign n6015 = pi10 ? n5954 : n6014;
  assign n6016 = pi09 ? n5865 : n6015;
  assign n6017 = pi08 ? n5850 : n6016;
  assign n6018 = pi20 ? n220 : n207;
  assign n6019 = pi19 ? n6018 : ~n32;
  assign n6020 = pi18 ? n32 : n6019;
  assign n6021 = pi17 ? n2531 : ~n6020;
  assign n6022 = pi16 ? n32 : n6021;
  assign n6023 = pi15 ? n32 : n6022;
  assign n6024 = pi17 ? n1933 : ~n2119;
  assign n6025 = pi16 ? n32 : n6024;
  assign n6026 = pi21 ? n173 : n313;
  assign n6027 = pi20 ? n6026 : ~n32;
  assign n6028 = pi19 ? n32 : ~n6027;
  assign n6029 = pi20 ? n501 : ~n207;
  assign n6030 = pi19 ? n6029 : n32;
  assign n6031 = pi18 ? n6028 : ~n6030;
  assign n6032 = pi17 ? n1933 : ~n6031;
  assign n6033 = pi16 ? n32 : n6032;
  assign n6034 = pi15 ? n6025 : n6033;
  assign n6035 = pi14 ? n6023 : n6034;
  assign n6036 = pi13 ? n32 : n6035;
  assign n6037 = pi12 ? n32 : n6036;
  assign n6038 = pi11 ? n32 : n6037;
  assign n6039 = pi10 ? n32 : n6038;
  assign n6040 = pi19 ? n2317 : ~n1818;
  assign n6041 = pi18 ? n32 : n6040;
  assign n6042 = pi20 ? n1324 : ~n32;
  assign n6043 = pi19 ? n507 : ~n6042;
  assign n6044 = pi18 ? n6043 : ~n32;
  assign n6045 = pi17 ? n6041 : ~n6044;
  assign n6046 = pi16 ? n32 : n6045;
  assign n6047 = pi19 ? n589 : ~n275;
  assign n6048 = pi18 ? n32 : n6047;
  assign n6049 = pi20 ? n357 : n342;
  assign n6050 = pi21 ? n206 : ~n174;
  assign n6051 = pi20 ? n6050 : ~n342;
  assign n6052 = pi19 ? n6049 : ~n6051;
  assign n6053 = pi18 ? n6052 : ~n32;
  assign n6054 = pi17 ? n6048 : ~n6053;
  assign n6055 = pi16 ? n32 : n6054;
  assign n6056 = pi15 ? n6046 : n6055;
  assign n6057 = pi20 ? n32 : n1331;
  assign n6058 = pi19 ? n6057 : n1165;
  assign n6059 = pi19 ? n1757 : n32;
  assign n6060 = pi18 ? n6058 : ~n6059;
  assign n6061 = pi17 ? n1807 : ~n6060;
  assign n6062 = pi16 ? n32 : n6061;
  assign n6063 = pi19 ? n1740 : ~n32;
  assign n6064 = pi18 ? n4380 : n6063;
  assign n6065 = pi17 ? n2136 : ~n6064;
  assign n6066 = pi16 ? n32 : n6065;
  assign n6067 = pi15 ? n6062 : n6066;
  assign n6068 = pi14 ? n6056 : n6067;
  assign n6069 = pi17 ? n2136 : ~n1933;
  assign n6070 = pi16 ? n32 : n6069;
  assign n6071 = pi19 ? n32 : n4491;
  assign n6072 = pi18 ? n1575 : ~n6071;
  assign n6073 = pi20 ? n32 : n3847;
  assign n6074 = pi20 ? n357 : n1368;
  assign n6075 = pi19 ? n6073 : n6074;
  assign n6076 = pi18 ? n6075 : n350;
  assign n6077 = pi17 ? n6072 : ~n6076;
  assign n6078 = pi16 ? n32 : n6077;
  assign n6079 = pi15 ? n6070 : n6078;
  assign n6080 = pi17 ? n1833 : ~n5696;
  assign n6081 = pi16 ? n32 : n6080;
  assign n6082 = pi20 ? n623 : n1331;
  assign n6083 = pi19 ? n32 : n6082;
  assign n6084 = pi18 ? n2142 : ~n6083;
  assign n6085 = pi21 ? n309 : n174;
  assign n6086 = pi20 ? n6085 : ~n32;
  assign n6087 = pi19 ? n4964 : n6086;
  assign n6088 = pi18 ? n6087 : ~n32;
  assign n6089 = pi17 ? n6084 : ~n6088;
  assign n6090 = pi16 ? n32 : n6089;
  assign n6091 = pi15 ? n6081 : n6090;
  assign n6092 = pi14 ? n6079 : n6091;
  assign n6093 = pi13 ? n6068 : n6092;
  assign n6094 = pi19 ? n4342 : n343;
  assign n6095 = pi18 ? n6094 : ~n32;
  assign n6096 = pi17 ? n1580 : ~n6095;
  assign n6097 = pi16 ? n32 : n6096;
  assign n6098 = pi18 ? n1509 : ~n5667;
  assign n6099 = pi17 ? n1593 : ~n6098;
  assign n6100 = pi16 ? n32 : n6099;
  assign n6101 = pi15 ? n6097 : n6100;
  assign n6102 = pi18 ? n32 : ~n5725;
  assign n6103 = pi17 ? n1213 : ~n6102;
  assign n6104 = pi16 ? n32 : n6103;
  assign n6105 = pi20 ? n428 : n448;
  assign n6106 = pi20 ? n175 : ~n339;
  assign n6107 = pi19 ? n6105 : n6106;
  assign n6108 = pi19 ? n519 : ~n236;
  assign n6109 = pi18 ? n6107 : ~n6108;
  assign n6110 = pi17 ? n1213 : ~n6109;
  assign n6111 = pi16 ? n32 : n6110;
  assign n6112 = pi15 ? n6104 : n6111;
  assign n6113 = pi14 ? n6101 : n6112;
  assign n6114 = pi19 ? n32 : n358;
  assign n6115 = pi18 ? n209 : ~n6114;
  assign n6116 = pi17 ? n6115 : ~n6095;
  assign n6117 = pi16 ? n32 : n6116;
  assign n6118 = pi19 ? n594 : n32;
  assign n6119 = pi18 ? n341 : ~n6118;
  assign n6120 = pi20 ? n339 : ~n207;
  assign n6121 = pi19 ? n6120 : n502;
  assign n6122 = pi18 ? n6121 : ~n32;
  assign n6123 = pi17 ? n6119 : ~n6122;
  assign n6124 = pi16 ? n32 : n6123;
  assign n6125 = pi15 ? n6117 : n6124;
  assign n6126 = pi17 ? n1232 : ~n5336;
  assign n6127 = pi16 ? n32 : n6126;
  assign n6128 = pi15 ? n5349 : n6127;
  assign n6129 = pi14 ? n6125 : n6128;
  assign n6130 = pi13 ? n6113 : n6129;
  assign n6131 = pi12 ? n6093 : n6130;
  assign n6132 = pi19 ? n349 : ~n236;
  assign n6133 = pi18 ? n32 : ~n6132;
  assign n6134 = pi17 ? n1232 : ~n6133;
  assign n6135 = pi16 ? n32 : n6134;
  assign n6136 = pi20 ? n765 : n32;
  assign n6137 = pi20 ? n1368 : n321;
  assign n6138 = pi19 ? n6136 : n6137;
  assign n6139 = pi20 ? n32 : n5854;
  assign n6140 = pi19 ? n6139 : n32;
  assign n6141 = pi18 ? n6138 : ~n6140;
  assign n6142 = pi17 ? n1966 : ~n6141;
  assign n6143 = pi16 ? n32 : n6142;
  assign n6144 = pi15 ? n6135 : n6143;
  assign n6145 = pi19 ? n507 : n32;
  assign n6146 = pi18 ? n1965 : ~n6145;
  assign n6147 = pi19 ? n208 : ~n617;
  assign n6148 = pi18 ? n6147 : n32;
  assign n6149 = pi17 ? n6146 : n6148;
  assign n6150 = pi16 ? n32 : n6149;
  assign n6151 = pi18 ? n2830 : ~n936;
  assign n6152 = pi19 ? n1885 : n349;
  assign n6153 = pi18 ? n6152 : ~n32;
  assign n6154 = pi17 ? n6151 : ~n6153;
  assign n6155 = pi16 ? n32 : n6154;
  assign n6156 = pi15 ? n6150 : n6155;
  assign n6157 = pi14 ? n6144 : n6156;
  assign n6158 = pi20 ? n321 : ~n428;
  assign n6159 = pi19 ? n6158 : n32;
  assign n6160 = pi18 ? n940 : ~n6159;
  assign n6161 = pi17 ? n1706 : ~n6160;
  assign n6162 = pi16 ? n32 : n6161;
  assign n6163 = pi19 ? n349 : n32;
  assign n6164 = pi18 ? n940 : ~n6163;
  assign n6165 = pi17 ? n1706 : ~n6164;
  assign n6166 = pi16 ? n32 : n6165;
  assign n6167 = pi15 ? n6162 : n6166;
  assign n6168 = pi18 ? n32 : ~n6163;
  assign n6169 = pi17 ? n1706 : ~n6168;
  assign n6170 = pi16 ? n32 : n6169;
  assign n6171 = pi20 ? n1324 : n32;
  assign n6172 = pi19 ? n6171 : ~n502;
  assign n6173 = pi20 ? n321 : n220;
  assign n6174 = pi19 ? n6173 : n32;
  assign n6175 = pi18 ? n6172 : ~n6174;
  assign n6176 = pi17 ? n1706 : ~n6175;
  assign n6177 = pi16 ? n32 : n6176;
  assign n6178 = pi15 ? n6170 : n6177;
  assign n6179 = pi14 ? n6167 : n6178;
  assign n6180 = pi13 ? n6157 : n6179;
  assign n6181 = pi19 ? n349 : ~n531;
  assign n6182 = pi18 ? n6181 : n32;
  assign n6183 = pi17 ? n1978 : n6182;
  assign n6184 = pi16 ? n32 : n6183;
  assign n6185 = pi18 ? n940 : ~n5357;
  assign n6186 = pi17 ? n4659 : ~n6185;
  assign n6187 = pi16 ? n32 : n6186;
  assign n6188 = pi15 ? n6184 : n6187;
  assign n6189 = pi17 ? n4659 : ~n2512;
  assign n6190 = pi16 ? n32 : n6189;
  assign n6191 = pi14 ? n6188 : n6190;
  assign n6192 = pi17 ? n4822 : ~n2512;
  assign n6193 = pi16 ? n32 : n6192;
  assign n6194 = pi14 ? n6190 : n6193;
  assign n6195 = pi13 ? n6191 : n6194;
  assign n6196 = pi12 ? n6180 : n6195;
  assign n6197 = pi11 ? n6131 : n6196;
  assign n6198 = pi15 ? n6193 : n5377;
  assign n6199 = pi14 ? n6193 : n6198;
  assign n6200 = pi17 ? n4341 : ~n2512;
  assign n6201 = pi16 ? n32 : n6200;
  assign n6202 = pi15 ? n5377 : n6201;
  assign n6203 = pi14 ? n6202 : n6201;
  assign n6204 = pi13 ? n6199 : n6203;
  assign n6205 = pi17 ? n1718 : ~n2512;
  assign n6206 = pi16 ? n32 : n6205;
  assign n6207 = pi15 ? n6206 : n6007;
  assign n6208 = pi17 ? n1718 : ~n2750;
  assign n6209 = pi16 ? n32 : n6208;
  assign n6210 = pi15 ? n6209 : n5773;
  assign n6211 = pi14 ? n6207 : n6210;
  assign n6212 = pi17 ? n1718 : ~n2519;
  assign n6213 = pi16 ? n32 : n6212;
  assign n6214 = pi17 ? n1215 : ~n2519;
  assign n6215 = pi16 ? n32 : n6214;
  assign n6216 = pi17 ? n4167 : ~n2512;
  assign n6217 = pi16 ? n32 : n6216;
  assign n6218 = pi15 ? n6215 : n6217;
  assign n6219 = pi14 ? n6213 : n6218;
  assign n6220 = pi13 ? n6211 : n6219;
  assign n6221 = pi12 ? n6204 : n6220;
  assign n6222 = pi19 ? n507 : ~n161;
  assign n6223 = pi18 ? n32 : n6222;
  assign n6224 = pi17 ? n4167 : ~n6223;
  assign n6225 = pi16 ? n32 : n6224;
  assign n6226 = pi15 ? n6217 : n6225;
  assign n6227 = pi15 ? n6009 : n6007;
  assign n6228 = pi14 ? n6226 : n6227;
  assign n6229 = pi21 ? n2076 : n32;
  assign n6230 = pi20 ? n6229 : n32;
  assign n6231 = pi19 ? n507 : ~n6230;
  assign n6232 = pi18 ? n32 : n6231;
  assign n6233 = pi17 ? n5765 : ~n6232;
  assign n6234 = pi16 ? n32 : n6233;
  assign n6235 = pi19 ? n507 : n236;
  assign n6236 = pi18 ? n32 : n6235;
  assign n6237 = pi17 ? n5765 : ~n6236;
  assign n6238 = pi16 ? n32 : n6237;
  assign n6239 = pi15 ? n6234 : n6238;
  assign n6240 = pi19 ? n507 : ~n53;
  assign n6241 = pi18 ? n32 : n6240;
  assign n6242 = pi17 ? n4682 : ~n6241;
  assign n6243 = pi16 ? n32 : n6242;
  assign n6244 = pi15 ? n6007 : n6243;
  assign n6245 = pi14 ? n6239 : n6244;
  assign n6246 = pi13 ? n6228 : n6245;
  assign n6247 = pi17 ? n4682 : ~n2750;
  assign n6248 = pi16 ? n32 : n6247;
  assign n6249 = pi19 ? n6057 : n617;
  assign n6250 = pi18 ? n32 : n6249;
  assign n6251 = pi17 ? n4682 : ~n6250;
  assign n6252 = pi16 ? n32 : n6251;
  assign n6253 = pi15 ? n6248 : n6252;
  assign n6254 = pi17 ? n1989 : ~n2750;
  assign n6255 = pi16 ? n32 : n6254;
  assign n6256 = pi17 ? n4341 : ~n2855;
  assign n6257 = pi16 ? n32 : n6256;
  assign n6258 = pi15 ? n6255 : n6257;
  assign n6259 = pi14 ? n6253 : n6258;
  assign n6260 = pi17 ? n4341 : ~n2623;
  assign n6261 = pi16 ? n32 : n6260;
  assign n6262 = pi17 ? n5930 : ~n2623;
  assign n6263 = pi16 ? n32 : n6262;
  assign n6264 = pi15 ? n6261 : n6263;
  assign n6265 = pi17 ? n5930 : ~n2618;
  assign n6266 = pi16 ? n32 : n6265;
  assign n6267 = pi17 ? n1480 : ~n3621;
  assign n6268 = pi16 ? n32 : n6267;
  assign n6269 = pi15 ? n6266 : n6268;
  assign n6270 = pi14 ? n6264 : n6269;
  assign n6271 = pi13 ? n6259 : n6270;
  assign n6272 = pi12 ? n6246 : n6271;
  assign n6273 = pi11 ? n6221 : n6272;
  assign n6274 = pi10 ? n6197 : n6273;
  assign n6275 = pi09 ? n6039 : n6274;
  assign n6276 = pi17 ? n2408 : ~n6020;
  assign n6277 = pi16 ? n32 : n6276;
  assign n6278 = pi15 ? n32 : n6277;
  assign n6279 = pi17 ? n2531 : ~n2119;
  assign n6280 = pi16 ? n32 : n6279;
  assign n6281 = pi20 ? n246 : n1817;
  assign n6282 = pi19 ? n531 : ~n6281;
  assign n6283 = pi18 ? n32 : n6282;
  assign n6284 = pi20 ? n3843 : n820;
  assign n6285 = pi19 ? n275 : ~n6284;
  assign n6286 = pi18 ? n6285 : ~n5749;
  assign n6287 = pi17 ? n6283 : ~n6286;
  assign n6288 = pi16 ? n32 : n6287;
  assign n6289 = pi15 ? n6280 : n6288;
  assign n6290 = pi14 ? n6278 : n6289;
  assign n6291 = pi13 ? n32 : n6290;
  assign n6292 = pi12 ? n32 : n6291;
  assign n6293 = pi11 ? n32 : n6292;
  assign n6294 = pi10 ? n32 : n6293;
  assign n6295 = pi20 ? n3523 : n1817;
  assign n6296 = pi19 ? n2297 : ~n6295;
  assign n6297 = pi18 ? n32 : n6296;
  assign n6298 = pi20 ? n246 : ~n32;
  assign n6299 = pi19 ? n507 : ~n6298;
  assign n6300 = pi18 ? n6299 : ~n32;
  assign n6301 = pi17 ? n6297 : ~n6300;
  assign n6302 = pi16 ? n32 : n6301;
  assign n6303 = pi21 ? n174 : ~n259;
  assign n6304 = pi20 ? n6303 : n266;
  assign n6305 = pi19 ? n429 : ~n6304;
  assign n6306 = pi18 ? n32 : n6305;
  assign n6307 = pi20 ? n207 : ~n342;
  assign n6308 = pi20 ? n220 : ~n342;
  assign n6309 = pi19 ? n6307 : n6308;
  assign n6310 = pi18 ? n6309 : n32;
  assign n6311 = pi17 ? n6306 : n6310;
  assign n6312 = pi16 ? n32 : n6311;
  assign n6313 = pi15 ? n6302 : n6312;
  assign n6314 = pi20 ? n310 : n32;
  assign n6315 = pi19 ? n6314 : n32;
  assign n6316 = pi18 ? n863 : ~n6315;
  assign n6317 = pi17 ? n1933 : ~n6316;
  assign n6318 = pi16 ? n32 : n6317;
  assign n6319 = pi17 ? n2319 : ~n6064;
  assign n6320 = pi16 ? n32 : n6319;
  assign n6321 = pi15 ? n6318 : n6320;
  assign n6322 = pi14 ? n6313 : n6321;
  assign n6323 = pi20 ? n749 : ~n428;
  assign n6324 = pi20 ? n2140 : n32;
  assign n6325 = pi19 ? n6323 : ~n6324;
  assign n6326 = pi18 ? n32 : n6325;
  assign n6327 = pi20 ? n274 : n207;
  assign n6328 = pi19 ? n6327 : ~n5163;
  assign n6329 = pi18 ? n6328 : n350;
  assign n6330 = pi17 ? n6326 : ~n6329;
  assign n6331 = pi16 ? n32 : n6330;
  assign n6332 = pi15 ? n6070 : n6331;
  assign n6333 = pi20 ? n1940 : ~n175;
  assign n6334 = pi19 ? n6333 : ~n32;
  assign n6335 = pi18 ? n32 : n6334;
  assign n6336 = pi17 ? n6335 : ~n5696;
  assign n6337 = pi16 ? n32 : n6336;
  assign n6338 = pi20 ? n207 : ~n1368;
  assign n6339 = pi20 ? n220 : n266;
  assign n6340 = pi19 ? n6338 : ~n6339;
  assign n6341 = pi18 ? n32 : n6340;
  assign n6342 = pi20 ? n6050 : n32;
  assign n6343 = pi19 ? n4964 : ~n6342;
  assign n6344 = pi18 ? n6343 : ~n32;
  assign n6345 = pi17 ? n6341 : ~n6344;
  assign n6346 = pi16 ? n32 : n6345;
  assign n6347 = pi15 ? n6337 : n6346;
  assign n6348 = pi14 ? n6332 : n6347;
  assign n6349 = pi13 ? n6322 : n6348;
  assign n6350 = pi20 ? n1076 : n32;
  assign n6351 = pi19 ? n6350 : n429;
  assign n6352 = pi18 ? n6351 : ~n32;
  assign n6353 = pi17 ? n3351 : ~n6352;
  assign n6354 = pi16 ? n32 : n6353;
  assign n6355 = pi20 ? n32 : ~n6050;
  assign n6356 = pi19 ? n32 : n6355;
  assign n6357 = pi18 ? n6356 : ~n5667;
  assign n6358 = pi17 ? n1576 : ~n6357;
  assign n6359 = pi16 ? n32 : n6358;
  assign n6360 = pi15 ? n6354 : n6359;
  assign n6361 = pi17 ? n1593 : ~n6102;
  assign n6362 = pi16 ? n32 : n6361;
  assign n6363 = pi19 ? n5741 : n5748;
  assign n6364 = pi18 ? n6363 : ~n5667;
  assign n6365 = pi17 ? n1593 : ~n6364;
  assign n6366 = pi16 ? n32 : n6365;
  assign n6367 = pi15 ? n6362 : n6366;
  assign n6368 = pi14 ? n6360 : n6367;
  assign n6369 = pi18 ? n1841 : ~n6114;
  assign n6370 = pi17 ? n6369 : ~n6095;
  assign n6371 = pi16 ? n32 : n6370;
  assign n6372 = pi20 ? n314 : ~n207;
  assign n6373 = pi19 ? n6372 : n589;
  assign n6374 = pi18 ? n6373 : ~n32;
  assign n6375 = pi17 ? n1478 : ~n6374;
  assign n6376 = pi16 ? n32 : n6375;
  assign n6377 = pi15 ? n6371 : n6376;
  assign n6378 = pi20 ? n32 : ~n3523;
  assign n6379 = pi19 ? n32 : n6378;
  assign n6380 = pi19 ? n594 : ~n617;
  assign n6381 = pi18 ? n6379 : ~n6380;
  assign n6382 = pi17 ? n1478 : ~n6381;
  assign n6383 = pi16 ? n32 : n6382;
  assign n6384 = pi19 ? n531 : ~n617;
  assign n6385 = pi18 ? n863 : ~n6384;
  assign n6386 = pi17 ? n1213 : ~n6385;
  assign n6387 = pi16 ? n32 : n6386;
  assign n6388 = pi15 ? n6383 : n6387;
  assign n6389 = pi14 ? n6377 : n6388;
  assign n6390 = pi13 ? n6368 : n6389;
  assign n6391 = pi12 ? n6349 : n6390;
  assign n6392 = pi17 ? n1213 : ~n6133;
  assign n6393 = pi16 ? n32 : n6392;
  assign n6394 = pi18 ? n209 : ~n4492;
  assign n6395 = pi20 ? n207 : ~n501;
  assign n6396 = pi20 ? n749 : n321;
  assign n6397 = pi19 ? n6395 : n6396;
  assign n6398 = pi20 ? n32 : n3523;
  assign n6399 = pi19 ? n6398 : n32;
  assign n6400 = pi18 ? n6397 : ~n6399;
  assign n6401 = pi17 ? n6394 : ~n6400;
  assign n6402 = pi16 ? n32 : n6401;
  assign n6403 = pi15 ? n6393 : n6402;
  assign n6404 = pi18 ? n245 : ~n6145;
  assign n6405 = pi19 ? n208 : ~n236;
  assign n6406 = pi18 ? n6405 : n32;
  assign n6407 = pi17 ? n6404 : n6406;
  assign n6408 = pi16 ? n32 : n6407;
  assign n6409 = pi17 ? n1041 : ~n6153;
  assign n6410 = pi16 ? n32 : n6409;
  assign n6411 = pi15 ? n6408 : n6410;
  assign n6412 = pi14 ? n6403 : n6411;
  assign n6413 = pi17 ? n1134 : ~n6160;
  assign n6414 = pi16 ? n32 : n6413;
  assign n6415 = pi17 ? n1134 : ~n6164;
  assign n6416 = pi16 ? n32 : n6415;
  assign n6417 = pi15 ? n6414 : n6416;
  assign n6418 = pi17 ? n4798 : ~n6168;
  assign n6419 = pi16 ? n32 : n6418;
  assign n6420 = pi20 ? n321 : ~n339;
  assign n6421 = pi19 ? n6420 : ~n349;
  assign n6422 = pi18 ? n6421 : ~n6174;
  assign n6423 = pi17 ? n4798 : ~n6422;
  assign n6424 = pi16 ? n32 : n6423;
  assign n6425 = pi15 ? n6419 : n6424;
  assign n6426 = pi14 ? n6417 : n6425;
  assign n6427 = pi13 ? n6412 : n6426;
  assign n6428 = pi17 ? n1966 : n6182;
  assign n6429 = pi16 ? n32 : n6428;
  assign n6430 = pi17 ? n4804 : ~n6185;
  assign n6431 = pi16 ? n32 : n6430;
  assign n6432 = pi15 ? n6429 : n6431;
  assign n6433 = pi17 ? n4804 : ~n2512;
  assign n6434 = pi16 ? n32 : n6433;
  assign n6435 = pi14 ? n6432 : n6434;
  assign n6436 = pi17 ? n1700 : ~n2512;
  assign n6437 = pi16 ? n32 : n6436;
  assign n6438 = pi15 ? n6434 : n6437;
  assign n6439 = pi18 ? n2849 : ~n32;
  assign n6440 = pi17 ? n6439 : ~n2512;
  assign n6441 = pi16 ? n32 : n6440;
  assign n6442 = pi14 ? n6438 : n6441;
  assign n6443 = pi13 ? n6435 : n6442;
  assign n6444 = pi12 ? n6427 : n6443;
  assign n6445 = pi11 ? n6391 : n6444;
  assign n6446 = pi15 ? n6441 : n5522;
  assign n6447 = pi14 ? n6441 : n6446;
  assign n6448 = pi19 ? n322 : ~n5597;
  assign n6449 = pi18 ? n32 : n6448;
  assign n6450 = pi17 ? n4497 : ~n6449;
  assign n6451 = pi16 ? n32 : n6450;
  assign n6452 = pi17 ? n4497 : ~n2512;
  assign n6453 = pi16 ? n32 : n6452;
  assign n6454 = pi15 ? n6451 : n6453;
  assign n6455 = pi14 ? n6454 : n6453;
  assign n6456 = pi13 ? n6447 : n6455;
  assign n6457 = pi17 ? n1984 : ~n2512;
  assign n6458 = pi16 ? n32 : n6457;
  assign n6459 = pi17 ? n1984 : ~n2750;
  assign n6460 = pi16 ? n32 : n6459;
  assign n6461 = pi17 ? n1984 : ~n2519;
  assign n6462 = pi16 ? n32 : n6461;
  assign n6463 = pi15 ? n6460 : n6462;
  assign n6464 = pi14 ? n6458 : n6463;
  assign n6465 = pi17 ? n1989 : ~n2519;
  assign n6466 = pi16 ? n32 : n6465;
  assign n6467 = pi15 ? n6462 : n6466;
  assign n6468 = pi17 ? n1989 : ~n5978;
  assign n6469 = pi16 ? n32 : n6468;
  assign n6470 = pi15 ? n6466 : n6469;
  assign n6471 = pi14 ? n6467 : n6470;
  assign n6472 = pi13 ? n6464 : n6471;
  assign n6473 = pi12 ? n6456 : n6472;
  assign n6474 = pi20 ? n140 : ~n32;
  assign n6475 = pi19 ? n507 : n6474;
  assign n6476 = pi18 ? n32 : n6475;
  assign n6477 = pi17 ? n4341 : ~n6476;
  assign n6478 = pi16 ? n32 : n6477;
  assign n6479 = pi15 ? n6201 : n6478;
  assign n6480 = pi17 ? n5930 : ~n2512;
  assign n6481 = pi16 ? n32 : n6480;
  assign n6482 = pi14 ? n6479 : n6481;
  assign n6483 = pi17 ? n5930 : ~n6236;
  assign n6484 = pi16 ? n32 : n6483;
  assign n6485 = pi15 ? n6481 : n6484;
  assign n6486 = pi15 ? n6481 : n6458;
  assign n6487 = pi14 ? n6485 : n6486;
  assign n6488 = pi13 ? n6482 : n6487;
  assign n6489 = pi17 ? n4822 : ~n2750;
  assign n6490 = pi16 ? n32 : n6489;
  assign n6491 = pi17 ? n4822 : ~n6250;
  assign n6492 = pi16 ? n32 : n6491;
  assign n6493 = pi15 ? n6490 : n6492;
  assign n6494 = pi17 ? n4497 : ~n2750;
  assign n6495 = pi16 ? n32 : n6494;
  assign n6496 = pi17 ? n4497 : ~n2855;
  assign n6497 = pi16 ? n32 : n6496;
  assign n6498 = pi15 ? n6495 : n6497;
  assign n6499 = pi14 ? n6493 : n6498;
  assign n6500 = pi19 ? n6057 : ~n32;
  assign n6501 = pi18 ? n32 : n6500;
  assign n6502 = pi17 ? n4497 : ~n6501;
  assign n6503 = pi16 ? n32 : n6502;
  assign n6504 = pi20 ? n3847 : n32;
  assign n6505 = pi19 ? n6504 : n1105;
  assign n6506 = pi18 ? n32 : n6505;
  assign n6507 = pi17 ? n2159 : ~n6506;
  assign n6508 = pi16 ? n32 : n6507;
  assign n6509 = pi15 ? n6503 : n6508;
  assign n6510 = pi17 ? n4659 : ~n2618;
  assign n6511 = pi16 ? n32 : n6510;
  assign n6512 = pi17 ? n2159 : ~n3621;
  assign n6513 = pi16 ? n32 : n6512;
  assign n6514 = pi15 ? n6511 : n6513;
  assign n6515 = pi14 ? n6509 : n6514;
  assign n6516 = pi13 ? n6499 : n6515;
  assign n6517 = pi12 ? n6488 : n6516;
  assign n6518 = pi11 ? n6473 : n6517;
  assign n6519 = pi10 ? n6445 : n6518;
  assign n6520 = pi09 ? n6294 : n6519;
  assign n6521 = pi08 ? n6275 : n6520;
  assign n6522 = pi07 ? n6017 : n6521;
  assign n6523 = pi06 ? n5651 : n6522;
  assign n6524 = pi05 ? n4963 : n6523;
  assign n6525 = pi04 ? n3691 : n6524;
  assign n6526 = pi03 ? n1675 : n6525;
  assign n6527 = pi02 ? n193 : n6526;
  assign n6528 = pi01 ? n32 : n6527;
  assign n6529 = pi17 ? n2414 : ~n2750;
  assign n6530 = pi16 ? n32 : n6529;
  assign n6531 = pi15 ? n32 : n6530;
  assign n6532 = pi17 ? n2414 : ~n3067;
  assign n6533 = pi16 ? n32 : n6532;
  assign n6534 = pi17 ? n2119 : ~n3067;
  assign n6535 = pi16 ? n32 : n6534;
  assign n6536 = pi15 ? n6533 : n6535;
  assign n6537 = pi14 ? n6531 : n6536;
  assign n6538 = pi13 ? n32 : n6537;
  assign n6539 = pi12 ? n32 : n6538;
  assign n6540 = pi11 ? n32 : n6539;
  assign n6541 = pi10 ? n32 : n6540;
  assign n6542 = pi17 ? n2425 : ~n2726;
  assign n6543 = pi16 ? n32 : n6542;
  assign n6544 = pi17 ? n2531 : ~n3067;
  assign n6545 = pi16 ? n32 : n6544;
  assign n6546 = pi15 ? n6543 : n6545;
  assign n6547 = pi17 ? n2299 : ~n3067;
  assign n6548 = pi16 ? n32 : n6547;
  assign n6549 = pi17 ? n2319 : ~n3067;
  assign n6550 = pi16 ? n32 : n6549;
  assign n6551 = pi15 ? n6548 : n6550;
  assign n6552 = pi14 ? n6546 : n6551;
  assign n6553 = pi17 ? n2537 : ~n3067;
  assign n6554 = pi16 ? n32 : n6553;
  assign n6555 = pi15 ? n6550 : n6554;
  assign n6556 = pi17 ? n3337 : ~n3067;
  assign n6557 = pi16 ? n32 : n6556;
  assign n6558 = pi17 ? n1807 : ~n3067;
  assign n6559 = pi16 ? n32 : n6558;
  assign n6560 = pi15 ? n6557 : n6559;
  assign n6561 = pi14 ? n6555 : n6560;
  assign n6562 = pi13 ? n6552 : n6561;
  assign n6563 = pi17 ? n2136 : ~n3067;
  assign n6564 = pi16 ? n32 : n6563;
  assign n6565 = pi17 ? n1576 : ~n3067;
  assign n6566 = pi16 ? n32 : n6565;
  assign n6567 = pi17 ? n1833 : ~n3067;
  assign n6568 = pi16 ? n32 : n6567;
  assign n6569 = pi15 ? n6566 : n6568;
  assign n6570 = pi14 ? n6564 : n6569;
  assign n6571 = pi17 ? n2143 : ~n3067;
  assign n6572 = pi16 ? n32 : n6571;
  assign n6573 = pi17 ? n1580 : ~n3067;
  assign n6574 = pi16 ? n32 : n6573;
  assign n6575 = pi15 ? n6572 : n6574;
  assign n6576 = pi17 ? n1593 : ~n3067;
  assign n6577 = pi16 ? n32 : n6576;
  assign n6578 = pi14 ? n6575 : n6577;
  assign n6579 = pi13 ? n6570 : n6578;
  assign n6580 = pi12 ? n6562 : n6579;
  assign n6581 = pi19 ? n322 : ~n349;
  assign n6582 = pi18 ? n32 : ~n6581;
  assign n6583 = pi17 ? n1842 : ~n6582;
  assign n6584 = pi16 ? n32 : n6583;
  assign n6585 = pi15 ? n6577 : n6584;
  assign n6586 = pi19 ? n358 : n349;
  assign n6587 = pi18 ? n32 : n6586;
  assign n6588 = pi17 ? n1470 : ~n6587;
  assign n6589 = pi16 ? n32 : n6588;
  assign n6590 = pi17 ? n1470 : ~n3067;
  assign n6591 = pi16 ? n32 : n6590;
  assign n6592 = pi15 ? n6589 : n6591;
  assign n6593 = pi14 ? n6585 : n6592;
  assign n6594 = pi17 ? n1971 : ~n3067;
  assign n6595 = pi16 ? n32 : n6594;
  assign n6596 = pi19 ? n5694 : n349;
  assign n6597 = pi18 ? n32 : n6596;
  assign n6598 = pi17 ? n1971 : ~n6597;
  assign n6599 = pi16 ? n32 : n6598;
  assign n6600 = pi19 ? n322 : n1757;
  assign n6601 = pi18 ? n1592 : ~n6600;
  assign n6602 = pi17 ? n1213 : ~n6601;
  assign n6603 = pi16 ? n32 : n6602;
  assign n6604 = pi15 ? n6599 : n6603;
  assign n6605 = pi14 ? n6595 : n6604;
  assign n6606 = pi13 ? n6593 : n6605;
  assign n6607 = pi18 ? n32 : ~n5747;
  assign n6608 = pi17 ? n930 : ~n6607;
  assign n6609 = pi16 ? n32 : n6608;
  assign n6610 = pi17 ? n930 : ~n3067;
  assign n6611 = pi16 ? n32 : n6610;
  assign n6612 = pi15 ? n6609 : n6611;
  assign n6613 = pi17 ? n1697 : ~n2736;
  assign n6614 = pi16 ? n32 : n6613;
  assign n6615 = pi15 ? n6611 : n6614;
  assign n6616 = pi14 ? n6612 : n6615;
  assign n6617 = pi21 ? n259 : n173;
  assign n6618 = pi20 ? n6617 : ~n207;
  assign n6619 = pi20 ? n5854 : ~n32;
  assign n6620 = pi19 ? n6618 : n6619;
  assign n6621 = pi21 ? n206 : n174;
  assign n6622 = pi20 ? n32 : n6621;
  assign n6623 = pi19 ? n6622 : n32;
  assign n6624 = pi18 ? n6620 : ~n6623;
  assign n6625 = pi17 ? n1697 : ~n6624;
  assign n6626 = pi16 ? n32 : n6625;
  assign n6627 = pi15 ? n6614 : n6626;
  assign n6628 = pi19 ? n349 : ~n502;
  assign n6629 = pi18 ? n32 : ~n6628;
  assign n6630 = pi17 ? n4798 : ~n6629;
  assign n6631 = pi16 ? n32 : n6630;
  assign n6632 = pi17 ? n4798 : ~n2736;
  assign n6633 = pi16 ? n32 : n6632;
  assign n6634 = pi15 ? n6631 : n6633;
  assign n6635 = pi14 ? n6627 : n6634;
  assign n6636 = pi13 ? n6616 : n6635;
  assign n6637 = pi12 ? n6606 : n6636;
  assign n6638 = pi11 ? n6580 : n6637;
  assign n6639 = pi17 ? n4798 : ~n3067;
  assign n6640 = pi16 ? n32 : n6639;
  assign n6641 = pi19 ? n4342 : n349;
  assign n6642 = pi18 ? n32 : n6641;
  assign n6643 = pi17 ? n1706 : ~n6642;
  assign n6644 = pi16 ? n32 : n6643;
  assign n6645 = pi19 ? n322 : ~n236;
  assign n6646 = pi18 ? n209 : ~n6645;
  assign n6647 = pi17 ? n4656 : ~n6646;
  assign n6648 = pi16 ? n32 : n6647;
  assign n6649 = pi15 ? n6644 : n6648;
  assign n6650 = pi14 ? n6640 : n6649;
  assign n6651 = pi21 ? n206 : ~n124;
  assign n6652 = pi20 ? n6651 : ~n32;
  assign n6653 = pi19 ? n32 : n6652;
  assign n6654 = pi18 ? n32 : n6653;
  assign n6655 = pi17 ? n4656 : ~n6654;
  assign n6656 = pi16 ? n32 : n6655;
  assign n6657 = pi17 ? n4656 : ~n3067;
  assign n6658 = pi16 ? n32 : n6657;
  assign n6659 = pi15 ? n6656 : n6658;
  assign n6660 = pi19 ? n1818 : n349;
  assign n6661 = pi18 ? n32 : n6660;
  assign n6662 = pi17 ? n4656 : ~n6661;
  assign n6663 = pi16 ? n32 : n6662;
  assign n6664 = pi15 ? n6663 : n6658;
  assign n6665 = pi14 ? n6659 : n6664;
  assign n6666 = pi13 ? n6650 : n6665;
  assign n6667 = pi17 ? n1978 : ~n3067;
  assign n6668 = pi16 ? n32 : n6667;
  assign n6669 = pi19 ? n531 : ~n349;
  assign n6670 = pi18 ? n32 : ~n6669;
  assign n6671 = pi17 ? n4659 : ~n6670;
  assign n6672 = pi16 ? n32 : n6671;
  assign n6673 = pi15 ? n6668 : n6672;
  assign n6674 = pi17 ? n4659 : ~n3067;
  assign n6675 = pi16 ? n32 : n6674;
  assign n6676 = pi15 ? n6668 : n6675;
  assign n6677 = pi14 ? n6673 : n6676;
  assign n6678 = pi17 ? n1472 : ~n3067;
  assign n6679 = pi16 ? n32 : n6678;
  assign n6680 = pi15 ? n6668 : n6679;
  assign n6681 = pi17 ? n1472 : ~n2733;
  assign n6682 = pi16 ? n32 : n6681;
  assign n6683 = pi20 ? n2358 : ~n32;
  assign n6684 = pi19 ? n32 : n6683;
  assign n6685 = pi18 ? n32 : n6684;
  assign n6686 = pi17 ? n4497 : ~n6685;
  assign n6687 = pi16 ? n32 : n6686;
  assign n6688 = pi15 ? n6682 : n6687;
  assign n6689 = pi14 ? n6680 : n6688;
  assign n6690 = pi13 ? n6677 : n6689;
  assign n6691 = pi12 ? n6666 : n6690;
  assign n6692 = pi21 ? n1009 : n140;
  assign n6693 = pi20 ? n6692 : ~n32;
  assign n6694 = pi19 ? n32 : n6693;
  assign n6695 = pi18 ? n32 : n6694;
  assign n6696 = pi17 ? n4497 : ~n6695;
  assign n6697 = pi16 ? n32 : n6696;
  assign n6698 = pi15 ? n6687 : n6697;
  assign n6699 = pi17 ? n2159 : ~n3067;
  assign n6700 = pi16 ? n32 : n6699;
  assign n6701 = pi15 ? n6700 : n6675;
  assign n6702 = pi14 ? n6698 : n6701;
  assign n6703 = pi17 ? n2159 : ~n2736;
  assign n6704 = pi16 ? n32 : n6703;
  assign n6705 = pi17 ? n4659 : ~n2736;
  assign n6706 = pi16 ? n32 : n6705;
  assign n6707 = pi15 ? n6704 : n6706;
  assign n6708 = pi17 ? n6439 : ~n2736;
  assign n6709 = pi16 ? n32 : n6708;
  assign n6710 = pi15 ? n6706 : n6709;
  assign n6711 = pi14 ? n6707 : n6710;
  assign n6712 = pi13 ? n6702 : n6711;
  assign n6713 = pi17 ? n6439 : ~n2855;
  assign n6714 = pi16 ? n32 : n6713;
  assign n6715 = pi15 ? n6709 : n6714;
  assign n6716 = pi17 ? n1700 : ~n2855;
  assign n6717 = pi16 ? n32 : n6716;
  assign n6718 = pi17 ? n4656 : ~n3812;
  assign n6719 = pi16 ? n32 : n6718;
  assign n6720 = pi15 ? n6717 : n6719;
  assign n6721 = pi14 ? n6715 : n6720;
  assign n6722 = pi20 ? n32 : n405;
  assign n6723 = pi19 ? n6722 : n1105;
  assign n6724 = pi18 ? n32 : n6723;
  assign n6725 = pi17 ? n4656 : ~n6724;
  assign n6726 = pi16 ? n32 : n6725;
  assign n6727 = pi20 ? n32 : ~n785;
  assign n6728 = pi19 ? n6727 : n1105;
  assign n6729 = pi18 ? n32 : n6728;
  assign n6730 = pi17 ? n4804 : ~n6729;
  assign n6731 = pi16 ? n32 : n6730;
  assign n6732 = pi15 ? n6726 : n6731;
  assign n6733 = pi17 ? n4804 : ~n3621;
  assign n6734 = pi16 ? n32 : n6733;
  assign n6735 = pi17 ? n1706 : ~n3621;
  assign n6736 = pi16 ? n32 : n6735;
  assign n6737 = pi15 ? n6734 : n6736;
  assign n6738 = pi14 ? n6732 : n6737;
  assign n6739 = pi13 ? n6721 : n6738;
  assign n6740 = pi12 ? n6712 : n6739;
  assign n6741 = pi11 ? n6691 : n6740;
  assign n6742 = pi10 ? n6638 : n6741;
  assign n6743 = pi09 ? n6541 : n6742;
  assign n6744 = pi17 ? n2512 : ~n2750;
  assign n6745 = pi16 ? n32 : n6744;
  assign n6746 = pi15 ? n32 : n6745;
  assign n6747 = pi17 ? n2512 : ~n3067;
  assign n6748 = pi16 ? n32 : n6747;
  assign n6749 = pi17 ? n2517 : ~n3067;
  assign n6750 = pi16 ? n32 : n6749;
  assign n6751 = pi15 ? n6748 : n6750;
  assign n6752 = pi14 ? n6746 : n6751;
  assign n6753 = pi13 ? n32 : n6752;
  assign n6754 = pi12 ? n32 : n6753;
  assign n6755 = pi11 ? n32 : n6754;
  assign n6756 = pi10 ? n32 : n6755;
  assign n6757 = pi17 ? n2755 : ~n2726;
  assign n6758 = pi16 ? n32 : n6757;
  assign n6759 = pi17 ? n2408 : ~n3067;
  assign n6760 = pi16 ? n32 : n6759;
  assign n6761 = pi15 ? n6758 : n6760;
  assign n6762 = pi15 ? n6533 : n6548;
  assign n6763 = pi14 ? n6761 : n6762;
  assign n6764 = pi17 ? n2410 : ~n3067;
  assign n6765 = pi16 ? n32 : n6764;
  assign n6766 = pi15 ? n6548 : n6765;
  assign n6767 = pi19 ? n32 : n6042;
  assign n6768 = pi18 ? n32 : n6767;
  assign n6769 = pi17 ? n2305 : ~n6768;
  assign n6770 = pi16 ? n32 : n6769;
  assign n6771 = pi17 ? n1933 : ~n3067;
  assign n6772 = pi16 ? n32 : n6771;
  assign n6773 = pi15 ? n6770 : n6772;
  assign n6774 = pi14 ? n6766 : n6773;
  assign n6775 = pi13 ? n6763 : n6774;
  assign n6776 = pi15 ? n6550 : n6564;
  assign n6777 = pi17 ? n1943 : ~n3067;
  assign n6778 = pi16 ? n32 : n6777;
  assign n6779 = pi15 ? n6564 : n6778;
  assign n6780 = pi14 ? n6776 : n6779;
  assign n6781 = pi17 ? n2325 : ~n3067;
  assign n6782 = pi16 ? n32 : n6781;
  assign n6783 = pi17 ? n3351 : ~n3067;
  assign n6784 = pi16 ? n32 : n6783;
  assign n6785 = pi15 ? n6782 : n6784;
  assign n6786 = pi14 ? n6785 : n6566;
  assign n6787 = pi13 ? n6780 : n6786;
  assign n6788 = pi12 ? n6775 : n6787;
  assign n6789 = pi20 ? n820 : ~n321;
  assign n6790 = pi19 ? n6789 : n349;
  assign n6791 = pi18 ? n32 : n6790;
  assign n6792 = pi17 ? n1833 : ~n6791;
  assign n6793 = pi16 ? n32 : n6792;
  assign n6794 = pi15 ? n6566 : n6793;
  assign n6795 = pi14 ? n6794 : n6572;
  assign n6796 = pi17 ? n1322 : ~n3067;
  assign n6797 = pi16 ? n32 : n6796;
  assign n6798 = pi17 ? n1322 : ~n6597;
  assign n6799 = pi16 ? n32 : n6798;
  assign n6800 = pi20 ? n339 : ~n321;
  assign n6801 = pi19 ? n6800 : n6683;
  assign n6802 = pi18 ? n32 : n6801;
  assign n6803 = pi17 ? n1593 : ~n6802;
  assign n6804 = pi16 ? n32 : n6803;
  assign n6805 = pi15 ? n6799 : n6804;
  assign n6806 = pi14 ? n6797 : n6805;
  assign n6807 = pi13 ? n6795 : n6806;
  assign n6808 = pi18 ? n32 : n6152;
  assign n6809 = pi17 ? n1842 : ~n6808;
  assign n6810 = pi16 ? n32 : n6809;
  assign n6811 = pi17 ? n1842 : ~n3067;
  assign n6812 = pi16 ? n32 : n6811;
  assign n6813 = pi15 ? n6810 : n6812;
  assign n6814 = pi17 ? n1704 : ~n3067;
  assign n6815 = pi16 ? n32 : n6814;
  assign n6816 = pi17 ? n1704 : ~n2736;
  assign n6817 = pi16 ? n32 : n6816;
  assign n6818 = pi15 ? n6815 : n6817;
  assign n6819 = pi14 ? n6813 : n6818;
  assign n6820 = pi17 ? n1704 : ~n2852;
  assign n6821 = pi16 ? n32 : n6820;
  assign n6822 = pi21 ? n174 : n173;
  assign n6823 = pi20 ? n6822 : n357;
  assign n6824 = pi20 ? n3523 : ~n2256;
  assign n6825 = pi19 ? n6823 : n6824;
  assign n6826 = pi19 ? n4126 : n5614;
  assign n6827 = pi18 ? n6825 : ~n6826;
  assign n6828 = pi17 ? n1971 : ~n6827;
  assign n6829 = pi16 ? n32 : n6828;
  assign n6830 = pi15 ? n6821 : n6829;
  assign n6831 = pi17 ? n1971 : ~n6607;
  assign n6832 = pi16 ? n32 : n6831;
  assign n6833 = pi17 ? n1971 : ~n2736;
  assign n6834 = pi16 ? n32 : n6833;
  assign n6835 = pi15 ? n6832 : n6834;
  assign n6836 = pi14 ? n6830 : n6835;
  assign n6837 = pi13 ? n6819 : n6836;
  assign n6838 = pi12 ? n6807 : n6837;
  assign n6839 = pi11 ? n6788 : n6838;
  assign n6840 = pi17 ? n1134 : ~n3067;
  assign n6841 = pi16 ? n32 : n6840;
  assign n6842 = pi15 ? n6595 : n6841;
  assign n6843 = pi17 ? n1134 : ~n6642;
  assign n6844 = pi16 ? n32 : n6843;
  assign n6845 = pi18 ? n1957 : ~n6645;
  assign n6846 = pi17 ? n1232 : ~n6845;
  assign n6847 = pi16 ? n32 : n6846;
  assign n6848 = pi15 ? n6844 : n6847;
  assign n6849 = pi14 ? n6842 : n6848;
  assign n6850 = pi17 ? n1232 : ~n2736;
  assign n6851 = pi16 ? n32 : n6850;
  assign n6852 = pi17 ? n1232 : ~n3067;
  assign n6853 = pi16 ? n32 : n6852;
  assign n6854 = pi15 ? n6851 : n6853;
  assign n6855 = pi17 ? n1232 : ~n6661;
  assign n6856 = pi16 ? n32 : n6855;
  assign n6857 = pi17 ? n1966 : ~n3067;
  assign n6858 = pi16 ? n32 : n6857;
  assign n6859 = pi15 ? n6856 : n6858;
  assign n6860 = pi14 ? n6854 : n6859;
  assign n6861 = pi13 ? n6849 : n6860;
  assign n6862 = pi19 ? n531 : ~n1077;
  assign n6863 = pi18 ? n32 : ~n6862;
  assign n6864 = pi17 ? n1966 : ~n6863;
  assign n6865 = pi16 ? n32 : n6864;
  assign n6866 = pi15 ? n6858 : n6865;
  assign n6867 = pi19 ? n1844 : n32;
  assign n6868 = pi18 ? n1965 : ~n6867;
  assign n6869 = pi17 ? n6868 : ~n3067;
  assign n6870 = pi16 ? n32 : n6869;
  assign n6871 = pi15 ? n6870 : n6858;
  assign n6872 = pi14 ? n6866 : n6871;
  assign n6873 = pi17 ? n1700 : ~n3067;
  assign n6874 = pi16 ? n32 : n6873;
  assign n6875 = pi15 ? n6870 : n6874;
  assign n6876 = pi17 ? n1700 : ~n2733;
  assign n6877 = pi16 ? n32 : n6876;
  assign n6878 = pi17 ? n1700 : ~n6685;
  assign n6879 = pi16 ? n32 : n6878;
  assign n6880 = pi15 ? n6877 : n6879;
  assign n6881 = pi14 ? n6875 : n6880;
  assign n6882 = pi13 ? n6872 : n6881;
  assign n6883 = pi12 ? n6861 : n6882;
  assign n6884 = pi17 ? n4656 : ~n6685;
  assign n6885 = pi16 ? n32 : n6884;
  assign n6886 = pi21 ? n309 : n140;
  assign n6887 = pi20 ? n6886 : ~n32;
  assign n6888 = pi19 ? n32 : n6887;
  assign n6889 = pi18 ? n32 : n6888;
  assign n6890 = pi17 ? n4656 : ~n6889;
  assign n6891 = pi16 ? n32 : n6890;
  assign n6892 = pi15 ? n6885 : n6891;
  assign n6893 = pi17 ? n4804 : ~n3067;
  assign n6894 = pi16 ? n32 : n6893;
  assign n6895 = pi14 ? n6892 : n6894;
  assign n6896 = pi17 ? n4804 : ~n2736;
  assign n6897 = pi16 ? n32 : n6896;
  assign n6898 = pi22 ? n173 : ~n84;
  assign n6899 = pi21 ? n6898 : ~n32;
  assign n6900 = pi20 ? n6899 : ~n32;
  assign n6901 = pi19 ? n32 : n6900;
  assign n6902 = pi18 ? n32 : n6901;
  assign n6903 = pi17 ? n4804 : ~n6902;
  assign n6904 = pi16 ? n32 : n6903;
  assign n6905 = pi15 ? n6897 : n6904;
  assign n6906 = pi17 ? n1966 : ~n2736;
  assign n6907 = pi16 ? n32 : n6906;
  assign n6908 = pi15 ? n6897 : n6907;
  assign n6909 = pi14 ? n6905 : n6908;
  assign n6910 = pi13 ? n6895 : n6909;
  assign n6911 = pi17 ? n4798 : ~n2731;
  assign n6912 = pi16 ? n32 : n6911;
  assign n6913 = pi17 ? n4798 : ~n2855;
  assign n6914 = pi16 ? n32 : n6913;
  assign n6915 = pi15 ? n6912 : n6914;
  assign n6916 = pi17 ? n1232 : ~n2855;
  assign n6917 = pi16 ? n32 : n6916;
  assign n6918 = pi19 ? n594 : n1105;
  assign n6919 = pi18 ? n32 : n6918;
  assign n6920 = pi17 ? n1232 : ~n6919;
  assign n6921 = pi16 ? n32 : n6920;
  assign n6922 = pi15 ? n6917 : n6921;
  assign n6923 = pi14 ? n6915 : n6922;
  assign n6924 = pi17 ? n1232 : ~n6724;
  assign n6925 = pi16 ? n32 : n6924;
  assign n6926 = pi19 ? n6727 : ~n32;
  assign n6927 = pi18 ? n32 : n6926;
  assign n6928 = pi17 ? n1134 : ~n6927;
  assign n6929 = pi16 ? n32 : n6928;
  assign n6930 = pi15 ? n6925 : n6929;
  assign n6931 = pi17 ? n930 : ~n3621;
  assign n6932 = pi16 ? n32 : n6931;
  assign n6933 = pi17 ? n1134 : ~n3621;
  assign n6934 = pi16 ? n32 : n6933;
  assign n6935 = pi15 ? n6932 : n6934;
  assign n6936 = pi14 ? n6930 : n6935;
  assign n6937 = pi13 ? n6923 : n6936;
  assign n6938 = pi12 ? n6910 : n6937;
  assign n6939 = pi11 ? n6883 : n6938;
  assign n6940 = pi10 ? n6839 : n6939;
  assign n6941 = pi09 ? n6756 : n6940;
  assign n6942 = pi08 ? n6743 : n6941;
  assign n6943 = pi17 ? n2623 : ~n2750;
  assign n6944 = pi16 ? n32 : n6943;
  assign n6945 = pi15 ? n32 : n6944;
  assign n6946 = pi17 ? n2623 : ~n3067;
  assign n6947 = pi16 ? n32 : n6946;
  assign n6948 = pi17 ? n4099 : ~n3067;
  assign n6949 = pi16 ? n32 : n6948;
  assign n6950 = pi15 ? n6947 : n6949;
  assign n6951 = pi14 ? n6945 : n6950;
  assign n6952 = pi13 ? n32 : n6951;
  assign n6953 = pi12 ? n32 : n6952;
  assign n6954 = pi11 ? n32 : n6953;
  assign n6955 = pi10 ? n32 : n6954;
  assign n6956 = pi17 ? n2618 : ~n2726;
  assign n6957 = pi16 ? n32 : n6956;
  assign n6958 = pi15 ? n6957 : n6748;
  assign n6959 = pi17 ? n2748 : ~n3067;
  assign n6960 = pi16 ? n32 : n6959;
  assign n6961 = pi15 ? n6960 : n6535;
  assign n6962 = pi14 ? n6958 : n6961;
  assign n6963 = pi17 ? n2425 : ~n3067;
  assign n6964 = pi16 ? n32 : n6963;
  assign n6965 = pi15 ? n6535 : n6964;
  assign n6966 = pi17 ? n2653 : ~n6768;
  assign n6967 = pi16 ? n32 : n6966;
  assign n6968 = pi15 ? n6967 : n6548;
  assign n6969 = pi14 ? n6965 : n6968;
  assign n6970 = pi13 ? n6962 : n6969;
  assign n6971 = pi14 ? n6551 : n6555;
  assign n6972 = pi17 ? n3337 : ~n6768;
  assign n6973 = pi16 ? n32 : n6972;
  assign n6974 = pi15 ? n6973 : n6559;
  assign n6975 = pi14 ? n6974 : n6564;
  assign n6976 = pi13 ? n6971 : n6975;
  assign n6977 = pi12 ? n6970 : n6976;
  assign n6978 = pi19 ? n267 : n349;
  assign n6979 = pi18 ? n32 : n6978;
  assign n6980 = pi17 ? n1943 : ~n6979;
  assign n6981 = pi16 ? n32 : n6980;
  assign n6982 = pi15 ? n6564 : n6981;
  assign n6983 = pi14 ? n6982 : n6782;
  assign n6984 = pi17 ? n1682 : ~n3067;
  assign n6985 = pi16 ? n32 : n6984;
  assign n6986 = pi17 ? n1682 : ~n6597;
  assign n6987 = pi16 ? n32 : n6986;
  assign n6988 = pi20 ? n342 : ~n321;
  assign n6989 = pi19 ? n6988 : n349;
  assign n6990 = pi18 ? n32 : n6989;
  assign n6991 = pi17 ? n1576 : ~n6990;
  assign n6992 = pi16 ? n32 : n6991;
  assign n6993 = pi15 ? n6987 : n6992;
  assign n6994 = pi14 ? n6985 : n6993;
  assign n6995 = pi13 ? n6983 : n6994;
  assign n6996 = pi14 ? n6568 : n6574;
  assign n6997 = pi20 ? n321 : ~n206;
  assign n6998 = pi19 ? n6997 : n349;
  assign n6999 = pi18 ? n32 : n6998;
  assign n7000 = pi17 ? n1322 : ~n6999;
  assign n7001 = pi16 ? n32 : n7000;
  assign n7002 = pi15 ? n6574 : n7001;
  assign n7003 = pi14 ? n7002 : n6797;
  assign n7004 = pi13 ? n6996 : n7003;
  assign n7005 = pi12 ? n6995 : n7004;
  assign n7006 = pi11 ? n6977 : n7005;
  assign n7007 = pi21 ? n32 : ~n124;
  assign n7008 = pi20 ? n7007 : ~n32;
  assign n7009 = pi19 ? n4342 : n7008;
  assign n7010 = pi18 ? n32 : n7009;
  assign n7011 = pi17 ? n1470 : ~n7010;
  assign n7012 = pi16 ? n32 : n7011;
  assign n7013 = pi21 ? n206 : n140;
  assign n7014 = pi20 ? n7013 : ~n32;
  assign n7015 = pi19 ? n4964 : n7014;
  assign n7016 = pi18 ? n32 : n7015;
  assign n7017 = pi17 ? n1478 : ~n7016;
  assign n7018 = pi16 ? n32 : n7017;
  assign n7019 = pi15 ? n7012 : n7018;
  assign n7020 = pi14 ? n6591 : n7019;
  assign n7021 = pi17 ? n1478 : ~n2850;
  assign n7022 = pi16 ? n32 : n7021;
  assign n7023 = pi20 ? n1839 : n339;
  assign n7024 = pi19 ? n1464 : n7023;
  assign n7025 = pi18 ? n32 : n7024;
  assign n7026 = pi17 ? n1478 : ~n7025;
  assign n7027 = pi16 ? n32 : n7026;
  assign n7028 = pi15 ? n7022 : n7027;
  assign n7029 = pi19 ? n1464 : n2848;
  assign n7030 = pi18 ? n32 : n7029;
  assign n7031 = pi17 ? n1478 : ~n7030;
  assign n7032 = pi16 ? n32 : n7031;
  assign n7033 = pi17 ? n1213 : ~n3067;
  assign n7034 = pi16 ? n32 : n7033;
  assign n7035 = pi15 ? n7032 : n7034;
  assign n7036 = pi14 ? n7028 : n7035;
  assign n7037 = pi13 ? n7020 : n7036;
  assign n7038 = pi19 ? n32 : n6298;
  assign n7039 = pi18 ? n32 : n7038;
  assign n7040 = pi17 ? n1213 : ~n7039;
  assign n7041 = pi16 ? n32 : n7040;
  assign n7042 = pi19 ? n531 : ~n343;
  assign n7043 = pi18 ? n32 : ~n7042;
  assign n7044 = pi17 ? n1213 : ~n7043;
  assign n7045 = pi16 ? n32 : n7044;
  assign n7046 = pi15 ? n7041 : n7045;
  assign n7047 = pi17 ? n1213 : ~n6768;
  assign n7048 = pi16 ? n32 : n7047;
  assign n7049 = pi14 ? n7046 : n7048;
  assign n7050 = pi17 ? n1697 : ~n3067;
  assign n7051 = pi16 ? n32 : n7050;
  assign n7052 = pi15 ? n7034 : n7051;
  assign n7053 = pi17 ? n1697 : ~n2733;
  assign n7054 = pi16 ? n32 : n7053;
  assign n7055 = pi19 ? n594 : n349;
  assign n7056 = pi18 ? n32 : n7055;
  assign n7057 = pi17 ? n1232 : ~n7056;
  assign n7058 = pi16 ? n32 : n7057;
  assign n7059 = pi15 ? n7054 : n7058;
  assign n7060 = pi14 ? n7052 : n7059;
  assign n7061 = pi13 ? n7049 : n7060;
  assign n7062 = pi12 ? n7037 : n7061;
  assign n7063 = pi17 ? n1232 : ~n2839;
  assign n7064 = pi16 ? n32 : n7063;
  assign n7065 = pi17 ? n1232 : ~n2850;
  assign n7066 = pi16 ? n32 : n7065;
  assign n7067 = pi15 ? n7064 : n7066;
  assign n7068 = pi17 ? n1134 : ~n7056;
  assign n7069 = pi16 ? n32 : n7068;
  assign n7070 = pi15 ? n7069 : n6611;
  assign n7071 = pi14 ? n7067 : n7070;
  assign n7072 = pi17 ? n1134 : ~n3798;
  assign n7073 = pi16 ? n32 : n7072;
  assign n7074 = pi17 ? n930 : ~n4245;
  assign n7075 = pi16 ? n32 : n7074;
  assign n7076 = pi15 ? n7073 : n7075;
  assign n7077 = pi17 ? n930 : ~n3967;
  assign n7078 = pi16 ? n32 : n7077;
  assign n7079 = pi15 ? n7078 : n6834;
  assign n7080 = pi14 ? n7076 : n7079;
  assign n7081 = pi13 ? n7071 : n7080;
  assign n7082 = pi17 ? n1971 : ~n2731;
  assign n7083 = pi16 ? n32 : n7082;
  assign n7084 = pi17 ? n1971 : ~n2750;
  assign n7085 = pi16 ? n32 : n7084;
  assign n7086 = pi15 ? n7083 : n7085;
  assign n7087 = pi17 ? n1704 : ~n2855;
  assign n7088 = pi16 ? n32 : n7087;
  assign n7089 = pi20 ? n342 : ~n220;
  assign n7090 = pi19 ? n7089 : ~n32;
  assign n7091 = pi18 ? n32 : n7090;
  assign n7092 = pi17 ? n1478 : ~n7091;
  assign n7093 = pi16 ? n32 : n7092;
  assign n7094 = pi15 ? n7088 : n7093;
  assign n7095 = pi14 ? n7086 : n7094;
  assign n7096 = pi20 ? n448 : n207;
  assign n7097 = pi19 ? n7096 : ~n1105;
  assign n7098 = pi18 ? n32 : ~n7097;
  assign n7099 = pi17 ? n1478 : ~n7098;
  assign n7100 = pi16 ? n32 : n7099;
  assign n7101 = pi20 ? n32 : ~n5854;
  assign n7102 = pi19 ? n7101 : ~n32;
  assign n7103 = pi18 ? n32 : n7102;
  assign n7104 = pi17 ? n1842 : ~n7103;
  assign n7105 = pi16 ? n32 : n7104;
  assign n7106 = pi15 ? n7100 : n7105;
  assign n7107 = pi22 ? n32 : ~n34;
  assign n7108 = pi21 ? n32 : ~n7107;
  assign n7109 = pi20 ? n207 : n7108;
  assign n7110 = pi19 ? n7109 : ~n32;
  assign n7111 = pi18 ? n6071 : n7110;
  assign n7112 = pi17 ? n1842 : ~n7111;
  assign n7113 = pi16 ? n32 : n7112;
  assign n7114 = pi17 ? n1842 : ~n2618;
  assign n7115 = pi16 ? n32 : n7114;
  assign n7116 = pi15 ? n7113 : n7115;
  assign n7117 = pi14 ? n7106 : n7116;
  assign n7118 = pi13 ? n7095 : n7117;
  assign n7119 = pi12 ? n7081 : n7118;
  assign n7120 = pi11 ? n7062 : n7119;
  assign n7121 = pi10 ? n7006 : n7120;
  assign n7122 = pi09 ? n6955 : n7121;
  assign n7123 = pi17 ? n3067 : ~n2750;
  assign n7124 = pi16 ? n32 : n7123;
  assign n7125 = pi15 ? n32 : n7124;
  assign n7126 = pi17 ? n4245 : ~n3067;
  assign n7127 = pi16 ? n32 : n7126;
  assign n7128 = pi17 ? n2724 : ~n3067;
  assign n7129 = pi16 ? n32 : n7128;
  assign n7130 = pi15 ? n7127 : n7129;
  assign n7131 = pi14 ? n7125 : n7130;
  assign n7132 = pi13 ? n32 : n7131;
  assign n7133 = pi12 ? n32 : n7132;
  assign n7134 = pi11 ? n32 : n7133;
  assign n7135 = pi10 ? n32 : n7134;
  assign n7136 = pi17 ? n2731 : ~n2726;
  assign n7137 = pi16 ? n32 : n7136;
  assign n7138 = pi15 ? n7137 : n6947;
  assign n7139 = pi17 ? n2750 : ~n3067;
  assign n7140 = pi16 ? n32 : n7139;
  assign n7141 = pi15 ? n7140 : n6960;
  assign n7142 = pi14 ? n7138 : n7141;
  assign n7143 = pi17 ? n2755 : ~n3067;
  assign n7144 = pi16 ? n32 : n7143;
  assign n7145 = pi15 ? n6960 : n7144;
  assign n7146 = pi17 ? n2519 : ~n6768;
  assign n7147 = pi16 ? n32 : n7146;
  assign n7148 = pi15 ? n7147 : n6533;
  assign n7149 = pi14 ? n7145 : n7148;
  assign n7150 = pi13 ? n7142 : n7149;
  assign n7151 = pi14 ? n6762 : n6766;
  assign n7152 = pi14 ? n6773 : n6550;
  assign n7153 = pi13 ? n7151 : n7152;
  assign n7154 = pi12 ? n7150 : n7153;
  assign n7155 = pi17 ? n2537 : ~n6979;
  assign n7156 = pi16 ? n32 : n7155;
  assign n7157 = pi15 ? n6550 : n7156;
  assign n7158 = pi14 ? n7157 : n6557;
  assign n7159 = pi17 ? n1814 : ~n3067;
  assign n7160 = pi16 ? n32 : n7159;
  assign n7161 = pi17 ? n1814 : ~n6597;
  assign n7162 = pi16 ? n32 : n7161;
  assign n7163 = pi17 ? n2136 : ~n6990;
  assign n7164 = pi16 ? n32 : n7163;
  assign n7165 = pi15 ? n7162 : n7164;
  assign n7166 = pi14 ? n7160 : n7165;
  assign n7167 = pi13 ? n7158 : n7166;
  assign n7168 = pi20 ? n321 : ~n1331;
  assign n7169 = pi19 ? n32 : n7168;
  assign n7170 = pi18 ? n32 : n7169;
  assign n7171 = pi17 ? n1943 : ~n7170;
  assign n7172 = pi16 ? n32 : n7171;
  assign n7173 = pi15 ? n7172 : n6778;
  assign n7174 = pi17 ? n1677 : ~n3067;
  assign n7175 = pi16 ? n32 : n7174;
  assign n7176 = pi14 ? n7173 : n7175;
  assign n7177 = pi17 ? n1682 : ~n6999;
  assign n7178 = pi16 ? n32 : n7177;
  assign n7179 = pi15 ? n7175 : n7178;
  assign n7180 = pi14 ? n7179 : n6985;
  assign n7181 = pi13 ? n7176 : n7180;
  assign n7182 = pi12 ? n7167 : n7181;
  assign n7183 = pi11 ? n7154 : n7182;
  assign n7184 = pi17 ? n1833 : ~n2850;
  assign n7185 = pi16 ? n32 : n7184;
  assign n7186 = pi15 ? n6568 : n7185;
  assign n7187 = pi19 ? n4342 : n589;
  assign n7188 = pi18 ? n32 : n7187;
  assign n7189 = pi17 ? n1833 : ~n7188;
  assign n7190 = pi16 ? n32 : n7189;
  assign n7191 = pi20 ? n7013 : ~n481;
  assign n7192 = pi19 ? n4964 : n7191;
  assign n7193 = pi18 ? n32 : n7192;
  assign n7194 = pi17 ? n2143 : ~n7193;
  assign n7195 = pi16 ? n32 : n7194;
  assign n7196 = pi15 ? n7190 : n7195;
  assign n7197 = pi14 ? n7186 : n7196;
  assign n7198 = pi17 ? n2143 : ~n2850;
  assign n7199 = pi16 ? n32 : n7198;
  assign n7200 = pi17 ? n2143 : ~n7025;
  assign n7201 = pi16 ? n32 : n7200;
  assign n7202 = pi15 ? n7199 : n7201;
  assign n7203 = pi17 ? n1593 : ~n7030;
  assign n7204 = pi16 ? n32 : n7203;
  assign n7205 = pi21 ? n32 : ~n35;
  assign n7206 = pi20 ? n7205 : ~n32;
  assign n7207 = pi19 ? n32 : n7206;
  assign n7208 = pi18 ? n32 : n7207;
  assign n7209 = pi17 ? n1593 : ~n7208;
  assign n7210 = pi16 ? n32 : n7209;
  assign n7211 = pi15 ? n7204 : n7210;
  assign n7212 = pi14 ? n7202 : n7211;
  assign n7213 = pi13 ? n7197 : n7212;
  assign n7214 = pi17 ? n1593 : ~n7039;
  assign n7215 = pi16 ? n32 : n7214;
  assign n7216 = pi19 ? n531 : ~n2317;
  assign n7217 = pi18 ? n32 : ~n7216;
  assign n7218 = pi17 ? n1593 : ~n7217;
  assign n7219 = pi16 ? n32 : n7218;
  assign n7220 = pi15 ? n7215 : n7219;
  assign n7221 = pi19 ? n462 : n32;
  assign n7222 = pi18 ? n1592 : ~n7221;
  assign n7223 = pi17 ? n7222 : ~n6768;
  assign n7224 = pi16 ? n32 : n7223;
  assign n7225 = pi17 ? n1593 : ~n6768;
  assign n7226 = pi16 ? n32 : n7225;
  assign n7227 = pi15 ? n7224 : n7226;
  assign n7228 = pi14 ? n7220 : n7227;
  assign n7229 = pi21 ? n32 : ~n51;
  assign n7230 = pi20 ? n7229 : ~n32;
  assign n7231 = pi19 ? n32 : n7230;
  assign n7232 = pi18 ? n32 : n7231;
  assign n7233 = pi17 ? n7222 : ~n7232;
  assign n7234 = pi16 ? n32 : n7233;
  assign n7235 = pi17 ? n1704 : ~n7232;
  assign n7236 = pi16 ? n32 : n7235;
  assign n7237 = pi15 ? n7234 : n7236;
  assign n7238 = pi17 ? n1478 : ~n2733;
  assign n7239 = pi16 ? n32 : n7238;
  assign n7240 = pi15 ? n7239 : n6815;
  assign n7241 = pi14 ? n7237 : n7240;
  assign n7242 = pi13 ? n7228 : n7241;
  assign n7243 = pi12 ? n7213 : n7242;
  assign n7244 = pi17 ? n1478 : ~n2836;
  assign n7245 = pi16 ? n32 : n7244;
  assign n7246 = pi17 ? n1478 : ~n3067;
  assign n7247 = pi16 ? n32 : n7246;
  assign n7248 = pi15 ? n7245 : n7247;
  assign n7249 = pi17 ? n1842 : ~n7056;
  assign n7250 = pi16 ? n32 : n7249;
  assign n7251 = pi17 ? n1842 : ~n2724;
  assign n7252 = pi16 ? n32 : n7251;
  assign n7253 = pi15 ? n7250 : n7252;
  assign n7254 = pi14 ? n7248 : n7253;
  assign n7255 = pi17 ? n1842 : ~n3798;
  assign n7256 = pi16 ? n32 : n7255;
  assign n7257 = pi15 ? n7256 : n7252;
  assign n7258 = pi17 ? n1593 : ~n3967;
  assign n7259 = pi16 ? n32 : n7258;
  assign n7260 = pi17 ? n1593 : ~n2731;
  assign n7261 = pi16 ? n32 : n7260;
  assign n7262 = pi15 ? n7259 : n7261;
  assign n7263 = pi14 ? n7257 : n7262;
  assign n7264 = pi13 ? n7254 : n7263;
  assign n7265 = pi17 ? n1322 : ~n2855;
  assign n7266 = pi16 ? n32 : n7265;
  assign n7267 = pi17 ? n1322 : ~n2750;
  assign n7268 = pi16 ? n32 : n7267;
  assign n7269 = pi15 ? n7266 : n7268;
  assign n7270 = pi17 ? n2143 : ~n2855;
  assign n7271 = pi16 ? n32 : n7270;
  assign n7272 = pi17 ? n2143 : ~n7091;
  assign n7273 = pi16 ? n32 : n7272;
  assign n7274 = pi15 ? n7271 : n7273;
  assign n7275 = pi14 ? n7269 : n7274;
  assign n7276 = pi17 ? n1833 : ~n7098;
  assign n7277 = pi16 ? n32 : n7276;
  assign n7278 = pi19 ? n4721 : ~n32;
  assign n7279 = pi18 ? n32 : n7278;
  assign n7280 = pi17 ? n1833 : ~n7279;
  assign n7281 = pi16 ? n32 : n7280;
  assign n7282 = pi15 ? n7277 : n7281;
  assign n7283 = pi20 ? n749 : n7108;
  assign n7284 = pi19 ? n7283 : ~n32;
  assign n7285 = pi18 ? n32 : n7284;
  assign n7286 = pi17 ? n1576 : ~n7285;
  assign n7287 = pi16 ? n32 : n7286;
  assign n7288 = pi17 ? n1833 : ~n2512;
  assign n7289 = pi16 ? n32 : n7288;
  assign n7290 = pi15 ? n7287 : n7289;
  assign n7291 = pi14 ? n7282 : n7290;
  assign n7292 = pi13 ? n7275 : n7291;
  assign n7293 = pi12 ? n7264 : n7292;
  assign n7294 = pi11 ? n7243 : n7293;
  assign n7295 = pi10 ? n7183 : n7294;
  assign n7296 = pi09 ? n7135 : n7295;
  assign n7297 = pi08 ? n7122 : n7296;
  assign n7298 = pi07 ? n6942 : n7297;
  assign n7299 = pi17 ? n2733 : ~n3067;
  assign n7300 = pi16 ? n32 : n7299;
  assign n7301 = pi15 ? n32 : n7300;
  assign n7302 = pi17 ? n2836 : ~n3067;
  assign n7303 = pi16 ? n32 : n7302;
  assign n7304 = pi15 ? n7300 : n7303;
  assign n7305 = pi14 ? n7301 : n7304;
  assign n7306 = pi13 ? n32 : n7305;
  assign n7307 = pi12 ? n32 : n7306;
  assign n7308 = pi11 ? n32 : n7307;
  assign n7309 = pi10 ? n32 : n7308;
  assign n7310 = pi17 ? n2839 : ~n2726;
  assign n7311 = pi16 ? n32 : n7310;
  assign n7312 = pi17 ? n3067 : ~n2726;
  assign n7313 = pi16 ? n32 : n7312;
  assign n7314 = pi15 ? n7311 : n7313;
  assign n7315 = pi17 ? n2750 : ~n2726;
  assign n7316 = pi16 ? n32 : n7315;
  assign n7317 = pi14 ? n7314 : n7316;
  assign n7318 = pi17 ? n2618 : ~n3067;
  assign n7319 = pi16 ? n32 : n7318;
  assign n7320 = pi15 ? n7140 : n7319;
  assign n7321 = pi17 ? n2628 : ~n3067;
  assign n7322 = pi16 ? n32 : n7321;
  assign n7323 = pi17 ? n2748 : ~n2733;
  assign n7324 = pi16 ? n32 : n7323;
  assign n7325 = pi15 ? n7322 : n7324;
  assign n7326 = pi14 ? n7320 : n7325;
  assign n7327 = pi13 ? n7317 : n7326;
  assign n7328 = pi14 ? n6961 : n6965;
  assign n7329 = pi17 ? n2653 : ~n2726;
  assign n7330 = pi16 ? n32 : n7329;
  assign n7331 = pi15 ? n7330 : n6548;
  assign n7332 = pi14 ? n7331 : n6548;
  assign n7333 = pi13 ? n7328 : n7332;
  assign n7334 = pi12 ? n7327 : n7333;
  assign n7335 = pi17 ? n2305 : ~n3067;
  assign n7336 = pi16 ? n32 : n7335;
  assign n7337 = pi15 ? n6770 : n7336;
  assign n7338 = pi14 ? n6766 : n7337;
  assign n7339 = pi17 ? n1933 : ~n2750;
  assign n7340 = pi16 ? n32 : n7339;
  assign n7341 = pi17 ? n2319 : ~n2750;
  assign n7342 = pi16 ? n32 : n7341;
  assign n7343 = pi15 ? n7340 : n7342;
  assign n7344 = pi14 ? n6772 : n7343;
  assign n7345 = pi13 ? n7338 : n7344;
  assign n7346 = pi17 ? n2537 : ~n6768;
  assign n7347 = pi16 ? n32 : n7346;
  assign n7348 = pi15 ? n7347 : n6554;
  assign n7349 = pi20 ? n428 : ~n207;
  assign n7350 = pi19 ? n32 : ~n7349;
  assign n7351 = pi18 ? n32 : n7350;
  assign n7352 = pi17 ? n1807 : ~n7351;
  assign n7353 = pi16 ? n32 : n7352;
  assign n7354 = pi17 ? n1807 : ~n2750;
  assign n7355 = pi16 ? n32 : n7354;
  assign n7356 = pi15 ? n7353 : n7355;
  assign n7357 = pi14 ? n7348 : n7356;
  assign n7358 = pi17 ? n1807 : ~n2519;
  assign n7359 = pi16 ? n32 : n7358;
  assign n7360 = pi17 ? n1814 : ~n2519;
  assign n7361 = pi16 ? n32 : n7360;
  assign n7362 = pi15 ? n7359 : n7361;
  assign n7363 = pi20 ? n342 : ~n274;
  assign n7364 = pi19 ? n32 : n7363;
  assign n7365 = pi18 ? n32 : n7364;
  assign n7366 = pi17 ? n1814 : ~n7365;
  assign n7367 = pi16 ? n32 : n7366;
  assign n7368 = pi19 ? n32 : n5435;
  assign n7369 = pi18 ? n32 : n7368;
  assign n7370 = pi17 ? n1814 : ~n7369;
  assign n7371 = pi16 ? n32 : n7370;
  assign n7372 = pi15 ? n7367 : n7371;
  assign n7373 = pi14 ? n7362 : n7372;
  assign n7374 = pi13 ? n7357 : n7373;
  assign n7375 = pi12 ? n7345 : n7374;
  assign n7376 = pi11 ? n7334 : n7375;
  assign n7377 = pi21 ? n32 : n1009;
  assign n7378 = pi20 ? n7377 : n1940;
  assign n7379 = pi19 ? n32 : n7378;
  assign n7380 = pi18 ? n32 : n7379;
  assign n7381 = pi17 ? n3351 : ~n7380;
  assign n7382 = pi16 ? n32 : n7381;
  assign n7383 = pi15 ? n6784 : n7382;
  assign n7384 = pi19 ? n32 : n7023;
  assign n7385 = pi18 ? n32 : n7384;
  assign n7386 = pi17 ? n3351 : ~n7385;
  assign n7387 = pi16 ? n32 : n7386;
  assign n7388 = pi21 ? n206 : ~n140;
  assign n7389 = pi20 ? n7388 : n481;
  assign n7390 = pi19 ? n32 : ~n7389;
  assign n7391 = pi18 ? n32 : n7390;
  assign n7392 = pi17 ? n2123 : ~n7391;
  assign n7393 = pi16 ? n32 : n7392;
  assign n7394 = pi15 ? n7387 : n7393;
  assign n7395 = pi14 ? n7383 : n7394;
  assign n7396 = pi18 ? n32 : n1758;
  assign n7397 = pi17 ? n2123 : ~n7396;
  assign n7398 = pi16 ? n32 : n7397;
  assign n7399 = pi20 ? n266 : ~n339;
  assign n7400 = pi19 ? n32 : ~n7399;
  assign n7401 = pi18 ? n32 : n7400;
  assign n7402 = pi17 ? n2123 : ~n7401;
  assign n7403 = pi16 ? n32 : n7402;
  assign n7404 = pi15 ? n7398 : n7403;
  assign n7405 = pi20 ? n206 : ~n339;
  assign n7406 = pi19 ? n32 : ~n7405;
  assign n7407 = pi18 ? n32 : n7406;
  assign n7408 = pi17 ? n1682 : ~n7407;
  assign n7409 = pi16 ? n32 : n7408;
  assign n7410 = pi22 ? n84 : ~n32;
  assign n7411 = pi21 ? n206 : ~n7410;
  assign n7412 = pi20 ? n7411 : n32;
  assign n7413 = pi19 ? n32 : ~n7412;
  assign n7414 = pi18 ? n32 : n7413;
  assign n7415 = pi17 ? n1682 : ~n7414;
  assign n7416 = pi16 ? n32 : n7415;
  assign n7417 = pi15 ? n7409 : n7416;
  assign n7418 = pi14 ? n7404 : n7417;
  assign n7419 = pi13 ? n7395 : n7418;
  assign n7420 = pi21 ? n174 : ~n35;
  assign n7421 = pi20 ? n7420 : n32;
  assign n7422 = pi19 ? n32 : ~n7421;
  assign n7423 = pi18 ? n32 : n7422;
  assign n7424 = pi17 ? n1682 : ~n7423;
  assign n7425 = pi16 ? n32 : n7424;
  assign n7426 = pi21 ? n206 : ~n35;
  assign n7427 = pi20 ? n7426 : n32;
  assign n7428 = pi19 ? n32 : ~n7427;
  assign n7429 = pi18 ? n32 : n7428;
  assign n7430 = pi17 ? n1682 : ~n7429;
  assign n7431 = pi16 ? n32 : n7430;
  assign n7432 = pi15 ? n7425 : n7431;
  assign n7433 = pi17 ? n1682 : ~n6768;
  assign n7434 = pi16 ? n32 : n7433;
  assign n7435 = pi20 ? n6621 : n32;
  assign n7436 = pi19 ? n32 : ~n7435;
  assign n7437 = pi18 ? n32 : n7436;
  assign n7438 = pi17 ? n1682 : ~n7437;
  assign n7439 = pi16 ? n32 : n7438;
  assign n7440 = pi15 ? n7434 : n7439;
  assign n7441 = pi14 ? n7432 : n7440;
  assign n7442 = pi21 ? n206 : ~n1939;
  assign n7443 = pi20 ? n7442 : n32;
  assign n7444 = pi19 ? n32 : ~n7443;
  assign n7445 = pi18 ? n32 : n7444;
  assign n7446 = pi17 ? n1580 : ~n7445;
  assign n7447 = pi16 ? n32 : n7446;
  assign n7448 = pi21 ? n206 : n51;
  assign n7449 = pi20 ? n7448 : n32;
  assign n7450 = pi19 ? n1464 : ~n7449;
  assign n7451 = pi18 ? n32 : n7450;
  assign n7452 = pi17 ? n1580 : ~n7451;
  assign n7453 = pi16 ? n32 : n7452;
  assign n7454 = pi15 ? n7447 : n7453;
  assign n7455 = pi19 ? n322 : ~n3692;
  assign n7456 = pi18 ? n32 : n7455;
  assign n7457 = pi17 ? n2143 : ~n7456;
  assign n7458 = pi16 ? n32 : n7457;
  assign n7459 = pi19 ? n1464 : n2317;
  assign n7460 = pi18 ? n32 : n7459;
  assign n7461 = pi17 ? n2143 : ~n7460;
  assign n7462 = pi16 ? n32 : n7461;
  assign n7463 = pi15 ? n7458 : n7462;
  assign n7464 = pi14 ? n7454 : n7463;
  assign n7465 = pi13 ? n7441 : n7464;
  assign n7466 = pi12 ? n7419 : n7465;
  assign n7467 = pi21 ? n206 : ~n242;
  assign n7468 = pi20 ? n7467 : n32;
  assign n7469 = pi19 ? n32 : ~n7468;
  assign n7470 = pi18 ? n32 : n7469;
  assign n7471 = pi17 ? n2143 : ~n7470;
  assign n7472 = pi16 ? n32 : n7471;
  assign n7473 = pi15 ? n7472 : n7185;
  assign n7474 = pi19 ? n1464 : ~n1757;
  assign n7475 = pi18 ? n32 : n7474;
  assign n7476 = pi17 ? n1833 : ~n7475;
  assign n7477 = pi16 ? n32 : n7476;
  assign n7478 = pi22 ? n173 : n34;
  assign n7479 = pi21 ? n7478 : ~n32;
  assign n7480 = pi20 ? n7479 : ~n32;
  assign n7481 = pi19 ? n32 : n7480;
  assign n7482 = pi18 ? n32 : n7481;
  assign n7483 = pi17 ? n6072 : ~n7482;
  assign n7484 = pi16 ? n32 : n7483;
  assign n7485 = pi15 ? n7477 : n7484;
  assign n7486 = pi14 ? n7473 : n7485;
  assign n7487 = pi21 ? n7107 : n32;
  assign n7488 = pi20 ? n7487 : n32;
  assign n7489 = pi19 ? n1464 : ~n7488;
  assign n7490 = pi18 ? n32 : n7489;
  assign n7491 = pi17 ? n1576 : ~n7490;
  assign n7492 = pi16 ? n32 : n7491;
  assign n7493 = pi19 ? n507 : ~n440;
  assign n7494 = pi18 ? n32 : n7493;
  assign n7495 = pi17 ? n1576 : ~n7494;
  assign n7496 = pi16 ? n32 : n7495;
  assign n7497 = pi15 ? n7492 : n7496;
  assign n7498 = pi17 ? n1682 : ~n7494;
  assign n7499 = pi16 ? n32 : n7498;
  assign n7500 = pi22 ? n173 : ~n50;
  assign n7501 = pi21 ? n7500 : n32;
  assign n7502 = pi20 ? n7501 : n32;
  assign n7503 = pi19 ? n507 : ~n7502;
  assign n7504 = pi18 ? n32 : n7503;
  assign n7505 = pi17 ? n1677 : ~n7504;
  assign n7506 = pi16 ? n32 : n7505;
  assign n7507 = pi15 ? n7499 : n7506;
  assign n7508 = pi14 ? n7497 : n7507;
  assign n7509 = pi13 ? n7486 : n7508;
  assign n7510 = pi19 ? n507 : ~n5626;
  assign n7511 = pi18 ? n32 : n7510;
  assign n7512 = pi17 ? n1677 : ~n7511;
  assign n7513 = pi16 ? n32 : n7512;
  assign n7514 = pi19 ? n1464 : n2614;
  assign n7515 = pi18 ? n32 : n7514;
  assign n7516 = pi17 ? n2123 : ~n7515;
  assign n7517 = pi16 ? n32 : n7516;
  assign n7518 = pi15 ? n7513 : n7517;
  assign n7519 = pi19 ? n507 : n1105;
  assign n7520 = pi18 ? n32 : n7519;
  assign n7521 = pi17 ? n2123 : ~n7520;
  assign n7522 = pi16 ? n32 : n7521;
  assign n7523 = pi17 ? n3351 : ~n2623;
  assign n7524 = pi16 ? n32 : n7523;
  assign n7525 = pi15 ? n7522 : n7524;
  assign n7526 = pi14 ? n7518 : n7525;
  assign n7527 = pi17 ? n3351 : ~n2750;
  assign n7528 = pi16 ? n32 : n7527;
  assign n7529 = pi17 ? n2325 : ~n2750;
  assign n7530 = pi16 ? n32 : n7529;
  assign n7531 = pi15 ? n7528 : n7530;
  assign n7532 = pi17 ? n1943 : ~n2512;
  assign n7533 = pi16 ? n32 : n7532;
  assign n7534 = pi19 ? n4280 : ~n32;
  assign n7535 = pi18 ? n32 : n7534;
  assign n7536 = pi17 ? n1943 : ~n7535;
  assign n7537 = pi16 ? n32 : n7536;
  assign n7538 = pi15 ? n7533 : n7537;
  assign n7539 = pi14 ? n7531 : n7538;
  assign n7540 = pi13 ? n7526 : n7539;
  assign n7541 = pi12 ? n7509 : n7540;
  assign n7542 = pi11 ? n7466 : n7541;
  assign n7543 = pi10 ? n7376 : n7542;
  assign n7544 = pi09 ? n7309 : n7543;
  assign n7545 = pi17 ? n3175 : ~n3067;
  assign n7546 = pi16 ? n32 : n7545;
  assign n7547 = pi15 ? n32 : n7546;
  assign n7548 = pi17 ? n2963 : ~n3067;
  assign n7549 = pi16 ? n32 : n7548;
  assign n7550 = pi15 ? n7546 : n7549;
  assign n7551 = pi14 ? n7547 : n7550;
  assign n7552 = pi13 ? n32 : n7551;
  assign n7553 = pi12 ? n32 : n7552;
  assign n7554 = pi11 ? n32 : n7553;
  assign n7555 = pi10 ? n32 : n7554;
  assign n7556 = pi17 ? n2831 : ~n2726;
  assign n7557 = pi16 ? n32 : n7556;
  assign n7558 = pi17 ? n2733 : ~n2726;
  assign n7559 = pi16 ? n32 : n7558;
  assign n7560 = pi15 ? n7557 : n7559;
  assign n7561 = pi17 ? n4245 : ~n2726;
  assign n7562 = pi16 ? n32 : n7561;
  assign n7563 = pi14 ? n7560 : n7562;
  assign n7564 = pi17 ? n2731 : ~n3067;
  assign n7565 = pi16 ? n32 : n7564;
  assign n7566 = pi15 ? n7129 : n7565;
  assign n7567 = pi17 ? n2736 : ~n3067;
  assign n7568 = pi16 ? n32 : n7567;
  assign n7569 = pi17 ? n2750 : ~n2733;
  assign n7570 = pi16 ? n32 : n7569;
  assign n7571 = pi15 ? n7568 : n7570;
  assign n7572 = pi14 ? n7566 : n7571;
  assign n7573 = pi13 ? n7563 : n7572;
  assign n7574 = pi14 ? n7141 : n7145;
  assign n7575 = pi17 ? n2519 : ~n2726;
  assign n7576 = pi16 ? n32 : n7575;
  assign n7577 = pi15 ? n7576 : n6533;
  assign n7578 = pi14 ? n7577 : n6536;
  assign n7579 = pi13 ? n7574 : n7578;
  assign n7580 = pi12 ? n7573 : n7579;
  assign n7581 = pi15 ? n6967 : n6545;
  assign n7582 = pi14 ? n6965 : n7581;
  assign n7583 = pi17 ? n2531 : ~n2750;
  assign n7584 = pi16 ? n32 : n7583;
  assign n7585 = pi17 ? n2299 : ~n2750;
  assign n7586 = pi16 ? n32 : n7585;
  assign n7587 = pi15 ? n7584 : n7586;
  assign n7588 = pi14 ? n6545 : n7587;
  assign n7589 = pi13 ? n7582 : n7588;
  assign n7590 = pi17 ? n2410 : ~n6768;
  assign n7591 = pi16 ? n32 : n7590;
  assign n7592 = pi15 ? n7591 : n6765;
  assign n7593 = pi17 ? n2305 : ~n7351;
  assign n7594 = pi16 ? n32 : n7593;
  assign n7595 = pi17 ? n2305 : ~n2750;
  assign n7596 = pi16 ? n32 : n7595;
  assign n7597 = pi15 ? n7594 : n7596;
  assign n7598 = pi14 ? n7592 : n7597;
  assign n7599 = pi17 ? n2305 : ~n2519;
  assign n7600 = pi16 ? n32 : n7599;
  assign n7601 = pi17 ? n1933 : ~n2519;
  assign n7602 = pi16 ? n32 : n7601;
  assign n7603 = pi15 ? n7600 : n7602;
  assign n7604 = pi20 ? n428 : ~n274;
  assign n7605 = pi19 ? n32 : n7604;
  assign n7606 = pi18 ? n32 : n7605;
  assign n7607 = pi17 ? n1933 : ~n7606;
  assign n7608 = pi16 ? n32 : n7607;
  assign n7609 = pi17 ? n1933 : ~n7369;
  assign n7610 = pi16 ? n32 : n7609;
  assign n7611 = pi15 ? n7608 : n7610;
  assign n7612 = pi14 ? n7603 : n7611;
  assign n7613 = pi13 ? n7598 : n7612;
  assign n7614 = pi12 ? n7589 : n7613;
  assign n7615 = pi11 ? n7580 : n7614;
  assign n7616 = pi20 ? n3523 : n1940;
  assign n7617 = pi19 ? n32 : n7616;
  assign n7618 = pi18 ? n32 : n7617;
  assign n7619 = pi17 ? n2537 : ~n7618;
  assign n7620 = pi16 ? n32 : n7619;
  assign n7621 = pi15 ? n6973 : n7620;
  assign n7622 = pi20 ? n1324 : n339;
  assign n7623 = pi19 ? n32 : n7622;
  assign n7624 = pi18 ? n32 : n7623;
  assign n7625 = pi17 ? n2537 : ~n7624;
  assign n7626 = pi16 ? n32 : n7625;
  assign n7627 = pi20 ? n1685 : n481;
  assign n7628 = pi19 ? n32 : ~n7627;
  assign n7629 = pi18 ? n32 : n7628;
  assign n7630 = pi17 ? n3337 : ~n7629;
  assign n7631 = pi16 ? n32 : n7630;
  assign n7632 = pi15 ? n7626 : n7631;
  assign n7633 = pi14 ? n7621 : n7632;
  assign n7634 = pi17 ? n3337 : ~n7396;
  assign n7635 = pi16 ? n32 : n7634;
  assign n7636 = pi20 ? n1685 : ~n339;
  assign n7637 = pi19 ? n32 : ~n7636;
  assign n7638 = pi18 ? n32 : n7637;
  assign n7639 = pi17 ? n3337 : ~n7638;
  assign n7640 = pi16 ? n32 : n7639;
  assign n7641 = pi15 ? n7635 : n7640;
  assign n7642 = pi20 ? n206 : n32;
  assign n7643 = pi19 ? n32 : ~n7642;
  assign n7644 = pi18 ? n32 : n7643;
  assign n7645 = pi17 ? n1943 : ~n7644;
  assign n7646 = pi16 ? n32 : n7645;
  assign n7647 = pi19 ? n32 : ~n3692;
  assign n7648 = pi18 ? n32 : n7647;
  assign n7649 = pi17 ? n1943 : ~n7648;
  assign n7650 = pi16 ? n32 : n7649;
  assign n7651 = pi15 ? n7646 : n7650;
  assign n7652 = pi14 ? n7641 : n7651;
  assign n7653 = pi13 ? n7633 : n7652;
  assign n7654 = pi17 ? n1943 : ~n7423;
  assign n7655 = pi16 ? n32 : n7654;
  assign n7656 = pi20 ? n1940 : ~n428;
  assign n7657 = pi19 ? n7656 : ~n32;
  assign n7658 = pi18 ? n32 : n7657;
  assign n7659 = pi22 ? n34 : n173;
  assign n7660 = pi21 ? n206 : ~n7659;
  assign n7661 = pi20 ? n7660 : n32;
  assign n7662 = pi19 ? n32 : ~n7661;
  assign n7663 = pi18 ? n32 : n7662;
  assign n7664 = pi17 ? n7658 : ~n7663;
  assign n7665 = pi16 ? n32 : n7664;
  assign n7666 = pi15 ? n7655 : n7665;
  assign n7667 = pi20 ? n1940 : ~n342;
  assign n7668 = pi19 ? n7667 : ~n32;
  assign n7669 = pi18 ? n32 : n7668;
  assign n7670 = pi17 ? n7669 : ~n6768;
  assign n7671 = pi16 ? n32 : n7670;
  assign n7672 = pi19 ? n32 : ~n7449;
  assign n7673 = pi18 ? n32 : n7672;
  assign n7674 = pi17 ? n7658 : ~n7673;
  assign n7675 = pi16 ? n32 : n7674;
  assign n7676 = pi15 ? n7671 : n7675;
  assign n7677 = pi14 ? n7666 : n7676;
  assign n7678 = pi17 ? n1677 : ~n7445;
  assign n7679 = pi16 ? n32 : n7678;
  assign n7680 = pi17 ? n3351 : ~n7475;
  assign n7681 = pi16 ? n32 : n7680;
  assign n7682 = pi15 ? n7679 : n7681;
  assign n7683 = pi17 ? n3351 : ~n7456;
  assign n7684 = pi16 ? n32 : n7683;
  assign n7685 = pi19 ? n322 : n2317;
  assign n7686 = pi18 ? n32 : n7685;
  assign n7687 = pi17 ? n2123 : ~n7686;
  assign n7688 = pi16 ? n32 : n7687;
  assign n7689 = pi15 ? n7684 : n7688;
  assign n7690 = pi14 ? n7682 : n7689;
  assign n7691 = pi13 ? n7677 : n7690;
  assign n7692 = pi12 ? n7653 : n7691;
  assign n7693 = pi20 ? n7388 : n32;
  assign n7694 = pi19 ? n32 : ~n7693;
  assign n7695 = pi18 ? n32 : n7694;
  assign n7696 = pi17 ? n2123 : ~n7695;
  assign n7697 = pi16 ? n32 : n7696;
  assign n7698 = pi17 ? n3351 : ~n2850;
  assign n7699 = pi16 ? n32 : n7698;
  assign n7700 = pi15 ? n7697 : n7699;
  assign n7701 = pi19 ? n2614 : ~n4491;
  assign n7702 = pi18 ? n32 : n7701;
  assign n7703 = pi19 ? n32 : ~n7488;
  assign n7704 = pi18 ? n32 : n7703;
  assign n7705 = pi17 ? n7702 : ~n7704;
  assign n7706 = pi16 ? n32 : n7705;
  assign n7707 = pi15 ? n7681 : n7706;
  assign n7708 = pi14 ? n7700 : n7707;
  assign n7709 = pi17 ? n2325 : ~n7490;
  assign n7710 = pi16 ? n32 : n7709;
  assign n7711 = pi17 ? n2136 : ~n7494;
  assign n7712 = pi16 ? n32 : n7711;
  assign n7713 = pi15 ? n7710 : n7712;
  assign n7714 = pi17 ? n2136 : ~n7511;
  assign n7715 = pi16 ? n32 : n7714;
  assign n7716 = pi15 ? n7712 : n7715;
  assign n7717 = pi14 ? n7713 : n7716;
  assign n7718 = pi13 ? n7708 : n7717;
  assign n7719 = pi17 ? n1814 : ~n7515;
  assign n7720 = pi16 ? n32 : n7719;
  assign n7721 = pi15 ? n7715 : n7720;
  assign n7722 = pi17 ? n1814 : ~n7520;
  assign n7723 = pi16 ? n32 : n7722;
  assign n7724 = pi17 ? n1807 : ~n2623;
  assign n7725 = pi16 ? n32 : n7724;
  assign n7726 = pi15 ? n7723 : n7725;
  assign n7727 = pi14 ? n7721 : n7726;
  assign n7728 = pi17 ? n2537 : ~n2750;
  assign n7729 = pi16 ? n32 : n7728;
  assign n7730 = pi17 ? n2537 : ~n2512;
  assign n7731 = pi16 ? n32 : n7730;
  assign n7732 = pi17 ? n2537 : ~n7535;
  assign n7733 = pi16 ? n32 : n7732;
  assign n7734 = pi15 ? n7731 : n7733;
  assign n7735 = pi14 ? n7729 : n7734;
  assign n7736 = pi13 ? n7727 : n7735;
  assign n7737 = pi12 ? n7718 : n7736;
  assign n7738 = pi11 ? n7692 : n7737;
  assign n7739 = pi10 ? n7615 : n7738;
  assign n7740 = pi09 ? n7555 : n7739;
  assign n7741 = pi08 ? n7544 : n7740;
  assign n7742 = pi17 ? n3164 : ~n3067;
  assign n7743 = pi16 ? n32 : n7742;
  assign n7744 = pi15 ? n32 : n7743;
  assign n7745 = pi17 ? n3046 : ~n3067;
  assign n7746 = pi16 ? n32 : n7745;
  assign n7747 = pi17 ? n3292 : ~n3067;
  assign n7748 = pi16 ? n32 : n7747;
  assign n7749 = pi15 ? n7746 : n7748;
  assign n7750 = pi14 ? n7744 : n7749;
  assign n7751 = pi13 ? n32 : n7750;
  assign n7752 = pi12 ? n32 : n7751;
  assign n7753 = pi11 ? n32 : n7752;
  assign n7754 = pi10 ? n32 : n7753;
  assign n7755 = pi17 ? n2952 : ~n2726;
  assign n7756 = pi16 ? n32 : n7755;
  assign n7757 = pi17 ? n3175 : ~n2726;
  assign n7758 = pi16 ? n32 : n7757;
  assign n7759 = pi15 ? n7756 : n7758;
  assign n7760 = pi17 ? n2836 : ~n2726;
  assign n7761 = pi16 ? n32 : n7760;
  assign n7762 = pi14 ? n7759 : n7761;
  assign n7763 = pi17 ? n2839 : ~n3067;
  assign n7764 = pi16 ? n32 : n7763;
  assign n7765 = pi15 ? n7303 : n7764;
  assign n7766 = pi17 ? n2850 : ~n3067;
  assign n7767 = pi16 ? n32 : n7766;
  assign n7768 = pi17 ? n4245 : ~n2733;
  assign n7769 = pi16 ? n32 : n7768;
  assign n7770 = pi15 ? n7767 : n7769;
  assign n7771 = pi14 ? n7765 : n7770;
  assign n7772 = pi13 ? n7762 : n7771;
  assign n7773 = pi14 ? n7140 : n7320;
  assign n7774 = pi17 ? n2628 : ~n2726;
  assign n7775 = pi16 ? n32 : n7774;
  assign n7776 = pi15 ? n7775 : n6960;
  assign n7777 = pi14 ? n7776 : n6960;
  assign n7778 = pi13 ? n7773 : n7777;
  assign n7779 = pi12 ? n7772 : n7778;
  assign n7780 = pi17 ? n2519 : ~n3067;
  assign n7781 = pi16 ? n32 : n7780;
  assign n7782 = pi15 ? n7781 : n6760;
  assign n7783 = pi14 ? n7145 : n7782;
  assign n7784 = pi15 ? n6760 : n6533;
  assign n7785 = pi17 ? n2119 : ~n2750;
  assign n7786 = pi16 ? n32 : n7785;
  assign n7787 = pi15 ? n6530 : n7786;
  assign n7788 = pi14 ? n7784 : n7787;
  assign n7789 = pi13 ? n7783 : n7788;
  assign n7790 = pi17 ? n2425 : ~n7039;
  assign n7791 = pi16 ? n32 : n7790;
  assign n7792 = pi17 ? n3787 : ~n3067;
  assign n7793 = pi16 ? n32 : n7792;
  assign n7794 = pi15 ? n7791 : n7793;
  assign n7795 = pi20 ? n32 : ~n1839;
  assign n7796 = pi19 ? n32 : ~n7795;
  assign n7797 = pi18 ? n32 : n7796;
  assign n7798 = pi17 ? n3787 : ~n7797;
  assign n7799 = pi16 ? n32 : n7798;
  assign n7800 = pi17 ? n3787 : ~n2750;
  assign n7801 = pi16 ? n32 : n7800;
  assign n7802 = pi15 ? n7799 : n7801;
  assign n7803 = pi14 ? n7794 : n7802;
  assign n7804 = pi19 ? n322 : ~n275;
  assign n7805 = pi18 ? n32 : n7804;
  assign n7806 = pi17 ? n3787 : ~n7805;
  assign n7807 = pi16 ? n32 : n7806;
  assign n7808 = pi17 ? n2531 : ~n2519;
  assign n7809 = pi16 ? n32 : n7808;
  assign n7810 = pi15 ? n7807 : n7809;
  assign n7811 = pi17 ? n2531 : ~n7365;
  assign n7812 = pi16 ? n32 : n7811;
  assign n7813 = pi20 ? n246 : n749;
  assign n7814 = pi19 ? n32 : n7813;
  assign n7815 = pi18 ? n32 : n7814;
  assign n7816 = pi17 ? n2531 : ~n7815;
  assign n7817 = pi16 ? n32 : n7816;
  assign n7818 = pi15 ? n7812 : n7817;
  assign n7819 = pi14 ? n7810 : n7818;
  assign n7820 = pi13 ? n7803 : n7819;
  assign n7821 = pi12 ? n7789 : n7820;
  assign n7822 = pi11 ? n7779 : n7821;
  assign n7823 = pi20 ? n246 : n1940;
  assign n7824 = pi19 ? n32 : n7823;
  assign n7825 = pi18 ? n32 : n7824;
  assign n7826 = pi17 ? n2299 : ~n7825;
  assign n7827 = pi16 ? n32 : n7826;
  assign n7828 = pi15 ? n6548 : n7827;
  assign n7829 = pi20 ? n1331 : ~n243;
  assign n7830 = pi19 ? n32 : ~n7829;
  assign n7831 = pi18 ? n32 : n7830;
  assign n7832 = pi17 ? n2410 : ~n7831;
  assign n7833 = pi16 ? n32 : n7832;
  assign n7834 = pi15 ? n6548 : n7833;
  assign n7835 = pi14 ? n7828 : n7834;
  assign n7836 = pi18 ? n32 : n1845;
  assign n7837 = pi17 ? n2410 : ~n7836;
  assign n7838 = pi16 ? n32 : n7837;
  assign n7839 = pi21 ? n405 : ~n206;
  assign n7840 = pi20 ? n7839 : ~n339;
  assign n7841 = pi19 ? n32 : ~n7840;
  assign n7842 = pi18 ? n32 : n7841;
  assign n7843 = pi17 ? n2410 : ~n7842;
  assign n7844 = pi16 ? n32 : n7843;
  assign n7845 = pi15 ? n7838 : n7844;
  assign n7846 = pi21 ? n206 : n1392;
  assign n7847 = pi20 ? n7846 : n32;
  assign n7848 = pi19 ? n32 : ~n7847;
  assign n7849 = pi18 ? n32 : n7848;
  assign n7850 = pi17 ? n2537 : ~n7849;
  assign n7851 = pi16 ? n32 : n7850;
  assign n7852 = pi21 ? n405 : ~n242;
  assign n7853 = pi20 ? n7852 : n32;
  assign n7854 = pi19 ? n32 : ~n7853;
  assign n7855 = pi18 ? n32 : n7854;
  assign n7856 = pi17 ? n2319 : ~n7855;
  assign n7857 = pi16 ? n32 : n7856;
  assign n7858 = pi15 ? n7851 : n7857;
  assign n7859 = pi14 ? n7845 : n7858;
  assign n7860 = pi13 ? n7835 : n7859;
  assign n7861 = pi21 ? n206 : ~n1009;
  assign n7862 = pi20 ? n7861 : n32;
  assign n7863 = pi19 ? n32 : ~n7862;
  assign n7864 = pi18 ? n32 : n7863;
  assign n7865 = pi17 ? n2319 : ~n7864;
  assign n7866 = pi16 ? n32 : n7865;
  assign n7867 = pi17 ? n1933 : ~n7855;
  assign n7868 = pi16 ? n32 : n7867;
  assign n7869 = pi15 ? n7866 : n7868;
  assign n7870 = pi19 ? n2317 : ~n5614;
  assign n7871 = pi18 ? n32 : n7870;
  assign n7872 = pi17 ? n7871 : ~n6768;
  assign n7873 = pi16 ? n32 : n7872;
  assign n7874 = pi19 ? n343 : ~n5614;
  assign n7875 = pi18 ? n32 : n7874;
  assign n7876 = pi17 ? n7875 : ~n7836;
  assign n7877 = pi16 ? n32 : n7876;
  assign n7878 = pi15 ? n7873 : n7877;
  assign n7879 = pi14 ? n7869 : n7878;
  assign n7880 = pi21 ? n32 : ~n1939;
  assign n7881 = pi20 ? n7880 : n32;
  assign n7882 = pi19 ? n32 : ~n7881;
  assign n7883 = pi18 ? n32 : n7882;
  assign n7884 = pi17 ? n1807 : ~n7883;
  assign n7885 = pi16 ? n32 : n7884;
  assign n7886 = pi17 ? n1807 : ~n7475;
  assign n7887 = pi16 ? n32 : n7886;
  assign n7888 = pi15 ? n7885 : n7887;
  assign n7889 = pi19 ? n322 : ~n247;
  assign n7890 = pi18 ? n32 : n7889;
  assign n7891 = pi17 ? n1807 : ~n7890;
  assign n7892 = pi16 ? n32 : n7891;
  assign n7893 = pi17 ? n1814 : ~n7460;
  assign n7894 = pi16 ? n32 : n7893;
  assign n7895 = pi15 ? n7892 : n7894;
  assign n7896 = pi14 ? n7888 : n7895;
  assign n7897 = pi13 ? n7879 : n7896;
  assign n7898 = pi12 ? n7860 : n7897;
  assign n7899 = pi19 ? n857 : ~n1757;
  assign n7900 = pi18 ? n32 : n7899;
  assign n7901 = pi17 ? n1814 : ~n7900;
  assign n7902 = pi16 ? n32 : n7901;
  assign n7903 = pi17 ? n1807 : ~n2850;
  assign n7904 = pi16 ? n32 : n7903;
  assign n7905 = pi15 ? n7902 : n7904;
  assign n7906 = pi17 ? n2537 : ~n7490;
  assign n7907 = pi16 ? n32 : n7906;
  assign n7908 = pi17 ? n2537 : ~n4245;
  assign n7909 = pi16 ? n32 : n7908;
  assign n7910 = pi15 ? n7907 : n7909;
  assign n7911 = pi14 ? n7905 : n7910;
  assign n7912 = pi19 ? n1464 : ~n5614;
  assign n7913 = pi18 ? n32 : n7912;
  assign n7914 = pi17 ? n2319 : ~n7913;
  assign n7915 = pi16 ? n32 : n7914;
  assign n7916 = pi17 ? n2319 : ~n7494;
  assign n7917 = pi16 ? n32 : n7916;
  assign n7918 = pi15 ? n7915 : n7917;
  assign n7919 = pi17 ? n2319 : ~n2512;
  assign n7920 = pi16 ? n32 : n7919;
  assign n7921 = pi19 ? n507 : n617;
  assign n7922 = pi18 ? n32 : n7921;
  assign n7923 = pi17 ? n2319 : ~n7922;
  assign n7924 = pi16 ? n32 : n7923;
  assign n7925 = pi15 ? n7920 : n7924;
  assign n7926 = pi14 ? n7918 : n7925;
  assign n7927 = pi13 ? n7911 : n7926;
  assign n7928 = pi17 ? n2319 : ~n7511;
  assign n7929 = pi16 ? n32 : n7928;
  assign n7930 = pi19 ? n1464 : n617;
  assign n7931 = pi18 ? n32 : n7930;
  assign n7932 = pi17 ? n1933 : ~n7931;
  assign n7933 = pi16 ? n32 : n7932;
  assign n7934 = pi15 ? n7929 : n7933;
  assign n7935 = pi17 ? n2410 : ~n2512;
  assign n7936 = pi16 ? n32 : n7935;
  assign n7937 = pi15 ? n7936 : n7586;
  assign n7938 = pi14 ? n7934 : n7937;
  assign n7939 = pi21 ? n259 : n206;
  assign n7940 = pi20 ? n7939 : n207;
  assign n7941 = pi19 ? n32 : ~n7940;
  assign n7942 = pi21 ? n173 : ~n206;
  assign n7943 = pi20 ? n7942 : n342;
  assign n7944 = pi19 ? n7943 : ~n32;
  assign n7945 = pi18 ? n7941 : n7944;
  assign n7946 = pi17 ? n2299 : ~n7945;
  assign n7947 = pi16 ? n32 : n7946;
  assign n7948 = pi15 ? n7586 : n7947;
  assign n7949 = pi17 ? n2299 : ~n2512;
  assign n7950 = pi16 ? n32 : n7949;
  assign n7951 = pi14 ? n7948 : n7950;
  assign n7952 = pi13 ? n7938 : n7951;
  assign n7953 = pi12 ? n7927 : n7952;
  assign n7954 = pi11 ? n7898 : n7953;
  assign n7955 = pi10 ? n7822 : n7954;
  assign n7956 = pi09 ? n7754 : n7955;
  assign n7957 = pi17 ? n2954 : ~n3067;
  assign n7958 = pi16 ? n32 : n7957;
  assign n7959 = pi15 ? n32 : n7958;
  assign n7960 = pi17 ? n4111 : ~n3067;
  assign n7961 = pi16 ? n32 : n7960;
  assign n7962 = pi15 ? n7958 : n7961;
  assign n7963 = pi14 ? n7959 : n7962;
  assign n7964 = pi13 ? n32 : n7963;
  assign n7965 = pi12 ? n32 : n7964;
  assign n7966 = pi11 ? n32 : n7965;
  assign n7967 = pi10 ? n32 : n7966;
  assign n7968 = pi17 ? n3160 : ~n2726;
  assign n7969 = pi16 ? n32 : n7968;
  assign n7970 = pi17 ? n3164 : ~n2726;
  assign n7971 = pi16 ? n32 : n7970;
  assign n7972 = pi15 ? n7969 : n7971;
  assign n7973 = pi17 ? n2726 : ~n2726;
  assign n7974 = pi16 ? n32 : n7973;
  assign n7975 = pi14 ? n7972 : n7974;
  assign n7976 = pi17 ? n2726 : ~n3067;
  assign n7977 = pi16 ? n32 : n7976;
  assign n7978 = pi17 ? n3182 : ~n3067;
  assign n7979 = pi16 ? n32 : n7978;
  assign n7980 = pi15 ? n7977 : n7979;
  assign n7981 = pi17 ? n2836 : ~n2733;
  assign n7982 = pi16 ? n32 : n7981;
  assign n7983 = pi15 ? n7300 : n7982;
  assign n7984 = pi14 ? n7980 : n7983;
  assign n7985 = pi13 ? n7975 : n7984;
  assign n7986 = pi14 ? n7127 : n7566;
  assign n7987 = pi17 ? n2736 : ~n2726;
  assign n7988 = pi16 ? n32 : n7987;
  assign n7989 = pi15 ? n7988 : n7140;
  assign n7990 = pi14 ? n7989 : n7140;
  assign n7991 = pi13 ? n7986 : n7990;
  assign n7992 = pi12 ? n7985 : n7991;
  assign n7993 = pi20 ? n321 : n141;
  assign n7994 = pi19 ? n32 : n7993;
  assign n7995 = pi18 ? n32 : n7994;
  assign n7996 = pi17 ? n2618 : ~n7995;
  assign n7997 = pi16 ? n32 : n7996;
  assign n7998 = pi15 ? n7140 : n7997;
  assign n7999 = pi15 ? n7322 : n6748;
  assign n8000 = pi14 ? n7998 : n7999;
  assign n8001 = pi17 ? n2517 : ~n2750;
  assign n8002 = pi16 ? n32 : n8001;
  assign n8003 = pi15 ? n6745 : n8002;
  assign n8004 = pi14 ? n6748 : n8003;
  assign n8005 = pi13 ? n8000 : n8004;
  assign n8006 = pi20 ? n246 : ~n160;
  assign n8007 = pi19 ? n32 : n8006;
  assign n8008 = pi18 ? n32 : n8007;
  assign n8009 = pi17 ? n2755 : ~n8008;
  assign n8010 = pi16 ? n32 : n8009;
  assign n8011 = pi17 ? n2292 : ~n3067;
  assign n8012 = pi16 ? n32 : n8011;
  assign n8013 = pi15 ? n8010 : n8012;
  assign n8014 = pi17 ? n2292 : ~n7797;
  assign n8015 = pi16 ? n32 : n8014;
  assign n8016 = pi17 ? n2408 : ~n2750;
  assign n8017 = pi16 ? n32 : n8016;
  assign n8018 = pi15 ? n8015 : n8017;
  assign n8019 = pi14 ? n8013 : n8018;
  assign n8020 = pi17 ? n2408 : ~n7805;
  assign n8021 = pi16 ? n32 : n8020;
  assign n8022 = pi17 ? n2414 : ~n2519;
  assign n8023 = pi16 ? n32 : n8022;
  assign n8024 = pi15 ? n8021 : n8023;
  assign n8025 = pi17 ? n2414 : ~n7365;
  assign n8026 = pi16 ? n32 : n8025;
  assign n8027 = pi17 ? n2425 : ~n7825;
  assign n8028 = pi16 ? n32 : n8027;
  assign n8029 = pi15 ? n8026 : n8028;
  assign n8030 = pi14 ? n8024 : n8029;
  assign n8031 = pi13 ? n8019 : n8030;
  assign n8032 = pi12 ? n8005 : n8031;
  assign n8033 = pi11 ? n7992 : n8032;
  assign n8034 = pi15 ? n6964 : n8028;
  assign n8035 = pi20 ? n32 : ~n243;
  assign n8036 = pi19 ? n32 : ~n8035;
  assign n8037 = pi18 ? n32 : n8036;
  assign n8038 = pi17 ? n2653 : ~n8037;
  assign n8039 = pi16 ? n32 : n8038;
  assign n8040 = pi15 ? n6964 : n8039;
  assign n8041 = pi14 ? n8034 : n8040;
  assign n8042 = pi17 ? n2653 : ~n7836;
  assign n8043 = pi16 ? n32 : n8042;
  assign n8044 = pi20 ? n246 : ~n339;
  assign n8045 = pi19 ? n32 : ~n8044;
  assign n8046 = pi18 ? n32 : n8045;
  assign n8047 = pi17 ? n2653 : ~n8046;
  assign n8048 = pi16 ? n32 : n8047;
  assign n8049 = pi15 ? n8043 : n8048;
  assign n8050 = pi17 ? n3787 : ~n7849;
  assign n8051 = pi16 ? n32 : n8050;
  assign n8052 = pi19 ? n32 : ~n5597;
  assign n8053 = pi18 ? n32 : n8052;
  assign n8054 = pi17 ? n3787 : ~n8053;
  assign n8055 = pi16 ? n32 : n8054;
  assign n8056 = pi15 ? n8051 : n8055;
  assign n8057 = pi14 ? n8049 : n8056;
  assign n8058 = pi13 ? n8041 : n8057;
  assign n8059 = pi17 ? n3787 : ~n7864;
  assign n8060 = pi16 ? n32 : n8059;
  assign n8061 = pi17 ? n3787 : ~n7855;
  assign n8062 = pi16 ? n32 : n8061;
  assign n8063 = pi15 ? n8060 : n8062;
  assign n8064 = pi20 ? n6303 : n32;
  assign n8065 = pi19 ? n365 : ~n8064;
  assign n8066 = pi18 ? n32 : n8065;
  assign n8067 = pi17 ? n8066 : ~n6768;
  assign n8068 = pi16 ? n32 : n8067;
  assign n8069 = pi17 ? n8066 : ~n7836;
  assign n8070 = pi16 ? n32 : n8069;
  assign n8071 = pi15 ? n8068 : n8070;
  assign n8072 = pi14 ? n8063 : n8071;
  assign n8073 = pi17 ? n1933 : ~n7883;
  assign n8074 = pi16 ? n32 : n8073;
  assign n8075 = pi17 ? n2305 : ~n7475;
  assign n8076 = pi16 ? n32 : n8075;
  assign n8077 = pi15 ? n8074 : n8076;
  assign n8078 = pi17 ? n2305 : ~n7890;
  assign n8079 = pi16 ? n32 : n8078;
  assign n8080 = pi17 ? n2410 : ~n7030;
  assign n8081 = pi16 ? n32 : n8080;
  assign n8082 = pi15 ? n8079 : n8081;
  assign n8083 = pi14 ? n8077 : n8082;
  assign n8084 = pi13 ? n8072 : n8083;
  assign n8085 = pi12 ? n8058 : n8084;
  assign n8086 = pi19 ? n507 : ~n1757;
  assign n8087 = pi18 ? n32 : n8086;
  assign n8088 = pi17 ? n2299 : ~n8087;
  assign n8089 = pi16 ? n32 : n8088;
  assign n8090 = pi17 ? n2299 : ~n2850;
  assign n8091 = pi16 ? n32 : n8090;
  assign n8092 = pi15 ? n8089 : n8091;
  assign n8093 = pi17 ? n2299 : ~n7490;
  assign n8094 = pi16 ? n32 : n8093;
  assign n8095 = pi17 ? n2299 : ~n4245;
  assign n8096 = pi16 ? n32 : n8095;
  assign n8097 = pi15 ? n8094 : n8096;
  assign n8098 = pi14 ? n8092 : n8097;
  assign n8099 = pi17 ? n2299 : ~n7913;
  assign n8100 = pi16 ? n32 : n8099;
  assign n8101 = pi17 ? n2299 : ~n7494;
  assign n8102 = pi16 ? n32 : n8101;
  assign n8103 = pi15 ? n8100 : n8102;
  assign n8104 = pi17 ? n2531 : ~n7511;
  assign n8105 = pi16 ? n32 : n8104;
  assign n8106 = pi19 ? n857 : n32;
  assign n8107 = pi18 ? n8106 : n7921;
  assign n8108 = pi17 ? n2531 : ~n8107;
  assign n8109 = pi16 ? n32 : n8108;
  assign n8110 = pi15 ? n8105 : n8109;
  assign n8111 = pi14 ? n8103 : n8110;
  assign n8112 = pi13 ? n8098 : n8111;
  assign n8113 = pi17 ? n2653 : ~n7511;
  assign n8114 = pi16 ? n32 : n8113;
  assign n8115 = pi17 ? n2425 : ~n7931;
  assign n8116 = pi16 ? n32 : n8115;
  assign n8117 = pi15 ? n8114 : n8116;
  assign n8118 = pi17 ? n2653 : ~n2512;
  assign n8119 = pi16 ? n32 : n8118;
  assign n8120 = pi17 ? n2425 : ~n2750;
  assign n8121 = pi16 ? n32 : n8120;
  assign n8122 = pi15 ? n8119 : n8121;
  assign n8123 = pi14 ? n8117 : n8122;
  assign n8124 = pi17 ? n2425 : ~n2618;
  assign n8125 = pi16 ? n32 : n8124;
  assign n8126 = pi19 ? n208 : ~n4491;
  assign n8127 = pi18 ? n32 : n8126;
  assign n8128 = pi20 ? n7839 : n342;
  assign n8129 = pi19 ? n8128 : ~n32;
  assign n8130 = pi18 ? n7941 : n8129;
  assign n8131 = pi17 ? n8127 : ~n8130;
  assign n8132 = pi16 ? n32 : n8131;
  assign n8133 = pi15 ? n8125 : n8132;
  assign n8134 = pi17 ? n2119 : ~n7535;
  assign n8135 = pi16 ? n32 : n8134;
  assign n8136 = pi17 ? n2408 : ~n2512;
  assign n8137 = pi16 ? n32 : n8136;
  assign n8138 = pi15 ? n8135 : n8137;
  assign n8139 = pi14 ? n8133 : n8138;
  assign n8140 = pi13 ? n8123 : n8139;
  assign n8141 = pi12 ? n8112 : n8140;
  assign n8142 = pi11 ? n8085 : n8141;
  assign n8143 = pi10 ? n8033 : n8142;
  assign n8144 = pi09 ? n7967 : n8143;
  assign n8145 = pi08 ? n7956 : n8144;
  assign n8146 = pi07 ? n7741 : n8145;
  assign n8147 = pi06 ? n7298 : n8146;
  assign n8148 = pi18 ? n1676 : ~n6978;
  assign n8149 = pi17 ? n32 : n8148;
  assign n8150 = pi16 ? n32 : n8149;
  assign n8151 = pi15 ? n32 : n8150;
  assign n8152 = pi17 ? n3569 : ~n3067;
  assign n8153 = pi16 ? n32 : n8152;
  assign n8154 = pi19 ? n267 : n236;
  assign n8155 = pi18 ? n32 : n8154;
  assign n8156 = pi17 ? n3569 : ~n8155;
  assign n8157 = pi16 ? n32 : n8156;
  assign n8158 = pi15 ? n8153 : n8157;
  assign n8159 = pi14 ? n8151 : n8158;
  assign n8160 = pi13 ? n32 : n8159;
  assign n8161 = pi12 ? n32 : n8160;
  assign n8162 = pi11 ? n32 : n8161;
  assign n8163 = pi10 ? n32 : n8162;
  assign n8164 = pi17 ? n3282 : ~n3067;
  assign n8165 = pi16 ? n32 : n8164;
  assign n8166 = pi17 ? n3155 : ~n3067;
  assign n8167 = pi16 ? n32 : n8166;
  assign n8168 = pi15 ? n8165 : n8167;
  assign n8169 = pi17 ? n3046 : ~n2726;
  assign n8170 = pi16 ? n32 : n8169;
  assign n8171 = pi14 ? n8168 : n8170;
  assign n8172 = pi17 ? n3587 : ~n3067;
  assign n8173 = pi16 ? n32 : n8172;
  assign n8174 = pi15 ? n7748 : n8173;
  assign n8175 = pi15 ? n7546 : n7977;
  assign n8176 = pi14 ? n8174 : n8175;
  assign n8177 = pi13 ? n8171 : n8176;
  assign n8178 = pi14 ? n7761 : n7765;
  assign n8179 = pi17 ? n2850 : ~n2726;
  assign n8180 = pi16 ? n32 : n8179;
  assign n8181 = pi15 ? n8180 : n7562;
  assign n8182 = pi14 ? n8181 : n7562;
  assign n8183 = pi13 ? n8178 : n8182;
  assign n8184 = pi12 ? n8177 : n8183;
  assign n8185 = pi20 ? n1324 : ~n1817;
  assign n8186 = pi19 ? n32 : n8185;
  assign n8187 = pi18 ? n32 : n8186;
  assign n8188 = pi17 ? n2623 : ~n8187;
  assign n8189 = pi16 ? n32 : n8188;
  assign n8190 = pi15 ? n7568 : n8189;
  assign n8191 = pi14 ? n7566 : n8190;
  assign n8192 = pi19 ? n32 : n321;
  assign n8193 = pi18 ? n32 : n8192;
  assign n8194 = pi17 ? n2623 : ~n8193;
  assign n8195 = pi16 ? n32 : n8194;
  assign n8196 = pi20 ? n321 : n518;
  assign n8197 = pi19 ? n32 : n8196;
  assign n8198 = pi18 ? n32 : n8197;
  assign n8199 = pi17 ? n2623 : ~n8198;
  assign n8200 = pi16 ? n32 : n8199;
  assign n8201 = pi15 ? n8195 : n8200;
  assign n8202 = pi20 ? n1385 : n321;
  assign n8203 = pi19 ? n32 : n8202;
  assign n8204 = pi18 ? n32 : n8203;
  assign n8205 = pi17 ? n2623 : ~n8204;
  assign n8206 = pi16 ? n32 : n8205;
  assign n8207 = pi17 ? n4099 : ~n8198;
  assign n8208 = pi16 ? n32 : n8207;
  assign n8209 = pi15 ? n8206 : n8208;
  assign n8210 = pi14 ? n8201 : n8209;
  assign n8211 = pi13 ? n8191 : n8210;
  assign n8212 = pi20 ? n321 : n1839;
  assign n8213 = pi19 ? n32 : n8212;
  assign n8214 = pi18 ? n32 : n8213;
  assign n8215 = pi17 ? n2618 : ~n8214;
  assign n8216 = pi16 ? n32 : n8215;
  assign n8217 = pi17 ? n2628 : ~n8193;
  assign n8218 = pi16 ? n32 : n8217;
  assign n8219 = pi15 ? n8216 : n8218;
  assign n8220 = pi20 ? n321 : ~n274;
  assign n8221 = pi19 ? n32 : n8220;
  assign n8222 = pi18 ? n32 : n8221;
  assign n8223 = pi17 ? n2628 : ~n8222;
  assign n8224 = pi16 ? n32 : n8223;
  assign n8225 = pi15 ? n8224 : n7322;
  assign n8226 = pi14 ? n8219 : n8225;
  assign n8227 = pi17 ? n2748 : ~n2959;
  assign n8228 = pi16 ? n32 : n8227;
  assign n8229 = pi15 ? n8224 : n8228;
  assign n8230 = pi20 ? n1324 : n207;
  assign n8231 = pi19 ? n32 : n8230;
  assign n8232 = pi18 ? n32 : n8231;
  assign n8233 = pi17 ? n2748 : ~n8232;
  assign n8234 = pi16 ? n32 : n8233;
  assign n8235 = pi20 ? n32 : ~n52;
  assign n8236 = pi19 ? n32 : n8235;
  assign n8237 = pi18 ? n32 : n8236;
  assign n8238 = pi17 ? n2755 : ~n8237;
  assign n8239 = pi16 ? n32 : n8238;
  assign n8240 = pi15 ? n8234 : n8239;
  assign n8241 = pi14 ? n8229 : n8240;
  assign n8242 = pi13 ? n8226 : n8241;
  assign n8243 = pi12 ? n8211 : n8242;
  assign n8244 = pi11 ? n8184 : n8243;
  assign n8245 = pi17 ? n2755 : ~n7369;
  assign n8246 = pi16 ? n32 : n8245;
  assign n8247 = pi20 ? n321 : n243;
  assign n8248 = pi19 ? n32 : n8247;
  assign n8249 = pi18 ? n32 : n8248;
  assign n8250 = pi17 ? n2519 : ~n8249;
  assign n8251 = pi16 ? n32 : n8250;
  assign n8252 = pi15 ? n8246 : n8251;
  assign n8253 = pi19 ? n32 : ~n6420;
  assign n8254 = pi18 ? n32 : n8253;
  assign n8255 = pi17 ? n2292 : ~n8254;
  assign n8256 = pi16 ? n32 : n8255;
  assign n8257 = pi15 ? n7576 : n8256;
  assign n8258 = pi14 ? n8252 : n8257;
  assign n8259 = pi19 ? n32 : ~n5614;
  assign n8260 = pi18 ? n32 : n8259;
  assign n8261 = pi17 ? n2292 : ~n8260;
  assign n8262 = pi16 ? n32 : n8261;
  assign n8263 = pi17 ? n2414 : ~n2726;
  assign n8264 = pi16 ? n32 : n8263;
  assign n8265 = pi15 ? n8262 : n8264;
  assign n8266 = pi19 ? n32 : n7008;
  assign n8267 = pi18 ? n32 : n8266;
  assign n8268 = pi17 ? n2414 : ~n8267;
  assign n8269 = pi16 ? n32 : n8268;
  assign n8270 = pi17 ? n2414 : ~n7039;
  assign n8271 = pi16 ? n32 : n8270;
  assign n8272 = pi15 ? n8269 : n8271;
  assign n8273 = pi14 ? n8265 : n8272;
  assign n8274 = pi13 ? n8258 : n8273;
  assign n8275 = pi22 ? n50 : n173;
  assign n8276 = pi21 ? n32 : n8275;
  assign n8277 = pi20 ? n8276 : ~n32;
  assign n8278 = pi19 ? n32 : n8277;
  assign n8279 = pi18 ? n32 : n8278;
  assign n8280 = pi17 ? n2414 : ~n8279;
  assign n8281 = pi16 ? n32 : n8280;
  assign n8282 = pi15 ? n8281 : n6533;
  assign n8283 = pi17 ? n2414 : ~n2831;
  assign n8284 = pi16 ? n32 : n8283;
  assign n8285 = pi21 ? n206 : n1939;
  assign n8286 = pi20 ? n8285 : ~n32;
  assign n8287 = pi19 ? n32 : n8286;
  assign n8288 = pi18 ? n32 : n8287;
  assign n8289 = pi17 ? n2414 : ~n8288;
  assign n8290 = pi16 ? n32 : n8289;
  assign n8291 = pi15 ? n8284 : n8290;
  assign n8292 = pi14 ? n8282 : n8291;
  assign n8293 = pi15 ? n7793 : n6535;
  assign n8294 = pi17 ? n2425 : ~n2850;
  assign n8295 = pi16 ? n32 : n8294;
  assign n8296 = pi15 ? n6535 : n8295;
  assign n8297 = pi14 ? n8293 : n8296;
  assign n8298 = pi13 ? n8292 : n8297;
  assign n8299 = pi12 ? n8274 : n8298;
  assign n8300 = pi19 ? n857 : n813;
  assign n8301 = pi18 ? n32 : n8300;
  assign n8302 = pi17 ? n2119 : ~n8301;
  assign n8303 = pi16 ? n32 : n8302;
  assign n8304 = pi17 ? n2425 : ~n2736;
  assign n8305 = pi16 ? n32 : n8304;
  assign n8306 = pi15 ? n8303 : n8305;
  assign n8307 = pi14 ? n6964 : n8306;
  assign n8308 = pi17 ? n2119 : ~n2724;
  assign n8309 = pi16 ? n32 : n8308;
  assign n8310 = pi17 ? n2119 : ~n2855;
  assign n8311 = pi16 ? n32 : n8310;
  assign n8312 = pi15 ? n8309 : n8311;
  assign n8313 = pi17 ? n2292 : ~n2616;
  assign n8314 = pi16 ? n32 : n8313;
  assign n8315 = pi17 ? n2292 : ~n2855;
  assign n8316 = pi16 ? n32 : n8315;
  assign n8317 = pi15 ? n8314 : n8316;
  assign n8318 = pi14 ? n8312 : n8317;
  assign n8319 = pi13 ? n8307 : n8318;
  assign n8320 = pi17 ? n2292 : ~n2750;
  assign n8321 = pi16 ? n32 : n8320;
  assign n8322 = pi15 ? n8316 : n8321;
  assign n8323 = pi18 ? n32 : n4581;
  assign n8324 = pi17 ? n2292 : ~n8323;
  assign n8325 = pi16 ? n32 : n8324;
  assign n8326 = pi17 ? n2519 : ~n2512;
  assign n8327 = pi16 ? n32 : n8326;
  assign n8328 = pi15 ? n8325 : n8327;
  assign n8329 = pi14 ? n8322 : n8328;
  assign n8330 = pi17 ? n2748 : ~n2512;
  assign n8331 = pi16 ? n32 : n8330;
  assign n8332 = pi15 ? n8327 : n8331;
  assign n8333 = pi17 ? n2517 : ~n2512;
  assign n8334 = pi16 ? n32 : n8333;
  assign n8335 = pi17 ? n2517 : ~n2637;
  assign n8336 = pi16 ? n32 : n8335;
  assign n8337 = pi15 ? n8334 : n8336;
  assign n8338 = pi14 ? n8332 : n8337;
  assign n8339 = pi13 ? n8329 : n8338;
  assign n8340 = pi12 ? n8319 : n8339;
  assign n8341 = pi11 ? n8299 : n8340;
  assign n8342 = pi10 ? n8244 : n8341;
  assign n8343 = pi09 ? n8163 : n8342;
  assign n8344 = pi18 ? n3350 : ~n6978;
  assign n8345 = pi17 ? n32 : n8344;
  assign n8346 = pi16 ? n32 : n8345;
  assign n8347 = pi15 ? n32 : n8346;
  assign n8348 = pi18 ? n3350 : ~n496;
  assign n8349 = pi17 ? n32 : n8348;
  assign n8350 = pi16 ? n32 : n8349;
  assign n8351 = pi18 ? n3350 : ~n8154;
  assign n8352 = pi17 ? n32 : n8351;
  assign n8353 = pi16 ? n32 : n8352;
  assign n8354 = pi15 ? n8350 : n8353;
  assign n8355 = pi14 ? n8347 : n8354;
  assign n8356 = pi13 ? n32 : n8355;
  assign n8357 = pi12 ? n32 : n8356;
  assign n8358 = pi11 ? n32 : n8357;
  assign n8359 = pi10 ? n32 : n8358;
  assign n8360 = pi18 ? n618 : ~n496;
  assign n8361 = pi17 ? n32 : n8360;
  assign n8362 = pi16 ? n32 : n8361;
  assign n8363 = pi15 ? n8362 : n8167;
  assign n8364 = pi17 ? n2954 : ~n2726;
  assign n8365 = pi16 ? n32 : n8364;
  assign n8366 = pi17 ? n3728 : ~n2726;
  assign n8367 = pi16 ? n32 : n8366;
  assign n8368 = pi15 ? n8365 : n8367;
  assign n8369 = pi14 ? n8363 : n8368;
  assign n8370 = pi17 ? n3728 : ~n3067;
  assign n8371 = pi16 ? n32 : n8370;
  assign n8372 = pi17 ? n3160 : ~n3067;
  assign n8373 = pi16 ? n32 : n8372;
  assign n8374 = pi15 ? n8371 : n8373;
  assign n8375 = pi15 ? n7743 : n7746;
  assign n8376 = pi14 ? n8374 : n8375;
  assign n8377 = pi13 ? n8369 : n8376;
  assign n8378 = pi14 ? n7974 : n7980;
  assign n8379 = pi15 ? n7559 : n7761;
  assign n8380 = pi14 ? n8379 : n7761;
  assign n8381 = pi13 ? n8378 : n8380;
  assign n8382 = pi12 ? n8377 : n8381;
  assign n8383 = pi20 ? n321 : ~n111;
  assign n8384 = pi19 ? n32 : n8383;
  assign n8385 = pi18 ? n32 : n8384;
  assign n8386 = pi17 ? n2836 : ~n8385;
  assign n8387 = pi16 ? n32 : n8386;
  assign n8388 = pi20 ? n321 : ~n125;
  assign n8389 = pi19 ? n32 : n8388;
  assign n8390 = pi18 ? n32 : n8389;
  assign n8391 = pi17 ? n2839 : ~n8390;
  assign n8392 = pi16 ? n32 : n8391;
  assign n8393 = pi15 ? n8387 : n8392;
  assign n8394 = pi17 ? n3067 : ~n8187;
  assign n8395 = pi16 ? n32 : n8394;
  assign n8396 = pi15 ? n7767 : n8395;
  assign n8397 = pi14 ? n8393 : n8396;
  assign n8398 = pi17 ? n3067 : ~n8193;
  assign n8399 = pi16 ? n32 : n8398;
  assign n8400 = pi17 ? n3067 : ~n8198;
  assign n8401 = pi16 ? n32 : n8400;
  assign n8402 = pi15 ? n8399 : n8401;
  assign n8403 = pi17 ? n4245 : ~n8204;
  assign n8404 = pi16 ? n32 : n8403;
  assign n8405 = pi17 ? n2724 : ~n8198;
  assign n8406 = pi16 ? n32 : n8405;
  assign n8407 = pi15 ? n8404 : n8406;
  assign n8408 = pi14 ? n8402 : n8407;
  assign n8409 = pi13 ? n8397 : n8408;
  assign n8410 = pi17 ? n2731 : ~n8214;
  assign n8411 = pi16 ? n32 : n8410;
  assign n8412 = pi17 ? n2855 : ~n8193;
  assign n8413 = pi16 ? n32 : n8412;
  assign n8414 = pi15 ? n8411 : n8413;
  assign n8415 = pi17 ? n2855 : ~n8222;
  assign n8416 = pi16 ? n32 : n8415;
  assign n8417 = pi17 ? n2855 : ~n3067;
  assign n8418 = pi16 ? n32 : n8417;
  assign n8419 = pi15 ? n8416 : n8418;
  assign n8420 = pi14 ? n8414 : n8419;
  assign n8421 = pi17 ? n2750 : ~n2959;
  assign n8422 = pi16 ? n32 : n8421;
  assign n8423 = pi15 ? n8416 : n8422;
  assign n8424 = pi17 ? n2750 : ~n8232;
  assign n8425 = pi16 ? n32 : n8424;
  assign n8426 = pi17 ? n4099 : ~n8237;
  assign n8427 = pi16 ? n32 : n8426;
  assign n8428 = pi15 ? n8425 : n8427;
  assign n8429 = pi14 ? n8423 : n8428;
  assign n8430 = pi13 ? n8420 : n8429;
  assign n8431 = pi12 ? n8409 : n8430;
  assign n8432 = pi11 ? n8382 : n8431;
  assign n8433 = pi17 ? n4099 : ~n7369;
  assign n8434 = pi16 ? n32 : n8433;
  assign n8435 = pi17 ? n4099 : ~n8249;
  assign n8436 = pi16 ? n32 : n8435;
  assign n8437 = pi15 ? n8434 : n8436;
  assign n8438 = pi17 ? n4099 : ~n2726;
  assign n8439 = pi16 ? n32 : n8438;
  assign n8440 = pi17 ? n2628 : ~n8254;
  assign n8441 = pi16 ? n32 : n8440;
  assign n8442 = pi15 ? n8439 : n8441;
  assign n8443 = pi14 ? n8437 : n8442;
  assign n8444 = pi17 ? n2628 : ~n8260;
  assign n8445 = pi16 ? n32 : n8444;
  assign n8446 = pi17 ? n2517 : ~n3175;
  assign n8447 = pi16 ? n32 : n8446;
  assign n8448 = pi15 ? n8445 : n8447;
  assign n8449 = pi17 ? n2748 : ~n2850;
  assign n8450 = pi16 ? n32 : n8449;
  assign n8451 = pi17 ? n2517 : ~n7039;
  assign n8452 = pi16 ? n32 : n8451;
  assign n8453 = pi15 ? n8450 : n8452;
  assign n8454 = pi14 ? n8448 : n8453;
  assign n8455 = pi13 ? n8443 : n8454;
  assign n8456 = pi17 ? n2517 : ~n6768;
  assign n8457 = pi16 ? n32 : n8456;
  assign n8458 = pi15 ? n8457 : n6750;
  assign n8459 = pi17 ? n2517 : ~n2831;
  assign n8460 = pi16 ? n32 : n8459;
  assign n8461 = pi17 ? n2519 : ~n8288;
  assign n8462 = pi16 ? n32 : n8461;
  assign n8463 = pi15 ? n8460 : n8462;
  assign n8464 = pi14 ? n8458 : n8463;
  assign n8465 = pi17 ? n2292 : ~n2850;
  assign n8466 = pi16 ? n32 : n8465;
  assign n8467 = pi15 ? n7781 : n8466;
  assign n8468 = pi14 ? n7781 : n8467;
  assign n8469 = pi13 ? n8464 : n8468;
  assign n8470 = pi12 ? n8455 : n8469;
  assign n8471 = pi19 ? n507 : n813;
  assign n8472 = pi18 ? n32 : n8471;
  assign n8473 = pi17 ? n2519 : ~n8472;
  assign n8474 = pi16 ? n32 : n8473;
  assign n8475 = pi17 ? n2519 : ~n2736;
  assign n8476 = pi16 ? n32 : n8475;
  assign n8477 = pi15 ? n8474 : n8476;
  assign n8478 = pi14 ? n7781 : n8477;
  assign n8479 = pi17 ? n2748 : ~n2736;
  assign n8480 = pi16 ? n32 : n8479;
  assign n8481 = pi17 ? n2748 : ~n2855;
  assign n8482 = pi16 ? n32 : n8481;
  assign n8483 = pi15 ? n8480 : n8482;
  assign n8484 = pi17 ? n2748 : ~n2616;
  assign n8485 = pi16 ? n32 : n8484;
  assign n8486 = pi15 ? n8485 : n8482;
  assign n8487 = pi14 ? n8483 : n8486;
  assign n8488 = pi13 ? n8478 : n8487;
  assign n8489 = pi15 ? n8482 : n6745;
  assign n8490 = pi17 ? n2748 : ~n8323;
  assign n8491 = pi16 ? n32 : n8490;
  assign n8492 = pi17 ? n4099 : ~n2512;
  assign n8493 = pi16 ? n32 : n8492;
  assign n8494 = pi15 ? n8491 : n8493;
  assign n8495 = pi14 ? n8489 : n8494;
  assign n8496 = pi17 ? n4099 : ~n2628;
  assign n8497 = pi16 ? n32 : n8496;
  assign n8498 = pi15 ? n8497 : n8493;
  assign n8499 = pi17 ? n4099 : ~n2519;
  assign n8500 = pi16 ? n32 : n8499;
  assign n8501 = pi15 ? n8493 : n8500;
  assign n8502 = pi14 ? n8498 : n8501;
  assign n8503 = pi13 ? n8495 : n8502;
  assign n8504 = pi12 ? n8488 : n8503;
  assign n8505 = pi11 ? n8470 : n8504;
  assign n8506 = pi10 ? n8432 : n8505;
  assign n8507 = pi09 ? n8359 : n8506;
  assign n8508 = pi08 ? n8343 : n8507;
  assign n8509 = pi18 ? n1813 : ~n6978;
  assign n8510 = pi17 ? n32 : n8509;
  assign n8511 = pi16 ? n32 : n8510;
  assign n8512 = pi15 ? n32 : n8511;
  assign n8513 = pi18 ? n1813 : ~n496;
  assign n8514 = pi17 ? n32 : n8513;
  assign n8515 = pi16 ? n32 : n8514;
  assign n8516 = pi19 ? n267 : n813;
  assign n8517 = pi18 ? n814 : ~n8516;
  assign n8518 = pi17 ? n32 : n8517;
  assign n8519 = pi16 ? n32 : n8518;
  assign n8520 = pi15 ? n8515 : n8519;
  assign n8521 = pi14 ? n8512 : n8520;
  assign n8522 = pi13 ? n32 : n8521;
  assign n8523 = pi12 ? n32 : n8522;
  assign n8524 = pi11 ? n32 : n8523;
  assign n8525 = pi10 ? n32 : n8524;
  assign n8526 = pi18 ? n814 : ~n496;
  assign n8527 = pi17 ? n32 : n8526;
  assign n8528 = pi16 ? n32 : n8527;
  assign n8529 = pi18 ? n1676 : ~n496;
  assign n8530 = pi17 ? n32 : n8529;
  assign n8531 = pi16 ? n32 : n8530;
  assign n8532 = pi15 ? n8528 : n8531;
  assign n8533 = pi17 ? n32 : ~n2726;
  assign n8534 = pi16 ? n32 : n8533;
  assign n8535 = pi19 ? n5694 : n531;
  assign n8536 = pi18 ? n32 : n8535;
  assign n8537 = pi17 ? n32 : ~n8536;
  assign n8538 = pi16 ? n32 : n8537;
  assign n8539 = pi15 ? n8534 : n8538;
  assign n8540 = pi14 ? n8532 : n8539;
  assign n8541 = pi15 ? n8167 : n7958;
  assign n8542 = pi14 ? n8165 : n8541;
  assign n8543 = pi13 ? n8540 : n8542;
  assign n8544 = pi14 ? n8170 : n8174;
  assign n8545 = pi15 ? n7758 : n7974;
  assign n8546 = pi20 ? n32 : ~n1010;
  assign n8547 = pi19 ? n32 : n8546;
  assign n8548 = pi18 ? n32 : n8547;
  assign n8549 = pi17 ? n2726 : ~n8548;
  assign n8550 = pi16 ? n32 : n8549;
  assign n8551 = pi15 ? n7974 : n8550;
  assign n8552 = pi14 ? n8545 : n8551;
  assign n8553 = pi13 ? n8544 : n8552;
  assign n8554 = pi12 ? n8543 : n8553;
  assign n8555 = pi17 ? n2726 : ~n8385;
  assign n8556 = pi16 ? n32 : n8555;
  assign n8557 = pi15 ? n8556 : n7979;
  assign n8558 = pi17 ? n2733 : ~n8187;
  assign n8559 = pi16 ? n32 : n8558;
  assign n8560 = pi15 ? n7300 : n8559;
  assign n8561 = pi14 ? n8557 : n8560;
  assign n8562 = pi20 ? n1324 : n321;
  assign n8563 = pi19 ? n32 : n8562;
  assign n8564 = pi18 ? n32 : n8563;
  assign n8565 = pi17 ? n2733 : ~n8564;
  assign n8566 = pi16 ? n32 : n8565;
  assign n8567 = pi17 ? n2733 : ~n8193;
  assign n8568 = pi16 ? n32 : n8567;
  assign n8569 = pi15 ? n8566 : n8568;
  assign n8570 = pi17 ? n2836 : ~n8193;
  assign n8571 = pi16 ? n32 : n8570;
  assign n8572 = pi15 ? n8568 : n8571;
  assign n8573 = pi14 ? n8569 : n8572;
  assign n8574 = pi13 ? n8561 : n8573;
  assign n8575 = pi17 ? n2839 : ~n8193;
  assign n8576 = pi16 ? n32 : n8575;
  assign n8577 = pi17 ? n2850 : ~n8564;
  assign n8578 = pi16 ? n32 : n8577;
  assign n8579 = pi15 ? n8576 : n8578;
  assign n8580 = pi17 ? n2850 : ~n8222;
  assign n8581 = pi16 ? n32 : n8580;
  assign n8582 = pi17 ? n2850 : ~n6768;
  assign n8583 = pi16 ? n32 : n8582;
  assign n8584 = pi15 ? n8581 : n8583;
  assign n8585 = pi14 ? n8579 : n8584;
  assign n8586 = pi17 ? n3067 : ~n3067;
  assign n8587 = pi16 ? n32 : n8586;
  assign n8588 = pi18 ? n32 : n4546;
  assign n8589 = pi17 ? n4245 : ~n8588;
  assign n8590 = pi16 ? n32 : n8589;
  assign n8591 = pi15 ? n8587 : n8590;
  assign n8592 = pi20 ? n1385 : n207;
  assign n8593 = pi19 ? n32 : n8592;
  assign n8594 = pi18 ? n32 : n8593;
  assign n8595 = pi17 ? n4245 : ~n8594;
  assign n8596 = pi16 ? n32 : n8595;
  assign n8597 = pi17 ? n2736 : ~n2733;
  assign n8598 = pi16 ? n32 : n8597;
  assign n8599 = pi15 ? n8596 : n8598;
  assign n8600 = pi14 ? n8591 : n8599;
  assign n8601 = pi13 ? n8585 : n8600;
  assign n8602 = pi12 ? n8574 : n8601;
  assign n8603 = pi11 ? n8554 : n8602;
  assign n8604 = pi17 ? n2736 : ~n7369;
  assign n8605 = pi16 ? n32 : n8604;
  assign n8606 = pi19 ? n32 : n1600;
  assign n8607 = pi18 ? n32 : n8606;
  assign n8608 = pi17 ? n2736 : ~n8607;
  assign n8609 = pi16 ? n32 : n8608;
  assign n8610 = pi15 ? n8605 : n8609;
  assign n8611 = pi20 ? n274 : ~n32;
  assign n8612 = pi19 ? n32 : n8611;
  assign n8613 = pi18 ? n32 : n8612;
  assign n8614 = pi17 ? n2736 : ~n8613;
  assign n8615 = pi16 ? n32 : n8614;
  assign n8616 = pi19 ? n32 : ~n5707;
  assign n8617 = pi18 ? n32 : n8616;
  assign n8618 = pi17 ? n2855 : ~n8617;
  assign n8619 = pi16 ? n32 : n8618;
  assign n8620 = pi15 ? n8615 : n8619;
  assign n8621 = pi14 ? n8610 : n8620;
  assign n8622 = pi20 ? n32 : ~n339;
  assign n8623 = pi19 ? n32 : ~n8622;
  assign n8624 = pi18 ? n32 : n8623;
  assign n8625 = pi17 ? n2855 : ~n8624;
  assign n8626 = pi16 ? n32 : n8625;
  assign n8627 = pi17 ? n2623 : ~n2726;
  assign n8628 = pi16 ? n32 : n8627;
  assign n8629 = pi15 ? n8626 : n8628;
  assign n8630 = pi21 ? n32 : n1392;
  assign n8631 = pi20 ? n8630 : ~n32;
  assign n8632 = pi19 ? n32 : n8631;
  assign n8633 = pi18 ? n32 : n8632;
  assign n8634 = pi17 ? n2623 : ~n8633;
  assign n8635 = pi16 ? n32 : n8634;
  assign n8636 = pi15 ? n8635 : n6947;
  assign n8637 = pi14 ? n8629 : n8636;
  assign n8638 = pi13 ? n8621 : n8637;
  assign n8639 = pi18 ? n32 : n1156;
  assign n8640 = pi17 ? n2623 : ~n8639;
  assign n8641 = pi16 ? n32 : n8640;
  assign n8642 = pi19 ? n32 : ~n1818;
  assign n8643 = pi18 ? n32 : n8642;
  assign n8644 = pi21 ? n405 : ~n309;
  assign n8645 = pi20 ? n8644 : ~n32;
  assign n8646 = pi19 ? n32 : n8645;
  assign n8647 = pi18 ? n32 : n8646;
  assign n8648 = pi17 ? n8643 : ~n8647;
  assign n8649 = pi16 ? n32 : n8648;
  assign n8650 = pi15 ? n8641 : n8649;
  assign n8651 = pi17 ? n8643 : ~n2831;
  assign n8652 = pi16 ? n32 : n8651;
  assign n8653 = pi18 ? n32 : n4407;
  assign n8654 = pi17 ? n2512 : ~n8653;
  assign n8655 = pi16 ? n32 : n8654;
  assign n8656 = pi15 ? n8652 : n8655;
  assign n8657 = pi14 ? n8650 : n8656;
  assign n8658 = pi17 ? n2628 : ~n8639;
  assign n8659 = pi16 ? n32 : n8658;
  assign n8660 = pi15 ? n6748 : n8659;
  assign n8661 = pi21 ? n32 : ~n7410;
  assign n8662 = pi20 ? n32 : n8661;
  assign n8663 = pi19 ? n8662 : n2848;
  assign n8664 = pi18 ? n32 : n8663;
  assign n8665 = pi17 ? n2618 : ~n8664;
  assign n8666 = pi16 ? n32 : n8665;
  assign n8667 = pi15 ? n7322 : n8666;
  assign n8668 = pi14 ? n8660 : n8667;
  assign n8669 = pi13 ? n8657 : n8668;
  assign n8670 = pi12 ? n8638 : n8669;
  assign n8671 = pi17 ? n4099 : ~n2724;
  assign n8672 = pi16 ? n32 : n8671;
  assign n8673 = pi15 ? n8672 : n6949;
  assign n8674 = pi19 ? n857 : n236;
  assign n8675 = pi18 ? n32 : n8674;
  assign n8676 = pi17 ? n4099 : ~n8675;
  assign n8677 = pi16 ? n32 : n8676;
  assign n8678 = pi17 ? n4099 : ~n8301;
  assign n8679 = pi16 ? n32 : n8678;
  assign n8680 = pi15 ? n8677 : n8679;
  assign n8681 = pi14 ? n8673 : n8680;
  assign n8682 = pi17 ? n4099 : ~n2736;
  assign n8683 = pi16 ? n32 : n8682;
  assign n8684 = pi17 ? n4099 : ~n2616;
  assign n8685 = pi16 ? n32 : n8684;
  assign n8686 = pi15 ? n8683 : n8685;
  assign n8687 = pi17 ? n2750 : ~n2616;
  assign n8688 = pi16 ? n32 : n8687;
  assign n8689 = pi17 ? n2750 : ~n2855;
  assign n8690 = pi16 ? n32 : n8689;
  assign n8691 = pi15 ? n8688 : n8690;
  assign n8692 = pi14 ? n8686 : n8691;
  assign n8693 = pi13 ? n8681 : n8692;
  assign n8694 = pi17 ? n2855 : ~n2750;
  assign n8695 = pi16 ? n32 : n8694;
  assign n8696 = pi18 ? n7221 : n702;
  assign n8697 = pi17 ? n2616 : ~n8696;
  assign n8698 = pi16 ? n32 : n8697;
  assign n8699 = pi15 ? n8695 : n8698;
  assign n8700 = pi17 ? n2855 : ~n2512;
  assign n8701 = pi16 ? n32 : n8700;
  assign n8702 = pi17 ? n2616 : ~n2512;
  assign n8703 = pi16 ? n32 : n8702;
  assign n8704 = pi15 ? n8701 : n8703;
  assign n8705 = pi14 ? n8699 : n8704;
  assign n8706 = pi17 ? n2616 : ~n2628;
  assign n8707 = pi16 ? n32 : n8706;
  assign n8708 = pi17 ? n2736 : ~n2512;
  assign n8709 = pi16 ? n32 : n8708;
  assign n8710 = pi15 ? n8707 : n8709;
  assign n8711 = pi19 ? n6049 : ~n32;
  assign n8712 = pi18 ? n32 : n8711;
  assign n8713 = pi17 ? n2736 : ~n8712;
  assign n8714 = pi16 ? n32 : n8713;
  assign n8715 = pi17 ? n2724 : ~n2517;
  assign n8716 = pi16 ? n32 : n8715;
  assign n8717 = pi15 ? n8714 : n8716;
  assign n8718 = pi14 ? n8710 : n8717;
  assign n8719 = pi13 ? n8705 : n8718;
  assign n8720 = pi12 ? n8693 : n8719;
  assign n8721 = pi11 ? n8670 : n8720;
  assign n8722 = pi10 ? n8603 : n8721;
  assign n8723 = pi09 ? n8525 : n8722;
  assign n8724 = pi18 ? n2298 : ~n6978;
  assign n8725 = pi17 ? n32 : n8724;
  assign n8726 = pi16 ? n32 : n8725;
  assign n8727 = pi15 ? n32 : n8726;
  assign n8728 = pi18 ? n430 : ~n496;
  assign n8729 = pi17 ? n32 : n8728;
  assign n8730 = pi16 ? n32 : n8729;
  assign n8731 = pi18 ? n430 : ~n8516;
  assign n8732 = pi17 ? n32 : n8731;
  assign n8733 = pi16 ? n32 : n8732;
  assign n8734 = pi15 ? n8730 : n8733;
  assign n8735 = pi14 ? n8727 : n8734;
  assign n8736 = pi13 ? n32 : n8735;
  assign n8737 = pi12 ? n32 : n8736;
  assign n8738 = pi11 ? n32 : n8737;
  assign n8739 = pi10 ? n32 : n8738;
  assign n8740 = pi18 ? n2304 : ~n496;
  assign n8741 = pi17 ? n32 : n8740;
  assign n8742 = pi16 ? n32 : n8741;
  assign n8743 = pi18 ? n1942 : ~n496;
  assign n8744 = pi17 ? n32 : n8743;
  assign n8745 = pi16 ? n32 : n8744;
  assign n8746 = pi15 ? n8742 : n8745;
  assign n8747 = pi18 ? n237 : ~n880;
  assign n8748 = pi17 ? n32 : n8747;
  assign n8749 = pi16 ? n32 : n8748;
  assign n8750 = pi18 ? n618 : ~n8535;
  assign n8751 = pi17 ? n32 : n8750;
  assign n8752 = pi16 ? n32 : n8751;
  assign n8753 = pi15 ? n8749 : n8752;
  assign n8754 = pi14 ? n8746 : n8753;
  assign n8755 = pi15 ? n8531 : n7958;
  assign n8756 = pi14 ? n8362 : n8755;
  assign n8757 = pi13 ? n8754 : n8756;
  assign n8758 = pi14 ? n8368 : n8374;
  assign n8759 = pi15 ? n7971 : n8170;
  assign n8760 = pi21 ? n1009 : n51;
  assign n8761 = pi20 ? n32 : ~n8760;
  assign n8762 = pi19 ? n32 : n8761;
  assign n8763 = pi18 ? n32 : n8762;
  assign n8764 = pi17 ? n3046 : ~n8763;
  assign n8765 = pi16 ? n32 : n8764;
  assign n8766 = pi15 ? n8170 : n8765;
  assign n8767 = pi14 ? n8759 : n8766;
  assign n8768 = pi13 ? n8758 : n8767;
  assign n8769 = pi12 ? n8757 : n8768;
  assign n8770 = pi17 ? n3292 : ~n8385;
  assign n8771 = pi16 ? n32 : n8770;
  assign n8772 = pi15 ? n8771 : n8173;
  assign n8773 = pi17 ? n3175 : ~n8187;
  assign n8774 = pi16 ? n32 : n8773;
  assign n8775 = pi15 ? n7546 : n8774;
  assign n8776 = pi14 ? n8772 : n8775;
  assign n8777 = pi17 ? n3175 : ~n8564;
  assign n8778 = pi16 ? n32 : n8777;
  assign n8779 = pi17 ? n3175 : ~n8193;
  assign n8780 = pi16 ? n32 : n8779;
  assign n8781 = pi15 ? n8778 : n8780;
  assign n8782 = pi17 ? n2963 : ~n8193;
  assign n8783 = pi16 ? n32 : n8782;
  assign n8784 = pi15 ? n8780 : n8783;
  assign n8785 = pi14 ? n8781 : n8784;
  assign n8786 = pi13 ? n8776 : n8785;
  assign n8787 = pi17 ? n2831 : ~n8193;
  assign n8788 = pi16 ? n32 : n8787;
  assign n8789 = pi17 ? n2831 : ~n8564;
  assign n8790 = pi16 ? n32 : n8789;
  assign n8791 = pi15 ? n8788 : n8790;
  assign n8792 = pi17 ? n2831 : ~n8222;
  assign n8793 = pi16 ? n32 : n8792;
  assign n8794 = pi17 ? n2831 : ~n6768;
  assign n8795 = pi16 ? n32 : n8794;
  assign n8796 = pi15 ? n8793 : n8795;
  assign n8797 = pi14 ? n8791 : n8796;
  assign n8798 = pi17 ? n2831 : ~n3067;
  assign n8799 = pi16 ? n32 : n8798;
  assign n8800 = pi17 ? n2733 : ~n8588;
  assign n8801 = pi16 ? n32 : n8800;
  assign n8802 = pi15 ? n8799 : n8801;
  assign n8803 = pi20 ? n1385 : n1940;
  assign n8804 = pi19 ? n32 : n8803;
  assign n8805 = pi18 ? n32 : n8804;
  assign n8806 = pi17 ? n2733 : ~n8805;
  assign n8807 = pi16 ? n32 : n8806;
  assign n8808 = pi15 ? n8807 : n7982;
  assign n8809 = pi14 ? n8802 : n8808;
  assign n8810 = pi13 ? n8797 : n8809;
  assign n8811 = pi12 ? n8786 : n8810;
  assign n8812 = pi11 ? n8769 : n8811;
  assign n8813 = pi17 ? n2836 : ~n7825;
  assign n8814 = pi16 ? n32 : n8813;
  assign n8815 = pi17 ? n2836 : ~n8607;
  assign n8816 = pi16 ? n32 : n8815;
  assign n8817 = pi15 ? n8814 : n8816;
  assign n8818 = pi20 ? n266 : ~n32;
  assign n8819 = pi19 ? n32 : n8818;
  assign n8820 = pi18 ? n32 : n8819;
  assign n8821 = pi17 ? n2839 : ~n8820;
  assign n8822 = pi16 ? n32 : n8821;
  assign n8823 = pi17 ? n2850 : ~n8617;
  assign n8824 = pi16 ? n32 : n8823;
  assign n8825 = pi15 ? n8822 : n8824;
  assign n8826 = pi14 ? n8817 : n8825;
  assign n8827 = pi17 ? n2850 : ~n8624;
  assign n8828 = pi16 ? n32 : n8827;
  assign n8829 = pi17 ? n2724 : ~n2726;
  assign n8830 = pi16 ? n32 : n8829;
  assign n8831 = pi15 ? n8828 : n8830;
  assign n8832 = pi17 ? n2724 : ~n8633;
  assign n8833 = pi16 ? n32 : n8832;
  assign n8834 = pi15 ? n8833 : n7129;
  assign n8835 = pi14 ? n8831 : n8834;
  assign n8836 = pi13 ? n8826 : n8835;
  assign n8837 = pi17 ? n2724 : ~n8639;
  assign n8838 = pi16 ? n32 : n8837;
  assign n8839 = pi20 ? n1940 : ~n1076;
  assign n8840 = pi19 ? n32 : n8839;
  assign n8841 = pi18 ? n32 : n8840;
  assign n8842 = pi17 ? n8841 : ~n8647;
  assign n8843 = pi16 ? n32 : n8842;
  assign n8844 = pi15 ? n8838 : n8843;
  assign n8845 = pi17 ? n8841 : ~n2733;
  assign n8846 = pi16 ? n32 : n8845;
  assign n8847 = pi17 ? n2623 : ~n8653;
  assign n8848 = pi16 ? n32 : n8847;
  assign n8849 = pi15 ? n8846 : n8848;
  assign n8850 = pi14 ? n8844 : n8849;
  assign n8851 = pi19 ? n1785 : n349;
  assign n8852 = pi18 ? n32 : n8851;
  assign n8853 = pi17 ? n2623 : ~n8852;
  assign n8854 = pi16 ? n32 : n8853;
  assign n8855 = pi17 ? n2736 : ~n8852;
  assign n8856 = pi16 ? n32 : n8855;
  assign n8857 = pi15 ? n8854 : n8856;
  assign n8858 = pi19 ? n1464 : n349;
  assign n8859 = pi18 ? n32 : n8858;
  assign n8860 = pi17 ? n2616 : ~n8859;
  assign n8861 = pi16 ? n32 : n8860;
  assign n8862 = pi15 ? n8856 : n8861;
  assign n8863 = pi14 ? n8857 : n8862;
  assign n8864 = pi13 ? n8850 : n8863;
  assign n8865 = pi12 ? n8836 : n8864;
  assign n8866 = pi19 ? n1785 : n813;
  assign n8867 = pi18 ? n32 : n8866;
  assign n8868 = pi17 ? n2616 : ~n8867;
  assign n8869 = pi16 ? n32 : n8868;
  assign n8870 = pi17 ? n2616 : ~n3067;
  assign n8871 = pi16 ? n32 : n8870;
  assign n8872 = pi15 ? n8869 : n8871;
  assign n8873 = pi17 ? n2616 : ~n8675;
  assign n8874 = pi16 ? n32 : n8873;
  assign n8875 = pi17 ? n2616 : ~n8301;
  assign n8876 = pi16 ? n32 : n8875;
  assign n8877 = pi15 ? n8874 : n8876;
  assign n8878 = pi14 ? n8872 : n8877;
  assign n8879 = pi17 ? n2736 : ~n2736;
  assign n8880 = pi16 ? n32 : n8879;
  assign n8881 = pi17 ? n2736 : ~n2616;
  assign n8882 = pi16 ? n32 : n8881;
  assign n8883 = pi15 ? n8880 : n8882;
  assign n8884 = pi19 ? n32 : ~n5626;
  assign n8885 = pi18 ? n32 : n8884;
  assign n8886 = pi17 ? n4245 : ~n8885;
  assign n8887 = pi16 ? n32 : n8886;
  assign n8888 = pi17 ? n4245 : ~n2616;
  assign n8889 = pi16 ? n32 : n8888;
  assign n8890 = pi15 ? n8887 : n8889;
  assign n8891 = pi14 ? n8883 : n8890;
  assign n8892 = pi13 ? n8878 : n8891;
  assign n8893 = pi17 ? n4245 : ~n2750;
  assign n8894 = pi16 ? n32 : n8893;
  assign n8895 = pi17 ? n4245 : ~n8696;
  assign n8896 = pi16 ? n32 : n8895;
  assign n8897 = pi15 ? n8894 : n8896;
  assign n8898 = pi17 ? n4245 : ~n2512;
  assign n8899 = pi16 ? n32 : n8898;
  assign n8900 = pi17 ? n3067 : ~n2512;
  assign n8901 = pi16 ? n32 : n8900;
  assign n8902 = pi15 ? n8899 : n8901;
  assign n8903 = pi14 ? n8897 : n8902;
  assign n8904 = pi17 ? n2836 : ~n2628;
  assign n8905 = pi16 ? n32 : n8904;
  assign n8906 = pi15 ? n8901 : n8905;
  assign n8907 = pi20 ? n207 : ~n518;
  assign n8908 = pi19 ? n8907 : n32;
  assign n8909 = pi18 ? n32 : ~n8908;
  assign n8910 = pi17 ? n2836 : ~n8909;
  assign n8911 = pi16 ? n32 : n8910;
  assign n8912 = pi17 ? n2836 : ~n2517;
  assign n8913 = pi16 ? n32 : n8912;
  assign n8914 = pi15 ? n8911 : n8913;
  assign n8915 = pi14 ? n8906 : n8914;
  assign n8916 = pi13 ? n8903 : n8915;
  assign n8917 = pi12 ? n8892 : n8916;
  assign n8918 = pi11 ? n8865 : n8917;
  assign n8919 = pi10 ? n8812 : n8918;
  assign n8920 = pi09 ? n8739 : n8919;
  assign n8921 = pi08 ? n8723 : n8920;
  assign n8922 = pi07 ? n8508 : n8921;
  assign n8923 = pi18 ? n418 : ~n8086;
  assign n8924 = pi17 ? n32 : n8923;
  assign n8925 = pi16 ? n32 : n8924;
  assign n8926 = pi15 ? n32 : n8925;
  assign n8927 = pi19 ? n6398 : ~n7488;
  assign n8928 = pi18 ? n418 : ~n8927;
  assign n8929 = pi17 ? n32 : n8928;
  assign n8930 = pi16 ? n32 : n8929;
  assign n8931 = pi19 ? n340 : ~n857;
  assign n8932 = pi20 ? n3847 : ~n915;
  assign n8933 = pi19 ? n8932 : ~n7488;
  assign n8934 = pi18 ? n8931 : ~n8933;
  assign n8935 = pi17 ? n32 : n8934;
  assign n8936 = pi16 ? n32 : n8935;
  assign n8937 = pi15 ? n8930 : n8936;
  assign n8938 = pi14 ? n8926 : n8937;
  assign n8939 = pi13 ? n32 : n8938;
  assign n8940 = pi12 ? n32 : n8939;
  assign n8941 = pi11 ? n32 : n8940;
  assign n8942 = pi10 ? n32 : n8941;
  assign n8943 = pi21 ? n405 : ~n174;
  assign n8944 = pi20 ? n1685 : n8943;
  assign n8945 = pi19 ? n365 : ~n8944;
  assign n8946 = pi20 ? n1611 : ~n32;
  assign n8947 = pi19 ? n8946 : n813;
  assign n8948 = pi18 ? n8945 : ~n8947;
  assign n8949 = pi17 ? n32 : n8948;
  assign n8950 = pi16 ? n32 : n8949;
  assign n8951 = pi19 ? n208 : n349;
  assign n8952 = pi18 ? n1813 : ~n8951;
  assign n8953 = pi17 ? n32 : n8952;
  assign n8954 = pi16 ? n32 : n8953;
  assign n8955 = pi15 ? n8950 : n8954;
  assign n8956 = pi19 ? n267 : n321;
  assign n8957 = pi18 ? n814 : ~n8956;
  assign n8958 = pi17 ? n32 : n8957;
  assign n8959 = pi16 ? n32 : n8958;
  assign n8960 = pi19 ? n221 : n321;
  assign n8961 = pi18 ? n814 : ~n8960;
  assign n8962 = pi17 ? n32 : n8961;
  assign n8963 = pi16 ? n32 : n8962;
  assign n8964 = pi15 ? n8959 : n8963;
  assign n8965 = pi14 ? n8955 : n8964;
  assign n8966 = pi19 ? n531 : n236;
  assign n8967 = pi18 ? n814 : ~n8966;
  assign n8968 = pi17 ? n32 : n8967;
  assign n8969 = pi16 ? n32 : n8968;
  assign n8970 = pi19 ? n916 : n236;
  assign n8971 = pi18 ? n1942 : ~n8970;
  assign n8972 = pi17 ? n32 : n8971;
  assign n8973 = pi16 ? n32 : n8972;
  assign n8974 = pi15 ? n8969 : n8973;
  assign n8975 = pi19 ? n221 : n236;
  assign n8976 = pi18 ? n1942 : ~n8975;
  assign n8977 = pi17 ? n32 : n8976;
  assign n8978 = pi16 ? n32 : n8977;
  assign n8979 = pi17 ? n32 : ~n6979;
  assign n8980 = pi16 ? n32 : n8979;
  assign n8981 = pi15 ? n8978 : n8980;
  assign n8982 = pi14 ? n8974 : n8981;
  assign n8983 = pi13 ? n8965 : n8982;
  assign n8984 = pi19 ? n5694 : n321;
  assign n8985 = pi18 ? n32 : n8984;
  assign n8986 = pi17 ? n32 : ~n8985;
  assign n8987 = pi16 ? n32 : n8986;
  assign n8988 = pi19 ? n5694 : n236;
  assign n8989 = pi18 ? n32 : n8988;
  assign n8990 = pi17 ? n3282 : ~n8989;
  assign n8991 = pi16 ? n32 : n8990;
  assign n8992 = pi19 ? n5694 : n617;
  assign n8993 = pi18 ? n32 : n8992;
  assign n8994 = pi17 ? n3282 : ~n8993;
  assign n8995 = pi16 ? n32 : n8994;
  assign n8996 = pi15 ? n8991 : n8995;
  assign n8997 = pi14 ? n8987 : n8996;
  assign n8998 = pi17 ? n3155 : ~n2726;
  assign n8999 = pi16 ? n32 : n8998;
  assign n9000 = pi21 ? n140 : ~n1939;
  assign n9001 = pi20 ? n32 : ~n9000;
  assign n9002 = pi19 ? n32 : n9001;
  assign n9003 = pi18 ? n32 : n9002;
  assign n9004 = pi17 ? n2954 : ~n9003;
  assign n9005 = pi16 ? n32 : n9004;
  assign n9006 = pi15 ? n8999 : n9005;
  assign n9007 = pi20 ? n32 : ~n207;
  assign n9008 = pi19 ? n9007 : n349;
  assign n9009 = pi18 ? n32 : n9008;
  assign n9010 = pi17 ? n2954 : ~n9009;
  assign n9011 = pi16 ? n32 : n9010;
  assign n9012 = pi19 ? n267 : n32;
  assign n9013 = pi21 ? n124 : n51;
  assign n9014 = pi20 ? n321 : ~n9013;
  assign n9015 = pi19 ? n5694 : n9014;
  assign n9016 = pi18 ? n9012 : n9015;
  assign n9017 = pi17 ? n3728 : ~n9016;
  assign n9018 = pi16 ? n32 : n9017;
  assign n9019 = pi15 ? n9011 : n9018;
  assign n9020 = pi14 ? n9006 : n9019;
  assign n9021 = pi13 ? n8997 : n9020;
  assign n9022 = pi12 ? n8983 : n9021;
  assign n9023 = pi17 ? n3728 : ~n8385;
  assign n9024 = pi16 ? n32 : n9023;
  assign n9025 = pi17 ? n3160 : ~n2736;
  assign n9026 = pi16 ? n32 : n9025;
  assign n9027 = pi15 ? n9024 : n9026;
  assign n9028 = pi20 ? n321 : ~n220;
  assign n9029 = pi19 ? n32 : n9028;
  assign n9030 = pi18 ? n32 : n9029;
  assign n9031 = pi17 ? n3164 : ~n9030;
  assign n9032 = pi16 ? n32 : n9031;
  assign n9033 = pi17 ? n3164 : ~n8193;
  assign n9034 = pi16 ? n32 : n9033;
  assign n9035 = pi15 ? n9032 : n9034;
  assign n9036 = pi14 ? n9027 : n9035;
  assign n9037 = pi20 ? n246 : n321;
  assign n9038 = pi19 ? n32 : n9037;
  assign n9039 = pi18 ? n32 : n9038;
  assign n9040 = pi17 ? n3164 : ~n9039;
  assign n9041 = pi16 ? n32 : n9040;
  assign n9042 = pi17 ? n3046 : ~n8193;
  assign n9043 = pi16 ? n32 : n9042;
  assign n9044 = pi17 ? n3292 : ~n8204;
  assign n9045 = pi16 ? n32 : n9044;
  assign n9046 = pi15 ? n9043 : n9045;
  assign n9047 = pi14 ? n9041 : n9046;
  assign n9048 = pi13 ? n9036 : n9047;
  assign n9049 = pi17 ? n2952 : ~n8193;
  assign n9050 = pi16 ? n32 : n9049;
  assign n9051 = pi17 ? n2952 : ~n8204;
  assign n9052 = pi16 ? n32 : n9051;
  assign n9053 = pi15 ? n9050 : n9052;
  assign n9054 = pi17 ? n2952 : ~n7369;
  assign n9055 = pi16 ? n32 : n9054;
  assign n9056 = pi18 ? n32 : n1387;
  assign n9057 = pi17 ? n2952 : ~n9056;
  assign n9058 = pi16 ? n32 : n9057;
  assign n9059 = pi15 ? n9055 : n9058;
  assign n9060 = pi14 ? n9053 : n9059;
  assign n9061 = pi19 ? n4670 : n422;
  assign n9062 = pi18 ? n32 : n9061;
  assign n9063 = pi17 ? n2952 : ~n9062;
  assign n9064 = pi16 ? n32 : n9063;
  assign n9065 = pi17 ? n2726 : ~n8232;
  assign n9066 = pi16 ? n32 : n9065;
  assign n9067 = pi15 ? n9064 : n9066;
  assign n9068 = pi20 ? n342 : n1940;
  assign n9069 = pi19 ? n32 : n9068;
  assign n9070 = pi18 ? n32 : n9069;
  assign n9071 = pi17 ? n2963 : ~n9070;
  assign n9072 = pi16 ? n32 : n9071;
  assign n9073 = pi18 ? n32 : n2026;
  assign n9074 = pi17 ? n2963 : ~n9073;
  assign n9075 = pi16 ? n32 : n9074;
  assign n9076 = pi15 ? n9072 : n9075;
  assign n9077 = pi14 ? n9067 : n9076;
  assign n9078 = pi13 ? n9060 : n9077;
  assign n9079 = pi12 ? n9048 : n9078;
  assign n9080 = pi11 ? n9022 : n9079;
  assign n9081 = pi17 ? n2963 : ~n7825;
  assign n9082 = pi16 ? n32 : n9081;
  assign n9083 = pi18 ? n32 : n4559;
  assign n9084 = pi17 ? n2963 : ~n9083;
  assign n9085 = pi16 ? n32 : n9084;
  assign n9086 = pi15 ? n9082 : n9085;
  assign n9087 = pi15 ? n7549 : n7979;
  assign n9088 = pi14 ? n9086 : n9087;
  assign n9089 = pi20 ? n5854 : n339;
  assign n9090 = pi19 ? n32 : n9089;
  assign n9091 = pi18 ? n32 : n9090;
  assign n9092 = pi17 ? n3182 : ~n9091;
  assign n9093 = pi16 ? n32 : n9092;
  assign n9094 = pi19 ? n32 : n6619;
  assign n9095 = pi18 ? n32 : n9094;
  assign n9096 = pi17 ? n2831 : ~n9095;
  assign n9097 = pi16 ? n32 : n9096;
  assign n9098 = pi15 ? n9093 : n9097;
  assign n9099 = pi17 ? n2839 : ~n3175;
  assign n9100 = pi16 ? n32 : n9099;
  assign n9101 = pi20 ? n785 : ~n32;
  assign n9102 = pi19 ? n32 : n9101;
  assign n9103 = pi18 ? n32 : n9102;
  assign n9104 = pi17 ? n2831 : ~n9103;
  assign n9105 = pi16 ? n32 : n9104;
  assign n9106 = pi15 ? n9100 : n9105;
  assign n9107 = pi14 ? n9098 : n9106;
  assign n9108 = pi13 ? n9088 : n9107;
  assign n9109 = pi17 ? n2839 : ~n8647;
  assign n9110 = pi16 ? n32 : n9109;
  assign n9111 = pi17 ? n2733 : ~n2852;
  assign n9112 = pi16 ? n32 : n9111;
  assign n9113 = pi15 ? n9110 : n9112;
  assign n9114 = pi21 ? n174 : ~n51;
  assign n9115 = pi20 ? n9114 : ~n32;
  assign n9116 = pi19 ? n32 : n9115;
  assign n9117 = pi18 ? n32 : n9116;
  assign n9118 = pi17 ? n2733 : ~n9117;
  assign n9119 = pi16 ? n32 : n9118;
  assign n9120 = pi17 ? n3067 : ~n2733;
  assign n9121 = pi16 ? n32 : n9120;
  assign n9122 = pi15 ? n9119 : n9121;
  assign n9123 = pi14 ? n9113 : n9122;
  assign n9124 = pi17 ? n2850 : ~n2724;
  assign n9125 = pi16 ? n32 : n9124;
  assign n9126 = pi15 ? n9121 : n9125;
  assign n9127 = pi17 ? n2850 : ~n8852;
  assign n9128 = pi16 ? n32 : n9127;
  assign n9129 = pi17 ? n3067 : ~n2724;
  assign n9130 = pi16 ? n32 : n9129;
  assign n9131 = pi15 ? n9128 : n9130;
  assign n9132 = pi14 ? n9126 : n9131;
  assign n9133 = pi13 ? n9123 : n9132;
  assign n9134 = pi12 ? n9108 : n9133;
  assign n9135 = pi19 ? n1785 : n236;
  assign n9136 = pi18 ? n32 : n9135;
  assign n9137 = pi17 ? n3067 : ~n9136;
  assign n9138 = pi16 ? n32 : n9137;
  assign n9139 = pi15 ? n8587 : n9138;
  assign n9140 = pi17 ? n3067 : ~n2736;
  assign n9141 = pi16 ? n32 : n9140;
  assign n9142 = pi15 ? n9130 : n9141;
  assign n9143 = pi14 ? n9139 : n9142;
  assign n9144 = pi17 ? n2836 : ~n2736;
  assign n9145 = pi16 ? n32 : n9144;
  assign n9146 = pi17 ? n2836 : ~n8885;
  assign n9147 = pi16 ? n32 : n9146;
  assign n9148 = pi15 ? n9145 : n9147;
  assign n9149 = pi17 ? n2733 : ~n2855;
  assign n9150 = pi16 ? n32 : n9149;
  assign n9151 = pi17 ? n2733 : ~n2616;
  assign n9152 = pi16 ? n32 : n9151;
  assign n9153 = pi15 ? n9150 : n9152;
  assign n9154 = pi14 ? n9148 : n9153;
  assign n9155 = pi13 ? n9143 : n9154;
  assign n9156 = pi17 ? n2733 : ~n2750;
  assign n9157 = pi16 ? n32 : n9156;
  assign n9158 = pi17 ? n2733 : ~n2618;
  assign n9159 = pi16 ? n32 : n9158;
  assign n9160 = pi17 ? n2963 : ~n2618;
  assign n9161 = pi16 ? n32 : n9160;
  assign n9162 = pi15 ? n9159 : n9161;
  assign n9163 = pi14 ? n9157 : n9162;
  assign n9164 = pi17 ? n2963 : ~n2628;
  assign n9165 = pi16 ? n32 : n9164;
  assign n9166 = pi17 ? n2726 : ~n2628;
  assign n9167 = pi16 ? n32 : n9166;
  assign n9168 = pi15 ? n9165 : n9167;
  assign n9169 = pi20 ? n3523 : n32;
  assign n9170 = pi19 ? n9169 : n32;
  assign n9171 = pi20 ? n274 : n518;
  assign n9172 = pi19 ? n9171 : ~n32;
  assign n9173 = pi18 ? n9170 : n9172;
  assign n9174 = pi17 ? n2726 : ~n9173;
  assign n9175 = pi16 ? n32 : n9174;
  assign n9176 = pi17 ? n2963 : ~n2517;
  assign n9177 = pi16 ? n32 : n9176;
  assign n9178 = pi15 ? n9175 : n9177;
  assign n9179 = pi14 ? n9168 : n9178;
  assign n9180 = pi13 ? n9163 : n9179;
  assign n9181 = pi12 ? n9155 : n9180;
  assign n9182 = pi11 ? n9134 : n9181;
  assign n9183 = pi10 ? n9080 : n9182;
  assign n9184 = pi09 ? n8942 : n9183;
  assign n9185 = pi18 ? n797 : ~n8086;
  assign n9186 = pi17 ? n32 : n9185;
  assign n9187 = pi16 ? n32 : n9186;
  assign n9188 = pi15 ? n32 : n9187;
  assign n9189 = pi19 ? n750 : ~n8622;
  assign n9190 = pi19 ? n6398 : ~n1757;
  assign n9191 = pi18 ? n9189 : ~n9190;
  assign n9192 = pi17 ? n32 : n9191;
  assign n9193 = pi16 ? n32 : n9192;
  assign n9194 = pi21 ? n309 : ~n173;
  assign n9195 = pi20 ? n9194 : ~n623;
  assign n9196 = pi19 ? n792 : ~n9195;
  assign n9197 = pi20 ? n6050 : ~n266;
  assign n9198 = pi19 ? n9197 : ~n32;
  assign n9199 = pi18 ? n9196 : ~n9198;
  assign n9200 = pi17 ? n32 : n9199;
  assign n9201 = pi16 ? n32 : n9200;
  assign n9202 = pi15 ? n9193 : n9201;
  assign n9203 = pi14 ? n9188 : n9202;
  assign n9204 = pi13 ? n32 : n9203;
  assign n9205 = pi12 ? n32 : n9204;
  assign n9206 = pi11 ? n32 : n9205;
  assign n9207 = pi10 ? n32 : n9206;
  assign n9208 = pi20 ? n220 : n749;
  assign n9209 = pi19 ? n208 : ~n9208;
  assign n9210 = pi18 ? n9209 : ~n8947;
  assign n9211 = pi17 ? n32 : n9210;
  assign n9212 = pi16 ? n32 : n9211;
  assign n9213 = pi18 ? n430 : ~n8951;
  assign n9214 = pi17 ? n32 : n9213;
  assign n9215 = pi16 ? n32 : n9214;
  assign n9216 = pi15 ? n9212 : n9215;
  assign n9217 = pi18 ? n430 : ~n8956;
  assign n9218 = pi17 ? n32 : n9217;
  assign n9219 = pi16 ? n32 : n9218;
  assign n9220 = pi20 ? n32 : n7839;
  assign n9221 = pi19 ? n9220 : n321;
  assign n9222 = pi18 ? n430 : ~n9221;
  assign n9223 = pi17 ? n32 : n9222;
  assign n9224 = pi16 ? n32 : n9223;
  assign n9225 = pi15 ? n9219 : n9224;
  assign n9226 = pi14 ? n9216 : n9225;
  assign n9227 = pi18 ? n2304 : ~n8966;
  assign n9228 = pi17 ? n32 : n9227;
  assign n9229 = pi16 ? n32 : n9228;
  assign n9230 = pi18 ? n2304 : ~n8970;
  assign n9231 = pi17 ? n32 : n9230;
  assign n9232 = pi16 ? n32 : n9231;
  assign n9233 = pi15 ? n9229 : n9232;
  assign n9234 = pi18 ? n344 : ~n8975;
  assign n9235 = pi17 ? n32 : n9234;
  assign n9236 = pi16 ? n32 : n9235;
  assign n9237 = pi18 ? n237 : ~n6978;
  assign n9238 = pi17 ? n32 : n9237;
  assign n9239 = pi16 ? n32 : n9238;
  assign n9240 = pi15 ? n9236 : n9239;
  assign n9241 = pi14 ? n9233 : n9240;
  assign n9242 = pi13 ? n9226 : n9241;
  assign n9243 = pi18 ? n237 : ~n8984;
  assign n9244 = pi17 ? n32 : n9243;
  assign n9245 = pi16 ? n32 : n9244;
  assign n9246 = pi18 ? n618 : ~n8984;
  assign n9247 = pi17 ? n32 : n9246;
  assign n9248 = pi16 ? n32 : n9247;
  assign n9249 = pi15 ? n9245 : n9248;
  assign n9250 = pi18 ? n618 : ~n8988;
  assign n9251 = pi17 ? n32 : n9250;
  assign n9252 = pi16 ? n32 : n9251;
  assign n9253 = pi18 ? n618 : ~n8992;
  assign n9254 = pi17 ? n32 : n9253;
  assign n9255 = pi16 ? n32 : n9254;
  assign n9256 = pi15 ? n9252 : n9255;
  assign n9257 = pi14 ? n9249 : n9256;
  assign n9258 = pi18 ? n1676 : ~n880;
  assign n9259 = pi17 ? n32 : n9258;
  assign n9260 = pi16 ? n32 : n9259;
  assign n9261 = pi17 ? n32 : ~n9003;
  assign n9262 = pi16 ? n32 : n9261;
  assign n9263 = pi15 ? n9260 : n9262;
  assign n9264 = pi17 ? n32 : ~n9009;
  assign n9265 = pi16 ? n32 : n9264;
  assign n9266 = pi19 ? n5694 : n8383;
  assign n9267 = pi18 ? n9012 : n9266;
  assign n9268 = pi17 ? n32 : ~n9267;
  assign n9269 = pi16 ? n32 : n9268;
  assign n9270 = pi15 ? n9265 : n9269;
  assign n9271 = pi14 ? n9263 : n9270;
  assign n9272 = pi13 ? n9257 : n9271;
  assign n9273 = pi12 ? n9242 : n9272;
  assign n9274 = pi17 ? n3282 : ~n2736;
  assign n9275 = pi16 ? n32 : n9274;
  assign n9276 = pi15 ? n8165 : n9275;
  assign n9277 = pi17 ? n3155 : ~n9030;
  assign n9278 = pi16 ? n32 : n9277;
  assign n9279 = pi17 ? n3155 : ~n8193;
  assign n9280 = pi16 ? n32 : n9279;
  assign n9281 = pi15 ? n9278 : n9280;
  assign n9282 = pi14 ? n9276 : n9281;
  assign n9283 = pi17 ? n3155 : ~n9039;
  assign n9284 = pi16 ? n32 : n9283;
  assign n9285 = pi17 ? n2954 : ~n9039;
  assign n9286 = pi16 ? n32 : n9285;
  assign n9287 = pi15 ? n9284 : n9286;
  assign n9288 = pi17 ? n2954 : ~n8193;
  assign n9289 = pi16 ? n32 : n9288;
  assign n9290 = pi17 ? n4111 : ~n8204;
  assign n9291 = pi16 ? n32 : n9290;
  assign n9292 = pi15 ? n9289 : n9291;
  assign n9293 = pi14 ? n9287 : n9292;
  assign n9294 = pi13 ? n9282 : n9293;
  assign n9295 = pi17 ? n3160 : ~n8193;
  assign n9296 = pi16 ? n32 : n9295;
  assign n9297 = pi17 ? n3160 : ~n8204;
  assign n9298 = pi16 ? n32 : n9297;
  assign n9299 = pi15 ? n9296 : n9298;
  assign n9300 = pi17 ? n3160 : ~n7369;
  assign n9301 = pi16 ? n32 : n9300;
  assign n9302 = pi17 ? n3160 : ~n9056;
  assign n9303 = pi16 ? n32 : n9302;
  assign n9304 = pi15 ? n9301 : n9303;
  assign n9305 = pi14 ? n9299 : n9304;
  assign n9306 = pi17 ? n3164 : ~n9062;
  assign n9307 = pi16 ? n32 : n9306;
  assign n9308 = pi17 ? n3046 : ~n8232;
  assign n9309 = pi16 ? n32 : n9308;
  assign n9310 = pi15 ? n9307 : n9309;
  assign n9311 = pi18 ? n32 : n1741;
  assign n9312 = pi17 ? n2959 : ~n9311;
  assign n9313 = pi16 ? n32 : n9312;
  assign n9314 = pi17 ? n2959 : ~n9073;
  assign n9315 = pi16 ? n32 : n9314;
  assign n9316 = pi15 ? n9313 : n9315;
  assign n9317 = pi14 ? n9310 : n9316;
  assign n9318 = pi13 ? n9305 : n9317;
  assign n9319 = pi12 ? n9294 : n9318;
  assign n9320 = pi11 ? n9273 : n9319;
  assign n9321 = pi20 ? n246 : n339;
  assign n9322 = pi19 ? n32 : n9321;
  assign n9323 = pi18 ? n32 : n9322;
  assign n9324 = pi17 ? n2959 : ~n9323;
  assign n9325 = pi16 ? n32 : n9324;
  assign n9326 = pi22 ? n32 : ~n84;
  assign n9327 = pi21 ? n9326 : n206;
  assign n9328 = pi20 ? n9327 : ~n32;
  assign n9329 = pi19 ? n32 : n9328;
  assign n9330 = pi18 ? n32 : n9329;
  assign n9331 = pi17 ? n2959 : ~n9330;
  assign n9332 = pi16 ? n32 : n9331;
  assign n9333 = pi15 ? n9325 : n9332;
  assign n9334 = pi17 ? n2959 : ~n3067;
  assign n9335 = pi16 ? n32 : n9334;
  assign n9336 = pi17 ? n2952 : ~n2736;
  assign n9337 = pi16 ? n32 : n9336;
  assign n9338 = pi15 ? n9335 : n9337;
  assign n9339 = pi14 ? n9333 : n9338;
  assign n9340 = pi20 ? n5854 : n141;
  assign n9341 = pi19 ? n32 : n9340;
  assign n9342 = pi18 ? n32 : n9341;
  assign n9343 = pi17 ? n3175 : ~n9342;
  assign n9344 = pi16 ? n32 : n9343;
  assign n9345 = pi20 ? n220 : ~n32;
  assign n9346 = pi19 ? n32 : n9345;
  assign n9347 = pi18 ? n32 : n9346;
  assign n9348 = pi17 ? n3175 : ~n9347;
  assign n9349 = pi16 ? n32 : n9348;
  assign n9350 = pi15 ? n9344 : n9349;
  assign n9351 = pi20 ? n653 : n141;
  assign n9352 = pi19 ? n32 : n9351;
  assign n9353 = pi18 ? n32 : n9352;
  assign n9354 = pi17 ? n3175 : ~n9353;
  assign n9355 = pi16 ? n32 : n9354;
  assign n9356 = pi17 ? n3175 : ~n9103;
  assign n9357 = pi16 ? n32 : n9356;
  assign n9358 = pi15 ? n9355 : n9357;
  assign n9359 = pi14 ? n9350 : n9358;
  assign n9360 = pi13 ? n9339 : n9359;
  assign n9361 = pi21 ? n405 : ~n1009;
  assign n9362 = pi20 ? n9361 : ~n32;
  assign n9363 = pi19 ? n32 : n9362;
  assign n9364 = pi18 ? n32 : n9363;
  assign n9365 = pi17 ? n3175 : ~n9364;
  assign n9366 = pi16 ? n32 : n9365;
  assign n9367 = pi21 ? n174 : n140;
  assign n9368 = pi20 ? n9367 : ~n32;
  assign n9369 = pi19 ? n32 : n9368;
  assign n9370 = pi18 ? n32 : n9369;
  assign n9371 = pi17 ? n3175 : ~n9370;
  assign n9372 = pi16 ? n32 : n9371;
  assign n9373 = pi15 ? n9366 : n9372;
  assign n9374 = pi21 ? n174 : ~n7500;
  assign n9375 = pi20 ? n9374 : ~n32;
  assign n9376 = pi19 ? n32 : n9375;
  assign n9377 = pi18 ? n32 : n9376;
  assign n9378 = pi17 ? n3175 : ~n9377;
  assign n9379 = pi16 ? n32 : n9378;
  assign n9380 = pi17 ? n2831 : ~n2733;
  assign n9381 = pi16 ? n32 : n9380;
  assign n9382 = pi15 ? n9379 : n9381;
  assign n9383 = pi14 ? n9373 : n9382;
  assign n9384 = pi17 ? n2831 : ~n2724;
  assign n9385 = pi16 ? n32 : n9384;
  assign n9386 = pi15 ? n9381 : n9385;
  assign n9387 = pi17 ? n2726 : ~n2850;
  assign n9388 = pi16 ? n32 : n9387;
  assign n9389 = pi17 ? n2963 : ~n2724;
  assign n9390 = pi16 ? n32 : n9389;
  assign n9391 = pi15 ? n9388 : n9390;
  assign n9392 = pi14 ? n9386 : n9391;
  assign n9393 = pi13 ? n9383 : n9392;
  assign n9394 = pi12 ? n9360 : n9393;
  assign n9395 = pi17 ? n2963 : ~n2850;
  assign n9396 = pi16 ? n32 : n9395;
  assign n9397 = pi17 ? n2963 : ~n2736;
  assign n9398 = pi16 ? n32 : n9397;
  assign n9399 = pi15 ? n9396 : n9398;
  assign n9400 = pi15 ? n9390 : n9398;
  assign n9401 = pi14 ? n9399 : n9400;
  assign n9402 = pi17 ? n2726 : ~n2736;
  assign n9403 = pi16 ? n32 : n9402;
  assign n9404 = pi17 ? n2726 : ~n2750;
  assign n9405 = pi16 ? n32 : n9404;
  assign n9406 = pi15 ? n9403 : n9405;
  assign n9407 = pi17 ? n2726 : ~n2855;
  assign n9408 = pi16 ? n32 : n9407;
  assign n9409 = pi17 ? n3050 : ~n2750;
  assign n9410 = pi16 ? n32 : n9409;
  assign n9411 = pi15 ? n9408 : n9410;
  assign n9412 = pi14 ? n9406 : n9411;
  assign n9413 = pi13 ? n9401 : n9412;
  assign n9414 = pi17 ? n3050 : ~n2623;
  assign n9415 = pi16 ? n32 : n9414;
  assign n9416 = pi17 ? n3050 : ~n2618;
  assign n9417 = pi16 ? n32 : n9416;
  assign n9418 = pi15 ? n9415 : n9417;
  assign n9419 = pi17 ? n2959 : ~n2618;
  assign n9420 = pi16 ? n32 : n9419;
  assign n9421 = pi15 ? n9417 : n9420;
  assign n9422 = pi14 ? n9418 : n9421;
  assign n9423 = pi17 ? n2959 : ~n2628;
  assign n9424 = pi16 ? n32 : n9423;
  assign n9425 = pi21 ? n405 : n1939;
  assign n9426 = pi20 ? n32 : n9425;
  assign n9427 = pi19 ? n9426 : ~n32;
  assign n9428 = pi18 ? n32 : n9427;
  assign n9429 = pi17 ? n2959 : ~n9428;
  assign n9430 = pi16 ? n32 : n9429;
  assign n9431 = pi15 ? n9424 : n9430;
  assign n9432 = pi17 ? n3046 : ~n9173;
  assign n9433 = pi16 ? n32 : n9432;
  assign n9434 = pi17 ? n2959 : ~n2519;
  assign n9435 = pi16 ? n32 : n9434;
  assign n9436 = pi15 ? n9433 : n9435;
  assign n9437 = pi14 ? n9431 : n9436;
  assign n9438 = pi13 ? n9422 : n9437;
  assign n9439 = pi12 ? n9413 : n9438;
  assign n9440 = pi11 ? n9394 : n9439;
  assign n9441 = pi10 ? n9320 : n9440;
  assign n9442 = pi09 ? n9207 : n9441;
  assign n9443 = pi08 ? n9184 : n9442;
  assign n9444 = pi18 ? n2627 : ~n7647;
  assign n9445 = pi17 ? n32 : n9444;
  assign n9446 = pi16 ? n32 : n9445;
  assign n9447 = pi15 ? n32 : n9446;
  assign n9448 = pi18 ? n605 : ~n8086;
  assign n9449 = pi17 ? n32 : n9448;
  assign n9450 = pi16 ? n32 : n9449;
  assign n9451 = pi15 ? n9446 : n9450;
  assign n9452 = pi14 ? n9447 : n9451;
  assign n9453 = pi13 ? n32 : n9452;
  assign n9454 = pi12 ? n32 : n9453;
  assign n9455 = pi11 ? n32 : n9454;
  assign n9456 = pi10 ? n32 : n9455;
  assign n9457 = pi19 ? n6398 : n343;
  assign n9458 = pi18 ? n2424 : ~n9457;
  assign n9459 = pi17 ? n32 : n9458;
  assign n9460 = pi16 ? n32 : n9459;
  assign n9461 = pi19 ? n507 : n349;
  assign n9462 = pi18 ? n418 : ~n9461;
  assign n9463 = pi17 ? n32 : n9462;
  assign n9464 = pi16 ? n32 : n9463;
  assign n9465 = pi15 ? n9460 : n9464;
  assign n9466 = pi18 ? n418 : ~n8192;
  assign n9467 = pi17 ? n32 : n9466;
  assign n9468 = pi16 ? n32 : n9467;
  assign n9469 = pi19 ? n1464 : n6396;
  assign n9470 = pi18 ? n3786 : ~n9469;
  assign n9471 = pi17 ? n32 : n9470;
  assign n9472 = pi16 ? n32 : n9471;
  assign n9473 = pi15 ? n9468 : n9472;
  assign n9474 = pi14 ? n9465 : n9473;
  assign n9475 = pi19 ? n750 : n813;
  assign n9476 = pi18 ? n3786 : ~n9475;
  assign n9477 = pi17 ? n32 : n9476;
  assign n9478 = pi16 ? n32 : n9477;
  assign n9479 = pi20 ? n1817 : n7839;
  assign n9480 = pi19 ? n365 : ~n9479;
  assign n9481 = pi18 ? n9480 : ~n496;
  assign n9482 = pi17 ? n32 : n9481;
  assign n9483 = pi16 ? n32 : n9482;
  assign n9484 = pi15 ? n9478 : n9483;
  assign n9485 = pi22 ? n173 : ~n65;
  assign n9486 = pi21 ? n7659 : ~n9485;
  assign n9487 = pi20 ? n32 : ~n9486;
  assign n9488 = pi21 ? n173 : n174;
  assign n9489 = pi20 ? n9488 : n6050;
  assign n9490 = pi19 ? n9487 : ~n9489;
  assign n9491 = pi21 ? n309 : ~n309;
  assign n9492 = pi20 ? n9491 : n207;
  assign n9493 = pi19 ? n9492 : ~n32;
  assign n9494 = pi18 ? n9490 : ~n9493;
  assign n9495 = pi17 ? n32 : n9494;
  assign n9496 = pi16 ? n32 : n9495;
  assign n9497 = pi19 ? n1812 : n236;
  assign n9498 = pi18 ? n9497 : ~n8951;
  assign n9499 = pi17 ? n32 : n9498;
  assign n9500 = pi16 ? n32 : n9499;
  assign n9501 = pi15 ? n9496 : n9500;
  assign n9502 = pi14 ? n9484 : n9501;
  assign n9503 = pi13 ? n9474 : n9502;
  assign n9504 = pi18 ? n814 : ~n8192;
  assign n9505 = pi17 ? n32 : n9504;
  assign n9506 = pi16 ? n32 : n9505;
  assign n9507 = pi15 ? n8959 : n9506;
  assign n9508 = pi19 ? n813 : n617;
  assign n9509 = pi19 ? n340 : n236;
  assign n9510 = pi18 ? n9508 : ~n9509;
  assign n9511 = pi17 ? n32 : n9510;
  assign n9512 = pi16 ? n32 : n9511;
  assign n9513 = pi15 ? n9512 : n8973;
  assign n9514 = pi14 ? n9507 : n9513;
  assign n9515 = pi19 ? n1941 : n617;
  assign n9516 = pi18 ? n9515 : ~n880;
  assign n9517 = pi17 ? n32 : n9516;
  assign n9518 = pi16 ? n32 : n9517;
  assign n9519 = pi18 ? n237 : ~n9002;
  assign n9520 = pi17 ? n32 : n9519;
  assign n9521 = pi16 ? n32 : n9520;
  assign n9522 = pi15 ? n9518 : n9521;
  assign n9523 = pi19 ? n6307 : ~n176;
  assign n9524 = pi20 ? n1331 : ~n342;
  assign n9525 = pi19 ? n9524 : n349;
  assign n9526 = pi18 ? n9523 : ~n9525;
  assign n9527 = pi17 ? n32 : n9526;
  assign n9528 = pi16 ? n32 : n9527;
  assign n9529 = pi18 ? n618 : ~n9266;
  assign n9530 = pi17 ? n32 : n9529;
  assign n9531 = pi16 ? n32 : n9530;
  assign n9532 = pi15 ? n9528 : n9531;
  assign n9533 = pi14 ? n9522 : n9532;
  assign n9534 = pi13 ? n9514 : n9533;
  assign n9535 = pi12 ? n9503 : n9534;
  assign n9536 = pi20 ? n339 : ~n175;
  assign n9537 = pi19 ? n9536 : ~n9169;
  assign n9538 = pi19 ? n261 : n617;
  assign n9539 = pi18 ? n9537 : ~n9538;
  assign n9540 = pi17 ? n32 : n9539;
  assign n9541 = pi16 ? n32 : n9540;
  assign n9542 = pi15 ? n8362 : n9541;
  assign n9543 = pi20 ? n321 : ~n260;
  assign n9544 = pi19 ? n32 : n9543;
  assign n9545 = pi18 ? n1676 : ~n9544;
  assign n9546 = pi17 ? n32 : n9545;
  assign n9547 = pi16 ? n32 : n9546;
  assign n9548 = pi20 ? n141 : ~n175;
  assign n9549 = pi19 ? n9548 : ~n32;
  assign n9550 = pi18 ? n9549 : ~n8192;
  assign n9551 = pi17 ? n32 : n9550;
  assign n9552 = pi16 ? n32 : n9551;
  assign n9553 = pi15 ? n9547 : n9552;
  assign n9554 = pi14 ? n9542 : n9553;
  assign n9555 = pi18 ? n1676 : ~n8192;
  assign n9556 = pi17 ? n32 : n9555;
  assign n9557 = pi16 ? n32 : n9556;
  assign n9558 = pi20 ? n141 : ~n3843;
  assign n9559 = pi20 ? n246 : n357;
  assign n9560 = pi19 ? n9558 : ~n9559;
  assign n9561 = pi19 ? n261 : n321;
  assign n9562 = pi18 ? n9560 : ~n9561;
  assign n9563 = pi17 ? n32 : n9562;
  assign n9564 = pi16 ? n32 : n9563;
  assign n9565 = pi15 ? n9557 : n9564;
  assign n9566 = pi17 ? n3569 : ~n8198;
  assign n9567 = pi16 ? n32 : n9566;
  assign n9568 = pi17 ? n3569 : ~n8214;
  assign n9569 = pi16 ? n32 : n9568;
  assign n9570 = pi15 ? n9567 : n9569;
  assign n9571 = pi14 ? n9565 : n9570;
  assign n9572 = pi13 ? n9554 : n9571;
  assign n9573 = pi17 ? n3282 : ~n8204;
  assign n9574 = pi16 ? n32 : n9573;
  assign n9575 = pi17 ? n3282 : ~n8214;
  assign n9576 = pi16 ? n32 : n9575;
  assign n9577 = pi15 ? n9574 : n9576;
  assign n9578 = pi19 ? n1818 : n32;
  assign n9579 = pi18 ? n9578 : n7368;
  assign n9580 = pi17 ? n3282 : ~n9579;
  assign n9581 = pi16 ? n32 : n9580;
  assign n9582 = pi20 ? n1324 : ~n274;
  assign n9583 = pi19 ? n32 : n9582;
  assign n9584 = pi18 ? n32 : n9583;
  assign n9585 = pi17 ? n3155 : ~n9584;
  assign n9586 = pi16 ? n32 : n9585;
  assign n9587 = pi15 ? n9581 : n9586;
  assign n9588 = pi14 ? n9577 : n9587;
  assign n9589 = pi20 ? n1331 : ~n339;
  assign n9590 = pi19 ? n5350 : n9589;
  assign n9591 = pi20 ? n428 : ~n321;
  assign n9592 = pi20 ? n220 : n274;
  assign n9593 = pi19 ? n9591 : ~n9592;
  assign n9594 = pi18 ? n9590 : n9593;
  assign n9595 = pi17 ? n3155 : ~n9594;
  assign n9596 = pi16 ? n32 : n9595;
  assign n9597 = pi20 ? n1385 : n749;
  assign n9598 = pi19 ? n32 : n9597;
  assign n9599 = pi18 ? n32 : n9598;
  assign n9600 = pi17 ? n3728 : ~n9599;
  assign n9601 = pi16 ? n32 : n9600;
  assign n9602 = pi15 ? n9596 : n9601;
  assign n9603 = pi17 ? n3728 : ~n8588;
  assign n9604 = pi16 ? n32 : n9603;
  assign n9605 = pi14 ? n9602 : n9604;
  assign n9606 = pi13 ? n9588 : n9605;
  assign n9607 = pi12 ? n9572 : n9606;
  assign n9608 = pi11 ? n9535 : n9607;
  assign n9609 = pi17 ? n3728 : ~n7039;
  assign n9610 = pi16 ? n32 : n9609;
  assign n9611 = pi19 ? n176 : n4406;
  assign n9612 = pi18 ? n7221 : n9611;
  assign n9613 = pi17 ? n3728 : ~n9612;
  assign n9614 = pi16 ? n32 : n9613;
  assign n9615 = pi15 ? n9610 : n9614;
  assign n9616 = pi17 ? n4111 : ~n8607;
  assign n9617 = pi16 ? n32 : n9616;
  assign n9618 = pi21 ? n7107 : ~n32;
  assign n9619 = pi20 ? n9618 : n339;
  assign n9620 = pi19 ? n32 : n9619;
  assign n9621 = pi18 ? n32 : n9620;
  assign n9622 = pi17 ? n3160 : ~n9621;
  assign n9623 = pi16 ? n32 : n9622;
  assign n9624 = pi15 ? n9617 : n9623;
  assign n9625 = pi14 ? n9615 : n9624;
  assign n9626 = pi17 ? n3292 : ~n7039;
  assign n9627 = pi16 ? n32 : n9626;
  assign n9628 = pi21 ? n100 : n206;
  assign n9629 = pi20 ? n9628 : ~n32;
  assign n9630 = pi19 ? n32 : n9629;
  assign n9631 = pi18 ? n32 : n9630;
  assign n9632 = pi17 ? n3292 : ~n9631;
  assign n9633 = pi16 ? n32 : n9632;
  assign n9634 = pi17 ? n3292 : ~n2850;
  assign n9635 = pi16 ? n32 : n9634;
  assign n9636 = pi15 ? n9633 : n9635;
  assign n9637 = pi14 ? n9627 : n9636;
  assign n9638 = pi13 ? n9625 : n9637;
  assign n9639 = pi21 ? n259 : ~n7659;
  assign n9640 = pi20 ? n175 : ~n9639;
  assign n9641 = pi21 ? n32 : ~n313;
  assign n9642 = pi20 ? n9641 : n1331;
  assign n9643 = pi19 ? n9640 : n9642;
  assign n9644 = pi20 ? n7942 : n32;
  assign n9645 = pi21 ? n206 : ~n454;
  assign n9646 = pi20 ? n9645 : ~n32;
  assign n9647 = pi19 ? n9644 : n9646;
  assign n9648 = pi18 ? n9643 : n9647;
  assign n9649 = pi17 ? n3292 : ~n9648;
  assign n9650 = pi16 ? n32 : n9649;
  assign n9651 = pi21 ? n405 : n8275;
  assign n9652 = pi20 ? n9651 : ~n32;
  assign n9653 = pi19 ? n32 : n9652;
  assign n9654 = pi18 ? n32 : n9653;
  assign n9655 = pi17 ? n3587 : ~n9654;
  assign n9656 = pi16 ? n32 : n9655;
  assign n9657 = pi15 ? n9650 : n9656;
  assign n9658 = pi17 ? n3175 : ~n3781;
  assign n9659 = pi16 ? n32 : n9658;
  assign n9660 = pi15 ? n7546 : n9659;
  assign n9661 = pi14 ? n9657 : n9660;
  assign n9662 = pi17 ? n2959 : ~n2724;
  assign n9663 = pi16 ? n32 : n9662;
  assign n9664 = pi17 ? n2959 : ~n3763;
  assign n9665 = pi16 ? n32 : n9664;
  assign n9666 = pi15 ? n9663 : n9665;
  assign n9667 = pi21 ? n405 : n140;
  assign n9668 = pi20 ? n9667 : ~n32;
  assign n9669 = pi19 ? n32 : n9668;
  assign n9670 = pi18 ? n32 : n9669;
  assign n9671 = pi17 ? n3587 : ~n9670;
  assign n9672 = pi16 ? n32 : n9671;
  assign n9673 = pi15 ? n9672 : n9335;
  assign n9674 = pi14 ? n9666 : n9673;
  assign n9675 = pi13 ? n9661 : n9674;
  assign n9676 = pi12 ? n9638 : n9675;
  assign n9677 = pi17 ? n2959 : ~n2850;
  assign n9678 = pi16 ? n32 : n9677;
  assign n9679 = pi15 ? n9678 : n9663;
  assign n9680 = pi17 ? n2959 : ~n2736;
  assign n9681 = pi16 ? n32 : n9680;
  assign n9682 = pi15 ? n9663 : n9681;
  assign n9683 = pi14 ? n9679 : n9682;
  assign n9684 = pi17 ? n3046 : ~n2855;
  assign n9685 = pi16 ? n32 : n9684;
  assign n9686 = pi15 ? n9681 : n9685;
  assign n9687 = pi17 ? n3046 : ~n2616;
  assign n9688 = pi16 ? n32 : n9687;
  assign n9689 = pi17 ? n3164 : ~n2623;
  assign n9690 = pi16 ? n32 : n9689;
  assign n9691 = pi15 ? n9688 : n9690;
  assign n9692 = pi14 ? n9686 : n9691;
  assign n9693 = pi13 ? n9683 : n9692;
  assign n9694 = pi17 ? n3164 : ~n3621;
  assign n9695 = pi16 ? n32 : n9694;
  assign n9696 = pi15 ? n9690 : n9695;
  assign n9697 = pi17 ? n3164 : ~n2618;
  assign n9698 = pi16 ? n32 : n9697;
  assign n9699 = pi15 ? n9698 : n9695;
  assign n9700 = pi14 ? n9696 : n9699;
  assign n9701 = pi17 ? n3728 : ~n2628;
  assign n9702 = pi16 ? n32 : n9701;
  assign n9703 = pi17 ? n3728 : ~n2748;
  assign n9704 = pi16 ? n32 : n9703;
  assign n9705 = pi15 ? n9702 : n9704;
  assign n9706 = pi17 ? n2954 : ~n2519;
  assign n9707 = pi16 ? n32 : n9706;
  assign n9708 = pi17 ? n3728 : ~n2519;
  assign n9709 = pi16 ? n32 : n9708;
  assign n9710 = pi15 ? n9707 : n9709;
  assign n9711 = pi14 ? n9705 : n9710;
  assign n9712 = pi13 ? n9700 : n9711;
  assign n9713 = pi12 ? n9693 : n9712;
  assign n9714 = pi11 ? n9676 : n9713;
  assign n9715 = pi10 ? n9608 : n9714;
  assign n9716 = pi09 ? n9456 : n9715;
  assign n9717 = pi18 ? n1750 : ~n7647;
  assign n9718 = pi17 ? n32 : n9717;
  assign n9719 = pi16 ? n32 : n9718;
  assign n9720 = pi15 ? n32 : n9719;
  assign n9721 = pi18 ? n2622 : ~n7647;
  assign n9722 = pi17 ? n32 : n9721;
  assign n9723 = pi16 ? n32 : n9722;
  assign n9724 = pi20 ? n1685 : n32;
  assign n9725 = pi19 ? n507 : ~n9724;
  assign n9726 = pi18 ? n323 : ~n9725;
  assign n9727 = pi17 ? n32 : n9726;
  assign n9728 = pi16 ? n32 : n9727;
  assign n9729 = pi15 ? n9723 : n9728;
  assign n9730 = pi14 ? n9720 : n9729;
  assign n9731 = pi13 ? n32 : n9730;
  assign n9732 = pi12 ? n32 : n9731;
  assign n9733 = pi11 ? n32 : n9732;
  assign n9734 = pi10 ? n32 : n9733;
  assign n9735 = pi18 ? n2291 : ~n684;
  assign n9736 = pi17 ? n32 : n9735;
  assign n9737 = pi16 ? n32 : n9736;
  assign n9738 = pi18 ? n797 : ~n9461;
  assign n9739 = pi17 ? n32 : n9738;
  assign n9740 = pi16 ? n32 : n9739;
  assign n9741 = pi15 ? n9737 : n9740;
  assign n9742 = pi18 ? n797 : ~n8192;
  assign n9743 = pi17 ? n32 : n9742;
  assign n9744 = pi16 ? n32 : n9743;
  assign n9745 = pi19 ? n6398 : n321;
  assign n9746 = pi18 ? n2413 : ~n9745;
  assign n9747 = pi17 ? n32 : n9746;
  assign n9748 = pi16 ? n32 : n9747;
  assign n9749 = pi15 ? n9744 : n9748;
  assign n9750 = pi14 ? n9741 : n9749;
  assign n9751 = pi19 ? n322 : n813;
  assign n9752 = pi18 ? n2413 : ~n9751;
  assign n9753 = pi17 ? n32 : n9752;
  assign n9754 = pi16 ? n32 : n9753;
  assign n9755 = pi19 ? n1969 : ~n1818;
  assign n9756 = pi18 ? n9755 : ~n496;
  assign n9757 = pi17 ? n32 : n9756;
  assign n9758 = pi16 ? n32 : n9757;
  assign n9759 = pi15 ? n9754 : n9758;
  assign n9760 = pi20 ? n1331 : n7839;
  assign n9761 = pi19 ? n244 : ~n9760;
  assign n9762 = pi20 ? n1611 : n749;
  assign n9763 = pi19 ? n9762 : ~n5614;
  assign n9764 = pi18 ? n9761 : ~n9763;
  assign n9765 = pi17 ? n32 : n9764;
  assign n9766 = pi16 ? n32 : n9765;
  assign n9767 = pi19 ? n429 : n617;
  assign n9768 = pi19 ? n750 : n349;
  assign n9769 = pi18 ? n9767 : ~n9768;
  assign n9770 = pi17 ? n32 : n9769;
  assign n9771 = pi16 ? n32 : n9770;
  assign n9772 = pi15 ? n9766 : n9771;
  assign n9773 = pi14 ? n9759 : n9772;
  assign n9774 = pi13 ? n9750 : n9773;
  assign n9775 = pi19 ? n6057 : n321;
  assign n9776 = pi18 ? n430 : ~n9775;
  assign n9777 = pi17 ? n32 : n9776;
  assign n9778 = pi16 ? n32 : n9777;
  assign n9779 = pi18 ? n430 : ~n8192;
  assign n9780 = pi17 ? n32 : n9779;
  assign n9781 = pi16 ? n32 : n9780;
  assign n9782 = pi15 ? n9778 : n9781;
  assign n9783 = pi19 ? n208 : n813;
  assign n9784 = pi18 ? n2304 : ~n9783;
  assign n9785 = pi17 ? n32 : n9784;
  assign n9786 = pi16 ? n32 : n9785;
  assign n9787 = pi18 ? n2304 : ~n8516;
  assign n9788 = pi17 ? n32 : n9787;
  assign n9789 = pi16 ? n32 : n9788;
  assign n9790 = pi15 ? n9786 : n9789;
  assign n9791 = pi14 ? n9782 : n9790;
  assign n9792 = pi18 ? n344 : ~n880;
  assign n9793 = pi17 ? n32 : n9792;
  assign n9794 = pi16 ? n32 : n9793;
  assign n9795 = pi18 ? n1813 : ~n9002;
  assign n9796 = pi17 ? n32 : n9795;
  assign n9797 = pi16 ? n32 : n9796;
  assign n9798 = pi15 ? n9794 : n9797;
  assign n9799 = pi20 ? n749 : ~n175;
  assign n9800 = pi19 ? n9799 : ~n32;
  assign n9801 = pi19 ? n261 : n349;
  assign n9802 = pi18 ? n9800 : ~n9801;
  assign n9803 = pi17 ? n32 : n9802;
  assign n9804 = pi16 ? n32 : n9803;
  assign n9805 = pi19 ? n916 : n8383;
  assign n9806 = pi18 ? n814 : ~n9805;
  assign n9807 = pi17 ? n32 : n9806;
  assign n9808 = pi16 ? n32 : n9807;
  assign n9809 = pi15 ? n9804 : n9808;
  assign n9810 = pi14 ? n9798 : n9809;
  assign n9811 = pi13 ? n9791 : n9810;
  assign n9812 = pi12 ? n9774 : n9811;
  assign n9813 = pi18 ? n814 : ~n7994;
  assign n9814 = pi17 ? n32 : n9813;
  assign n9815 = pi16 ? n32 : n9814;
  assign n9816 = pi20 ? n207 : n141;
  assign n9817 = pi19 ? n261 : n9816;
  assign n9818 = pi18 ? n1942 : ~n9817;
  assign n9819 = pi17 ? n32 : n9818;
  assign n9820 = pi16 ? n32 : n9819;
  assign n9821 = pi15 ? n9815 : n9820;
  assign n9822 = pi20 ? n321 : n342;
  assign n9823 = pi19 ? n32 : n9822;
  assign n9824 = pi18 ? n1942 : ~n9823;
  assign n9825 = pi17 ? n32 : n9824;
  assign n9826 = pi16 ? n32 : n9825;
  assign n9827 = pi18 ? n1942 : ~n8192;
  assign n9828 = pi17 ? n32 : n9827;
  assign n9829 = pi16 ? n32 : n9828;
  assign n9830 = pi15 ? n9826 : n9829;
  assign n9831 = pi14 ? n9821 : n9830;
  assign n9832 = pi19 ? n2614 : ~n9169;
  assign n9833 = pi18 ? n9832 : ~n9561;
  assign n9834 = pi17 ? n32 : n9833;
  assign n9835 = pi16 ? n32 : n9834;
  assign n9836 = pi15 ? n9829 : n9835;
  assign n9837 = pi18 ? n3350 : ~n8197;
  assign n9838 = pi17 ? n32 : n9837;
  assign n9839 = pi16 ? n32 : n9838;
  assign n9840 = pi18 ? n3350 : ~n8213;
  assign n9841 = pi17 ? n32 : n9840;
  assign n9842 = pi16 ? n32 : n9841;
  assign n9843 = pi15 ? n9839 : n9842;
  assign n9844 = pi14 ? n9836 : n9843;
  assign n9845 = pi13 ? n9831 : n9844;
  assign n9846 = pi20 ? n1385 : n1839;
  assign n9847 = pi19 ? n32 : n9846;
  assign n9848 = pi18 ? n618 : ~n9847;
  assign n9849 = pi17 ? n32 : n9848;
  assign n9850 = pi16 ? n32 : n9849;
  assign n9851 = pi18 ? n618 : ~n8213;
  assign n9852 = pi17 ? n32 : n9851;
  assign n9853 = pi16 ? n32 : n9852;
  assign n9854 = pi15 ? n9850 : n9853;
  assign n9855 = pi18 ? n618 : ~n7368;
  assign n9856 = pi17 ? n32 : n9855;
  assign n9857 = pi16 ? n32 : n9856;
  assign n9858 = pi18 ? n618 : ~n9583;
  assign n9859 = pi17 ? n32 : n9858;
  assign n9860 = pi16 ? n32 : n9859;
  assign n9861 = pi15 ? n9857 : n9860;
  assign n9862 = pi14 ? n9854 : n9861;
  assign n9863 = pi21 ? n405 : ~n259;
  assign n9864 = pi20 ? n32 : n9863;
  assign n9865 = pi19 ? n9864 : n32;
  assign n9866 = pi20 ? n1611 : ~n274;
  assign n9867 = pi19 ? n5694 : n9866;
  assign n9868 = pi18 ? n9865 : n9867;
  assign n9869 = pi17 ? n32 : ~n9868;
  assign n9870 = pi16 ? n32 : n9869;
  assign n9871 = pi17 ? n32 : ~n9599;
  assign n9872 = pi16 ? n32 : n9871;
  assign n9873 = pi15 ? n9870 : n9872;
  assign n9874 = pi20 ? n175 : n1940;
  assign n9875 = pi19 ? n32 : n9874;
  assign n9876 = pi18 ? n32 : n9875;
  assign n9877 = pi17 ? n32 : ~n9876;
  assign n9878 = pi16 ? n32 : n9877;
  assign n9879 = pi14 ? n9873 : n9878;
  assign n9880 = pi13 ? n9862 : n9879;
  assign n9881 = pi12 ? n9845 : n9880;
  assign n9882 = pi11 ? n9812 : n9881;
  assign n9883 = pi17 ? n32 : ~n7039;
  assign n9884 = pi16 ? n32 : n9883;
  assign n9885 = pi17 ? n3569 : ~n9330;
  assign n9886 = pi16 ? n32 : n9885;
  assign n9887 = pi15 ? n9884 : n9886;
  assign n9888 = pi17 ? n3569 : ~n8249;
  assign n9889 = pi16 ? n32 : n9888;
  assign n9890 = pi20 ? n501 : n339;
  assign n9891 = pi19 ? n32 : n9890;
  assign n9892 = pi18 ? n32 : n9891;
  assign n9893 = pi17 ? n4111 : ~n9892;
  assign n9894 = pi16 ? n32 : n9893;
  assign n9895 = pi15 ? n9889 : n9894;
  assign n9896 = pi14 ? n9887 : n9895;
  assign n9897 = pi21 ? n100 : ~n206;
  assign n9898 = pi20 ? n9897 : n141;
  assign n9899 = pi19 ? n32 : n9898;
  assign n9900 = pi18 ? n32 : n9899;
  assign n9901 = pi17 ? n3155 : ~n9900;
  assign n9902 = pi16 ? n32 : n9901;
  assign n9903 = pi20 ? n246 : n141;
  assign n9904 = pi19 ? n32 : n9903;
  assign n9905 = pi18 ? n32 : n9904;
  assign n9906 = pi17 ? n4111 : ~n9905;
  assign n9907 = pi16 ? n32 : n9906;
  assign n9908 = pi15 ? n9902 : n9907;
  assign n9909 = pi17 ? n3155 : ~n3781;
  assign n9910 = pi16 ? n32 : n9909;
  assign n9911 = pi17 ? n3155 : ~n2850;
  assign n9912 = pi16 ? n32 : n9911;
  assign n9913 = pi15 ? n9910 : n9912;
  assign n9914 = pi14 ? n9908 : n9913;
  assign n9915 = pi13 ? n9896 : n9914;
  assign n9916 = pi19 ? n8622 : n4670;
  assign n9917 = pi19 ? n247 : n9646;
  assign n9918 = pi18 ? n9916 : n9917;
  assign n9919 = pi17 ? n2954 : ~n9918;
  assign n9920 = pi16 ? n32 : n9919;
  assign n9921 = pi20 ? n8943 : ~n32;
  assign n9922 = pi19 ? n32 : n9921;
  assign n9923 = pi18 ? n32 : n9922;
  assign n9924 = pi17 ? n2954 : ~n9923;
  assign n9925 = pi16 ? n32 : n9924;
  assign n9926 = pi15 ? n9920 : n9925;
  assign n9927 = pi17 ? n3164 : ~n3781;
  assign n9928 = pi16 ? n32 : n9927;
  assign n9929 = pi15 ? n7743 : n9928;
  assign n9930 = pi14 ? n9926 : n9929;
  assign n9931 = pi17 ? n3160 : ~n2724;
  assign n9932 = pi16 ? n32 : n9931;
  assign n9933 = pi17 ? n3160 : ~n3763;
  assign n9934 = pi16 ? n32 : n9933;
  assign n9935 = pi15 ? n9932 : n9934;
  assign n9936 = pi19 ? n1818 : n2848;
  assign n9937 = pi18 ? n32 : n9936;
  assign n9938 = pi17 ? n3164 : ~n9937;
  assign n9939 = pi16 ? n32 : n9938;
  assign n9940 = pi15 ? n9026 : n9939;
  assign n9941 = pi14 ? n9935 : n9940;
  assign n9942 = pi13 ? n9930 : n9941;
  assign n9943 = pi12 ? n9915 : n9942;
  assign n9944 = pi19 ? n472 : n1812;
  assign n9945 = pi18 ? n32 : n9944;
  assign n9946 = pi17 ? n3164 : ~n9945;
  assign n9947 = pi16 ? n32 : n9946;
  assign n9948 = pi17 ? n3164 : ~n4245;
  assign n9949 = pi16 ? n32 : n9948;
  assign n9950 = pi15 ? n9947 : n9949;
  assign n9951 = pi17 ? n3164 : ~n2736;
  assign n9952 = pi16 ? n32 : n9951;
  assign n9953 = pi17 ? n3728 : ~n2736;
  assign n9954 = pi16 ? n32 : n9953;
  assign n9955 = pi15 ? n9952 : n9954;
  assign n9956 = pi14 ? n9950 : n9955;
  assign n9957 = pi17 ? n2954 : ~n2616;
  assign n9958 = pi16 ? n32 : n9957;
  assign n9959 = pi15 ? n9954 : n9958;
  assign n9960 = pi19 ? n594 : n2614;
  assign n9961 = pi18 ? n32 : n9960;
  assign n9962 = pi17 ? n2954 : ~n9961;
  assign n9963 = pi16 ? n32 : n9962;
  assign n9964 = pi17 ? n2954 : ~n2623;
  assign n9965 = pi16 ? n32 : n9964;
  assign n9966 = pi15 ? n9963 : n9965;
  assign n9967 = pi14 ? n9959 : n9966;
  assign n9968 = pi13 ? n9956 : n9967;
  assign n9969 = pi17 ? n2954 : ~n2618;
  assign n9970 = pi16 ? n32 : n9969;
  assign n9971 = pi17 ? n2954 : ~n3621;
  assign n9972 = pi16 ? n32 : n9971;
  assign n9973 = pi15 ? n9970 : n9972;
  assign n9974 = pi18 ? n6071 : n595;
  assign n9975 = pi17 ? n3569 : ~n9974;
  assign n9976 = pi16 ? n32 : n9975;
  assign n9977 = pi17 ? n3569 : ~n3621;
  assign n9978 = pi16 ? n32 : n9977;
  assign n9979 = pi15 ? n9976 : n9978;
  assign n9980 = pi14 ? n9973 : n9979;
  assign n9981 = pi17 ? n32 : ~n2628;
  assign n9982 = pi16 ? n32 : n9981;
  assign n9983 = pi17 ? n32 : ~n2748;
  assign n9984 = pi16 ? n32 : n9983;
  assign n9985 = pi15 ? n9982 : n9984;
  assign n9986 = pi17 ? n32 : ~n2519;
  assign n9987 = pi16 ? n32 : n9986;
  assign n9988 = pi14 ? n9985 : n9987;
  assign n9989 = pi13 ? n9980 : n9988;
  assign n9990 = pi12 ? n9968 : n9989;
  assign n9991 = pi11 ? n9943 : n9990;
  assign n9992 = pi10 ? n9882 : n9991;
  assign n9993 = pi09 ? n9734 : n9992;
  assign n9994 = pi08 ? n9716 : n9993;
  assign n9995 = pi07 ? n9443 : n9994;
  assign n9996 = pi06 ? n8922 : n9995;
  assign n9997 = pi05 ? n8147 : n9996;
  assign n9998 = pi18 ? n962 : ~n880;
  assign n9999 = pi17 ? n32 : n9998;
  assign n10000 = pi16 ? n32 : n9999;
  assign n10001 = pi15 ? n32 : n10000;
  assign n10002 = pi18 ? n2730 : ~n940;
  assign n10003 = pi17 ? n32 : n10002;
  assign n10004 = pi16 ? n32 : n10003;
  assign n10005 = pi18 ? n702 : ~n940;
  assign n10006 = pi17 ? n32 : n10005;
  assign n10007 = pi16 ? n32 : n10006;
  assign n10008 = pi15 ? n10004 : n10007;
  assign n10009 = pi14 ? n10001 : n10008;
  assign n10010 = pi13 ? n32 : n10009;
  assign n10011 = pi12 ? n32 : n10010;
  assign n10012 = pi11 ? n32 : n10011;
  assign n10013 = pi10 ? n32 : n10012;
  assign n10014 = pi18 ? n4098 : ~n940;
  assign n10015 = pi17 ? n32 : n10014;
  assign n10016 = pi16 ? n32 : n10015;
  assign n10017 = pi18 ? n595 : ~n940;
  assign n10018 = pi17 ? n32 : n10017;
  assign n10019 = pi16 ? n32 : n10018;
  assign n10020 = pi15 ? n10016 : n10019;
  assign n10021 = pi18 ? n595 : ~n880;
  assign n10022 = pi17 ? n32 : n10021;
  assign n10023 = pi16 ? n32 : n10022;
  assign n10024 = pi18 ? n2627 : ~n880;
  assign n10025 = pi17 ? n32 : n10024;
  assign n10026 = pi16 ? n32 : n10025;
  assign n10027 = pi15 ? n10023 : n10026;
  assign n10028 = pi14 ? n10020 : n10027;
  assign n10029 = pi18 ? n508 : ~n880;
  assign n10030 = pi17 ? n32 : n10029;
  assign n10031 = pi16 ? n32 : n10030;
  assign n10032 = pi18 ? n2424 : ~n880;
  assign n10033 = pi17 ? n32 : n10032;
  assign n10034 = pi16 ? n32 : n10033;
  assign n10035 = pi18 ? n418 : ~n880;
  assign n10036 = pi17 ? n32 : n10035;
  assign n10037 = pi16 ? n32 : n10036;
  assign n10038 = pi15 ? n10034 : n10037;
  assign n10039 = pi14 ? n10031 : n10038;
  assign n10040 = pi13 ? n10028 : n10039;
  assign n10041 = pi18 ? n3786 : ~n940;
  assign n10042 = pi17 ? n32 : n10041;
  assign n10043 = pi16 ? n32 : n10042;
  assign n10044 = pi14 ? n10037 : n10043;
  assign n10045 = pi18 ? n532 : ~n880;
  assign n10046 = pi17 ? n32 : n10045;
  assign n10047 = pi16 ? n32 : n10046;
  assign n10048 = pi18 ? n2298 : ~n880;
  assign n10049 = pi17 ? n32 : n10048;
  assign n10050 = pi16 ? n32 : n10049;
  assign n10051 = pi15 ? n10047 : n10050;
  assign n10052 = pi20 ? n32 : ~n111;
  assign n10053 = pi19 ? n32 : n10052;
  assign n10054 = pi18 ? n430 : ~n10053;
  assign n10055 = pi17 ? n32 : n10054;
  assign n10056 = pi16 ? n32 : n10055;
  assign n10057 = pi20 ? n342 : ~n111;
  assign n10058 = pi19 ? n32 : n10057;
  assign n10059 = pi18 ? n430 : ~n10058;
  assign n10060 = pi17 ? n32 : n10059;
  assign n10061 = pi16 ? n32 : n10060;
  assign n10062 = pi15 ? n10056 : n10061;
  assign n10063 = pi14 ? n10051 : n10062;
  assign n10064 = pi13 ? n10044 : n10063;
  assign n10065 = pi12 ? n10040 : n10064;
  assign n10066 = pi21 ? n1009 : n206;
  assign n10067 = pi20 ? n342 : n10066;
  assign n10068 = pi19 ? n32 : n10067;
  assign n10069 = pi18 ? n430 : ~n10068;
  assign n10070 = pi17 ? n32 : n10069;
  assign n10071 = pi16 ? n32 : n10070;
  assign n10072 = pi20 ? n342 : n141;
  assign n10073 = pi19 ? n32 : n10072;
  assign n10074 = pi18 ? n2304 : ~n10073;
  assign n10075 = pi17 ? n32 : n10074;
  assign n10076 = pi16 ? n32 : n10075;
  assign n10077 = pi15 ? n10071 : n10076;
  assign n10078 = pi19 ? n32 : n342;
  assign n10079 = pi18 ? n2304 : ~n10078;
  assign n10080 = pi17 ? n32 : n10079;
  assign n10081 = pi16 ? n32 : n10080;
  assign n10082 = pi18 ? n344 : ~n684;
  assign n10083 = pi17 ? n32 : n10082;
  assign n10084 = pi16 ? n32 : n10083;
  assign n10085 = pi15 ? n10081 : n10084;
  assign n10086 = pi14 ? n10077 : n10085;
  assign n10087 = pi18 ? n350 : ~n684;
  assign n10088 = pi17 ? n32 : n10087;
  assign n10089 = pi16 ? n32 : n10088;
  assign n10090 = pi18 ? n1813 : ~n684;
  assign n10091 = pi17 ? n32 : n10090;
  assign n10092 = pi16 ? n32 : n10091;
  assign n10093 = pi15 ? n10089 : n10092;
  assign n10094 = pi20 ? n175 : ~n1817;
  assign n10095 = pi19 ? n32 : n10094;
  assign n10096 = pi18 ? n1813 : ~n10095;
  assign n10097 = pi17 ? n32 : n10096;
  assign n10098 = pi16 ? n32 : n10097;
  assign n10099 = pi18 ? n1813 : ~n2043;
  assign n10100 = pi17 ? n32 : n10099;
  assign n10101 = pi16 ? n32 : n10100;
  assign n10102 = pi15 ? n10098 : n10101;
  assign n10103 = pi14 ? n10093 : n10102;
  assign n10104 = pi13 ? n10086 : n10103;
  assign n10105 = pi18 ? n814 : ~n9847;
  assign n10106 = pi17 ? n32 : n10105;
  assign n10107 = pi16 ? n32 : n10106;
  assign n10108 = pi18 ? n814 : ~n7038;
  assign n10109 = pi17 ? n32 : n10108;
  assign n10110 = pi16 ? n32 : n10109;
  assign n10111 = pi15 ? n10107 : n10110;
  assign n10112 = pi18 ? n814 : ~n1965;
  assign n10113 = pi17 ? n32 : n10112;
  assign n10114 = pi16 ? n32 : n10113;
  assign n10115 = pi18 ? n814 : ~n880;
  assign n10116 = pi17 ? n32 : n10115;
  assign n10117 = pi16 ? n32 : n10116;
  assign n10118 = pi15 ? n10114 : n10117;
  assign n10119 = pi14 ? n10111 : n10118;
  assign n10120 = pi20 ? n1324 : n749;
  assign n10121 = pi19 ? n32 : n10120;
  assign n10122 = pi18 ? n237 : ~n10121;
  assign n10123 = pi17 ? n32 : n10122;
  assign n10124 = pi16 ? n32 : n10123;
  assign n10125 = pi20 ? n428 : ~n52;
  assign n10126 = pi19 ? n32 : n10125;
  assign n10127 = pi18 ? n237 : ~n10126;
  assign n10128 = pi17 ? n32 : n10127;
  assign n10129 = pi16 ? n32 : n10128;
  assign n10130 = pi15 ? n10124 : n10129;
  assign n10131 = pi18 ? n237 : ~n7824;
  assign n10132 = pi17 ? n32 : n10131;
  assign n10133 = pi16 ? n32 : n10132;
  assign n10134 = pi18 ? n237 : ~n1970;
  assign n10135 = pi17 ? n32 : n10134;
  assign n10136 = pi16 ? n32 : n10135;
  assign n10137 = pi15 ? n10133 : n10136;
  assign n10138 = pi14 ? n10130 : n10137;
  assign n10139 = pi13 ? n10119 : n10138;
  assign n10140 = pi12 ? n10104 : n10139;
  assign n10141 = pi11 ? n10065 : n10140;
  assign n10142 = pi18 ? n237 : ~n684;
  assign n10143 = pi17 ? n32 : n10142;
  assign n10144 = pi16 ? n32 : n10143;
  assign n10145 = pi18 ? n237 : ~n245;
  assign n10146 = pi17 ? n32 : n10145;
  assign n10147 = pi16 ? n32 : n10146;
  assign n10148 = pi20 ? n9628 : n339;
  assign n10149 = pi19 ? n32 : n10148;
  assign n10150 = pi18 ? n618 : ~n10149;
  assign n10151 = pi17 ? n32 : n10150;
  assign n10152 = pi16 ? n32 : n10151;
  assign n10153 = pi15 ? n10147 : n10152;
  assign n10154 = pi14 ? n10144 : n10153;
  assign n10155 = pi18 ? n618 : ~n366;
  assign n10156 = pi17 ? n32 : n10155;
  assign n10157 = pi16 ? n32 : n10156;
  assign n10158 = pi20 ? n1331 : n141;
  assign n10159 = pi19 ? n32 : n10158;
  assign n10160 = pi18 ? n618 : ~n10159;
  assign n10161 = pi17 ? n32 : n10160;
  assign n10162 = pi16 ? n32 : n10161;
  assign n10163 = pi15 ? n10157 : n10162;
  assign n10164 = pi18 ? n618 : ~n9630;
  assign n10165 = pi17 ? n32 : n10164;
  assign n10166 = pi16 ? n32 : n10165;
  assign n10167 = pi21 ? n2076 : n405;
  assign n10168 = pi20 ? n10167 : ~n32;
  assign n10169 = pi19 ? n267 : n10168;
  assign n10170 = pi18 ? n618 : ~n10169;
  assign n10171 = pi17 ? n32 : n10170;
  assign n10172 = pi16 ? n32 : n10171;
  assign n10173 = pi15 ? n10166 : n10172;
  assign n10174 = pi14 ? n10163 : n10173;
  assign n10175 = pi13 ? n10154 : n10174;
  assign n10176 = pi20 ? n141 : ~n246;
  assign n10177 = pi19 ? n10176 : ~n32;
  assign n10178 = pi19 ? n267 : n8277;
  assign n10179 = pi18 ? n10177 : ~n10178;
  assign n10180 = pi17 ? n32 : n10179;
  assign n10181 = pi16 ? n32 : n10180;
  assign n10182 = pi22 ? n65 : n173;
  assign n10183 = pi21 ? n32 : n10182;
  assign n10184 = pi20 ? n10183 : ~n32;
  assign n10185 = pi19 ? n32 : n10184;
  assign n10186 = pi18 ? n1676 : ~n10185;
  assign n10187 = pi17 ? n32 : n10186;
  assign n10188 = pi16 ? n32 : n10187;
  assign n10189 = pi15 ? n10181 : n10188;
  assign n10190 = pi17 ? n3155 : ~n8639;
  assign n10191 = pi16 ? n32 : n10190;
  assign n10192 = pi14 ? n10189 : n10191;
  assign n10193 = pi19 ? n472 : n589;
  assign n10194 = pi18 ? n32 : n10193;
  assign n10195 = pi17 ? n32 : ~n10194;
  assign n10196 = pi16 ? n32 : n10195;
  assign n10197 = pi15 ? n8167 : n10196;
  assign n10198 = pi17 ? n32 : ~n2850;
  assign n10199 = pi16 ? n32 : n10198;
  assign n10200 = pi17 ? n3569 : ~n9937;
  assign n10201 = pi16 ? n32 : n10200;
  assign n10202 = pi15 ? n10199 : n10201;
  assign n10203 = pi14 ? n10197 : n10202;
  assign n10204 = pi13 ? n10192 : n10203;
  assign n10205 = pi12 ? n10175 : n10204;
  assign n10206 = pi19 ? n1320 : n1812;
  assign n10207 = pi18 ? n32 : n10206;
  assign n10208 = pi17 ? n3569 : ~n10207;
  assign n10209 = pi16 ? n32 : n10208;
  assign n10210 = pi19 ? n1818 : n1812;
  assign n10211 = pi18 ? n32 : n10210;
  assign n10212 = pi17 ? n3569 : ~n10211;
  assign n10213 = pi16 ? n32 : n10212;
  assign n10214 = pi15 ? n10209 : n10213;
  assign n10215 = pi17 ? n3569 : ~n2736;
  assign n10216 = pi16 ? n32 : n10215;
  assign n10217 = pi17 ? n32 : ~n2736;
  assign n10218 = pi16 ? n32 : n10217;
  assign n10219 = pi15 ? n10216 : n10218;
  assign n10220 = pi14 ? n10214 : n10219;
  assign n10221 = pi17 ? n32 : ~n2616;
  assign n10222 = pi16 ? n32 : n10221;
  assign n10223 = pi15 ? n10218 : n10222;
  assign n10224 = pi18 ? n3350 : ~n2622;
  assign n10225 = pi17 ? n32 : n10224;
  assign n10226 = pi16 ? n32 : n10225;
  assign n10227 = pi18 ? n3350 : ~n595;
  assign n10228 = pi17 ? n32 : n10227;
  assign n10229 = pi16 ? n32 : n10228;
  assign n10230 = pi15 ? n10226 : n10229;
  assign n10231 = pi14 ? n10223 : n10230;
  assign n10232 = pi13 ? n10220 : n10231;
  assign n10233 = pi18 ? n3350 : ~n4098;
  assign n10234 = pi17 ? n32 : n10233;
  assign n10235 = pi16 ? n32 : n10234;
  assign n10236 = pi15 ? n10235 : n10229;
  assign n10237 = pi18 ? n237 : ~n595;
  assign n10238 = pi17 ? n32 : n10237;
  assign n10239 = pi16 ? n32 : n10238;
  assign n10240 = pi18 ? n237 : ~n508;
  assign n10241 = pi17 ? n32 : n10240;
  assign n10242 = pi16 ? n32 : n10241;
  assign n10243 = pi15 ? n10239 : n10242;
  assign n10244 = pi14 ? n10236 : n10243;
  assign n10245 = pi18 ? n237 : ~n323;
  assign n10246 = pi17 ? n32 : n10245;
  assign n10247 = pi16 ? n32 : n10246;
  assign n10248 = pi18 ? n1813 : ~n323;
  assign n10249 = pi17 ? n32 : n10248;
  assign n10250 = pi16 ? n32 : n10249;
  assign n10251 = pi15 ? n10247 : n10250;
  assign n10252 = pi14 ? n10251 : n10250;
  assign n10253 = pi13 ? n10244 : n10252;
  assign n10254 = pi12 ? n10232 : n10253;
  assign n10255 = pi11 ? n10205 : n10254;
  assign n10256 = pi10 ? n10141 : n10255;
  assign n10257 = pi09 ? n10013 : n10256;
  assign n10258 = pi18 ? n590 : ~n880;
  assign n10259 = pi17 ? n32 : n10258;
  assign n10260 = pi16 ? n32 : n10259;
  assign n10261 = pi15 ? n32 : n10260;
  assign n10262 = pi18 ? n2849 : ~n940;
  assign n10263 = pi17 ? n32 : n10262;
  assign n10264 = pi16 ? n32 : n10263;
  assign n10265 = pi18 ? n697 : ~n940;
  assign n10266 = pi17 ? n32 : n10265;
  assign n10267 = pi16 ? n32 : n10266;
  assign n10268 = pi15 ? n10264 : n10267;
  assign n10269 = pi14 ? n10261 : n10268;
  assign n10270 = pi13 ? n32 : n10269;
  assign n10271 = pi12 ? n32 : n10270;
  assign n10272 = pi11 ? n32 : n10271;
  assign n10273 = pi10 ? n32 : n10272;
  assign n10274 = pi18 ? n2615 : ~n940;
  assign n10275 = pi17 ? n32 : n10274;
  assign n10276 = pi16 ? n32 : n10275;
  assign n10277 = pi18 ? n1750 : ~n940;
  assign n10278 = pi17 ? n32 : n10277;
  assign n10279 = pi16 ? n32 : n10278;
  assign n10280 = pi15 ? n10276 : n10279;
  assign n10281 = pi18 ? n1750 : ~n880;
  assign n10282 = pi17 ? n32 : n10281;
  assign n10283 = pi16 ? n32 : n10282;
  assign n10284 = pi18 ? n2622 : ~n880;
  assign n10285 = pi17 ? n32 : n10284;
  assign n10286 = pi16 ? n32 : n10285;
  assign n10287 = pi15 ? n10283 : n10286;
  assign n10288 = pi14 ? n10280 : n10287;
  assign n10289 = pi18 ? n702 : ~n880;
  assign n10290 = pi17 ? n32 : n10289;
  assign n10291 = pi16 ? n32 : n10290;
  assign n10292 = pi15 ? n10286 : n10291;
  assign n10293 = pi18 ? n2291 : ~n880;
  assign n10294 = pi17 ? n32 : n10293;
  assign n10295 = pi16 ? n32 : n10294;
  assign n10296 = pi18 ? n797 : ~n880;
  assign n10297 = pi17 ? n32 : n10296;
  assign n10298 = pi16 ? n32 : n10297;
  assign n10299 = pi15 ? n10295 : n10298;
  assign n10300 = pi14 ? n10292 : n10299;
  assign n10301 = pi13 ? n10288 : n10300;
  assign n10302 = pi18 ? n2413 : ~n940;
  assign n10303 = pi17 ? n32 : n10302;
  assign n10304 = pi16 ? n32 : n10303;
  assign n10305 = pi14 ? n10298 : n10304;
  assign n10306 = pi18 ? n2413 : ~n880;
  assign n10307 = pi17 ? n32 : n10306;
  assign n10308 = pi16 ? n32 : n10307;
  assign n10309 = pi15 ? n10308 : n10034;
  assign n10310 = pi18 ? n418 : ~n10053;
  assign n10311 = pi17 ? n32 : n10310;
  assign n10312 = pi16 ? n32 : n10311;
  assign n10313 = pi18 ? n418 : ~n10073;
  assign n10314 = pi17 ? n32 : n10313;
  assign n10315 = pi16 ? n32 : n10314;
  assign n10316 = pi15 ? n10312 : n10315;
  assign n10317 = pi14 ? n10309 : n10316;
  assign n10318 = pi13 ? n10305 : n10317;
  assign n10319 = pi12 ? n10301 : n10318;
  assign n10320 = pi18 ? n418 : ~n10068;
  assign n10321 = pi17 ? n32 : n10320;
  assign n10322 = pi16 ? n32 : n10321;
  assign n10323 = pi18 ? n3786 : ~n10073;
  assign n10324 = pi17 ? n32 : n10323;
  assign n10325 = pi16 ? n32 : n10324;
  assign n10326 = pi15 ? n10322 : n10325;
  assign n10327 = pi20 ? n342 : ~n726;
  assign n10328 = pi19 ? n32 : n10327;
  assign n10329 = pi18 ? n3786 : ~n10328;
  assign n10330 = pi17 ? n32 : n10329;
  assign n10331 = pi16 ? n32 : n10330;
  assign n10332 = pi18 ? n532 : ~n684;
  assign n10333 = pi17 ? n32 : n10332;
  assign n10334 = pi16 ? n32 : n10333;
  assign n10335 = pi15 ? n10331 : n10334;
  assign n10336 = pi14 ? n10326 : n10335;
  assign n10337 = pi18 ? n2298 : ~n684;
  assign n10338 = pi17 ? n32 : n10337;
  assign n10339 = pi16 ? n32 : n10338;
  assign n10340 = pi15 ? n10334 : n10339;
  assign n10341 = pi18 ? n2298 : ~n10095;
  assign n10342 = pi17 ? n32 : n10341;
  assign n10343 = pi16 ? n32 : n10342;
  assign n10344 = pi18 ? n2298 : ~n2043;
  assign n10345 = pi17 ? n32 : n10344;
  assign n10346 = pi16 ? n32 : n10345;
  assign n10347 = pi15 ? n10343 : n10346;
  assign n10348 = pi14 ? n10340 : n10347;
  assign n10349 = pi13 ? n10336 : n10348;
  assign n10350 = pi18 ? n430 : ~n9847;
  assign n10351 = pi17 ? n32 : n10350;
  assign n10352 = pi16 ? n32 : n10351;
  assign n10353 = pi18 ? n430 : ~n7038;
  assign n10354 = pi17 ? n32 : n10353;
  assign n10355 = pi16 ? n32 : n10354;
  assign n10356 = pi15 ? n10352 : n10355;
  assign n10357 = pi18 ? n2304 : ~n1965;
  assign n10358 = pi17 ? n32 : n10357;
  assign n10359 = pi16 ? n32 : n10358;
  assign n10360 = pi18 ? n3336 : ~n880;
  assign n10361 = pi17 ? n32 : n10360;
  assign n10362 = pi16 ? n32 : n10361;
  assign n10363 = pi15 ? n10359 : n10362;
  assign n10364 = pi14 ? n10356 : n10363;
  assign n10365 = pi18 ? n350 : ~n10121;
  assign n10366 = pi17 ? n32 : n10365;
  assign n10367 = pi16 ? n32 : n10366;
  assign n10368 = pi18 ? n350 : ~n1965;
  assign n10369 = pi17 ? n32 : n10368;
  assign n10370 = pi16 ? n32 : n10369;
  assign n10371 = pi15 ? n10367 : n10370;
  assign n10372 = pi18 ? n350 : ~n7824;
  assign n10373 = pi17 ? n32 : n10372;
  assign n10374 = pi16 ? n32 : n10373;
  assign n10375 = pi18 ? n350 : ~n341;
  assign n10376 = pi17 ? n32 : n10375;
  assign n10377 = pi16 ? n32 : n10376;
  assign n10378 = pi15 ? n10374 : n10377;
  assign n10379 = pi14 ? n10371 : n10378;
  assign n10380 = pi13 ? n10364 : n10379;
  assign n10381 = pi12 ? n10349 : n10380;
  assign n10382 = pi11 ? n10319 : n10381;
  assign n10383 = pi18 ? n350 : ~n245;
  assign n10384 = pi17 ? n32 : n10383;
  assign n10385 = pi16 ? n32 : n10384;
  assign n10386 = pi18 ? n814 : ~n3780;
  assign n10387 = pi17 ? n32 : n10386;
  assign n10388 = pi16 ? n32 : n10387;
  assign n10389 = pi15 ? n10385 : n10388;
  assign n10390 = pi14 ? n10089 : n10389;
  assign n10391 = pi18 ? n814 : ~n366;
  assign n10392 = pi17 ? n32 : n10391;
  assign n10393 = pi16 ? n32 : n10392;
  assign n10394 = pi20 ? n405 : ~n32;
  assign n10395 = pi19 ? n32 : n10394;
  assign n10396 = pi18 ? n814 : ~n10395;
  assign n10397 = pi17 ? n32 : n10396;
  assign n10398 = pi16 ? n32 : n10397;
  assign n10399 = pi15 ? n10393 : n10398;
  assign n10400 = pi18 ? n814 : ~n684;
  assign n10401 = pi17 ? n32 : n10400;
  assign n10402 = pi16 ? n32 : n10401;
  assign n10403 = pi19 ? n267 : n429;
  assign n10404 = pi18 ? n814 : ~n10403;
  assign n10405 = pi17 ? n32 : n10404;
  assign n10406 = pi16 ? n32 : n10405;
  assign n10407 = pi15 ? n10402 : n10406;
  assign n10408 = pi14 ? n10399 : n10407;
  assign n10409 = pi13 ? n10390 : n10408;
  assign n10410 = pi20 ? n1940 : ~n246;
  assign n10411 = pi19 ? n10410 : ~n32;
  assign n10412 = pi18 ? n10411 : ~n10178;
  assign n10413 = pi17 ? n32 : n10412;
  assign n10414 = pi16 ? n32 : n10413;
  assign n10415 = pi18 ? n814 : ~n8632;
  assign n10416 = pi17 ? n32 : n10415;
  assign n10417 = pi16 ? n32 : n10416;
  assign n10418 = pi15 ? n10414 : n10417;
  assign n10419 = pi18 ? n1676 : ~n1156;
  assign n10420 = pi17 ? n32 : n10419;
  assign n10421 = pi16 ? n32 : n10420;
  assign n10422 = pi18 ? n237 : ~n496;
  assign n10423 = pi17 ? n32 : n10422;
  assign n10424 = pi16 ? n32 : n10423;
  assign n10425 = pi15 ? n10421 : n10424;
  assign n10426 = pi14 ? n10418 : n10425;
  assign n10427 = pi18 ? n1942 : ~n590;
  assign n10428 = pi17 ? n32 : n10427;
  assign n10429 = pi16 ? n32 : n10428;
  assign n10430 = pi15 ? n8745 : n10429;
  assign n10431 = pi18 ? n1942 : ~n2849;
  assign n10432 = pi17 ? n32 : n10431;
  assign n10433 = pi16 ? n32 : n10432;
  assign n10434 = pi18 ? n237 : ~n7029;
  assign n10435 = pi17 ? n32 : n10434;
  assign n10436 = pi16 ? n32 : n10435;
  assign n10437 = pi15 ? n10433 : n10436;
  assign n10438 = pi14 ? n10430 : n10437;
  assign n10439 = pi13 ? n10426 : n10438;
  assign n10440 = pi12 ? n10409 : n10439;
  assign n10441 = pi19 ? n507 : n1812;
  assign n10442 = pi18 ? n237 : ~n10441;
  assign n10443 = pi17 ? n32 : n10442;
  assign n10444 = pi16 ? n32 : n10443;
  assign n10445 = pi22 ? n173 : n50;
  assign n10446 = pi21 ? n10445 : ~n32;
  assign n10447 = pi20 ? n10446 : ~n32;
  assign n10448 = pi19 ? n1464 : n10447;
  assign n10449 = pi18 ? n237 : ~n10448;
  assign n10450 = pi17 ? n32 : n10449;
  assign n10451 = pi16 ? n32 : n10450;
  assign n10452 = pi15 ? n10444 : n10451;
  assign n10453 = pi18 ? n237 : ~n697;
  assign n10454 = pi17 ? n32 : n10453;
  assign n10455 = pi16 ? n32 : n10454;
  assign n10456 = pi14 ? n10452 : n10455;
  assign n10457 = pi18 ? n1813 : ~n697;
  assign n10458 = pi17 ? n32 : n10457;
  assign n10459 = pi16 ? n32 : n10458;
  assign n10460 = pi18 ? n350 : ~n2615;
  assign n10461 = pi17 ? n32 : n10460;
  assign n10462 = pi16 ? n32 : n10461;
  assign n10463 = pi15 ? n10459 : n10462;
  assign n10464 = pi18 ? n350 : ~n2622;
  assign n10465 = pi17 ? n32 : n10464;
  assign n10466 = pi16 ? n32 : n10465;
  assign n10467 = pi18 ? n350 : ~n595;
  assign n10468 = pi17 ? n32 : n10467;
  assign n10469 = pi16 ? n32 : n10468;
  assign n10470 = pi15 ? n10466 : n10469;
  assign n10471 = pi14 ? n10463 : n10470;
  assign n10472 = pi13 ? n10456 : n10471;
  assign n10473 = pi18 ? n350 : ~n4098;
  assign n10474 = pi17 ? n32 : n10473;
  assign n10475 = pi16 ? n32 : n10474;
  assign n10476 = pi15 ? n10475 : n10469;
  assign n10477 = pi18 ? n2318 : ~n508;
  assign n10478 = pi17 ? n32 : n10477;
  assign n10479 = pi16 ? n32 : n10478;
  assign n10480 = pi15 ? n10469 : n10479;
  assign n10481 = pi14 ? n10476 : n10480;
  assign n10482 = pi18 ? n344 : ~n323;
  assign n10483 = pi17 ? n32 : n10482;
  assign n10484 = pi16 ? n32 : n10483;
  assign n10485 = pi20 ? n428 : n321;
  assign n10486 = pi19 ? n10485 : ~n32;
  assign n10487 = pi18 ? n2318 : ~n10486;
  assign n10488 = pi17 ? n32 : n10487;
  assign n10489 = pi16 ? n32 : n10488;
  assign n10490 = pi15 ? n10484 : n10489;
  assign n10491 = pi14 ? n10484 : n10490;
  assign n10492 = pi13 ? n10481 : n10491;
  assign n10493 = pi12 ? n10472 : n10492;
  assign n10494 = pi11 ? n10440 : n10493;
  assign n10495 = pi10 ? n10382 : n10494;
  assign n10496 = pi09 ? n10273 : n10495;
  assign n10497 = pi08 ? n10257 : n10496;
  assign n10498 = pi16 ? n32 : n882;
  assign n10499 = pi15 ? n32 : n10498;
  assign n10500 = pi18 ? n2830 : ~n940;
  assign n10501 = pi17 ? n32 : n10500;
  assign n10502 = pi16 ? n32 : n10501;
  assign n10503 = pi18 ? n496 : ~n940;
  assign n10504 = pi17 ? n32 : n10503;
  assign n10505 = pi16 ? n32 : n10504;
  assign n10506 = pi15 ? n10502 : n10505;
  assign n10507 = pi14 ? n10499 : n10506;
  assign n10508 = pi13 ? n32 : n10507;
  assign n10509 = pi12 ? n32 : n10508;
  assign n10510 = pi11 ? n32 : n10509;
  assign n10511 = pi10 ? n32 : n10510;
  assign n10512 = pi18 ? n4244 : ~n940;
  assign n10513 = pi17 ? n32 : n10512;
  assign n10514 = pi16 ? n32 : n10513;
  assign n10515 = pi18 ? n962 : ~n940;
  assign n10516 = pi17 ? n32 : n10515;
  assign n10517 = pi16 ? n32 : n10516;
  assign n10518 = pi15 ? n10514 : n10517;
  assign n10519 = pi18 ? n2730 : ~n880;
  assign n10520 = pi17 ? n32 : n10519;
  assign n10521 = pi16 ? n32 : n10520;
  assign n10522 = pi15 ? n10000 : n10521;
  assign n10523 = pi14 ? n10518 : n10522;
  assign n10524 = pi18 ? n697 : ~n880;
  assign n10525 = pi17 ? n32 : n10524;
  assign n10526 = pi16 ? n32 : n10525;
  assign n10527 = pi15 ? n10521 : n10526;
  assign n10528 = pi18 ? n4098 : ~n880;
  assign n10529 = pi17 ? n32 : n10528;
  assign n10530 = pi16 ? n32 : n10529;
  assign n10531 = pi15 ? n10530 : n10023;
  assign n10532 = pi14 ? n10527 : n10531;
  assign n10533 = pi13 ? n10523 : n10532;
  assign n10534 = pi18 ? n2627 : ~n940;
  assign n10535 = pi17 ? n32 : n10534;
  assign n10536 = pi16 ? n32 : n10535;
  assign n10537 = pi18 ? n508 : ~n940;
  assign n10538 = pi17 ? n32 : n10537;
  assign n10539 = pi16 ? n32 : n10538;
  assign n10540 = pi15 ? n10536 : n10539;
  assign n10541 = pi14 ? n10023 : n10540;
  assign n10542 = pi15 ? n10031 : n10295;
  assign n10543 = pi18 ? n797 : ~n10053;
  assign n10544 = pi17 ? n32 : n10543;
  assign n10545 = pi16 ? n32 : n10544;
  assign n10546 = pi18 ? n797 : ~n10073;
  assign n10547 = pi17 ? n32 : n10546;
  assign n10548 = pi16 ? n32 : n10547;
  assign n10549 = pi15 ? n10545 : n10548;
  assign n10550 = pi14 ? n10542 : n10549;
  assign n10551 = pi13 ? n10541 : n10550;
  assign n10552 = pi12 ? n10533 : n10551;
  assign n10553 = pi18 ? n797 : ~n10078;
  assign n10554 = pi17 ? n32 : n10553;
  assign n10555 = pi16 ? n32 : n10554;
  assign n10556 = pi18 ? n2413 : ~n10073;
  assign n10557 = pi17 ? n32 : n10556;
  assign n10558 = pi16 ? n32 : n10557;
  assign n10559 = pi15 ? n10555 : n10558;
  assign n10560 = pi18 ? n2413 : ~n10328;
  assign n10561 = pi17 ? n32 : n10560;
  assign n10562 = pi16 ? n32 : n10561;
  assign n10563 = pi18 ? n2413 : ~n684;
  assign n10564 = pi17 ? n32 : n10563;
  assign n10565 = pi16 ? n32 : n10564;
  assign n10566 = pi15 ? n10562 : n10565;
  assign n10567 = pi14 ? n10559 : n10566;
  assign n10568 = pi20 ? n342 : ~n1817;
  assign n10569 = pi19 ? n32 : n10568;
  assign n10570 = pi18 ? n605 : ~n10569;
  assign n10571 = pi17 ? n32 : n10570;
  assign n10572 = pi16 ? n32 : n10571;
  assign n10573 = pi18 ? n2424 : ~n2043;
  assign n10574 = pi17 ? n32 : n10573;
  assign n10575 = pi16 ? n32 : n10574;
  assign n10576 = pi15 ? n10572 : n10575;
  assign n10577 = pi18 ? n2424 : ~n10569;
  assign n10578 = pi17 ? n32 : n10577;
  assign n10579 = pi16 ? n32 : n10578;
  assign n10580 = pi18 ? n2424 : ~n684;
  assign n10581 = pi17 ? n32 : n10580;
  assign n10582 = pi16 ? n32 : n10581;
  assign n10583 = pi15 ? n10579 : n10582;
  assign n10584 = pi14 ? n10576 : n10583;
  assign n10585 = pi13 ? n10567 : n10584;
  assign n10586 = pi18 ? n418 : ~n8213;
  assign n10587 = pi17 ? n32 : n10586;
  assign n10588 = pi16 ? n32 : n10587;
  assign n10589 = pi18 ? n418 : ~n496;
  assign n10590 = pi17 ? n32 : n10589;
  assign n10591 = pi16 ? n32 : n10590;
  assign n10592 = pi15 ? n10588 : n10591;
  assign n10593 = pi20 ? n342 : ~n6229;
  assign n10594 = pi19 ? n32 : n10593;
  assign n10595 = pi18 ? n3786 : ~n10594;
  assign n10596 = pi17 ? n32 : n10595;
  assign n10597 = pi16 ? n32 : n10596;
  assign n10598 = pi18 ? n3786 : ~n684;
  assign n10599 = pi17 ? n32 : n10598;
  assign n10600 = pi16 ? n32 : n10599;
  assign n10601 = pi15 ? n10597 : n10600;
  assign n10602 = pi14 ? n10592 : n10601;
  assign n10603 = pi18 ? n532 : ~n9598;
  assign n10604 = pi17 ? n32 : n10603;
  assign n10605 = pi16 ? n32 : n10604;
  assign n10606 = pi15 ? n10605 : n10334;
  assign n10607 = pi18 ? n532 : ~n8804;
  assign n10608 = pi17 ? n32 : n10607;
  assign n10609 = pi16 ? n32 : n10608;
  assign n10610 = pi15 ? n10609 : n10334;
  assign n10611 = pi14 ? n10606 : n10610;
  assign n10612 = pi13 ? n10602 : n10611;
  assign n10613 = pi12 ? n10585 : n10612;
  assign n10614 = pi11 ? n10552 : n10613;
  assign n10615 = pi20 ? n342 : n243;
  assign n10616 = pi19 ? n32 : n10615;
  assign n10617 = pi18 ? n532 : ~n10616;
  assign n10618 = pi17 ? n32 : n10617;
  assign n10619 = pi16 ? n32 : n10618;
  assign n10620 = pi15 ? n10619 : n10339;
  assign n10621 = pi18 ? n2318 : ~n245;
  assign n10622 = pi17 ? n32 : n10621;
  assign n10623 = pi16 ? n32 : n10622;
  assign n10624 = pi18 ? n1548 : ~n684;
  assign n10625 = pi17 ? n32 : n10624;
  assign n10626 = pi16 ? n32 : n10625;
  assign n10627 = pi15 ? n10623 : n10626;
  assign n10628 = pi14 ? n10620 : n10627;
  assign n10629 = pi18 ? n1548 : ~n366;
  assign n10630 = pi17 ? n32 : n10629;
  assign n10631 = pi16 ? n32 : n10630;
  assign n10632 = pi20 ? n260 : n32;
  assign n10633 = pi19 ? n32 : ~n10632;
  assign n10634 = pi18 ? n1548 : ~n10633;
  assign n10635 = pi17 ? n32 : n10634;
  assign n10636 = pi16 ? n32 : n10635;
  assign n10637 = pi15 ? n10631 : n10636;
  assign n10638 = pi18 ? n1548 : ~n1965;
  assign n10639 = pi17 ? n32 : n10638;
  assign n10640 = pi16 ? n32 : n10639;
  assign n10641 = pi15 ? n10640 : n10636;
  assign n10642 = pi14 ? n10637 : n10641;
  assign n10643 = pi13 ? n10628 : n10642;
  assign n10644 = pi21 ? n206 : ~n405;
  assign n10645 = pi20 ? n10644 : n32;
  assign n10646 = pi19 ? n32 : ~n10645;
  assign n10647 = pi18 ? n1548 : ~n10646;
  assign n10648 = pi17 ? n32 : n10647;
  assign n10649 = pi16 ? n32 : n10648;
  assign n10650 = pi18 ? n6047 : ~n684;
  assign n10651 = pi17 ? n32 : n10650;
  assign n10652 = pi16 ? n32 : n10651;
  assign n10653 = pi15 ? n10649 : n10652;
  assign n10654 = pi18 ? n3336 : ~n1156;
  assign n10655 = pi17 ? n32 : n10654;
  assign n10656 = pi16 ? n32 : n10655;
  assign n10657 = pi18 ? n3336 : ~n590;
  assign n10658 = pi17 ? n32 : n10657;
  assign n10659 = pi16 ? n32 : n10658;
  assign n10660 = pi15 ? n10656 : n10659;
  assign n10661 = pi14 ? n10653 : n10660;
  assign n10662 = pi20 ? n623 : n32;
  assign n10663 = pi19 ? n32 : ~n10662;
  assign n10664 = pi18 ? n3336 : ~n10663;
  assign n10665 = pi17 ? n32 : n10664;
  assign n10666 = pi16 ? n32 : n10665;
  assign n10667 = pi18 ? n3336 : ~n2849;
  assign n10668 = pi17 ? n32 : n10667;
  assign n10669 = pi16 ? n32 : n10668;
  assign n10670 = pi19 ? n507 : ~n7488;
  assign n10671 = pi18 ? n350 : ~n10670;
  assign n10672 = pi17 ? n32 : n10671;
  assign n10673 = pi16 ? n32 : n10672;
  assign n10674 = pi15 ? n10669 : n10673;
  assign n10675 = pi14 ? n10666 : n10674;
  assign n10676 = pi13 ? n10661 : n10675;
  assign n10677 = pi12 ? n10643 : n10676;
  assign n10678 = pi18 ? n350 : ~n508;
  assign n10679 = pi17 ? n32 : n10678;
  assign n10680 = pi16 ? n32 : n10679;
  assign n10681 = pi18 ? n350 : ~n2730;
  assign n10682 = pi17 ? n32 : n10681;
  assign n10683 = pi16 ? n32 : n10682;
  assign n10684 = pi15 ? n10680 : n10683;
  assign n10685 = pi18 ? n2318 : ~n697;
  assign n10686 = pi17 ? n32 : n10685;
  assign n10687 = pi16 ? n32 : n10686;
  assign n10688 = pi18 ? n344 : ~n697;
  assign n10689 = pi17 ? n32 : n10688;
  assign n10690 = pi16 ? n32 : n10689;
  assign n10691 = pi15 ? n10687 : n10690;
  assign n10692 = pi14 ? n10684 : n10691;
  assign n10693 = pi18 ? n344 : ~n1750;
  assign n10694 = pi17 ? n32 : n10693;
  assign n10695 = pi16 ? n32 : n10694;
  assign n10696 = pi18 ? n344 : ~n595;
  assign n10697 = pi17 ? n32 : n10696;
  assign n10698 = pi16 ? n32 : n10697;
  assign n10699 = pi15 ? n10695 : n10698;
  assign n10700 = pi18 ? n344 : ~n508;
  assign n10701 = pi17 ? n32 : n10700;
  assign n10702 = pi16 ? n32 : n10701;
  assign n10703 = pi15 ? n10698 : n10702;
  assign n10704 = pi14 ? n10699 : n10703;
  assign n10705 = pi13 ? n10692 : n10704;
  assign n10706 = pi18 ? n344 : ~n4098;
  assign n10707 = pi17 ? n32 : n10706;
  assign n10708 = pi16 ? n32 : n10707;
  assign n10709 = pi15 ? n10708 : n10698;
  assign n10710 = pi19 ? n1612 : ~n32;
  assign n10711 = pi18 ? n2298 : ~n10710;
  assign n10712 = pi17 ? n32 : n10711;
  assign n10713 = pi16 ? n32 : n10712;
  assign n10714 = pi18 ? n532 : ~n2754;
  assign n10715 = pi17 ? n32 : n10714;
  assign n10716 = pi16 ? n32 : n10715;
  assign n10717 = pi15 ? n10713 : n10716;
  assign n10718 = pi14 ? n10709 : n10717;
  assign n10719 = pi18 ? n532 : ~n1405;
  assign n10720 = pi17 ? n32 : n10719;
  assign n10721 = pi16 ? n32 : n10720;
  assign n10722 = pi15 ? n10721 : n10716;
  assign n10723 = pi18 ? n532 : ~n323;
  assign n10724 = pi17 ? n32 : n10723;
  assign n10725 = pi16 ? n32 : n10724;
  assign n10726 = pi18 ? n532 : ~n797;
  assign n10727 = pi17 ? n32 : n10726;
  assign n10728 = pi16 ? n32 : n10727;
  assign n10729 = pi15 ? n10725 : n10728;
  assign n10730 = pi14 ? n10722 : n10729;
  assign n10731 = pi13 ? n10718 : n10730;
  assign n10732 = pi12 ? n10705 : n10731;
  assign n10733 = pi11 ? n10677 : n10732;
  assign n10734 = pi10 ? n10614 : n10733;
  assign n10735 = pi09 ? n10511 : n10734;
  assign n10736 = pi18 ? n751 : ~n880;
  assign n10737 = pi17 ? n32 : n10736;
  assign n10738 = pi16 ? n32 : n10737;
  assign n10739 = pi15 ? n32 : n10738;
  assign n10740 = pi18 ? n684 : ~n940;
  assign n10741 = pi17 ? n32 : n10740;
  assign n10742 = pi16 ? n32 : n10741;
  assign n10743 = pi15 ? n10502 : n10742;
  assign n10744 = pi14 ? n10739 : n10743;
  assign n10745 = pi13 ? n32 : n10744;
  assign n10746 = pi12 ? n32 : n10745;
  assign n10747 = pi11 ? n32 : n10746;
  assign n10748 = pi10 ? n32 : n10747;
  assign n10749 = pi18 ? n2835 : ~n940;
  assign n10750 = pi17 ? n32 : n10749;
  assign n10751 = pi16 ? n32 : n10750;
  assign n10752 = pi18 ? n590 : ~n940;
  assign n10753 = pi17 ? n32 : n10752;
  assign n10754 = pi16 ? n32 : n10753;
  assign n10755 = pi15 ? n10751 : n10754;
  assign n10756 = pi18 ? n2849 : ~n880;
  assign n10757 = pi17 ? n32 : n10756;
  assign n10758 = pi16 ? n32 : n10757;
  assign n10759 = pi15 ? n10260 : n10758;
  assign n10760 = pi14 ? n10755 : n10759;
  assign n10761 = pi18 ? n496 : ~n880;
  assign n10762 = pi17 ? n32 : n10761;
  assign n10763 = pi16 ? n32 : n10762;
  assign n10764 = pi15 ? n10758 : n10763;
  assign n10765 = pi18 ? n2615 : ~n880;
  assign n10766 = pi17 ? n32 : n10765;
  assign n10767 = pi16 ? n32 : n10766;
  assign n10768 = pi15 ? n10767 : n10283;
  assign n10769 = pi14 ? n10764 : n10768;
  assign n10770 = pi13 ? n10760 : n10769;
  assign n10771 = pi18 ? n2622 : ~n940;
  assign n10772 = pi17 ? n32 : n10771;
  assign n10773 = pi16 ? n32 : n10772;
  assign n10774 = pi14 ? n10283 : n10773;
  assign n10775 = pi15 ? n10291 : n10530;
  assign n10776 = pi18 ? n595 : ~n10053;
  assign n10777 = pi17 ? n32 : n10776;
  assign n10778 = pi16 ? n32 : n10777;
  assign n10779 = pi18 ? n595 : ~n684;
  assign n10780 = pi17 ? n32 : n10779;
  assign n10781 = pi16 ? n32 : n10780;
  assign n10782 = pi15 ? n10778 : n10781;
  assign n10783 = pi14 ? n10775 : n10782;
  assign n10784 = pi13 ? n10774 : n10783;
  assign n10785 = pi12 ? n10770 : n10784;
  assign n10786 = pi18 ? n595 : ~n10328;
  assign n10787 = pi17 ? n32 : n10786;
  assign n10788 = pi16 ? n32 : n10787;
  assign n10789 = pi18 ? n2627 : ~n684;
  assign n10790 = pi17 ? n32 : n10789;
  assign n10791 = pi16 ? n32 : n10790;
  assign n10792 = pi15 ? n10788 : n10791;
  assign n10793 = pi20 ? n342 : ~n623;
  assign n10794 = pi19 ? n32 : n10793;
  assign n10795 = pi18 ? n508 : ~n10794;
  assign n10796 = pi17 ? n32 : n10795;
  assign n10797 = pi16 ? n32 : n10796;
  assign n10798 = pi18 ? n508 : ~n684;
  assign n10799 = pi17 ? n32 : n10798;
  assign n10800 = pi16 ? n32 : n10799;
  assign n10801 = pi15 ? n10797 : n10800;
  assign n10802 = pi14 ? n10792 : n10801;
  assign n10803 = pi18 ? n323 : ~n10569;
  assign n10804 = pi17 ? n32 : n10803;
  assign n10805 = pi16 ? n32 : n10804;
  assign n10806 = pi18 ? n2291 : ~n2043;
  assign n10807 = pi17 ? n32 : n10806;
  assign n10808 = pi16 ? n32 : n10807;
  assign n10809 = pi15 ? n10805 : n10808;
  assign n10810 = pi20 ? n342 : ~n160;
  assign n10811 = pi19 ? n32 : n10810;
  assign n10812 = pi18 ? n2291 : ~n10811;
  assign n10813 = pi17 ? n32 : n10812;
  assign n10814 = pi16 ? n32 : n10813;
  assign n10815 = pi15 ? n10814 : n9737;
  assign n10816 = pi14 ? n10809 : n10815;
  assign n10817 = pi13 ? n10802 : n10816;
  assign n10818 = pi18 ? n797 : ~n8213;
  assign n10819 = pi17 ? n32 : n10818;
  assign n10820 = pi16 ? n32 : n10819;
  assign n10821 = pi18 ? n797 : ~n496;
  assign n10822 = pi17 ? n32 : n10821;
  assign n10823 = pi16 ? n32 : n10822;
  assign n10824 = pi15 ? n10820 : n10823;
  assign n10825 = pi18 ? n797 : ~n10594;
  assign n10826 = pi17 ? n32 : n10825;
  assign n10827 = pi16 ? n32 : n10826;
  assign n10828 = pi15 ? n10827 : n10565;
  assign n10829 = pi14 ? n10824 : n10828;
  assign n10830 = pi18 ? n605 : ~n9598;
  assign n10831 = pi17 ? n32 : n10830;
  assign n10832 = pi16 ? n32 : n10831;
  assign n10833 = pi18 ? n605 : ~n684;
  assign n10834 = pi17 ? n32 : n10833;
  assign n10835 = pi16 ? n32 : n10834;
  assign n10836 = pi15 ? n10832 : n10835;
  assign n10837 = pi18 ? n605 : ~n8804;
  assign n10838 = pi17 ? n32 : n10837;
  assign n10839 = pi16 ? n32 : n10838;
  assign n10840 = pi15 ? n10839 : n10835;
  assign n10841 = pi14 ? n10836 : n10840;
  assign n10842 = pi13 ? n10829 : n10841;
  assign n10843 = pi12 ? n10817 : n10842;
  assign n10844 = pi11 ? n10785 : n10843;
  assign n10845 = pi18 ? n605 : ~n10616;
  assign n10846 = pi17 ? n32 : n10845;
  assign n10847 = pi16 ? n32 : n10846;
  assign n10848 = pi15 ? n10847 : n10582;
  assign n10849 = pi18 ? n2424 : ~n245;
  assign n10850 = pi17 ? n32 : n10849;
  assign n10851 = pi16 ? n32 : n10850;
  assign n10852 = pi18 ? n418 : ~n4559;
  assign n10853 = pi17 ? n32 : n10852;
  assign n10854 = pi16 ? n32 : n10853;
  assign n10855 = pi15 ? n10851 : n10854;
  assign n10856 = pi14 ? n10848 : n10855;
  assign n10857 = pi20 ? n52 : n141;
  assign n10858 = pi19 ? n32 : n10857;
  assign n10859 = pi18 ? n418 : ~n10858;
  assign n10860 = pi17 ? n32 : n10859;
  assign n10861 = pi16 ? n32 : n10860;
  assign n10862 = pi21 ? n1939 : ~n206;
  assign n10863 = pi20 ? n10862 : n32;
  assign n10864 = pi19 ? n32 : ~n10863;
  assign n10865 = pi18 ? n418 : ~n10864;
  assign n10866 = pi17 ? n32 : n10865;
  assign n10867 = pi16 ? n32 : n10866;
  assign n10868 = pi15 ? n10861 : n10867;
  assign n10869 = pi21 ? n51 : n405;
  assign n10870 = pi20 ? n10869 : ~n32;
  assign n10871 = pi19 ? n32 : n10870;
  assign n10872 = pi18 ? n418 : ~n10871;
  assign n10873 = pi17 ? n32 : n10872;
  assign n10874 = pi16 ? n32 : n10873;
  assign n10875 = pi15 ? n10874 : n10867;
  assign n10876 = pi14 ? n10868 : n10875;
  assign n10877 = pi13 ? n10856 : n10876;
  assign n10878 = pi21 ? n405 : ~n405;
  assign n10879 = pi20 ? n10878 : n32;
  assign n10880 = pi19 ? n32 : ~n10879;
  assign n10881 = pi18 ? n3786 : ~n10880;
  assign n10882 = pi17 ? n32 : n10881;
  assign n10883 = pi16 ? n32 : n10882;
  assign n10884 = pi19 ? n2303 : ~n267;
  assign n10885 = pi18 ? n10884 : ~n684;
  assign n10886 = pi17 ? n32 : n10885;
  assign n10887 = pi16 ? n32 : n10886;
  assign n10888 = pi15 ? n10883 : n10887;
  assign n10889 = pi21 ? n174 : n259;
  assign n10890 = pi20 ? n10889 : ~n32;
  assign n10891 = pi19 ? n32 : n10890;
  assign n10892 = pi18 ? n2304 : ~n10891;
  assign n10893 = pi17 ? n32 : n10892;
  assign n10894 = pi16 ? n32 : n10893;
  assign n10895 = pi20 ? n1377 : ~n32;
  assign n10896 = pi19 ? n32 : n10895;
  assign n10897 = pi18 ? n2304 : ~n10896;
  assign n10898 = pi17 ? n32 : n10897;
  assign n10899 = pi16 ? n32 : n10898;
  assign n10900 = pi15 ? n10894 : n10899;
  assign n10901 = pi14 ? n10888 : n10900;
  assign n10902 = pi19 ? n32 : ~n9724;
  assign n10903 = pi18 ? n2304 : ~n10902;
  assign n10904 = pi17 ? n32 : n10903;
  assign n10905 = pi16 ? n32 : n10904;
  assign n10906 = pi18 ? n532 : ~n6888;
  assign n10907 = pi17 ? n32 : n10906;
  assign n10908 = pi16 ? n32 : n10907;
  assign n10909 = pi18 ? n2298 : ~n10670;
  assign n10910 = pi17 ? n32 : n10909;
  assign n10911 = pi16 ? n32 : n10910;
  assign n10912 = pi15 ? n10908 : n10911;
  assign n10913 = pi14 ? n10905 : n10912;
  assign n10914 = pi13 ? n10901 : n10913;
  assign n10915 = pi12 ? n10877 : n10914;
  assign n10916 = pi18 ? n2298 : ~n6240;
  assign n10917 = pi17 ? n32 : n10916;
  assign n10918 = pi16 ? n32 : n10917;
  assign n10919 = pi18 ? n2298 : ~n2730;
  assign n10920 = pi17 ? n32 : n10919;
  assign n10921 = pi16 ? n32 : n10920;
  assign n10922 = pi15 ? n10918 : n10921;
  assign n10923 = pi19 ? n462 : n236;
  assign n10924 = pi18 ? n532 : ~n10923;
  assign n10925 = pi17 ? n32 : n10924;
  assign n10926 = pi16 ? n32 : n10925;
  assign n10927 = pi19 ? n275 : n236;
  assign n10928 = pi18 ? n532 : ~n10927;
  assign n10929 = pi17 ? n32 : n10928;
  assign n10930 = pi16 ? n32 : n10929;
  assign n10931 = pi15 ? n10926 : n10930;
  assign n10932 = pi14 ? n10922 : n10931;
  assign n10933 = pi18 ? n532 : ~n1750;
  assign n10934 = pi17 ? n32 : n10933;
  assign n10935 = pi16 ? n32 : n10934;
  assign n10936 = pi18 ? n532 : ~n595;
  assign n10937 = pi17 ? n32 : n10936;
  assign n10938 = pi16 ? n32 : n10937;
  assign n10939 = pi15 ? n10935 : n10938;
  assign n10940 = pi18 ? n532 : ~n4098;
  assign n10941 = pi17 ? n32 : n10940;
  assign n10942 = pi16 ? n32 : n10941;
  assign n10943 = pi18 ? n2424 : ~n508;
  assign n10944 = pi17 ? n32 : n10943;
  assign n10945 = pi16 ? n32 : n10944;
  assign n10946 = pi15 ? n10942 : n10945;
  assign n10947 = pi14 ? n10939 : n10946;
  assign n10948 = pi13 ? n10932 : n10947;
  assign n10949 = pi18 ? n2424 : ~n9427;
  assign n10950 = pi17 ? n32 : n10949;
  assign n10951 = pi16 ? n32 : n10950;
  assign n10952 = pi15 ? n10942 : n10951;
  assign n10953 = pi18 ? n605 : ~n418;
  assign n10954 = pi17 ? n32 : n10953;
  assign n10955 = pi16 ? n32 : n10954;
  assign n10956 = pi18 ? n605 : ~n2754;
  assign n10957 = pi17 ? n32 : n10956;
  assign n10958 = pi16 ? n32 : n10957;
  assign n10959 = pi15 ? n10955 : n10958;
  assign n10960 = pi14 ? n10952 : n10959;
  assign n10961 = pi18 ? n605 : ~n323;
  assign n10962 = pi17 ? n32 : n10961;
  assign n10963 = pi16 ? n32 : n10962;
  assign n10964 = pi18 ? n2291 : ~n797;
  assign n10965 = pi17 ? n32 : n10964;
  assign n10966 = pi16 ? n32 : n10965;
  assign n10967 = pi15 ? n10963 : n10966;
  assign n10968 = pi14 ? n10958 : n10967;
  assign n10969 = pi13 ? n10960 : n10968;
  assign n10970 = pi12 ? n10948 : n10969;
  assign n10971 = pi11 ? n10915 : n10970;
  assign n10972 = pi10 ? n10844 : n10971;
  assign n10973 = pi09 ? n10748 : n10972;
  assign n10974 = pi08 ? n10735 : n10973;
  assign n10975 = pi07 ? n10497 : n10974;
  assign n10976 = pi18 ? n1592 : ~n940;
  assign n10977 = pi17 ? n32 : n10976;
  assign n10978 = pi16 ? n32 : n10977;
  assign n10979 = pi15 ? n32 : n10978;
  assign n10980 = pi18 ? n1970 : ~n940;
  assign n10981 = pi17 ? n32 : n10980;
  assign n10982 = pi16 ? n32 : n10981;
  assign n10983 = pi18 ? n209 : ~n940;
  assign n10984 = pi17 ? n32 : n10983;
  assign n10985 = pi16 ? n32 : n10984;
  assign n10986 = pi15 ? n10982 : n10985;
  assign n10987 = pi14 ? n10979 : n10986;
  assign n10988 = pi13 ? n32 : n10987;
  assign n10989 = pi12 ? n32 : n10988;
  assign n10990 = pi11 ? n32 : n10989;
  assign n10991 = pi10 ? n32 : n10990;
  assign n10992 = pi16 ? n32 : n942;
  assign n10993 = pi16 ? n32 : n1046;
  assign n10994 = pi15 ? n10992 : n10993;
  assign n10995 = pi16 ? n32 : n1059;
  assign n10996 = pi15 ? n10498 : n10995;
  assign n10997 = pi14 ? n10994 : n10996;
  assign n10998 = pi18 ? n684 : ~n880;
  assign n10999 = pi17 ? n32 : n10998;
  assign n11000 = pi16 ? n32 : n10999;
  assign n11001 = pi15 ? n10995 : n11000;
  assign n11002 = pi18 ? n4244 : ~n880;
  assign n11003 = pi17 ? n32 : n11002;
  assign n11004 = pi16 ? n32 : n11003;
  assign n11005 = pi15 ? n11004 : n10000;
  assign n11006 = pi14 ? n11001 : n11005;
  assign n11007 = pi13 ? n10997 : n11006;
  assign n11008 = pi14 ? n10000 : n10004;
  assign n11009 = pi15 ? n10526 : n10767;
  assign n11010 = pi21 ? n124 : n1939;
  assign n11011 = pi20 ? n32 : n11010;
  assign n11012 = pi19 ? n32 : n11011;
  assign n11013 = pi18 ? n1750 : ~n11012;
  assign n11014 = pi17 ? n32 : n11013;
  assign n11015 = pi16 ? n32 : n11014;
  assign n11016 = pi15 ? n11015 : n10283;
  assign n11017 = pi14 ? n11009 : n11016;
  assign n11018 = pi13 ? n11008 : n11017;
  assign n11019 = pi12 ? n11007 : n11018;
  assign n11020 = pi18 ? n1750 : ~n8547;
  assign n11021 = pi17 ? n32 : n11020;
  assign n11022 = pi16 ? n32 : n11021;
  assign n11023 = pi18 ? n2622 : ~n684;
  assign n11024 = pi17 ? n32 : n11023;
  assign n11025 = pi16 ? n32 : n11024;
  assign n11026 = pi15 ? n11022 : n11025;
  assign n11027 = pi20 ? n32 : ~n1817;
  assign n11028 = pi19 ? n32 : n11027;
  assign n11029 = pi18 ? n2622 : ~n11028;
  assign n11030 = pi17 ? n32 : n11029;
  assign n11031 = pi16 ? n32 : n11030;
  assign n11032 = pi15 ? n11031 : n10291;
  assign n11033 = pi14 ? n11026 : n11032;
  assign n11034 = pi18 ? n702 : ~n11028;
  assign n11035 = pi17 ? n32 : n11034;
  assign n11036 = pi16 ? n32 : n11035;
  assign n11037 = pi15 ? n11036 : n10530;
  assign n11038 = pi18 ? n4098 : ~n10811;
  assign n11039 = pi17 ? n32 : n11038;
  assign n11040 = pi16 ? n32 : n11039;
  assign n11041 = pi18 ? n4098 : ~n684;
  assign n11042 = pi17 ? n32 : n11041;
  assign n11043 = pi16 ? n32 : n11042;
  assign n11044 = pi15 ? n11040 : n11043;
  assign n11045 = pi14 ? n11037 : n11044;
  assign n11046 = pi13 ? n11033 : n11045;
  assign n11047 = pi15 ? n10781 : n10791;
  assign n11048 = pi21 ? n9326 : ~n32;
  assign n11049 = pi20 ? n175 : n11048;
  assign n11050 = pi19 ? n32 : n11049;
  assign n11051 = pi18 ? n2627 : ~n11050;
  assign n11052 = pi17 ? n32 : n11051;
  assign n11053 = pi16 ? n32 : n11052;
  assign n11054 = pi18 ? n2754 : ~n1741;
  assign n11055 = pi17 ? n32 : n11054;
  assign n11056 = pi16 ? n32 : n11055;
  assign n11057 = pi15 ? n11053 : n11056;
  assign n11058 = pi14 ? n11047 : n11057;
  assign n11059 = pi20 ? n175 : ~n52;
  assign n11060 = pi19 ? n32 : n11059;
  assign n11061 = pi18 ? n323 : ~n11060;
  assign n11062 = pi17 ? n32 : n11061;
  assign n11063 = pi16 ? n32 : n11062;
  assign n11064 = pi18 ? n323 : ~n1741;
  assign n11065 = pi17 ? n32 : n11064;
  assign n11066 = pi16 ? n32 : n11065;
  assign n11067 = pi15 ? n11063 : n11066;
  assign n11068 = pi18 ? n323 : ~n341;
  assign n11069 = pi17 ? n32 : n11068;
  assign n11070 = pi16 ? n32 : n11069;
  assign n11071 = pi18 ? n323 : ~n880;
  assign n11072 = pi17 ? n32 : n11071;
  assign n11073 = pi16 ? n32 : n11072;
  assign n11074 = pi15 ? n11070 : n11073;
  assign n11075 = pi14 ? n11067 : n11074;
  assign n11076 = pi13 ? n11058 : n11075;
  assign n11077 = pi12 ? n11046 : n11076;
  assign n11078 = pi11 ? n11019 : n11077;
  assign n11079 = pi18 ? n323 : ~n245;
  assign n11080 = pi17 ? n32 : n11079;
  assign n11081 = pi16 ? n32 : n11080;
  assign n11082 = pi15 ? n11081 : n11073;
  assign n11083 = pi18 ? n2291 : ~n366;
  assign n11084 = pi17 ? n32 : n11083;
  assign n11085 = pi16 ? n32 : n11084;
  assign n11086 = pi21 ? n1939 : n32;
  assign n11087 = pi20 ? n11086 : n141;
  assign n11088 = pi19 ? n32 : n11087;
  assign n11089 = pi18 ? n797 : ~n11088;
  assign n11090 = pi17 ? n32 : n11089;
  assign n11091 = pi16 ? n32 : n11090;
  assign n11092 = pi15 ? n11085 : n11091;
  assign n11093 = pi14 ? n11082 : n11092;
  assign n11094 = pi18 ? n797 : ~n3780;
  assign n11095 = pi17 ? n32 : n11094;
  assign n11096 = pi16 ? n32 : n11095;
  assign n11097 = pi21 ? n51 : n206;
  assign n11098 = pi20 ? n11097 : ~n32;
  assign n11099 = pi19 ? n32 : n11098;
  assign n11100 = pi18 ? n797 : ~n11099;
  assign n11101 = pi17 ? n32 : n11100;
  assign n11102 = pi16 ? n32 : n11101;
  assign n11103 = pi15 ? n11096 : n11102;
  assign n11104 = pi18 ? n797 : ~n10646;
  assign n11105 = pi17 ? n32 : n11104;
  assign n11106 = pi16 ? n32 : n11105;
  assign n11107 = pi21 ? n206 : n405;
  assign n11108 = pi20 ? n11107 : ~n32;
  assign n11109 = pi19 ? n32 : n11108;
  assign n11110 = pi18 ? n797 : ~n11109;
  assign n11111 = pi17 ? n32 : n11110;
  assign n11112 = pi16 ? n32 : n11111;
  assign n11113 = pi15 ? n11106 : n11112;
  assign n11114 = pi14 ? n11103 : n11113;
  assign n11115 = pi13 ? n11093 : n11114;
  assign n11116 = pi21 ? n66 : n206;
  assign n11117 = pi20 ? n11116 : ~n32;
  assign n11118 = pi19 ? n32 : n11117;
  assign n11119 = pi18 ? n2413 : ~n11118;
  assign n11120 = pi17 ? n32 : n11119;
  assign n11121 = pi16 ? n32 : n11120;
  assign n11122 = pi21 ? n1939 : n259;
  assign n11123 = pi20 ? n11122 : ~n32;
  assign n11124 = pi19 ? n32 : n11123;
  assign n11125 = pi18 ? n3786 : ~n11124;
  assign n11126 = pi17 ? n32 : n11125;
  assign n11127 = pi16 ? n32 : n11126;
  assign n11128 = pi15 ? n11121 : n11127;
  assign n11129 = pi18 ? n3786 : ~n6653;
  assign n11130 = pi17 ? n32 : n11129;
  assign n11131 = pi16 ? n32 : n11130;
  assign n11132 = pi19 ? n32 : n288;
  assign n11133 = pi18 ? n2413 : ~n11132;
  assign n11134 = pi17 ? n32 : n11133;
  assign n11135 = pi16 ? n32 : n11134;
  assign n11136 = pi15 ? n11131 : n11135;
  assign n11137 = pi14 ? n11128 : n11136;
  assign n11138 = pi18 ? n2413 : ~n1758;
  assign n11139 = pi17 ? n32 : n11138;
  assign n11140 = pi16 ? n32 : n11139;
  assign n11141 = pi15 ? n11135 : n11140;
  assign n11142 = pi18 ? n2413 : ~n697;
  assign n11143 = pi17 ? n32 : n11142;
  assign n11144 = pi16 ? n32 : n11143;
  assign n11145 = pi20 ? n32 : ~n501;
  assign n11146 = pi19 ? n11145 : ~n53;
  assign n11147 = pi18 ? n605 : ~n11146;
  assign n11148 = pi17 ? n32 : n11147;
  assign n11149 = pi16 ? n32 : n11148;
  assign n11150 = pi15 ? n11144 : n11149;
  assign n11151 = pi14 ? n11141 : n11150;
  assign n11152 = pi13 ? n11137 : n11151;
  assign n11153 = pi12 ? n11115 : n11152;
  assign n11154 = pi19 ? n6057 : n1941;
  assign n11155 = pi18 ? n605 : ~n11154;
  assign n11156 = pi17 ? n32 : n11155;
  assign n11157 = pi16 ? n32 : n11156;
  assign n11158 = pi18 ? n605 : ~n2730;
  assign n11159 = pi17 ? n32 : n11158;
  assign n11160 = pi16 ? n32 : n11159;
  assign n11161 = pi15 ? n11157 : n11160;
  assign n11162 = pi18 ? n605 : ~n772;
  assign n11163 = pi17 ? n32 : n11162;
  assign n11164 = pi16 ? n32 : n11163;
  assign n11165 = pi18 ? n605 : ~n1750;
  assign n11166 = pi17 ? n32 : n11165;
  assign n11167 = pi16 ? n32 : n11166;
  assign n11168 = pi15 ? n11164 : n11167;
  assign n11169 = pi14 ? n11161 : n11168;
  assign n11170 = pi22 ? n65 : n34;
  assign n11171 = pi21 ? n32 : n11170;
  assign n11172 = pi20 ? n32 : n11171;
  assign n11173 = pi19 ? n11172 : ~n32;
  assign n11174 = pi18 ? n323 : ~n11173;
  assign n11175 = pi17 ? n32 : n11174;
  assign n11176 = pi16 ? n32 : n11175;
  assign n11177 = pi18 ? n323 : ~n4098;
  assign n11178 = pi17 ? n32 : n11177;
  assign n11179 = pi16 ? n32 : n11178;
  assign n11180 = pi15 ? n11176 : n11179;
  assign n11181 = pi14 ? n11176 : n11180;
  assign n11182 = pi13 ? n11169 : n11181;
  assign n11183 = pi20 ? n32 : n8630;
  assign n11184 = pi19 ? n11183 : ~n32;
  assign n11185 = pi18 ? n323 : ~n11184;
  assign n11186 = pi17 ? n32 : n11185;
  assign n11187 = pi16 ? n32 : n11186;
  assign n11188 = pi18 ? n323 : ~n323;
  assign n11189 = pi17 ? n32 : n11188;
  assign n11190 = pi16 ? n32 : n11189;
  assign n11191 = pi15 ? n11187 : n11190;
  assign n11192 = pi18 ? n323 : ~n2754;
  assign n11193 = pi17 ? n32 : n11192;
  assign n11194 = pi16 ? n32 : n11193;
  assign n11195 = pi14 ? n11191 : n11194;
  assign n11196 = pi18 ? n508 : ~n2754;
  assign n11197 = pi17 ? n32 : n11196;
  assign n11198 = pi16 ? n32 : n11197;
  assign n11199 = pi15 ? n11198 : n11194;
  assign n11200 = pi18 ? n508 : ~n323;
  assign n11201 = pi17 ? n32 : n11200;
  assign n11202 = pi16 ? n32 : n11201;
  assign n11203 = pi18 ? n508 : ~n797;
  assign n11204 = pi17 ? n32 : n11203;
  assign n11205 = pi16 ? n32 : n11204;
  assign n11206 = pi15 ? n11202 : n11205;
  assign n11207 = pi14 ? n11199 : n11206;
  assign n11208 = pi13 ? n11195 : n11207;
  assign n11209 = pi12 ? n11182 : n11208;
  assign n11210 = pi11 ? n11153 : n11209;
  assign n11211 = pi10 ? n11078 : n11210;
  assign n11212 = pi09 ? n10991 : n11211;
  assign n11213 = pi18 ? n2142 : ~n940;
  assign n11214 = pi17 ? n32 : n11213;
  assign n11215 = pi16 ? n32 : n11214;
  assign n11216 = pi15 ? n32 : n11215;
  assign n11217 = pi18 ? n1841 : ~n940;
  assign n11218 = pi17 ? n32 : n11217;
  assign n11219 = pi16 ? n32 : n11218;
  assign n11220 = pi18 ? n940 : ~n940;
  assign n11221 = pi17 ? n32 : n11220;
  assign n11222 = pi16 ? n32 : n11221;
  assign n11223 = pi15 ? n11219 : n11222;
  assign n11224 = pi14 ? n11216 : n11223;
  assign n11225 = pi13 ? n32 : n11224;
  assign n11226 = pi12 ? n32 : n11225;
  assign n11227 = pi11 ? n32 : n11226;
  assign n11228 = pi10 ? n32 : n11227;
  assign n11229 = pi18 ? n1477 : ~n940;
  assign n11230 = pi17 ? n32 : n11229;
  assign n11231 = pi16 ? n32 : n11230;
  assign n11232 = pi18 ? n751 : ~n940;
  assign n11233 = pi17 ? n32 : n11232;
  assign n11234 = pi16 ? n32 : n11233;
  assign n11235 = pi15 ? n11231 : n11234;
  assign n11236 = pi18 ? n1970 : ~n880;
  assign n11237 = pi17 ? n32 : n11236;
  assign n11238 = pi16 ? n32 : n11237;
  assign n11239 = pi15 ? n10738 : n11238;
  assign n11240 = pi14 ? n11235 : n11239;
  assign n11241 = pi15 ? n11238 : n11000;
  assign n11242 = pi18 ? n2835 : ~n880;
  assign n11243 = pi17 ? n32 : n11242;
  assign n11244 = pi16 ? n32 : n11243;
  assign n11245 = pi15 ? n11244 : n10260;
  assign n11246 = pi14 ? n11241 : n11245;
  assign n11247 = pi13 ? n11240 : n11246;
  assign n11248 = pi14 ? n10260 : n10264;
  assign n11249 = pi15 ? n10763 : n11004;
  assign n11250 = pi20 ? n32 : ~n726;
  assign n11251 = pi19 ? n32 : n11250;
  assign n11252 = pi18 ? n962 : ~n11251;
  assign n11253 = pi17 ? n32 : n11252;
  assign n11254 = pi16 ? n32 : n11253;
  assign n11255 = pi15 ? n11254 : n10000;
  assign n11256 = pi14 ? n11249 : n11255;
  assign n11257 = pi13 ? n11248 : n11256;
  assign n11258 = pi12 ? n11247 : n11257;
  assign n11259 = pi18 ? n962 : ~n8547;
  assign n11260 = pi17 ? n32 : n11259;
  assign n11261 = pi16 ? n32 : n11260;
  assign n11262 = pi18 ? n2730 : ~n684;
  assign n11263 = pi17 ? n32 : n11262;
  assign n11264 = pi16 ? n32 : n11263;
  assign n11265 = pi15 ? n11261 : n11264;
  assign n11266 = pi18 ? n2730 : ~n11028;
  assign n11267 = pi17 ? n32 : n11266;
  assign n11268 = pi16 ? n32 : n11267;
  assign n11269 = pi15 ? n11268 : n10526;
  assign n11270 = pi14 ? n11265 : n11269;
  assign n11271 = pi18 ? n697 : ~n11028;
  assign n11272 = pi17 ? n32 : n11271;
  assign n11273 = pi16 ? n32 : n11272;
  assign n11274 = pi15 ? n11273 : n10767;
  assign n11275 = pi18 ? n2615 : ~n10811;
  assign n11276 = pi17 ? n32 : n11275;
  assign n11277 = pi16 ? n32 : n11276;
  assign n11278 = pi18 ? n2615 : ~n684;
  assign n11279 = pi17 ? n32 : n11278;
  assign n11280 = pi16 ? n32 : n11279;
  assign n11281 = pi15 ? n11277 : n11280;
  assign n11282 = pi14 ? n11274 : n11281;
  assign n11283 = pi13 ? n11270 : n11282;
  assign n11284 = pi18 ? n1750 : ~n10594;
  assign n11285 = pi17 ? n32 : n11284;
  assign n11286 = pi16 ? n32 : n11285;
  assign n11287 = pi18 ? n1750 : ~n684;
  assign n11288 = pi17 ? n32 : n11287;
  assign n11289 = pi16 ? n32 : n11288;
  assign n11290 = pi15 ? n11286 : n11289;
  assign n11291 = pi18 ? n2622 : ~n11050;
  assign n11292 = pi17 ? n32 : n11291;
  assign n11293 = pi16 ? n32 : n11292;
  assign n11294 = pi18 ? n2622 : ~n1741;
  assign n11295 = pi17 ? n32 : n11294;
  assign n11296 = pi16 ? n32 : n11295;
  assign n11297 = pi15 ? n11293 : n11296;
  assign n11298 = pi14 ? n11290 : n11297;
  assign n11299 = pi18 ? n702 : ~n8236;
  assign n11300 = pi17 ? n32 : n11299;
  assign n11301 = pi16 ? n32 : n11300;
  assign n11302 = pi18 ? n702 : ~n1741;
  assign n11303 = pi17 ? n32 : n11302;
  assign n11304 = pi16 ? n32 : n11303;
  assign n11305 = pi15 ? n11301 : n11304;
  assign n11306 = pi18 ? n702 : ~n245;
  assign n11307 = pi17 ? n32 : n11306;
  assign n11308 = pi16 ? n32 : n11307;
  assign n11309 = pi15 ? n11308 : n10291;
  assign n11310 = pi14 ? n11305 : n11309;
  assign n11311 = pi13 ? n11298 : n11310;
  assign n11312 = pi12 ? n11283 : n11311;
  assign n11313 = pi11 ? n11258 : n11312;
  assign n11314 = pi18 ? n4098 : ~n245;
  assign n11315 = pi17 ? n32 : n11314;
  assign n11316 = pi16 ? n32 : n11315;
  assign n11317 = pi15 ? n11316 : n10530;
  assign n11318 = pi18 ? n2747 : ~n366;
  assign n11319 = pi17 ? n32 : n11318;
  assign n11320 = pi16 ? n32 : n11319;
  assign n11321 = pi20 ? n915 : n141;
  assign n11322 = pi19 ? n32 : n11321;
  assign n11323 = pi18 ? n520 : ~n11322;
  assign n11324 = pi17 ? n32 : n11323;
  assign n11325 = pi16 ? n32 : n11324;
  assign n11326 = pi15 ? n11320 : n11325;
  assign n11327 = pi14 ? n11317 : n11326;
  assign n11328 = pi21 ? n1939 : n9326;
  assign n11329 = pi20 ? n11328 : ~n32;
  assign n11330 = pi19 ? n32 : n11329;
  assign n11331 = pi18 ? n520 : ~n11330;
  assign n11332 = pi17 ? n32 : n11331;
  assign n11333 = pi16 ? n32 : n11332;
  assign n11334 = pi21 ? n51 : n9326;
  assign n11335 = pi20 ? n11334 : ~n32;
  assign n11336 = pi19 ? n32 : n11335;
  assign n11337 = pi18 ? n520 : ~n11336;
  assign n11338 = pi17 ? n32 : n11337;
  assign n11339 = pi16 ? n32 : n11338;
  assign n11340 = pi15 ? n11333 : n11339;
  assign n11341 = pi18 ? n520 : ~n10646;
  assign n11342 = pi17 ? n32 : n11341;
  assign n11343 = pi16 ? n32 : n11342;
  assign n11344 = pi18 ? n520 : ~n11109;
  assign n11345 = pi17 ? n32 : n11344;
  assign n11346 = pi16 ? n32 : n11345;
  assign n11347 = pi15 ? n11343 : n11346;
  assign n11348 = pi14 ? n11340 : n11347;
  assign n11349 = pi13 ? n11327 : n11348;
  assign n11350 = pi19 ? n519 : ~n8622;
  assign n11351 = pi18 ? n11350 : ~n684;
  assign n11352 = pi17 ? n32 : n11351;
  assign n11353 = pi16 ? n32 : n11352;
  assign n11354 = pi18 ? n2754 : ~n11124;
  assign n11355 = pi17 ? n32 : n11354;
  assign n11356 = pi16 ? n32 : n11355;
  assign n11357 = pi15 ? n11353 : n11356;
  assign n11358 = pi18 ? n2754 : ~n6653;
  assign n11359 = pi17 ? n32 : n11358;
  assign n11360 = pi16 ? n32 : n11359;
  assign n11361 = pi18 ? n2754 : ~n11132;
  assign n11362 = pi17 ? n32 : n11361;
  assign n11363 = pi16 ? n32 : n11362;
  assign n11364 = pi15 ? n11360 : n11363;
  assign n11365 = pi14 ? n11357 : n11364;
  assign n11366 = pi18 ? n2754 : ~n1758;
  assign n11367 = pi17 ? n32 : n11366;
  assign n11368 = pi16 ? n32 : n11367;
  assign n11369 = pi15 ? n11363 : n11368;
  assign n11370 = pi19 ? n654 : n236;
  assign n11371 = pi18 ? n2754 : ~n11370;
  assign n11372 = pi17 ? n32 : n11371;
  assign n11373 = pi16 ? n32 : n11372;
  assign n11374 = pi20 ? n32 : ~n314;
  assign n11375 = pi19 ? n11374 : ~n358;
  assign n11376 = pi18 ? n323 : ~n11375;
  assign n11377 = pi17 ? n32 : n11376;
  assign n11378 = pi16 ? n32 : n11377;
  assign n11379 = pi15 ? n11373 : n11378;
  assign n11380 = pi14 ? n11369 : n11379;
  assign n11381 = pi13 ? n11365 : n11380;
  assign n11382 = pi12 ? n11349 : n11381;
  assign n11383 = pi18 ? n323 : ~n2730;
  assign n11384 = pi17 ? n32 : n11383;
  assign n11385 = pi16 ? n32 : n11384;
  assign n11386 = pi19 ? n1818 : n236;
  assign n11387 = pi18 ? n323 : ~n11386;
  assign n11388 = pi17 ? n32 : n11387;
  assign n11389 = pi16 ? n32 : n11388;
  assign n11390 = pi15 ? n11385 : n11389;
  assign n11391 = pi18 ? n323 : ~n4581;
  assign n11392 = pi17 ? n32 : n11391;
  assign n11393 = pi16 ? n32 : n11392;
  assign n11394 = pi18 ? n508 : ~n11173;
  assign n11395 = pi17 ? n32 : n11394;
  assign n11396 = pi16 ? n32 : n11395;
  assign n11397 = pi15 ? n11393 : n11396;
  assign n11398 = pi14 ? n11390 : n11397;
  assign n11399 = pi18 ? n508 : ~n4098;
  assign n11400 = pi17 ? n32 : n11399;
  assign n11401 = pi16 ? n32 : n11400;
  assign n11402 = pi22 ? n32 : n33;
  assign n11403 = pi21 ? n32 : n11402;
  assign n11404 = pi20 ? n32 : n11403;
  assign n11405 = pi19 ? n11404 : ~n32;
  assign n11406 = pi18 ? n508 : ~n11405;
  assign n11407 = pi17 ? n32 : n11406;
  assign n11408 = pi16 ? n32 : n11407;
  assign n11409 = pi15 ? n11401 : n11408;
  assign n11410 = pi14 ? n11409 : n11401;
  assign n11411 = pi13 ? n11398 : n11410;
  assign n11412 = pi18 ? n508 : ~n2627;
  assign n11413 = pi17 ? n32 : n11412;
  assign n11414 = pi16 ? n32 : n11413;
  assign n11415 = pi15 ? n11414 : n11202;
  assign n11416 = pi18 ? n702 : ~n2754;
  assign n11417 = pi17 ? n32 : n11416;
  assign n11418 = pi16 ? n32 : n11417;
  assign n11419 = pi15 ? n11202 : n11418;
  assign n11420 = pi14 ? n11415 : n11419;
  assign n11421 = pi18 ? n702 : ~n323;
  assign n11422 = pi17 ? n32 : n11421;
  assign n11423 = pi16 ? n32 : n11422;
  assign n11424 = pi18 ? n702 : ~n605;
  assign n11425 = pi17 ? n32 : n11424;
  assign n11426 = pi16 ? n32 : n11425;
  assign n11427 = pi18 ? n702 : ~n418;
  assign n11428 = pi17 ? n32 : n11427;
  assign n11429 = pi16 ? n32 : n11428;
  assign n11430 = pi15 ? n11426 : n11429;
  assign n11431 = pi14 ? n11423 : n11430;
  assign n11432 = pi13 ? n11420 : n11431;
  assign n11433 = pi12 ? n11411 : n11432;
  assign n11434 = pi11 ? n11382 : n11433;
  assign n11435 = pi10 ? n11313 : n11434;
  assign n11436 = pi09 ? n11228 : n11435;
  assign n11437 = pi08 ? n11212 : n11436;
  assign n11438 = pi19 ? n1105 : ~n322;
  assign n11439 = pi18 ? n32 : n11438;
  assign n11440 = pi17 ? n32 : n11439;
  assign n11441 = pi16 ? n32 : n11440;
  assign n11442 = pi15 ? n32 : n11441;
  assign n11443 = pi18 ? n863 : ~n940;
  assign n11444 = pi17 ? n32 : n11443;
  assign n11445 = pi16 ? n32 : n11444;
  assign n11446 = pi15 ? n11215 : n11445;
  assign n11447 = pi14 ? n11442 : n11446;
  assign n11448 = pi13 ? n32 : n11447;
  assign n11449 = pi12 ? n32 : n11448;
  assign n11450 = pi11 ? n32 : n11449;
  assign n11451 = pi10 ? n32 : n11450;
  assign n11452 = pi15 ? n11445 : n10978;
  assign n11453 = pi18 ? n1592 : ~n880;
  assign n11454 = pi17 ? n32 : n11453;
  assign n11455 = pi16 ? n32 : n11454;
  assign n11456 = pi18 ? n1841 : ~n880;
  assign n11457 = pi17 ? n32 : n11456;
  assign n11458 = pi16 ? n32 : n11457;
  assign n11459 = pi15 ? n11455 : n11458;
  assign n11460 = pi14 ? n11452 : n11459;
  assign n11461 = pi18 ? n209 : ~n880;
  assign n11462 = pi17 ? n32 : n11461;
  assign n11463 = pi16 ? n32 : n11462;
  assign n11464 = pi15 ? n11458 : n11463;
  assign n11465 = pi18 ? n245 : ~n880;
  assign n11466 = pi17 ? n32 : n11465;
  assign n11467 = pi16 ? n32 : n11466;
  assign n11468 = pi15 ? n11467 : n10498;
  assign n11469 = pi14 ? n11464 : n11468;
  assign n11470 = pi13 ? n11460 : n11469;
  assign n11471 = pi16 ? n32 : n1243;
  assign n11472 = pi14 ? n10498 : n11471;
  assign n11473 = pi15 ? n11000 : n11244;
  assign n11474 = pi18 ? n590 : ~n11251;
  assign n11475 = pi17 ? n32 : n11474;
  assign n11476 = pi16 ? n32 : n11475;
  assign n11477 = pi15 ? n11476 : n10260;
  assign n11478 = pi14 ? n11473 : n11477;
  assign n11479 = pi13 ? n11472 : n11478;
  assign n11480 = pi12 ? n11470 : n11479;
  assign n11481 = pi18 ? n590 : ~n1965;
  assign n11482 = pi17 ? n32 : n11481;
  assign n11483 = pi16 ? n32 : n11482;
  assign n11484 = pi18 ? n2849 : ~n1965;
  assign n11485 = pi17 ? n32 : n11484;
  assign n11486 = pi16 ? n32 : n11485;
  assign n11487 = pi15 ? n11483 : n11486;
  assign n11488 = pi20 ? n428 : ~n1817;
  assign n11489 = pi19 ? n32 : n11488;
  assign n11490 = pi18 ? n2849 : ~n11489;
  assign n11491 = pi17 ? n32 : n11490;
  assign n11492 = pi16 ? n32 : n11491;
  assign n11493 = pi15 ? n11492 : n10763;
  assign n11494 = pi14 ? n11487 : n11493;
  assign n11495 = pi18 ? n496 : ~n1965;
  assign n11496 = pi17 ? n32 : n11495;
  assign n11497 = pi16 ? n32 : n11496;
  assign n11498 = pi18 ? n4244 : ~n1965;
  assign n11499 = pi17 ? n32 : n11498;
  assign n11500 = pi16 ? n32 : n11499;
  assign n11501 = pi15 ? n11497 : n11500;
  assign n11502 = pi14 ? n11501 : n11500;
  assign n11503 = pi13 ? n11494 : n11502;
  assign n11504 = pi20 ? n428 : ~n6229;
  assign n11505 = pi19 ? n32 : n11504;
  assign n11506 = pi18 ? n962 : ~n11505;
  assign n11507 = pi17 ? n32 : n11506;
  assign n11508 = pi16 ? n32 : n11507;
  assign n11509 = pi18 ? n962 : ~n1965;
  assign n11510 = pi17 ? n32 : n11509;
  assign n11511 = pi16 ? n32 : n11510;
  assign n11512 = pi15 ? n11508 : n11511;
  assign n11513 = pi18 ? n2730 : ~n209;
  assign n11514 = pi17 ? n32 : n11513;
  assign n11515 = pi16 ? n32 : n11514;
  assign n11516 = pi18 ? n2730 : ~n11050;
  assign n11517 = pi17 ? n32 : n11516;
  assign n11518 = pi16 ? n32 : n11517;
  assign n11519 = pi15 ? n11515 : n11518;
  assign n11520 = pi14 ? n11512 : n11519;
  assign n11521 = pi18 ? n697 : ~n1965;
  assign n11522 = pi17 ? n32 : n11521;
  assign n11523 = pi16 ? n32 : n11522;
  assign n11524 = pi18 ? n697 : ~n209;
  assign n11525 = pi17 ? n32 : n11524;
  assign n11526 = pi16 ? n32 : n11525;
  assign n11527 = pi15 ? n11523 : n11526;
  assign n11528 = pi18 ? n697 : ~n245;
  assign n11529 = pi17 ? n32 : n11528;
  assign n11530 = pi16 ? n32 : n11529;
  assign n11531 = pi20 ? n1817 : ~n32;
  assign n11532 = pi19 ? n32 : n11531;
  assign n11533 = pi18 ? n697 : ~n11532;
  assign n11534 = pi17 ? n32 : n11533;
  assign n11535 = pi16 ? n32 : n11534;
  assign n11536 = pi15 ? n11530 : n11535;
  assign n11537 = pi14 ? n11527 : n11536;
  assign n11538 = pi13 ? n11520 : n11537;
  assign n11539 = pi12 ? n11503 : n11538;
  assign n11540 = pi11 ? n11480 : n11539;
  assign n11541 = pi20 ? n9641 : ~n481;
  assign n11542 = pi19 ? n32 : n11541;
  assign n11543 = pi18 ? n697 : ~n11542;
  assign n11544 = pi17 ? n32 : n11543;
  assign n11545 = pi16 ? n32 : n11544;
  assign n11546 = pi20 ? n9641 : ~n32;
  assign n11547 = pi19 ? n32 : n11546;
  assign n11548 = pi18 ? n2615 : ~n11547;
  assign n11549 = pi17 ? n32 : n11548;
  assign n11550 = pi16 ? n32 : n11549;
  assign n11551 = pi15 ? n11545 : n11550;
  assign n11552 = pi18 ? n2615 : ~n366;
  assign n11553 = pi17 ? n32 : n11552;
  assign n11554 = pi16 ? n32 : n11553;
  assign n11555 = pi18 ? n1750 : ~n2962;
  assign n11556 = pi17 ? n32 : n11555;
  assign n11557 = pi16 ? n32 : n11556;
  assign n11558 = pi15 ? n11554 : n11557;
  assign n11559 = pi14 ? n11551 : n11558;
  assign n11560 = pi21 ? n206 : n100;
  assign n11561 = pi20 ? n11560 : ~n32;
  assign n11562 = pi19 ? n32 : n11561;
  assign n11563 = pi18 ? n1750 : ~n11562;
  assign n11564 = pi17 ? n32 : n11563;
  assign n11565 = pi16 ? n32 : n11564;
  assign n11566 = pi15 ? n11557 : n11565;
  assign n11567 = pi22 ? n32 : ~n65;
  assign n11568 = pi21 ? n11567 : ~n313;
  assign n11569 = pi20 ? n11568 : ~n32;
  assign n11570 = pi19 ? n32 : n11569;
  assign n11571 = pi18 ? n1750 : ~n11570;
  assign n11572 = pi17 ? n32 : n11571;
  assign n11573 = pi16 ? n32 : n11572;
  assign n11574 = pi21 ? n206 : ~n7500;
  assign n11575 = pi20 ? n11574 : ~n32;
  assign n11576 = pi19 ? n32 : n11575;
  assign n11577 = pi18 ? n595 : ~n11576;
  assign n11578 = pi17 ? n32 : n11577;
  assign n11579 = pi16 ? n32 : n11578;
  assign n11580 = pi15 ? n11573 : n11579;
  assign n11581 = pi14 ? n11566 : n11580;
  assign n11582 = pi13 ? n11559 : n11581;
  assign n11583 = pi21 ? n11567 : n259;
  assign n11584 = pi20 ? n11583 : ~n32;
  assign n11585 = pi19 ? n3495 : n11584;
  assign n11586 = pi18 ? n2622 : ~n11585;
  assign n11587 = pi17 ? n32 : n11586;
  assign n11588 = pi16 ? n32 : n11587;
  assign n11589 = pi21 ? n51 : ~n32;
  assign n11590 = pi20 ? n11589 : ~n32;
  assign n11591 = pi19 ? n32 : n11590;
  assign n11592 = pi18 ? n2627 : ~n11591;
  assign n11593 = pi17 ? n32 : n11592;
  assign n11594 = pi16 ? n32 : n11593;
  assign n11595 = pi15 ? n11588 : n11594;
  assign n11596 = pi18 ? n2627 : ~n6653;
  assign n11597 = pi17 ? n32 : n11596;
  assign n11598 = pi16 ? n32 : n11597;
  assign n11599 = pi18 ? n2627 : ~n697;
  assign n11600 = pi17 ? n32 : n11599;
  assign n11601 = pi16 ? n32 : n11600;
  assign n11602 = pi15 ? n11598 : n11601;
  assign n11603 = pi14 ? n11595 : n11602;
  assign n11604 = pi18 ? n2627 : ~n11132;
  assign n11605 = pi17 ? n32 : n11604;
  assign n11606 = pi16 ? n32 : n11605;
  assign n11607 = pi18 ? n2627 : ~n496;
  assign n11608 = pi17 ? n32 : n11607;
  assign n11609 = pi16 ? n32 : n11608;
  assign n11610 = pi15 ? n11606 : n11609;
  assign n11611 = pi18 ? n2627 : ~n2730;
  assign n11612 = pi17 ? n32 : n11611;
  assign n11613 = pi16 ? n32 : n11612;
  assign n11614 = pi18 ? n508 : ~n697;
  assign n11615 = pi17 ? n32 : n11614;
  assign n11616 = pi16 ? n32 : n11615;
  assign n11617 = pi15 ? n11613 : n11616;
  assign n11618 = pi14 ? n11610 : n11617;
  assign n11619 = pi13 ? n11603 : n11618;
  assign n11620 = pi12 ? n11582 : n11619;
  assign n11621 = pi19 ? n857 : n1941;
  assign n11622 = pi18 ? n508 : ~n11621;
  assign n11623 = pi17 ? n32 : n11622;
  assign n11624 = pi16 ? n32 : n11623;
  assign n11625 = pi15 ? n11624 : n11616;
  assign n11626 = pi18 ? n702 : ~n2615;
  assign n11627 = pi17 ? n32 : n11626;
  assign n11628 = pi16 ? n32 : n11627;
  assign n11629 = pi18 ? n702 : ~n4098;
  assign n11630 = pi17 ? n32 : n11629;
  assign n11631 = pi16 ? n32 : n11630;
  assign n11632 = pi15 ? n11628 : n11631;
  assign n11633 = pi14 ? n11625 : n11632;
  assign n11634 = pi18 ? n702 : ~n11405;
  assign n11635 = pi17 ? n32 : n11634;
  assign n11636 = pi16 ? n32 : n11635;
  assign n11637 = pi15 ? n11631 : n11636;
  assign n11638 = pi14 ? n11637 : n11631;
  assign n11639 = pi13 ? n11633 : n11638;
  assign n11640 = pi18 ? n702 : ~n2627;
  assign n11641 = pi17 ? n32 : n11640;
  assign n11642 = pi16 ? n32 : n11641;
  assign n11643 = pi15 ? n11642 : n11418;
  assign n11644 = pi18 ? n697 : ~n2754;
  assign n11645 = pi17 ? n32 : n11644;
  assign n11646 = pi16 ? n32 : n11645;
  assign n11647 = pi14 ? n11643 : n11646;
  assign n11648 = pi18 ? n697 : ~n323;
  assign n11649 = pi17 ? n32 : n11648;
  assign n11650 = pi16 ? n32 : n11649;
  assign n11651 = pi15 ? n11646 : n11650;
  assign n11652 = pi18 ? n697 : ~n605;
  assign n11653 = pi17 ? n32 : n11652;
  assign n11654 = pi16 ? n32 : n11653;
  assign n11655 = pi18 ? n697 : ~n418;
  assign n11656 = pi17 ? n32 : n11655;
  assign n11657 = pi16 ? n32 : n11656;
  assign n11658 = pi15 ? n11654 : n11657;
  assign n11659 = pi14 ? n11651 : n11658;
  assign n11660 = pi13 ? n11647 : n11659;
  assign n11661 = pi12 ? n11639 : n11660;
  assign n11662 = pi11 ? n11620 : n11661;
  assign n11663 = pi10 ? n11540 : n11662;
  assign n11664 = pi09 ? n11451 : n11663;
  assign n11665 = pi19 ? n1941 : ~n322;
  assign n11666 = pi18 ? n32 : n11665;
  assign n11667 = pi17 ? n32 : n11666;
  assign n11668 = pi16 ? n32 : n11667;
  assign n11669 = pi15 ? n32 : n11668;
  assign n11670 = pi18 ? n32 : ~n940;
  assign n11671 = pi17 ? n32 : n11670;
  assign n11672 = pi16 ? n32 : n11671;
  assign n11673 = pi15 ? n11441 : n11672;
  assign n11674 = pi14 ? n11669 : n11673;
  assign n11675 = pi13 ? n32 : n11674;
  assign n11676 = pi12 ? n32 : n11675;
  assign n11677 = pi11 ? n32 : n11676;
  assign n11678 = pi10 ? n32 : n11677;
  assign n11679 = pi18 ? n1575 : ~n940;
  assign n11680 = pi17 ? n32 : n11679;
  assign n11681 = pi16 ? n32 : n11680;
  assign n11682 = pi15 ? n11672 : n11681;
  assign n11683 = pi18 ? n1575 : ~n880;
  assign n11684 = pi17 ? n32 : n11683;
  assign n11685 = pi16 ? n32 : n11684;
  assign n11686 = pi18 ? n2142 : ~n880;
  assign n11687 = pi17 ? n32 : n11686;
  assign n11688 = pi16 ? n32 : n11687;
  assign n11689 = pi15 ? n11685 : n11688;
  assign n11690 = pi14 ? n11682 : n11689;
  assign n11691 = pi18 ? n863 : ~n880;
  assign n11692 = pi17 ? n32 : n11691;
  assign n11693 = pi16 ? n32 : n11692;
  assign n11694 = pi18 ? n940 : ~n880;
  assign n11695 = pi17 ? n32 : n11694;
  assign n11696 = pi16 ? n32 : n11695;
  assign n11697 = pi15 ? n11693 : n11696;
  assign n11698 = pi18 ? n1477 : ~n880;
  assign n11699 = pi17 ? n32 : n11698;
  assign n11700 = pi16 ? n32 : n11699;
  assign n11701 = pi15 ? n11700 : n10738;
  assign n11702 = pi14 ? n11697 : n11701;
  assign n11703 = pi13 ? n11690 : n11702;
  assign n11704 = pi14 ? n10738 : n10982;
  assign n11705 = pi15 ? n11463 : n11467;
  assign n11706 = pi18 ? n341 : ~n11251;
  assign n11707 = pi17 ? n32 : n11706;
  assign n11708 = pi16 ? n32 : n11707;
  assign n11709 = pi15 ? n11708 : n10498;
  assign n11710 = pi14 ? n11705 : n11709;
  assign n11711 = pi13 ? n11704 : n11710;
  assign n11712 = pi12 ? n11703 : n11711;
  assign n11713 = pi18 ? n341 : ~n1965;
  assign n11714 = pi17 ? n32 : n11713;
  assign n11715 = pi16 ? n32 : n11714;
  assign n11716 = pi16 ? n32 : n2101;
  assign n11717 = pi15 ? n11715 : n11716;
  assign n11718 = pi18 ? n366 : ~n11489;
  assign n11719 = pi17 ? n32 : n11718;
  assign n11720 = pi16 ? n32 : n11719;
  assign n11721 = pi15 ? n11720 : n11000;
  assign n11722 = pi14 ? n11717 : n11721;
  assign n11723 = pi18 ? n684 : ~n1965;
  assign n11724 = pi17 ? n32 : n11723;
  assign n11725 = pi16 ? n32 : n11724;
  assign n11726 = pi18 ? n2835 : ~n1965;
  assign n11727 = pi17 ? n32 : n11726;
  assign n11728 = pi16 ? n32 : n11727;
  assign n11729 = pi15 ? n11725 : n11728;
  assign n11730 = pi14 ? n11729 : n11728;
  assign n11731 = pi13 ? n11722 : n11730;
  assign n11732 = pi18 ? n590 : ~n11505;
  assign n11733 = pi17 ? n32 : n11732;
  assign n11734 = pi16 ? n32 : n11733;
  assign n11735 = pi15 ? n11734 : n11483;
  assign n11736 = pi18 ? n2849 : ~n209;
  assign n11737 = pi17 ? n32 : n11736;
  assign n11738 = pi16 ? n32 : n11737;
  assign n11739 = pi18 ? n2849 : ~n11050;
  assign n11740 = pi17 ? n32 : n11739;
  assign n11741 = pi16 ? n32 : n11740;
  assign n11742 = pi15 ? n11738 : n11741;
  assign n11743 = pi14 ? n11735 : n11742;
  assign n11744 = pi18 ? n496 : ~n1970;
  assign n11745 = pi17 ? n32 : n11744;
  assign n11746 = pi16 ? n32 : n11745;
  assign n11747 = pi15 ? n11497 : n11746;
  assign n11748 = pi18 ? n496 : ~n245;
  assign n11749 = pi17 ? n32 : n11748;
  assign n11750 = pi16 ? n32 : n11749;
  assign n11751 = pi18 ? n496 : ~n7038;
  assign n11752 = pi17 ? n32 : n11751;
  assign n11753 = pi16 ? n32 : n11752;
  assign n11754 = pi15 ? n11750 : n11753;
  assign n11755 = pi14 ? n11747 : n11754;
  assign n11756 = pi13 ? n11743 : n11755;
  assign n11757 = pi12 ? n11731 : n11756;
  assign n11758 = pi11 ? n11712 : n11757;
  assign n11759 = pi18 ? n496 : ~n7231;
  assign n11760 = pi17 ? n32 : n11759;
  assign n11761 = pi16 ? n32 : n11760;
  assign n11762 = pi20 ? n1324 : ~n481;
  assign n11763 = pi19 ? n32 : n11762;
  assign n11764 = pi18 ? n4244 : ~n11763;
  assign n11765 = pi17 ? n32 : n11764;
  assign n11766 = pi16 ? n32 : n11765;
  assign n11767 = pi15 ? n11761 : n11766;
  assign n11768 = pi20 ? n111 : n141;
  assign n11769 = pi19 ? n32 : n11768;
  assign n11770 = pi18 ? n4244 : ~n11769;
  assign n11771 = pi17 ? n32 : n11770;
  assign n11772 = pi16 ? n32 : n11771;
  assign n11773 = pi18 ? n962 : ~n2962;
  assign n11774 = pi17 ? n32 : n11773;
  assign n11775 = pi16 ? n32 : n11774;
  assign n11776 = pi15 ? n11772 : n11775;
  assign n11777 = pi14 ? n11767 : n11776;
  assign n11778 = pi18 ? n962 : ~n11109;
  assign n11779 = pi17 ? n32 : n11778;
  assign n11780 = pi16 ? n32 : n11779;
  assign n11781 = pi15 ? n11511 : n11780;
  assign n11782 = pi21 ? n206 : ~n7107;
  assign n11783 = pi20 ? n11782 : ~n32;
  assign n11784 = pi19 ? n32 : n11783;
  assign n11785 = pi18 ? n962 : ~n11784;
  assign n11786 = pi17 ? n32 : n11785;
  assign n11787 = pi16 ? n32 : n11786;
  assign n11788 = pi21 ? n1939 : ~n7500;
  assign n11789 = pi20 ? n11788 : ~n32;
  assign n11790 = pi19 ? n32 : n11789;
  assign n11791 = pi18 ? n962 : ~n11790;
  assign n11792 = pi17 ? n32 : n11791;
  assign n11793 = pi16 ? n32 : n11792;
  assign n11794 = pi15 ? n11787 : n11793;
  assign n11795 = pi14 ? n11781 : n11794;
  assign n11796 = pi13 ? n11777 : n11795;
  assign n11797 = pi19 ? n32 : n6333;
  assign n11798 = pi19 ? n247 : n288;
  assign n11799 = pi18 ? n11797 : ~n11798;
  assign n11800 = pi17 ? n32 : n11799;
  assign n11801 = pi16 ? n32 : n11800;
  assign n11802 = pi18 ? n2622 : ~n11591;
  assign n11803 = pi17 ? n32 : n11802;
  assign n11804 = pi16 ? n32 : n11803;
  assign n11805 = pi15 ? n11801 : n11804;
  assign n11806 = pi18 ? n2622 : ~n697;
  assign n11807 = pi17 ? n32 : n11806;
  assign n11808 = pi16 ? n32 : n11807;
  assign n11809 = pi14 ? n11805 : n11808;
  assign n11810 = pi18 ? n2730 : ~n697;
  assign n11811 = pi17 ? n32 : n11810;
  assign n11812 = pi16 ? n32 : n11811;
  assign n11813 = pi18 ? n2730 : ~n2730;
  assign n11814 = pi17 ? n32 : n11813;
  assign n11815 = pi16 ? n32 : n11814;
  assign n11816 = pi15 ? n11812 : n11815;
  assign n11817 = pi18 ? n697 : ~n2730;
  assign n11818 = pi17 ? n32 : n11817;
  assign n11819 = pi16 ? n32 : n11818;
  assign n11820 = pi15 ? n11815 : n11819;
  assign n11821 = pi14 ? n11816 : n11820;
  assign n11822 = pi13 ? n11809 : n11821;
  assign n11823 = pi12 ? n11796 : n11822;
  assign n11824 = pi19 ? n507 : n1941;
  assign n11825 = pi18 ? n697 : ~n11824;
  assign n11826 = pi17 ? n32 : n11825;
  assign n11827 = pi16 ? n32 : n11826;
  assign n11828 = pi15 ? n11827 : n11819;
  assign n11829 = pi18 ? n697 : ~n697;
  assign n11830 = pi17 ? n32 : n11829;
  assign n11831 = pi16 ? n32 : n11830;
  assign n11832 = pi18 ? n697 : ~n4098;
  assign n11833 = pi17 ? n32 : n11832;
  assign n11834 = pi16 ? n32 : n11833;
  assign n11835 = pi15 ? n11831 : n11834;
  assign n11836 = pi14 ? n11828 : n11835;
  assign n11837 = pi18 ? n697 : ~n595;
  assign n11838 = pi17 ? n32 : n11837;
  assign n11839 = pi16 ? n32 : n11838;
  assign n11840 = pi18 ? n496 : ~n595;
  assign n11841 = pi17 ? n32 : n11840;
  assign n11842 = pi16 ? n32 : n11841;
  assign n11843 = pi15 ? n11842 : n11839;
  assign n11844 = pi14 ? n11839 : n11843;
  assign n11845 = pi13 ? n11836 : n11844;
  assign n11846 = pi18 ? n496 : ~n2747;
  assign n11847 = pi17 ? n32 : n11846;
  assign n11848 = pi16 ? n32 : n11847;
  assign n11849 = pi18 ? n496 : ~n2754;
  assign n11850 = pi17 ? n32 : n11849;
  assign n11851 = pi16 ? n32 : n11850;
  assign n11852 = pi15 ? n11848 : n11851;
  assign n11853 = pi14 ? n11852 : n11851;
  assign n11854 = pi18 ? n496 : ~n797;
  assign n11855 = pi17 ? n32 : n11854;
  assign n11856 = pi16 ? n32 : n11855;
  assign n11857 = pi15 ? n11851 : n11856;
  assign n11858 = pi18 ? n684 : ~n605;
  assign n11859 = pi17 ? n32 : n11858;
  assign n11860 = pi16 ? n32 : n11859;
  assign n11861 = pi18 ? n684 : ~n418;
  assign n11862 = pi17 ? n32 : n11861;
  assign n11863 = pi16 ? n32 : n11862;
  assign n11864 = pi15 ? n11860 : n11863;
  assign n11865 = pi14 ? n11857 : n11864;
  assign n11866 = pi13 ? n11853 : n11865;
  assign n11867 = pi12 ? n11845 : n11866;
  assign n11868 = pi11 ? n11823 : n11867;
  assign n11869 = pi10 ? n11758 : n11868;
  assign n11870 = pi09 ? n11678 : n11869;
  assign n11871 = pi08 ? n11664 : n11870;
  assign n11872 = pi07 ? n11437 : n11871;
  assign n11873 = pi06 ? n10975 : n11872;
  assign n11874 = pi19 ? n1941 : ~n343;
  assign n11875 = pi18 ? n32 : n11874;
  assign n11876 = pi17 ? n32 : n11875;
  assign n11877 = pi16 ? n32 : n11876;
  assign n11878 = pi15 ? n32 : n11877;
  assign n11879 = pi20 ? n266 : ~n207;
  assign n11880 = pi19 ? n1941 : n11879;
  assign n11881 = pi18 ? n32 : n11880;
  assign n11882 = pi17 ? n32 : n11881;
  assign n11883 = pi16 ? n32 : n11882;
  assign n11884 = pi19 ? n236 : ~n531;
  assign n11885 = pi18 ? n32 : n11884;
  assign n11886 = pi17 ? n32 : n11885;
  assign n11887 = pi16 ? n32 : n11886;
  assign n11888 = pi15 ? n11883 : n11887;
  assign n11889 = pi14 ? n11878 : n11888;
  assign n11890 = pi13 ? n32 : n11889;
  assign n11891 = pi12 ? n32 : n11890;
  assign n11892 = pi11 ? n32 : n11891;
  assign n11893 = pi10 ? n32 : n11892;
  assign n11894 = pi19 ? n2614 : n4342;
  assign n11895 = pi18 ? n32 : n11894;
  assign n11896 = pi17 ? n32 : n11895;
  assign n11897 = pi16 ? n32 : n11896;
  assign n11898 = pi15 ? n11887 : n11897;
  assign n11899 = pi20 ? n339 : ~n342;
  assign n11900 = pi19 ? n11899 : n4342;
  assign n11901 = pi18 ? n32 : n11900;
  assign n11902 = pi17 ? n32 : n11901;
  assign n11903 = pi16 ? n32 : n11902;
  assign n11904 = pi18 ? n32 : ~n880;
  assign n11905 = pi17 ? n32 : n11904;
  assign n11906 = pi16 ? n32 : n11905;
  assign n11907 = pi15 ? n11903 : n11906;
  assign n11908 = pi14 ? n11898 : n11907;
  assign n11909 = pi15 ? n11672 : n11445;
  assign n11910 = pi18 ? n1321 : ~n880;
  assign n11911 = pi17 ? n32 : n11910;
  assign n11912 = pi16 ? n32 : n11911;
  assign n11913 = pi14 ? n11909 : n11912;
  assign n11914 = pi13 ? n11908 : n11913;
  assign n11915 = pi18 ? n1592 : ~n2043;
  assign n11916 = pi17 ? n32 : n11915;
  assign n11917 = pi16 ? n32 : n11916;
  assign n11918 = pi18 ? n1592 : ~n1387;
  assign n11919 = pi17 ? n32 : n11918;
  assign n11920 = pi16 ? n32 : n11919;
  assign n11921 = pi15 ? n11917 : n11920;
  assign n11922 = pi20 ? n175 : n321;
  assign n11923 = pi19 ? n32 : n11922;
  assign n11924 = pi18 ? n1841 : ~n11923;
  assign n11925 = pi17 ? n32 : n11924;
  assign n11926 = pi16 ? n32 : n11925;
  assign n11927 = pi15 ? n11926 : n11219;
  assign n11928 = pi14 ? n11921 : n11927;
  assign n11929 = pi20 ? n32 : ~n260;
  assign n11930 = pi19 ? n32 : n11929;
  assign n11931 = pi18 ? n940 : ~n11930;
  assign n11932 = pi17 ? n32 : n11931;
  assign n11933 = pi16 ? n32 : n11932;
  assign n11934 = pi18 ? n1477 : ~n7038;
  assign n11935 = pi17 ? n32 : n11934;
  assign n11936 = pi16 ? n32 : n11935;
  assign n11937 = pi15 ? n11933 : n11936;
  assign n11938 = pi20 ? n32 : ~n125;
  assign n11939 = pi19 ? n32 : n11938;
  assign n11940 = pi18 ? n751 : ~n11939;
  assign n11941 = pi17 ? n32 : n11940;
  assign n11942 = pi16 ? n32 : n11941;
  assign n11943 = pi18 ? n751 : ~n7038;
  assign n11944 = pi17 ? n32 : n11943;
  assign n11945 = pi16 ? n32 : n11944;
  assign n11946 = pi15 ? n11942 : n11945;
  assign n11947 = pi14 ? n11937 : n11946;
  assign n11948 = pi13 ? n11928 : n11947;
  assign n11949 = pi12 ? n11914 : n11948;
  assign n11950 = pi18 ? n751 : ~n6767;
  assign n11951 = pi17 ? n32 : n11950;
  assign n11952 = pi16 ? n32 : n11951;
  assign n11953 = pi18 ? n1970 : ~n1509;
  assign n11954 = pi17 ? n32 : n11953;
  assign n11955 = pi16 ? n32 : n11954;
  assign n11956 = pi15 ? n11952 : n11955;
  assign n11957 = pi14 ? n11956 : n10986;
  assign n11958 = pi14 ? n11705 : n10992;
  assign n11959 = pi13 ? n11957 : n11958;
  assign n11960 = pi20 ? n246 : n1475;
  assign n11961 = pi19 ? n32 : n11960;
  assign n11962 = pi18 ? n341 : ~n11961;
  assign n11963 = pi17 ? n32 : n11962;
  assign n11964 = pi16 ? n32 : n11963;
  assign n11965 = pi18 ? n341 : ~n1054;
  assign n11966 = pi17 ? n32 : n11965;
  assign n11967 = pi16 ? n32 : n11966;
  assign n11968 = pi15 ? n11964 : n11967;
  assign n11969 = pi18 ? n2830 : ~n209;
  assign n11970 = pi17 ? n32 : n11969;
  assign n11971 = pi16 ? n32 : n11970;
  assign n11972 = pi20 ? n32 : n11048;
  assign n11973 = pi19 ? n32 : n11972;
  assign n11974 = pi18 ? n2830 : ~n11973;
  assign n11975 = pi17 ? n32 : n11974;
  assign n11976 = pi16 ? n32 : n11975;
  assign n11977 = pi15 ? n11971 : n11976;
  assign n11978 = pi14 ? n11968 : n11977;
  assign n11979 = pi18 ? n684 : ~n7368;
  assign n11980 = pi17 ? n32 : n11979;
  assign n11981 = pi16 ? n32 : n11980;
  assign n11982 = pi18 ? n684 : ~n1970;
  assign n11983 = pi17 ? n32 : n11982;
  assign n11984 = pi16 ? n32 : n11983;
  assign n11985 = pi15 ? n11981 : n11984;
  assign n11986 = pi20 ? n246 : ~n481;
  assign n11987 = pi19 ? n32 : n11986;
  assign n11988 = pi18 ? n684 : ~n11987;
  assign n11989 = pi17 ? n32 : n11988;
  assign n11990 = pi16 ? n32 : n11989;
  assign n11991 = pi20 ? n32 : ~n481;
  assign n11992 = pi19 ? n32 : n11991;
  assign n11993 = pi18 ? n684 : ~n11992;
  assign n11994 = pi17 ? n32 : n11993;
  assign n11995 = pi16 ? n32 : n11994;
  assign n11996 = pi15 ? n11990 : n11995;
  assign n11997 = pi14 ? n11985 : n11996;
  assign n11998 = pi13 ? n11978 : n11997;
  assign n11999 = pi12 ? n11959 : n11998;
  assign n12000 = pi11 ? n11949 : n11999;
  assign n12001 = pi18 ? n2835 : ~n11992;
  assign n12002 = pi17 ? n32 : n12001;
  assign n12003 = pi16 ? n32 : n12002;
  assign n12004 = pi15 ? n11000 : n12003;
  assign n12005 = pi18 ? n2835 : ~n366;
  assign n12006 = pi17 ? n32 : n12005;
  assign n12007 = pi16 ? n32 : n12006;
  assign n12008 = pi20 ? n7108 : ~n32;
  assign n12009 = pi19 ? n32 : n12008;
  assign n12010 = pi18 ? n590 : ~n12009;
  assign n12011 = pi17 ? n32 : n12010;
  assign n12012 = pi16 ? n32 : n12011;
  assign n12013 = pi15 ? n12007 : n12012;
  assign n12014 = pi14 ? n12004 : n12013;
  assign n12015 = pi18 ? n590 : ~n2962;
  assign n12016 = pi17 ? n32 : n12015;
  assign n12017 = pi16 ? n32 : n12016;
  assign n12018 = pi15 ? n12017 : n11483;
  assign n12019 = pi21 ? n32 : n9326;
  assign n12020 = pi20 ? n12019 : ~n32;
  assign n12021 = pi19 ? n32 : n12020;
  assign n12022 = pi18 ? n590 : ~n12021;
  assign n12023 = pi17 ? n32 : n12022;
  assign n12024 = pi16 ? n32 : n12023;
  assign n12025 = pi18 ? n590 : ~n2830;
  assign n12026 = pi17 ? n32 : n12025;
  assign n12027 = pi16 ? n32 : n12026;
  assign n12028 = pi15 ? n12024 : n12027;
  assign n12029 = pi14 ? n12018 : n12028;
  assign n12030 = pi13 ? n12014 : n12029;
  assign n12031 = pi18 ? n2730 : ~n590;
  assign n12032 = pi17 ? n32 : n12031;
  assign n12033 = pi16 ? n32 : n12032;
  assign n12034 = pi18 ? n2849 : ~n590;
  assign n12035 = pi17 ? n32 : n12034;
  assign n12036 = pi16 ? n32 : n12035;
  assign n12037 = pi15 ? n12033 : n12036;
  assign n12038 = pi18 ? n2849 : ~n2730;
  assign n12039 = pi17 ? n32 : n12038;
  assign n12040 = pi16 ? n32 : n12039;
  assign n12041 = pi15 ? n12040 : n12036;
  assign n12042 = pi14 ? n12037 : n12041;
  assign n12043 = pi18 ? n2849 : ~n496;
  assign n12044 = pi17 ? n32 : n12043;
  assign n12045 = pi16 ? n32 : n12044;
  assign n12046 = pi15 ? n12045 : n12040;
  assign n12047 = pi18 ? n496 : ~n2730;
  assign n12048 = pi17 ? n32 : n12047;
  assign n12049 = pi16 ? n32 : n12048;
  assign n12050 = pi15 ? n12040 : n12049;
  assign n12051 = pi14 ? n12046 : n12050;
  assign n12052 = pi13 ? n12042 : n12051;
  assign n12053 = pi12 ? n12030 : n12052;
  assign n12054 = pi18 ? n496 : ~n697;
  assign n12055 = pi17 ? n32 : n12054;
  assign n12056 = pi16 ? n32 : n12055;
  assign n12057 = pi18 ? n684 : ~n4098;
  assign n12058 = pi17 ? n32 : n12057;
  assign n12059 = pi16 ? n32 : n12058;
  assign n12060 = pi15 ? n12056 : n12059;
  assign n12061 = pi14 ? n12049 : n12060;
  assign n12062 = pi21 ? n32 : n7478;
  assign n12063 = pi20 ? n32 : n12062;
  assign n12064 = pi19 ? n12063 : ~n32;
  assign n12065 = pi18 ? n684 : ~n12064;
  assign n12066 = pi17 ? n32 : n12065;
  assign n12067 = pi16 ? n32 : n12066;
  assign n12068 = pi18 ? n684 : ~n595;
  assign n12069 = pi17 ? n32 : n12068;
  assign n12070 = pi16 ? n32 : n12069;
  assign n12071 = pi15 ? n12067 : n12070;
  assign n12072 = pi14 ? n12059 : n12071;
  assign n12073 = pi13 ? n12061 : n12072;
  assign n12074 = pi18 ? n684 : ~n520;
  assign n12075 = pi17 ? n32 : n12074;
  assign n12076 = pi16 ? n32 : n12075;
  assign n12077 = pi18 ? n684 : ~n2754;
  assign n12078 = pi17 ? n32 : n12077;
  assign n12079 = pi16 ? n32 : n12078;
  assign n12080 = pi15 ? n12076 : n12079;
  assign n12081 = pi18 ? n880 : ~n2754;
  assign n12082 = pi17 ? n32 : n12081;
  assign n12083 = pi16 ? n32 : n12082;
  assign n12084 = pi15 ? n12079 : n12083;
  assign n12085 = pi14 ? n12080 : n12084;
  assign n12086 = pi18 ? n684 : ~n797;
  assign n12087 = pi17 ? n32 : n12086;
  assign n12088 = pi16 ? n32 : n12087;
  assign n12089 = pi18 ? n880 : ~n2413;
  assign n12090 = pi17 ? n32 : n12089;
  assign n12091 = pi16 ? n32 : n12090;
  assign n12092 = pi15 ? n12088 : n12091;
  assign n12093 = pi18 ? n880 : ~n605;
  assign n12094 = pi17 ? n32 : n12093;
  assign n12095 = pi16 ? n32 : n12094;
  assign n12096 = pi18 ? n880 : ~n418;
  assign n12097 = pi17 ? n32 : n12096;
  assign n12098 = pi16 ? n32 : n12097;
  assign n12099 = pi15 ? n12095 : n12098;
  assign n12100 = pi14 ? n12092 : n12099;
  assign n12101 = pi13 ? n12085 : n12100;
  assign n12102 = pi12 ? n12073 : n12101;
  assign n12103 = pi11 ? n12053 : n12102;
  assign n12104 = pi10 ? n12000 : n12103;
  assign n12105 = pi09 ? n11893 : n12104;
  assign n12106 = pi19 ? n2848 : ~n343;
  assign n12107 = pi18 ? n32 : n12106;
  assign n12108 = pi17 ? n32 : n12107;
  assign n12109 = pi16 ? n32 : n12108;
  assign n12110 = pi15 ? n32 : n12109;
  assign n12111 = pi19 ? n2848 : n11879;
  assign n12112 = pi18 ? n32 : n12111;
  assign n12113 = pi17 ? n32 : n12112;
  assign n12114 = pi16 ? n32 : n12113;
  assign n12115 = pi18 ? n32 : n6181;
  assign n12116 = pi17 ? n32 : n12115;
  assign n12117 = pi16 ? n32 : n12116;
  assign n12118 = pi15 ? n12114 : n12117;
  assign n12119 = pi14 ? n12110 : n12118;
  assign n12120 = pi13 ? n32 : n12119;
  assign n12121 = pi12 ? n32 : n12120;
  assign n12122 = pi11 ? n32 : n12121;
  assign n12123 = pi10 ? n32 : n12122;
  assign n12124 = pi19 ? n813 : n4342;
  assign n12125 = pi18 ? n32 : n12124;
  assign n12126 = pi17 ? n32 : n12125;
  assign n12127 = pi16 ? n32 : n12126;
  assign n12128 = pi15 ? n12117 : n12127;
  assign n12129 = pi19 ? n7667 : n4342;
  assign n12130 = pi18 ? n32 : n12129;
  assign n12131 = pi17 ? n32 : n12130;
  assign n12132 = pi16 ? n32 : n12131;
  assign n12133 = pi15 ? n12132 : n11887;
  assign n12134 = pi14 ? n12128 : n12133;
  assign n12135 = pi19 ? n236 : ~n322;
  assign n12136 = pi18 ? n32 : n12135;
  assign n12137 = pi17 ? n32 : n12136;
  assign n12138 = pi16 ? n32 : n12137;
  assign n12139 = pi15 ? n12138 : n11672;
  assign n12140 = pi14 ? n12139 : n11685;
  assign n12141 = pi13 ? n12134 : n12140;
  assign n12142 = pi18 ? n1575 : ~n2043;
  assign n12143 = pi17 ? n32 : n12142;
  assign n12144 = pi16 ? n32 : n12143;
  assign n12145 = pi18 ? n1575 : ~n1387;
  assign n12146 = pi17 ? n32 : n12145;
  assign n12147 = pi16 ? n32 : n12146;
  assign n12148 = pi15 ? n12144 : n12147;
  assign n12149 = pi18 ? n2142 : ~n11923;
  assign n12150 = pi17 ? n32 : n12149;
  assign n12151 = pi16 ? n32 : n12150;
  assign n12152 = pi15 ? n12151 : n11445;
  assign n12153 = pi14 ? n12148 : n12152;
  assign n12154 = pi18 ? n863 : ~n9002;
  assign n12155 = pi17 ? n32 : n12154;
  assign n12156 = pi16 ? n32 : n12155;
  assign n12157 = pi18 ? n1321 : ~n9904;
  assign n12158 = pi17 ? n32 : n12157;
  assign n12159 = pi16 ? n32 : n12158;
  assign n12160 = pi15 ? n12156 : n12159;
  assign n12161 = pi18 ? n1592 : ~n9904;
  assign n12162 = pi17 ? n32 : n12161;
  assign n12163 = pi16 ? n32 : n12162;
  assign n12164 = pi15 ? n11912 : n12163;
  assign n12165 = pi14 ? n12160 : n12164;
  assign n12166 = pi13 ? n12153 : n12165;
  assign n12167 = pi12 ? n12141 : n12166;
  assign n12168 = pi18 ? n1592 : ~n6767;
  assign n12169 = pi17 ? n32 : n12168;
  assign n12170 = pi16 ? n32 : n12169;
  assign n12171 = pi20 ? n32 : n10066;
  assign n12172 = pi19 ? n32 : n12171;
  assign n12173 = pi18 ? n1841 : ~n12172;
  assign n12174 = pi17 ? n32 : n12173;
  assign n12175 = pi16 ? n32 : n12174;
  assign n12176 = pi15 ? n12170 : n12175;
  assign n12177 = pi14 ? n12176 : n11223;
  assign n12178 = pi15 ? n11696 : n11700;
  assign n12179 = pi14 ? n12178 : n11231;
  assign n12180 = pi13 ? n12177 : n12179;
  assign n12181 = pi18 ? n751 : ~n7814;
  assign n12182 = pi17 ? n32 : n12181;
  assign n12183 = pi16 ? n32 : n12182;
  assign n12184 = pi18 ? n751 : ~n1054;
  assign n12185 = pi17 ? n32 : n12184;
  assign n12186 = pi16 ? n32 : n12185;
  assign n12187 = pi15 ? n12183 : n12186;
  assign n12188 = pi18 ? n1970 : ~n209;
  assign n12189 = pi17 ? n32 : n12188;
  assign n12190 = pi16 ? n32 : n12189;
  assign n12191 = pi20 ? n101 : n11048;
  assign n12192 = pi19 ? n32 : n12191;
  assign n12193 = pi18 ? n1970 : ~n12192;
  assign n12194 = pi17 ? n32 : n12193;
  assign n12195 = pi16 ? n32 : n12194;
  assign n12196 = pi15 ? n12190 : n12195;
  assign n12197 = pi14 ? n12187 : n12196;
  assign n12198 = pi18 ? n209 : ~n7368;
  assign n12199 = pi17 ? n32 : n12198;
  assign n12200 = pi16 ? n32 : n12199;
  assign n12201 = pi18 ? n209 : ~n245;
  assign n12202 = pi17 ? n32 : n12201;
  assign n12203 = pi16 ? n32 : n12202;
  assign n12204 = pi15 ? n12200 : n12203;
  assign n12205 = pi18 ? n209 : ~n7038;
  assign n12206 = pi17 ? n32 : n12205;
  assign n12207 = pi16 ? n32 : n12206;
  assign n12208 = pi15 ? n12207 : n11463;
  assign n12209 = pi14 ? n12204 : n12208;
  assign n12210 = pi13 ? n12197 : n12209;
  assign n12211 = pi12 ? n12180 : n12210;
  assign n12212 = pi11 ? n12167 : n12211;
  assign n12213 = pi18 ? n2962 : ~n880;
  assign n12214 = pi17 ? n32 : n12213;
  assign n12215 = pi16 ? n32 : n12214;
  assign n12216 = pi15 ? n11463 : n12215;
  assign n12217 = pi18 ? n2962 : ~n2962;
  assign n12218 = pi17 ? n32 : n12217;
  assign n12219 = pi16 ? n32 : n12218;
  assign n12220 = pi18 ? n1965 : ~n12009;
  assign n12221 = pi17 ? n32 : n12220;
  assign n12222 = pi16 ? n32 : n12221;
  assign n12223 = pi15 ? n12219 : n12222;
  assign n12224 = pi14 ? n12216 : n12223;
  assign n12225 = pi18 ? n1965 : ~n2962;
  assign n12226 = pi17 ? n32 : n12225;
  assign n12227 = pi16 ? n32 : n12226;
  assign n12228 = pi18 ? n1965 : ~n1965;
  assign n12229 = pi17 ? n32 : n12228;
  assign n12230 = pi16 ? n32 : n12229;
  assign n12231 = pi15 ? n12227 : n12230;
  assign n12232 = pi18 ? n1965 : ~n684;
  assign n12233 = pi17 ? n32 : n12232;
  assign n12234 = pi16 ? n32 : n12233;
  assign n12235 = pi18 ? n1965 : ~n590;
  assign n12236 = pi17 ? n32 : n12235;
  assign n12237 = pi16 ? n32 : n12236;
  assign n12238 = pi15 ? n12234 : n12237;
  assign n12239 = pi14 ? n12231 : n12238;
  assign n12240 = pi13 ? n12224 : n12239;
  assign n12241 = pi18 ? n2830 : ~n590;
  assign n12242 = pi17 ? n32 : n12241;
  assign n12243 = pi16 ? n32 : n12242;
  assign n12244 = pi21 ? n66 : ~n32;
  assign n12245 = pi20 ? n12244 : ~n32;
  assign n12246 = pi19 ? n32 : n12245;
  assign n12247 = pi18 ? n2830 : ~n12246;
  assign n12248 = pi17 ? n32 : n12247;
  assign n12249 = pi16 ? n32 : n12248;
  assign n12250 = pi15 ? n12249 : n12243;
  assign n12251 = pi14 ? n12243 : n12250;
  assign n12252 = pi18 ? n2830 : ~n2849;
  assign n12253 = pi17 ? n32 : n12252;
  assign n12254 = pi16 ? n32 : n12253;
  assign n12255 = pi18 ? n2830 : ~n2730;
  assign n12256 = pi17 ? n32 : n12255;
  assign n12257 = pi16 ? n32 : n12256;
  assign n12258 = pi15 ? n12254 : n12257;
  assign n12259 = pi18 ? n684 : ~n697;
  assign n12260 = pi17 ? n32 : n12259;
  assign n12261 = pi16 ? n32 : n12260;
  assign n12262 = pi15 ? n12257 : n12261;
  assign n12263 = pi14 ? n12258 : n12262;
  assign n12264 = pi13 ? n12251 : n12263;
  assign n12265 = pi12 ? n12240 : n12264;
  assign n12266 = pi18 ? n880 : ~n2622;
  assign n12267 = pi17 ? n32 : n12266;
  assign n12268 = pi16 ? n32 : n12267;
  assign n12269 = pi18 ? n880 : ~n4098;
  assign n12270 = pi17 ? n32 : n12269;
  assign n12271 = pi16 ? n32 : n12270;
  assign n12272 = pi15 ? n12268 : n12271;
  assign n12273 = pi14 ? n12261 : n12272;
  assign n12274 = pi22 ? n50 : n34;
  assign n12275 = pi21 ? n32 : n12274;
  assign n12276 = pi20 ? n32 : n12275;
  assign n12277 = pi19 ? n12276 : ~n32;
  assign n12278 = pi18 ? n880 : ~n12277;
  assign n12279 = pi17 ? n32 : n12278;
  assign n12280 = pi16 ? n32 : n12279;
  assign n12281 = pi18 ? n880 : ~n508;
  assign n12282 = pi17 ? n32 : n12281;
  assign n12283 = pi16 ? n32 : n12282;
  assign n12284 = pi15 ? n12280 : n12283;
  assign n12285 = pi14 ? n12271 : n12284;
  assign n12286 = pi13 ? n12273 : n12285;
  assign n12287 = pi18 ? n880 : ~n520;
  assign n12288 = pi17 ? n32 : n12287;
  assign n12289 = pi16 ? n32 : n12288;
  assign n12290 = pi15 ? n12289 : n12083;
  assign n12291 = pi18 ? n209 : ~n2754;
  assign n12292 = pi17 ? n32 : n12291;
  assign n12293 = pi16 ? n32 : n12292;
  assign n12294 = pi14 ? n12290 : n12293;
  assign n12295 = pi18 ? n209 : ~n797;
  assign n12296 = pi17 ? n32 : n12295;
  assign n12297 = pi16 ? n32 : n12296;
  assign n12298 = pi18 ? n209 : ~n2413;
  assign n12299 = pi17 ? n32 : n12298;
  assign n12300 = pi16 ? n32 : n12299;
  assign n12301 = pi15 ? n12297 : n12300;
  assign n12302 = pi18 ? n209 : ~n605;
  assign n12303 = pi17 ? n32 : n12302;
  assign n12304 = pi16 ? n32 : n12303;
  assign n12305 = pi18 ? n209 : ~n3786;
  assign n12306 = pi17 ? n32 : n12305;
  assign n12307 = pi16 ? n32 : n12306;
  assign n12308 = pi15 ? n12304 : n12307;
  assign n12309 = pi14 ? n12301 : n12308;
  assign n12310 = pi13 ? n12294 : n12309;
  assign n12311 = pi12 ? n12286 : n12310;
  assign n12312 = pi11 ? n12265 : n12311;
  assign n12313 = pi10 ? n12212 : n12312;
  assign n12314 = pi09 ? n12123 : n12313;
  assign n12315 = pi08 ? n12105 : n12314;
  assign n12316 = pi19 ? n2303 : ~n349;
  assign n12317 = pi18 ? n32 : n12316;
  assign n12318 = pi17 ? n32 : n12317;
  assign n12319 = pi16 ? n32 : n12318;
  assign n12320 = pi15 ? n32 : n12319;
  assign n12321 = pi19 ? n2303 : n1757;
  assign n12322 = pi18 ? n32 : n12321;
  assign n12323 = pi17 ? n32 : n12322;
  assign n12324 = pi16 ? n32 : n12323;
  assign n12325 = pi19 ? n2317 : ~n531;
  assign n12326 = pi18 ? n32 : n12325;
  assign n12327 = pi17 ? n32 : n12326;
  assign n12328 = pi16 ? n32 : n12327;
  assign n12329 = pi15 ? n12324 : n12328;
  assign n12330 = pi14 ? n12320 : n12329;
  assign n12331 = pi13 ? n32 : n12330;
  assign n12332 = pi12 ? n32 : n12331;
  assign n12333 = pi11 ? n32 : n12332;
  assign n12334 = pi10 ? n32 : n12333;
  assign n12335 = pi20 ? n1839 : ~n11107;
  assign n12336 = pi19 ? n12335 : n4342;
  assign n12337 = pi18 ? n32 : n12336;
  assign n12338 = pi17 ? n32 : n12337;
  assign n12339 = pi16 ? n32 : n12338;
  assign n12340 = pi15 ? n12328 : n12339;
  assign n12341 = pi19 ? n6158 : n4342;
  assign n12342 = pi18 ? n32 : n12341;
  assign n12343 = pi17 ? n32 : n12342;
  assign n12344 = pi16 ? n32 : n12343;
  assign n12345 = pi15 ? n12344 : n12117;
  assign n12346 = pi14 ? n12340 : n12345;
  assign n12347 = pi19 ? n236 : ~n11922;
  assign n12348 = pi18 ? n32 : n12347;
  assign n12349 = pi17 ? n32 : n12348;
  assign n12350 = pi16 ? n32 : n12349;
  assign n12351 = pi15 ? n12138 : n12350;
  assign n12352 = pi19 ? n2614 : ~n531;
  assign n12353 = pi18 ? n32 : n12352;
  assign n12354 = pi17 ? n32 : n12353;
  assign n12355 = pi16 ? n32 : n12354;
  assign n12356 = pi14 ? n12351 : n12355;
  assign n12357 = pi13 ? n12346 : n12356;
  assign n12358 = pi19 ? n2614 : ~n343;
  assign n12359 = pi18 ? n32 : n12358;
  assign n12360 = pi17 ? n32 : n12359;
  assign n12361 = pi16 ? n32 : n12360;
  assign n12362 = pi20 ? n339 : ~n1611;
  assign n12363 = pi19 ? n12362 : n4670;
  assign n12364 = pi18 ? n32 : n12363;
  assign n12365 = pi17 ? n32 : n12364;
  assign n12366 = pi16 ? n32 : n12365;
  assign n12367 = pi15 ? n12361 : n12366;
  assign n12368 = pi19 ? n32 : n1490;
  assign n12369 = pi18 ? n32 : ~n12368;
  assign n12370 = pi17 ? n32 : n12369;
  assign n12371 = pi16 ? n32 : n12370;
  assign n12372 = pi14 ? n12367 : n12371;
  assign n12373 = pi20 ? n175 : ~n9000;
  assign n12374 = pi19 ? n32 : n12373;
  assign n12375 = pi18 ? n32 : ~n12374;
  assign n12376 = pi17 ? n32 : n12375;
  assign n12377 = pi16 ? n32 : n12376;
  assign n12378 = pi18 ? n1575 : ~n9904;
  assign n12379 = pi17 ? n32 : n12378;
  assign n12380 = pi16 ? n32 : n12379;
  assign n12381 = pi15 ? n12377 : n12380;
  assign n12382 = pi15 ? n11685 : n12380;
  assign n12383 = pi14 ? n12381 : n12382;
  assign n12384 = pi13 ? n12372 : n12383;
  assign n12385 = pi12 ? n12357 : n12384;
  assign n12386 = pi18 ? n2142 : ~n11930;
  assign n12387 = pi17 ? n32 : n12386;
  assign n12388 = pi16 ? n32 : n12387;
  assign n12389 = pi15 ? n12380 : n12388;
  assign n12390 = pi18 ? n863 : ~n11923;
  assign n12391 = pi17 ? n32 : n12390;
  assign n12392 = pi16 ? n32 : n12391;
  assign n12393 = pi15 ? n12392 : n11445;
  assign n12394 = pi14 ? n12389 : n12393;
  assign n12395 = pi18 ? n863 : ~n2043;
  assign n12396 = pi17 ? n32 : n12395;
  assign n12397 = pi16 ? n32 : n12396;
  assign n12398 = pi18 ? n863 : ~n10095;
  assign n12399 = pi17 ? n32 : n12398;
  assign n12400 = pi16 ? n32 : n12399;
  assign n12401 = pi15 ? n12397 : n12400;
  assign n12402 = pi18 ? n1321 : ~n11923;
  assign n12403 = pi17 ? n32 : n12402;
  assign n12404 = pi16 ? n32 : n12403;
  assign n12405 = pi20 ? n175 : n1839;
  assign n12406 = pi19 ? n32 : n12405;
  assign n12407 = pi18 ? n1321 : ~n12406;
  assign n12408 = pi17 ? n32 : n12407;
  assign n12409 = pi16 ? n32 : n12408;
  assign n12410 = pi15 ? n12404 : n12409;
  assign n12411 = pi14 ? n12401 : n12410;
  assign n12412 = pi13 ? n12394 : n12411;
  assign n12413 = pi18 ? n1592 : ~n9598;
  assign n12414 = pi17 ? n32 : n12413;
  assign n12415 = pi16 ? n32 : n12414;
  assign n12416 = pi20 ? n9641 : ~n6229;
  assign n12417 = pi19 ? n32 : n12416;
  assign n12418 = pi18 ? n1592 : ~n12417;
  assign n12419 = pi17 ? n32 : n12418;
  assign n12420 = pi16 ? n32 : n12419;
  assign n12421 = pi15 ? n12415 : n12420;
  assign n12422 = pi18 ? n1841 : ~n751;
  assign n12423 = pi17 ? n32 : n12422;
  assign n12424 = pi16 ? n32 : n12423;
  assign n12425 = pi20 ? n428 : n1475;
  assign n12426 = pi19 ? n32 : n12425;
  assign n12427 = pi18 ? n1841 : ~n12426;
  assign n12428 = pi17 ? n32 : n12427;
  assign n12429 = pi16 ? n32 : n12428;
  assign n12430 = pi15 ? n12424 : n12429;
  assign n12431 = pi14 ? n12421 : n12430;
  assign n12432 = pi18 ? n940 : ~n8804;
  assign n12433 = pi17 ? n32 : n12432;
  assign n12434 = pi16 ? n32 : n12433;
  assign n12435 = pi20 ? n175 : n339;
  assign n12436 = pi19 ? n32 : n12435;
  assign n12437 = pi18 ? n940 : ~n12436;
  assign n12438 = pi17 ? n32 : n12437;
  assign n12439 = pi16 ? n32 : n12438;
  assign n12440 = pi15 ? n12434 : n12439;
  assign n12441 = pi18 ? n940 : ~n496;
  assign n12442 = pi17 ? n32 : n12441;
  assign n12443 = pi16 ? n32 : n12442;
  assign n12444 = pi18 ? n940 : ~n341;
  assign n12445 = pi17 ? n32 : n12444;
  assign n12446 = pi16 ? n32 : n12445;
  assign n12447 = pi15 ? n12443 : n12446;
  assign n12448 = pi14 ? n12440 : n12447;
  assign n12449 = pi13 ? n12431 : n12448;
  assign n12450 = pi12 ? n12412 : n12449;
  assign n12451 = pi11 ? n12385 : n12450;
  assign n12452 = pi18 ? n940 : ~n245;
  assign n12453 = pi17 ? n32 : n12452;
  assign n12454 = pi16 ? n32 : n12453;
  assign n12455 = pi18 ? n1477 : ~n341;
  assign n12456 = pi17 ? n32 : n12455;
  assign n12457 = pi16 ? n32 : n12456;
  assign n12458 = pi15 ? n12454 : n12457;
  assign n12459 = pi18 ? n1477 : ~n684;
  assign n12460 = pi17 ? n32 : n12459;
  assign n12461 = pi16 ? n32 : n12460;
  assign n12462 = pi18 ? n751 : ~n496;
  assign n12463 = pi17 ? n32 : n12462;
  assign n12464 = pi16 ? n32 : n12463;
  assign n12465 = pi15 ? n12461 : n12464;
  assign n12466 = pi14 ? n12458 : n12465;
  assign n12467 = pi18 ? n751 : ~n684;
  assign n12468 = pi17 ? n32 : n12467;
  assign n12469 = pi16 ? n32 : n12468;
  assign n12470 = pi18 ? n751 : ~n1965;
  assign n12471 = pi17 ? n32 : n12470;
  assign n12472 = pi16 ? n32 : n12471;
  assign n12473 = pi15 ? n12469 : n12472;
  assign n12474 = pi15 ? n12472 : n12464;
  assign n12475 = pi14 ? n12473 : n12474;
  assign n12476 = pi13 ? n12466 : n12475;
  assign n12477 = pi16 ? n32 : n960;
  assign n12478 = pi18 ? n366 : ~n10891;
  assign n12479 = pi17 ? n32 : n12478;
  assign n12480 = pi16 ? n32 : n12479;
  assign n12481 = pi16 ? n32 : n1881;
  assign n12482 = pi15 ? n12480 : n12481;
  assign n12483 = pi14 ? n12477 : n12482;
  assign n12484 = pi18 ? n366 : ~n2849;
  assign n12485 = pi17 ? n32 : n12484;
  assign n12486 = pi16 ? n32 : n12485;
  assign n12487 = pi16 ? n32 : n893;
  assign n12488 = pi15 ? n12486 : n12487;
  assign n12489 = pi18 ? n1970 : ~n2730;
  assign n12490 = pi17 ? n32 : n12489;
  assign n12491 = pi16 ? n32 : n12490;
  assign n12492 = pi19 ? n1574 : n236;
  assign n12493 = pi18 ? n366 : ~n12492;
  assign n12494 = pi17 ? n32 : n12493;
  assign n12495 = pi16 ? n32 : n12494;
  assign n12496 = pi15 ? n12491 : n12495;
  assign n12497 = pi14 ? n12488 : n12496;
  assign n12498 = pi13 ? n12483 : n12497;
  assign n12499 = pi12 ? n12476 : n12498;
  assign n12500 = pi18 ? n209 : ~n2730;
  assign n12501 = pi17 ? n32 : n12500;
  assign n12502 = pi16 ? n32 : n12501;
  assign n12503 = pi18 ? n209 : ~n697;
  assign n12504 = pi17 ? n32 : n12503;
  assign n12505 = pi16 ? n32 : n12504;
  assign n12506 = pi15 ? n12502 : n12505;
  assign n12507 = pi18 ? n209 : ~n2622;
  assign n12508 = pi17 ? n32 : n12507;
  assign n12509 = pi16 ? n32 : n12508;
  assign n12510 = pi18 ? n209 : ~n4098;
  assign n12511 = pi17 ? n32 : n12510;
  assign n12512 = pi16 ? n32 : n12511;
  assign n12513 = pi15 ? n12509 : n12512;
  assign n12514 = pi14 ? n12506 : n12513;
  assign n12515 = pi16 ? n32 : n1257;
  assign n12516 = pi18 ? n209 : ~n2747;
  assign n12517 = pi17 ? n32 : n12516;
  assign n12518 = pi16 ? n32 : n12517;
  assign n12519 = pi15 ? n12515 : n12518;
  assign n12520 = pi14 ? n12512 : n12519;
  assign n12521 = pi13 ? n12514 : n12520;
  assign n12522 = pi18 ? n940 : ~n2747;
  assign n12523 = pi17 ? n32 : n12522;
  assign n12524 = pi16 ? n32 : n12523;
  assign n12525 = pi18 ? n940 : ~n2754;
  assign n12526 = pi17 ? n32 : n12525;
  assign n12527 = pi16 ? n32 : n12526;
  assign n12528 = pi15 ? n12524 : n12527;
  assign n12529 = pi18 ? n940 : ~n797;
  assign n12530 = pi17 ? n32 : n12529;
  assign n12531 = pi16 ? n32 : n12530;
  assign n12532 = pi14 ? n12528 : n12531;
  assign n12533 = pi18 ? n940 : ~n2413;
  assign n12534 = pi17 ? n32 : n12533;
  assign n12535 = pi16 ? n32 : n12534;
  assign n12536 = pi18 ? n940 : ~n605;
  assign n12537 = pi17 ? n32 : n12536;
  assign n12538 = pi16 ? n32 : n12537;
  assign n12539 = pi15 ? n12535 : n12538;
  assign n12540 = pi18 ? n863 : ~n532;
  assign n12541 = pi17 ? n32 : n12540;
  assign n12542 = pi16 ? n32 : n12541;
  assign n12543 = pi18 ? n863 : ~n430;
  assign n12544 = pi17 ? n32 : n12543;
  assign n12545 = pi16 ? n32 : n12544;
  assign n12546 = pi15 ? n12542 : n12545;
  assign n12547 = pi14 ? n12539 : n12546;
  assign n12548 = pi13 ? n12532 : n12547;
  assign n12549 = pi12 ? n12521 : n12548;
  assign n12550 = pi11 ? n12499 : n12549;
  assign n12551 = pi10 ? n12451 : n12550;
  assign n12552 = pi09 ? n12334 : n12551;
  assign n12553 = pi19 ? n429 : ~n349;
  assign n12554 = pi18 ? n32 : n12553;
  assign n12555 = pi17 ? n32 : n12554;
  assign n12556 = pi16 ? n32 : n12555;
  assign n12557 = pi15 ? n32 : n12556;
  assign n12558 = pi19 ? n429 : n1757;
  assign n12559 = pi18 ? n32 : n12558;
  assign n12560 = pi17 ? n32 : n12559;
  assign n12561 = pi16 ? n32 : n12560;
  assign n12562 = pi19 ? n429 : ~n531;
  assign n12563 = pi18 ? n32 : n12562;
  assign n12564 = pi17 ? n32 : n12563;
  assign n12565 = pi16 ? n32 : n12564;
  assign n12566 = pi15 ? n12561 : n12565;
  assign n12567 = pi14 ? n12557 : n12566;
  assign n12568 = pi13 ? n32 : n12567;
  assign n12569 = pi12 ? n32 : n12568;
  assign n12570 = pi11 ? n32 : n12569;
  assign n12571 = pi10 ? n32 : n12570;
  assign n12572 = pi20 ? n342 : ~n11107;
  assign n12573 = pi19 ? n12572 : n4342;
  assign n12574 = pi18 ? n32 : n12573;
  assign n12575 = pi17 ? n32 : n12574;
  assign n12576 = pi16 ? n32 : n12575;
  assign n12577 = pi15 ? n12565 : n12576;
  assign n12578 = pi20 ? n342 : ~n428;
  assign n12579 = pi19 ? n12578 : n4342;
  assign n12580 = pi18 ? n32 : n12579;
  assign n12581 = pi17 ? n32 : n12580;
  assign n12582 = pi16 ? n32 : n12581;
  assign n12583 = pi19 ? n343 : ~n531;
  assign n12584 = pi18 ? n32 : n12583;
  assign n12585 = pi17 ? n32 : n12584;
  assign n12586 = pi16 ? n32 : n12585;
  assign n12587 = pi15 ? n12582 : n12586;
  assign n12588 = pi14 ? n12577 : n12587;
  assign n12589 = pi19 ? n349 : ~n322;
  assign n12590 = pi18 ? n32 : n12589;
  assign n12591 = pi17 ? n32 : n12590;
  assign n12592 = pi16 ? n32 : n12591;
  assign n12593 = pi19 ? n349 : ~n11922;
  assign n12594 = pi18 ? n32 : n12593;
  assign n12595 = pi17 ? n32 : n12594;
  assign n12596 = pi16 ? n32 : n12595;
  assign n12597 = pi15 ? n12592 : n12596;
  assign n12598 = pi19 ? n1812 : ~n531;
  assign n12599 = pi18 ? n32 : n12598;
  assign n12600 = pi17 ? n32 : n12599;
  assign n12601 = pi16 ? n32 : n12600;
  assign n12602 = pi14 ? n12597 : n12601;
  assign n12603 = pi13 ? n12588 : n12602;
  assign n12604 = pi19 ? n813 : ~n343;
  assign n12605 = pi18 ? n32 : n12604;
  assign n12606 = pi17 ? n32 : n12605;
  assign n12607 = pi16 ? n32 : n12606;
  assign n12608 = pi20 ? n1940 : ~n1611;
  assign n12609 = pi19 ? n12608 : n4670;
  assign n12610 = pi18 ? n32 : n12609;
  assign n12611 = pi17 ? n32 : n12610;
  assign n12612 = pi16 ? n32 : n12611;
  assign n12613 = pi15 ? n12607 : n12612;
  assign n12614 = pi19 ? n236 : ~n1490;
  assign n12615 = pi18 ? n32 : n12614;
  assign n12616 = pi17 ? n32 : n12615;
  assign n12617 = pi16 ? n32 : n12616;
  assign n12618 = pi14 ? n12613 : n12617;
  assign n12619 = pi19 ? n236 : ~n12373;
  assign n12620 = pi18 ? n32 : n12619;
  assign n12621 = pi17 ? n32 : n12620;
  assign n12622 = pi16 ? n32 : n12621;
  assign n12623 = pi19 ? n2614 : ~n6298;
  assign n12624 = pi18 ? n32 : n12623;
  assign n12625 = pi17 ? n32 : n12624;
  assign n12626 = pi16 ? n32 : n12625;
  assign n12627 = pi15 ? n12622 : n12626;
  assign n12628 = pi15 ? n12355 : n12626;
  assign n12629 = pi14 ? n12627 : n12628;
  assign n12630 = pi13 ? n12618 : n12629;
  assign n12631 = pi12 ? n12603 : n12630;
  assign n12632 = pi19 ? n617 : ~n9903;
  assign n12633 = pi18 ? n32 : n12632;
  assign n12634 = pi17 ? n32 : n12633;
  assign n12635 = pi16 ? n32 : n12634;
  assign n12636 = pi18 ? n32 : ~n863;
  assign n12637 = pi17 ? n32 : n12636;
  assign n12638 = pi16 ? n32 : n12637;
  assign n12639 = pi15 ? n12635 : n12638;
  assign n12640 = pi15 ? n12371 : n11672;
  assign n12641 = pi14 ? n12639 : n12640;
  assign n12642 = pi18 ? n32 : ~n2043;
  assign n12643 = pi17 ? n32 : n12642;
  assign n12644 = pi16 ? n32 : n12643;
  assign n12645 = pi18 ? n32 : ~n10095;
  assign n12646 = pi17 ? n32 : n12645;
  assign n12647 = pi16 ? n32 : n12646;
  assign n12648 = pi15 ? n12644 : n12647;
  assign n12649 = pi18 ? n32 : ~n12406;
  assign n12650 = pi17 ? n32 : n12649;
  assign n12651 = pi16 ? n32 : n12650;
  assign n12652 = pi14 ? n12648 : n12651;
  assign n12653 = pi13 ? n12641 : n12652;
  assign n12654 = pi18 ? n936 : ~n9598;
  assign n12655 = pi17 ? n32 : n12654;
  assign n12656 = pi16 ? n32 : n12655;
  assign n12657 = pi20 ? n321 : ~n6229;
  assign n12658 = pi19 ? n32 : n12657;
  assign n12659 = pi18 ? n2142 : ~n12658;
  assign n12660 = pi17 ? n32 : n12659;
  assign n12661 = pi16 ? n32 : n12660;
  assign n12662 = pi15 ? n12656 : n12661;
  assign n12663 = pi18 ? n2142 : ~n1477;
  assign n12664 = pi17 ? n32 : n12663;
  assign n12665 = pi16 ? n32 : n12664;
  assign n12666 = pi20 ? n175 : n1475;
  assign n12667 = pi19 ? n32 : n12666;
  assign n12668 = pi18 ? n2142 : ~n12667;
  assign n12669 = pi17 ? n32 : n12668;
  assign n12670 = pi16 ? n32 : n12669;
  assign n12671 = pi15 ? n12665 : n12670;
  assign n12672 = pi14 ? n12662 : n12671;
  assign n12673 = pi18 ? n2142 : ~n8804;
  assign n12674 = pi17 ? n32 : n12673;
  assign n12675 = pi16 ? n32 : n12674;
  assign n12676 = pi18 ? n863 : ~n12436;
  assign n12677 = pi17 ? n32 : n12676;
  assign n12678 = pi16 ? n32 : n12677;
  assign n12679 = pi15 ? n12675 : n12678;
  assign n12680 = pi20 ? n321 : ~n481;
  assign n12681 = pi19 ? n32 : n12680;
  assign n12682 = pi18 ? n863 : ~n12681;
  assign n12683 = pi17 ? n32 : n12682;
  assign n12684 = pi16 ? n32 : n12683;
  assign n12685 = pi18 ? n863 : ~n245;
  assign n12686 = pi17 ? n32 : n12685;
  assign n12687 = pi16 ? n32 : n12686;
  assign n12688 = pi15 ? n12684 : n12687;
  assign n12689 = pi14 ? n12679 : n12688;
  assign n12690 = pi13 ? n12672 : n12689;
  assign n12691 = pi12 ? n12653 : n12690;
  assign n12692 = pi11 ? n12631 : n12691;
  assign n12693 = pi18 ? n1321 : ~n341;
  assign n12694 = pi17 ? n32 : n12693;
  assign n12695 = pi16 ? n32 : n12694;
  assign n12696 = pi15 ? n12687 : n12695;
  assign n12697 = pi18 ? n1321 : ~n684;
  assign n12698 = pi17 ? n32 : n12697;
  assign n12699 = pi16 ? n32 : n12698;
  assign n12700 = pi18 ? n1592 : ~n496;
  assign n12701 = pi17 ? n32 : n12700;
  assign n12702 = pi16 ? n32 : n12701;
  assign n12703 = pi15 ? n12699 : n12702;
  assign n12704 = pi14 ? n12696 : n12703;
  assign n12705 = pi18 ? n1592 : ~n12021;
  assign n12706 = pi17 ? n32 : n12705;
  assign n12707 = pi16 ? n32 : n12706;
  assign n12708 = pi19 ? n4491 : n2297;
  assign n12709 = pi18 ? n1592 : ~n12708;
  assign n12710 = pi17 ? n32 : n12709;
  assign n12711 = pi16 ? n32 : n12710;
  assign n12712 = pi15 ? n12707 : n12711;
  assign n12713 = pi18 ? n1592 : ~n1965;
  assign n12714 = pi17 ? n32 : n12713;
  assign n12715 = pi16 ? n32 : n12714;
  assign n12716 = pi15 ? n12715 : n12702;
  assign n12717 = pi14 ? n12712 : n12716;
  assign n12718 = pi13 ? n12704 : n12717;
  assign n12719 = pi18 ? n1970 : ~n496;
  assign n12720 = pi17 ? n32 : n12719;
  assign n12721 = pi16 ? n32 : n12720;
  assign n12722 = pi18 ? n1841 : ~n10891;
  assign n12723 = pi17 ? n32 : n12722;
  assign n12724 = pi16 ? n32 : n12723;
  assign n12725 = pi18 ? n1841 : ~n2849;
  assign n12726 = pi17 ? n32 : n12725;
  assign n12727 = pi16 ? n32 : n12726;
  assign n12728 = pi15 ? n12724 : n12727;
  assign n12729 = pi14 ? n12721 : n12728;
  assign n12730 = pi18 ? n1841 : ~n962;
  assign n12731 = pi17 ? n32 : n12730;
  assign n12732 = pi16 ? n32 : n12731;
  assign n12733 = pi18 ? n1841 : ~n697;
  assign n12734 = pi17 ? n32 : n12733;
  assign n12735 = pi16 ? n32 : n12734;
  assign n12736 = pi15 ? n12732 : n12735;
  assign n12737 = pi18 ? n1841 : ~n2730;
  assign n12738 = pi17 ? n32 : n12737;
  assign n12739 = pi16 ? n32 : n12738;
  assign n12740 = pi18 ? n940 : ~n2730;
  assign n12741 = pi17 ? n32 : n12740;
  assign n12742 = pi16 ? n32 : n12741;
  assign n12743 = pi15 ? n12739 : n12742;
  assign n12744 = pi14 ? n12736 : n12743;
  assign n12745 = pi13 ? n12729 : n12744;
  assign n12746 = pi12 ? n12718 : n12745;
  assign n12747 = pi18 ? n940 : ~n1750;
  assign n12748 = pi17 ? n32 : n12747;
  assign n12749 = pi16 ? n32 : n12748;
  assign n12750 = pi15 ? n12742 : n12749;
  assign n12751 = pi18 ? n940 : ~n2622;
  assign n12752 = pi17 ? n32 : n12751;
  assign n12753 = pi16 ? n32 : n12752;
  assign n12754 = pi18 ? n940 : ~n4098;
  assign n12755 = pi17 ? n32 : n12754;
  assign n12756 = pi16 ? n32 : n12755;
  assign n12757 = pi15 ? n12753 : n12756;
  assign n12758 = pi14 ? n12750 : n12757;
  assign n12759 = pi18 ? n863 : ~n4098;
  assign n12760 = pi17 ? n32 : n12759;
  assign n12761 = pi16 ? n32 : n12760;
  assign n12762 = pi18 ? n863 : ~n508;
  assign n12763 = pi17 ? n32 : n12762;
  assign n12764 = pi16 ? n32 : n12763;
  assign n12765 = pi18 ? n863 : ~n2747;
  assign n12766 = pi17 ? n32 : n12765;
  assign n12767 = pi16 ? n32 : n12766;
  assign n12768 = pi15 ? n12764 : n12767;
  assign n12769 = pi14 ? n12761 : n12768;
  assign n12770 = pi13 ? n12758 : n12769;
  assign n12771 = pi18 ? n863 : ~n323;
  assign n12772 = pi17 ? n32 : n12771;
  assign n12773 = pi16 ? n32 : n12772;
  assign n12774 = pi15 ? n12767 : n12773;
  assign n12775 = pi18 ? n863 : ~n797;
  assign n12776 = pi17 ? n32 : n12775;
  assign n12777 = pi16 ? n32 : n12776;
  assign n12778 = pi14 ? n12774 : n12777;
  assign n12779 = pi18 ? n32 : ~n2413;
  assign n12780 = pi17 ? n32 : n12779;
  assign n12781 = pi16 ? n32 : n12780;
  assign n12782 = pi18 ? n32 : ~n605;
  assign n12783 = pi17 ? n32 : n12782;
  assign n12784 = pi16 ? n32 : n12783;
  assign n12785 = pi15 ? n12781 : n12784;
  assign n12786 = pi18 ? n32 : ~n532;
  assign n12787 = pi17 ? n32 : n12786;
  assign n12788 = pi16 ? n32 : n12787;
  assign n12789 = pi18 ? n32 : ~n2298;
  assign n12790 = pi17 ? n32 : n12789;
  assign n12791 = pi16 ? n32 : n12790;
  assign n12792 = pi15 ? n12788 : n12791;
  assign n12793 = pi14 ? n12785 : n12792;
  assign n12794 = pi13 ? n12778 : n12793;
  assign n12795 = pi12 ? n12770 : n12794;
  assign n12796 = pi11 ? n12746 : n12795;
  assign n12797 = pi10 ? n12692 : n12796;
  assign n12798 = pi09 ? n12571 : n12797;
  assign n12799 = pi08 ? n12552 : n12798;
  assign n12800 = pi07 ? n12315 : n12799;
  assign n12801 = pi20 ? n7939 : ~n32;
  assign n12802 = pi19 ? n531 : ~n12801;
  assign n12803 = pi18 ? n32 : n12802;
  assign n12804 = pi17 ? n32 : n12803;
  assign n12805 = pi16 ? n32 : n12804;
  assign n12806 = pi15 ? n32 : n12805;
  assign n12807 = pi19 ? n531 : ~n8946;
  assign n12808 = pi18 ? n32 : n12807;
  assign n12809 = pi17 ? n32 : n12808;
  assign n12810 = pi16 ? n32 : n12809;
  assign n12811 = pi19 ? n531 : ~n531;
  assign n12812 = pi18 ? n32 : n12811;
  assign n12813 = pi17 ? n32 : n12812;
  assign n12814 = pi16 ? n32 : n12813;
  assign n12815 = pi15 ? n12810 : n12814;
  assign n12816 = pi14 ? n12806 : n12815;
  assign n12817 = pi13 ? n32 : n12816;
  assign n12818 = pi12 ? n32 : n12817;
  assign n12819 = pi11 ? n32 : n12818;
  assign n12820 = pi10 ? n32 : n12819;
  assign n12821 = pi20 ? n32 : ~n175;
  assign n12822 = pi20 ? n564 : ~n32;
  assign n12823 = pi19 ? n12821 : ~n12822;
  assign n12824 = pi18 ? n32 : n12823;
  assign n12825 = pi17 ? n32 : n12824;
  assign n12826 = pi16 ? n32 : n12825;
  assign n12827 = pi19 ? n2297 : n5707;
  assign n12828 = pi18 ? n32 : n12827;
  assign n12829 = pi17 ? n32 : n12828;
  assign n12830 = pi16 ? n32 : n12829;
  assign n12831 = pi15 ? n12826 : n12830;
  assign n12832 = pi19 ? n2297 : ~n531;
  assign n12833 = pi18 ? n32 : n12832;
  assign n12834 = pi17 ? n32 : n12833;
  assign n12835 = pi16 ? n32 : n12834;
  assign n12836 = pi14 ? n12831 : n12835;
  assign n12837 = pi19 ? n12578 : n5694;
  assign n12838 = pi18 ? n32 : n12837;
  assign n12839 = pi17 ? n32 : n12838;
  assign n12840 = pi16 ? n32 : n12839;
  assign n12841 = pi20 ? n342 : ~n405;
  assign n12842 = pi19 ? n12841 : n5694;
  assign n12843 = pi18 ? n32 : n12842;
  assign n12844 = pi17 ? n32 : n12843;
  assign n12845 = pi16 ? n32 : n12844;
  assign n12846 = pi15 ? n12840 : n12845;
  assign n12847 = pi19 ? n589 : ~n531;
  assign n12848 = pi18 ? n32 : n12847;
  assign n12849 = pi17 ? n32 : n12848;
  assign n12850 = pi16 ? n32 : n12849;
  assign n12851 = pi14 ? n12846 : n12850;
  assign n12852 = pi13 ? n12836 : n12851;
  assign n12853 = pi20 ? n1839 : ~n405;
  assign n12854 = pi20 ? n501 : n32;
  assign n12855 = pi19 ? n12853 : n12854;
  assign n12856 = pi18 ? n32 : n12855;
  assign n12857 = pi17 ? n32 : n12856;
  assign n12858 = pi16 ? n32 : n12857;
  assign n12859 = pi19 ? n6158 : n5707;
  assign n12860 = pi18 ? n32 : n12859;
  assign n12861 = pi17 ? n32 : n12860;
  assign n12862 = pi16 ? n32 : n12861;
  assign n12863 = pi15 ? n12858 : n12862;
  assign n12864 = pi14 ? n12863 : n12117;
  assign n12865 = pi19 ? n349 : ~n10072;
  assign n12866 = pi18 ? n32 : n12865;
  assign n12867 = pi17 ? n32 : n12866;
  assign n12868 = pi16 ? n32 : n12867;
  assign n12869 = pi15 ? n12868 : n12601;
  assign n12870 = pi19 ? n1812 : ~n365;
  assign n12871 = pi18 ? n32 : n12870;
  assign n12872 = pi17 ? n32 : n12871;
  assign n12873 = pi16 ? n32 : n12872;
  assign n12874 = pi19 ? n813 : ~n12171;
  assign n12875 = pi18 ? n32 : n12874;
  assign n12876 = pi17 ? n32 : n12875;
  assign n12877 = pi16 ? n32 : n12876;
  assign n12878 = pi15 ? n12873 : n12877;
  assign n12879 = pi14 ? n12869 : n12878;
  assign n12880 = pi13 ? n12864 : n12879;
  assign n12881 = pi12 ? n12852 : n12880;
  assign n12882 = pi21 ? n259 : n405;
  assign n12883 = pi20 ? n1940 : ~n12882;
  assign n12884 = pi21 ? n309 : ~n206;
  assign n12885 = pi20 ? n12884 : n32;
  assign n12886 = pi19 ? n12883 : n12885;
  assign n12887 = pi18 ? n32 : n12886;
  assign n12888 = pi17 ? n32 : n12887;
  assign n12889 = pi16 ? n32 : n12888;
  assign n12890 = pi19 ? n236 : ~n507;
  assign n12891 = pi18 ? n32 : n12890;
  assign n12892 = pi17 ? n32 : n12891;
  assign n12893 = pi16 ? n32 : n12892;
  assign n12894 = pi15 ? n12889 : n12893;
  assign n12895 = pi19 ? n236 : ~n343;
  assign n12896 = pi18 ? n32 : n12895;
  assign n12897 = pi17 ? n32 : n12896;
  assign n12898 = pi16 ? n32 : n12897;
  assign n12899 = pi20 ? n207 : ~n274;
  assign n12900 = pi19 ? n12899 : ~n422;
  assign n12901 = pi18 ? n32 : n12900;
  assign n12902 = pi17 ? n32 : n12901;
  assign n12903 = pi16 ? n32 : n12902;
  assign n12904 = pi15 ? n12898 : n12903;
  assign n12905 = pi14 ? n12894 : n12904;
  assign n12906 = pi19 ? n236 : ~n422;
  assign n12907 = pi18 ? n32 : n12906;
  assign n12908 = pi17 ? n32 : n12907;
  assign n12909 = pi16 ? n32 : n12908;
  assign n12910 = pi19 ? n236 : ~n10094;
  assign n12911 = pi18 ? n32 : n12910;
  assign n12912 = pi17 ? n32 : n12911;
  assign n12913 = pi16 ? n32 : n12912;
  assign n12914 = pi15 ? n12909 : n12913;
  assign n12915 = pi19 ? n236 : ~n1840;
  assign n12916 = pi18 ? n32 : n12915;
  assign n12917 = pi17 ? n32 : n12916;
  assign n12918 = pi16 ? n32 : n12917;
  assign n12919 = pi19 ? n2614 : ~n10593;
  assign n12920 = pi18 ? n32 : n12919;
  assign n12921 = pi17 ? n32 : n12920;
  assign n12922 = pi16 ? n32 : n12921;
  assign n12923 = pi15 ? n12918 : n12922;
  assign n12924 = pi14 ? n12914 : n12923;
  assign n12925 = pi13 ? n12905 : n12924;
  assign n12926 = pi19 ? n1105 : ~n531;
  assign n12927 = pi18 ? n32 : n12926;
  assign n12928 = pi17 ? n32 : n12927;
  assign n12929 = pi16 ? n32 : n12928;
  assign n12930 = pi20 ? n9641 : n207;
  assign n12931 = pi19 ? n1105 : ~n12930;
  assign n12932 = pi18 ? n32 : n12931;
  assign n12933 = pi17 ? n32 : n12932;
  assign n12934 = pi16 ? n32 : n12933;
  assign n12935 = pi15 ? n12929 : n12934;
  assign n12936 = pi19 ? n1105 : ~n10593;
  assign n12937 = pi18 ? n32 : n12936;
  assign n12938 = pi17 ? n32 : n12937;
  assign n12939 = pi16 ? n32 : n12938;
  assign n12940 = pi20 ? n141 : ~n357;
  assign n12941 = pi19 ? n12940 : ~n750;
  assign n12942 = pi18 ? n32 : n12941;
  assign n12943 = pi17 ? n32 : n12942;
  assign n12944 = pi16 ? n32 : n12943;
  assign n12945 = pi15 ? n12939 : n12944;
  assign n12946 = pi14 ? n12935 : n12945;
  assign n12947 = pi20 ? n342 : ~n481;
  assign n12948 = pi19 ? n1105 : ~n12947;
  assign n12949 = pi18 ? n32 : n12948;
  assign n12950 = pi17 ? n32 : n12949;
  assign n12951 = pi16 ? n32 : n12950;
  assign n12952 = pi19 ? n1105 : ~n429;
  assign n12953 = pi18 ? n32 : n12952;
  assign n12954 = pi17 ? n32 : n12953;
  assign n12955 = pi16 ? n32 : n12954;
  assign n12956 = pi15 ? n12951 : n12955;
  assign n12957 = pi20 ? n428 : ~n481;
  assign n12958 = pi19 ? n32 : n12957;
  assign n12959 = pi18 ? n32 : ~n12958;
  assign n12960 = pi17 ? n32 : n12959;
  assign n12961 = pi16 ? n32 : n12960;
  assign n12962 = pi15 ? n12955 : n12961;
  assign n12963 = pi14 ? n12956 : n12962;
  assign n12964 = pi13 ? n12946 : n12963;
  assign n12965 = pi12 ? n12925 : n12964;
  assign n12966 = pi11 ? n12881 : n12965;
  assign n12967 = pi18 ? n1575 : ~n341;
  assign n12968 = pi17 ? n32 : n12967;
  assign n12969 = pi16 ? n32 : n12968;
  assign n12970 = pi18 ? n1575 : ~n12021;
  assign n12971 = pi17 ? n32 : n12970;
  assign n12972 = pi16 ? n32 : n12971;
  assign n12973 = pi15 ? n12969 : n12972;
  assign n12974 = pi18 ? n1575 : ~n1965;
  assign n12975 = pi17 ? n32 : n12974;
  assign n12976 = pi16 ? n32 : n12975;
  assign n12977 = pi15 ? n12976 : n12972;
  assign n12978 = pi14 ? n12973 : n12977;
  assign n12979 = pi18 ? n936 : ~n2962;
  assign n12980 = pi17 ? n32 : n12979;
  assign n12981 = pi16 ? n32 : n12980;
  assign n12982 = pi21 ? n259 : ~n100;
  assign n12983 = pi20 ? n12982 : n32;
  assign n12984 = pi19 ? n32 : ~n12983;
  assign n12985 = pi18 ? n936 : ~n12984;
  assign n12986 = pi17 ? n32 : n12985;
  assign n12987 = pi16 ? n32 : n12986;
  assign n12988 = pi15 ? n12981 : n12987;
  assign n12989 = pi18 ? n936 : ~n1965;
  assign n12990 = pi17 ? n32 : n12989;
  assign n12991 = pi16 ? n32 : n12990;
  assign n12992 = pi18 ? n936 : ~n496;
  assign n12993 = pi17 ? n32 : n12992;
  assign n12994 = pi16 ? n32 : n12993;
  assign n12995 = pi15 ? n12991 : n12994;
  assign n12996 = pi14 ? n12988 : n12995;
  assign n12997 = pi13 ? n12978 : n12996;
  assign n12998 = pi18 ? n2142 : ~n590;
  assign n12999 = pi17 ? n32 : n12998;
  assign n13000 = pi16 ? n32 : n12999;
  assign n13001 = pi18 ? n2142 : ~n10891;
  assign n13002 = pi17 ? n32 : n13001;
  assign n13003 = pi16 ? n32 : n13002;
  assign n13004 = pi18 ? n2142 : ~n2849;
  assign n13005 = pi17 ? n32 : n13004;
  assign n13006 = pi16 ? n32 : n13005;
  assign n13007 = pi15 ? n13003 : n13006;
  assign n13008 = pi14 ? n13000 : n13007;
  assign n13009 = pi18 ? n2142 : ~n962;
  assign n13010 = pi17 ? n32 : n13009;
  assign n13011 = pi16 ? n32 : n13010;
  assign n13012 = pi18 ? n2142 : ~n2730;
  assign n13013 = pi17 ? n32 : n13012;
  assign n13014 = pi16 ? n32 : n13013;
  assign n13015 = pi15 ? n13011 : n13014;
  assign n13016 = pi18 ? n863 : ~n2730;
  assign n13017 = pi17 ? n32 : n13016;
  assign n13018 = pi16 ? n32 : n13017;
  assign n13019 = pi15 ? n13014 : n13018;
  assign n13020 = pi14 ? n13015 : n13019;
  assign n13021 = pi13 ? n13008 : n13020;
  assign n13022 = pi12 ? n12997 : n13021;
  assign n13023 = pi18 ? n863 : ~n1750;
  assign n13024 = pi17 ? n32 : n13023;
  assign n13025 = pi16 ? n32 : n13024;
  assign n13026 = pi18 ? n863 : ~n2622;
  assign n13027 = pi17 ? n32 : n13026;
  assign n13028 = pi16 ? n32 : n13027;
  assign n13029 = pi15 ? n13025 : n13028;
  assign n13030 = pi18 ? n32 : ~n2622;
  assign n13031 = pi17 ? n32 : n13030;
  assign n13032 = pi16 ? n32 : n13031;
  assign n13033 = pi18 ? n32 : ~n4098;
  assign n13034 = pi17 ? n32 : n13033;
  assign n13035 = pi16 ? n32 : n13034;
  assign n13036 = pi15 ? n13032 : n13035;
  assign n13037 = pi14 ? n13029 : n13036;
  assign n13038 = pi18 ? n32 : ~n508;
  assign n13039 = pi17 ? n32 : n13038;
  assign n13040 = pi16 ? n32 : n13039;
  assign n13041 = pi18 ? n32 : ~n2747;
  assign n13042 = pi17 ? n32 : n13041;
  assign n13043 = pi16 ? n32 : n13042;
  assign n13044 = pi18 ? n32 : ~n520;
  assign n13045 = pi17 ? n32 : n13044;
  assign n13046 = pi16 ? n32 : n13045;
  assign n13047 = pi15 ? n13043 : n13046;
  assign n13048 = pi14 ? n13040 : n13047;
  assign n13049 = pi13 ? n13037 : n13048;
  assign n13050 = pi18 ? n32 : ~n2291;
  assign n13051 = pi17 ? n32 : n13050;
  assign n13052 = pi16 ? n32 : n13051;
  assign n13053 = pi18 ? n32 : ~n797;
  assign n13054 = pi17 ? n32 : n13053;
  assign n13055 = pi16 ? n32 : n13054;
  assign n13056 = pi15 ? n13052 : n13055;
  assign n13057 = pi20 ? n207 : ~n749;
  assign n13058 = pi19 ? n13057 : n32;
  assign n13059 = pi18 ? n32 : n13058;
  assign n13060 = pi17 ? n32 : n13059;
  assign n13061 = pi16 ? n32 : n13060;
  assign n13062 = pi20 ? n207 : ~n1940;
  assign n13063 = pi19 ? n13062 : n32;
  assign n13064 = pi18 ? n32 : n13063;
  assign n13065 = pi17 ? n32 : n13064;
  assign n13066 = pi16 ? n32 : n13065;
  assign n13067 = pi15 ? n13061 : n13066;
  assign n13068 = pi14 ? n13056 : n13067;
  assign n13069 = pi20 ? n207 : ~n207;
  assign n13070 = pi19 ? n13069 : n32;
  assign n13071 = pi18 ? n32 : n13070;
  assign n13072 = pi17 ? n32 : n13071;
  assign n13073 = pi16 ? n32 : n13072;
  assign n13074 = pi20 ? n207 : ~n141;
  assign n13075 = pi19 ? n13074 : n32;
  assign n13076 = pi18 ? n32 : n13075;
  assign n13077 = pi17 ? n32 : n13076;
  assign n13078 = pi16 ? n32 : n13077;
  assign n13079 = pi15 ? n13073 : n13078;
  assign n13080 = pi19 ? n5707 : n32;
  assign n13081 = pi18 ? n32 : n13080;
  assign n13082 = pi17 ? n32 : n13081;
  assign n13083 = pi16 ? n32 : n13082;
  assign n13084 = pi21 ? n206 : ~n100;
  assign n13085 = pi20 ? n13084 : n32;
  assign n13086 = pi19 ? n13085 : n32;
  assign n13087 = pi18 ? n32 : n13086;
  assign n13088 = pi17 ? n32 : n13087;
  assign n13089 = pi16 ? n32 : n13088;
  assign n13090 = pi15 ? n13083 : n13089;
  assign n13091 = pi14 ? n13079 : n13090;
  assign n13092 = pi13 ? n13068 : n13091;
  assign n13093 = pi12 ? n13049 : n13092;
  assign n13094 = pi11 ? n13022 : n13093;
  assign n13095 = pi10 ? n12966 : n13094;
  assign n13096 = pi09 ? n12820 : n13095;
  assign n13097 = pi19 ? n340 : ~n4406;
  assign n13098 = pi18 ? n32 : n13097;
  assign n13099 = pi17 ? n32 : n13098;
  assign n13100 = pi16 ? n32 : n13099;
  assign n13101 = pi15 ? n32 : n13100;
  assign n13102 = pi19 ? n340 : ~n343;
  assign n13103 = pi18 ? n32 : n13102;
  assign n13104 = pi17 ? n32 : n13103;
  assign n13105 = pi16 ? n32 : n13104;
  assign n13106 = pi19 ? n340 : ~n531;
  assign n13107 = pi18 ? n32 : n13106;
  assign n13108 = pi17 ? n32 : n13107;
  assign n13109 = pi16 ? n32 : n13108;
  assign n13110 = pi15 ? n13105 : n13109;
  assign n13111 = pi14 ? n13101 : n13110;
  assign n13112 = pi13 ? n32 : n13111;
  assign n13113 = pi12 ? n32 : n13112;
  assign n13114 = pi11 ? n32 : n13113;
  assign n13115 = pi10 ? n32 : n13114;
  assign n13116 = pi19 ? n559 : ~n8818;
  assign n13117 = pi18 ? n32 : n13116;
  assign n13118 = pi17 ? n32 : n13117;
  assign n13119 = pi16 ? n32 : n13118;
  assign n13120 = pi19 ? n531 : n5707;
  assign n13121 = pi18 ? n32 : n13120;
  assign n13122 = pi17 ? n32 : n13121;
  assign n13123 = pi16 ? n32 : n13122;
  assign n13124 = pi15 ? n13119 : n13123;
  assign n13125 = pi14 ? n13124 : n12814;
  assign n13126 = pi20 ? n2140 : ~n101;
  assign n13127 = pi19 ? n13126 : n5694;
  assign n13128 = pi18 ? n32 : n13127;
  assign n13129 = pi17 ? n32 : n13128;
  assign n13130 = pi16 ? n32 : n13129;
  assign n13131 = pi20 ? n1331 : ~n321;
  assign n13132 = pi19 ? n2303 : n13131;
  assign n13133 = pi18 ? n32 : n13132;
  assign n13134 = pi17 ? n32 : n13133;
  assign n13135 = pi16 ? n32 : n13134;
  assign n13136 = pi15 ? n13130 : n13135;
  assign n13137 = pi19 ? n2303 : ~n531;
  assign n13138 = pi18 ? n32 : n13137;
  assign n13139 = pi17 ? n32 : n13138;
  assign n13140 = pi16 ? n32 : n13139;
  assign n13141 = pi14 ? n13136 : n13140;
  assign n13142 = pi13 ? n13125 : n13141;
  assign n13143 = pi19 ? n343 : n12854;
  assign n13144 = pi18 ? n32 : n13143;
  assign n13145 = pi17 ? n32 : n13144;
  assign n13146 = pi16 ? n32 : n13145;
  assign n13147 = pi19 ? n343 : n5707;
  assign n13148 = pi18 ? n32 : n13147;
  assign n13149 = pi17 ? n32 : n13148;
  assign n13150 = pi16 ? n32 : n13149;
  assign n13151 = pi15 ? n13146 : n13150;
  assign n13152 = pi14 ? n13151 : n12586;
  assign n13153 = pi19 ? n343 : ~n10072;
  assign n13154 = pi18 ? n32 : n13153;
  assign n13155 = pi17 ? n32 : n13154;
  assign n13156 = pi16 ? n32 : n13155;
  assign n13157 = pi15 ? n13156 : n12850;
  assign n13158 = pi19 ? n589 : ~n365;
  assign n13159 = pi18 ? n32 : n13158;
  assign n13160 = pi17 ? n32 : n13159;
  assign n13161 = pi16 ? n32 : n13160;
  assign n13162 = pi19 ? n2848 : ~n1508;
  assign n13163 = pi18 ? n32 : n13162;
  assign n13164 = pi17 ? n32 : n13163;
  assign n13165 = pi16 ? n32 : n13164;
  assign n13166 = pi15 ? n13161 : n13165;
  assign n13167 = pi14 ? n13157 : n13166;
  assign n13168 = pi13 ? n13152 : n13167;
  assign n13169 = pi12 ? n13142 : n13168;
  assign n13170 = pi20 ? n321 : ~n11107;
  assign n13171 = pi21 ? n313 : ~n206;
  assign n13172 = pi20 ? n13171 : n32;
  assign n13173 = pi19 ? n13170 : n13172;
  assign n13174 = pi18 ? n32 : n13173;
  assign n13175 = pi17 ? n32 : n13174;
  assign n13176 = pi16 ? n32 : n13175;
  assign n13177 = pi19 ? n349 : ~n11250;
  assign n13178 = pi18 ? n32 : n13177;
  assign n13179 = pi17 ? n32 : n13178;
  assign n13180 = pi16 ? n32 : n13179;
  assign n13181 = pi15 ? n13176 : n13180;
  assign n13182 = pi19 ? n349 : ~n343;
  assign n13183 = pi18 ? n32 : n13182;
  assign n13184 = pi17 ? n32 : n13183;
  assign n13185 = pi16 ? n32 : n13184;
  assign n13186 = pi15 ? n13185 : n12117;
  assign n13187 = pi14 ? n13181 : n13186;
  assign n13188 = pi19 ? n349 : ~n422;
  assign n13189 = pi18 ? n32 : n13188;
  assign n13190 = pi17 ? n32 : n13189;
  assign n13191 = pi16 ? n32 : n13190;
  assign n13192 = pi19 ? n349 : ~n10094;
  assign n13193 = pi18 ? n32 : n13192;
  assign n13194 = pi17 ? n32 : n13193;
  assign n13195 = pi16 ? n32 : n13194;
  assign n13196 = pi15 ? n13191 : n13195;
  assign n13197 = pi19 ? n1812 : ~n1840;
  assign n13198 = pi18 ? n32 : n13197;
  assign n13199 = pi17 ? n32 : n13198;
  assign n13200 = pi16 ? n32 : n13199;
  assign n13201 = pi15 ? n13200 : n12607;
  assign n13202 = pi14 ? n13196 : n13201;
  assign n13203 = pi13 ? n13187 : n13202;
  assign n13204 = pi19 ? n1941 : ~n531;
  assign n13205 = pi18 ? n32 : n13204;
  assign n13206 = pi17 ? n32 : n13205;
  assign n13207 = pi16 ? n32 : n13206;
  assign n13208 = pi19 ? n1941 : ~n12930;
  assign n13209 = pi18 ? n32 : n13208;
  assign n13210 = pi17 ? n32 : n13209;
  assign n13211 = pi16 ? n32 : n13210;
  assign n13212 = pi15 ? n13207 : n13211;
  assign n13213 = pi19 ? n1941 : ~n10593;
  assign n13214 = pi18 ? n32 : n13213;
  assign n13215 = pi17 ? n32 : n13214;
  assign n13216 = pi16 ? n32 : n13215;
  assign n13217 = pi19 ? n1941 : ~n750;
  assign n13218 = pi18 ? n32 : n13217;
  assign n13219 = pi17 ? n32 : n13218;
  assign n13220 = pi16 ? n32 : n13219;
  assign n13221 = pi15 ? n13216 : n13220;
  assign n13222 = pi14 ? n13212 : n13221;
  assign n13223 = pi19 ? n1941 : ~n429;
  assign n13224 = pi18 ? n32 : n13223;
  assign n13225 = pi17 ? n32 : n13224;
  assign n13226 = pi16 ? n32 : n13225;
  assign n13227 = pi15 ? n11877 : n13226;
  assign n13228 = pi19 ? n236 : ~n429;
  assign n13229 = pi18 ? n32 : n13228;
  assign n13230 = pi17 ? n32 : n13229;
  assign n13231 = pi16 ? n32 : n13230;
  assign n13232 = pi19 ? n2614 : ~n12957;
  assign n13233 = pi18 ? n32 : n13232;
  assign n13234 = pi17 ? n32 : n13233;
  assign n13235 = pi16 ? n32 : n13234;
  assign n13236 = pi15 ? n13231 : n13235;
  assign n13237 = pi14 ? n13227 : n13236;
  assign n13238 = pi13 ? n13222 : n13237;
  assign n13239 = pi12 ? n13203 : n13238;
  assign n13240 = pi11 ? n13169 : n13239;
  assign n13241 = pi19 ? n2614 : ~n340;
  assign n13242 = pi18 ? n32 : n13241;
  assign n13243 = pi17 ? n32 : n13242;
  assign n13244 = pi16 ? n32 : n13243;
  assign n13245 = pi21 ? n259 : ~n9326;
  assign n13246 = pi20 ? n13245 : n32;
  assign n13247 = pi19 ? n2614 : n13246;
  assign n13248 = pi18 ? n32 : n13247;
  assign n13249 = pi17 ? n32 : n13248;
  assign n13250 = pi16 ? n32 : n13249;
  assign n13251 = pi15 ? n13244 : n13250;
  assign n13252 = pi19 ? n2614 : ~n429;
  assign n13253 = pi18 ? n32 : n13252;
  assign n13254 = pi17 ? n32 : n13253;
  assign n13255 = pi16 ? n32 : n13254;
  assign n13256 = pi19 ? n2614 : ~n12020;
  assign n13257 = pi18 ? n32 : n13256;
  assign n13258 = pi17 ? n32 : n13257;
  assign n13259 = pi16 ? n32 : n13258;
  assign n13260 = pi15 ? n13255 : n13259;
  assign n13261 = pi14 ? n13251 : n13260;
  assign n13262 = pi21 ? n124 : n100;
  assign n13263 = pi20 ? n13262 : ~n32;
  assign n13264 = pi19 ? n2614 : ~n13263;
  assign n13265 = pi18 ? n32 : n13264;
  assign n13266 = pi17 ? n32 : n13265;
  assign n13267 = pi16 ? n32 : n13266;
  assign n13268 = pi15 ? n13267 : n13255;
  assign n13269 = pi21 ? n124 : n259;
  assign n13270 = pi20 ? n13269 : ~n32;
  assign n13271 = pi19 ? n617 : ~n13270;
  assign n13272 = pi18 ? n32 : n13271;
  assign n13273 = pi17 ? n32 : n13272;
  assign n13274 = pi16 ? n32 : n13273;
  assign n13275 = pi19 ? n1105 : ~n349;
  assign n13276 = pi18 ? n32 : n13275;
  assign n13277 = pi17 ? n32 : n13276;
  assign n13278 = pi16 ? n32 : n13277;
  assign n13279 = pi15 ? n13274 : n13278;
  assign n13280 = pi14 ? n13268 : n13279;
  assign n13281 = pi13 ? n13261 : n13280;
  assign n13282 = pi19 ? n1105 : ~n589;
  assign n13283 = pi18 ? n32 : n13282;
  assign n13284 = pi17 ? n32 : n13283;
  assign n13285 = pi16 ? n32 : n13284;
  assign n13286 = pi19 ? n1105 : ~n10890;
  assign n13287 = pi18 ? n32 : n13286;
  assign n13288 = pi17 ? n32 : n13287;
  assign n13289 = pi16 ? n32 : n13288;
  assign n13290 = pi19 ? n1105 : ~n1812;
  assign n13291 = pi18 ? n32 : n13290;
  assign n13292 = pi17 ? n32 : n13291;
  assign n13293 = pi16 ? n32 : n13292;
  assign n13294 = pi15 ? n13289 : n13293;
  assign n13295 = pi14 ? n13285 : n13294;
  assign n13296 = pi19 ? n1105 : ~n813;
  assign n13297 = pi18 ? n32 : n13296;
  assign n13298 = pi17 ? n32 : n13297;
  assign n13299 = pi16 ? n32 : n13298;
  assign n13300 = pi20 ? n243 : ~n428;
  assign n13301 = pi19 ? n13300 : ~n1941;
  assign n13302 = pi18 ? n32 : n13301;
  assign n13303 = pi17 ? n32 : n13302;
  assign n13304 = pi16 ? n32 : n13303;
  assign n13305 = pi15 ? n13299 : n13304;
  assign n13306 = pi19 ? n1105 : ~n1941;
  assign n13307 = pi18 ? n32 : n13306;
  assign n13308 = pi17 ? n32 : n13307;
  assign n13309 = pi16 ? n32 : n13308;
  assign n13310 = pi15 ? n13309 : n13304;
  assign n13311 = pi14 ? n13305 : n13310;
  assign n13312 = pi13 ? n13295 : n13311;
  assign n13313 = pi12 ? n13281 : n13312;
  assign n13314 = pi19 ? n2614 : ~n617;
  assign n13315 = pi18 ? n32 : n13314;
  assign n13316 = pi17 ? n32 : n13315;
  assign n13317 = pi16 ? n32 : n13316;
  assign n13318 = pi19 ? n236 : ~n1105;
  assign n13319 = pi18 ? n32 : n13318;
  assign n13320 = pi17 ? n32 : n13319;
  assign n13321 = pi16 ? n32 : n13320;
  assign n13322 = pi15 ? n13317 : n13321;
  assign n13323 = pi20 ? n207 : ~n428;
  assign n13324 = pi19 ? n13323 : n32;
  assign n13325 = pi18 ? n32 : n13324;
  assign n13326 = pi17 ? n32 : n13325;
  assign n13327 = pi16 ? n32 : n13326;
  assign n13328 = pi15 ? n13321 : n13327;
  assign n13329 = pi14 ? n13322 : n13328;
  assign n13330 = pi20 ? n207 : ~n2385;
  assign n13331 = pi19 ? n13330 : n32;
  assign n13332 = pi18 ? n32 : n13331;
  assign n13333 = pi17 ? n32 : n13332;
  assign n13334 = pi16 ? n32 : n13333;
  assign n13335 = pi19 ? n6307 : n32;
  assign n13336 = pi18 ? n32 : n13335;
  assign n13337 = pi17 ? n32 : n13336;
  assign n13338 = pi16 ? n32 : n13337;
  assign n13339 = pi15 ? n13334 : n13338;
  assign n13340 = pi20 ? n207 : ~n1319;
  assign n13341 = pi19 ? n13340 : n32;
  assign n13342 = pi18 ? n32 : n13341;
  assign n13343 = pi17 ? n32 : n13342;
  assign n13344 = pi16 ? n32 : n13343;
  assign n13345 = pi20 ? n749 : ~n518;
  assign n13346 = pi19 ? n13345 : n32;
  assign n13347 = pi18 ? n32 : n13346;
  assign n13348 = pi17 ? n32 : n13347;
  assign n13349 = pi16 ? n32 : n13348;
  assign n13350 = pi15 ? n13344 : n13349;
  assign n13351 = pi14 ? n13339 : n13350;
  assign n13352 = pi13 ? n13329 : n13351;
  assign n13353 = pi20 ? n1475 : ~n1475;
  assign n13354 = pi19 ? n13353 : n32;
  assign n13355 = pi18 ? n32 : n13354;
  assign n13356 = pi17 ? n32 : n13355;
  assign n13357 = pi16 ? n32 : n13356;
  assign n13358 = pi18 ? n32 : n5164;
  assign n13359 = pi17 ? n32 : n13358;
  assign n13360 = pi16 ? n32 : n13359;
  assign n13361 = pi15 ? n13357 : n13360;
  assign n13362 = pi20 ? n1475 : ~n749;
  assign n13363 = pi19 ? n13362 : n32;
  assign n13364 = pi18 ? n32 : n13363;
  assign n13365 = pi17 ? n32 : n13364;
  assign n13366 = pi16 ? n32 : n13365;
  assign n13367 = pi18 ? n32 : n5005;
  assign n13368 = pi17 ? n32 : n13367;
  assign n13369 = pi16 ? n32 : n13368;
  assign n13370 = pi15 ? n13366 : n13369;
  assign n13371 = pi14 ? n13361 : n13370;
  assign n13372 = pi19 ? n6420 : n32;
  assign n13373 = pi18 ? n32 : n13372;
  assign n13374 = pi17 ? n32 : n13373;
  assign n13375 = pi16 ? n32 : n13374;
  assign n13376 = pi20 ? n321 : ~n141;
  assign n13377 = pi19 ? n13376 : n32;
  assign n13378 = pi18 ? n32 : n13377;
  assign n13379 = pi17 ? n32 : n13378;
  assign n13380 = pi16 ? n32 : n13379;
  assign n13381 = pi15 ? n13375 : n13380;
  assign n13382 = pi20 ? n1319 : n32;
  assign n13383 = pi19 ? n13382 : n32;
  assign n13384 = pi18 ? n32 : n13383;
  assign n13385 = pi17 ? n32 : n13384;
  assign n13386 = pi16 ? n32 : n13385;
  assign n13387 = pi21 ? n32 : n7107;
  assign n13388 = pi20 ? n13387 : n32;
  assign n13389 = pi19 ? n13388 : n32;
  assign n13390 = pi18 ? n32 : n13389;
  assign n13391 = pi17 ? n32 : n13390;
  assign n13392 = pi16 ? n32 : n13391;
  assign n13393 = pi15 ? n13386 : n13392;
  assign n13394 = pi14 ? n13381 : n13393;
  assign n13395 = pi13 ? n13371 : n13394;
  assign n13396 = pi12 ? n13352 : n13395;
  assign n13397 = pi11 ? n13313 : n13396;
  assign n13398 = pi10 ? n13240 : n13397;
  assign n13399 = pi09 ? n13115 : n13398;
  assign n13400 = pi08 ? n13096 : n13399;
  assign n13401 = pi19 ? n1969 : ~n343;
  assign n13402 = pi18 ? n32 : n13401;
  assign n13403 = pi17 ? n32 : n13402;
  assign n13404 = pi16 ? n32 : n13403;
  assign n13405 = pi15 ? n32 : n13404;
  assign n13406 = pi19 ? n1969 : ~n531;
  assign n13407 = pi18 ? n32 : n13406;
  assign n13408 = pi17 ? n32 : n13407;
  assign n13409 = pi16 ? n32 : n13408;
  assign n13410 = pi15 ? n13404 : n13409;
  assign n13411 = pi14 ? n13405 : n13410;
  assign n13412 = pi13 ? n32 : n13411;
  assign n13413 = pi12 ? n32 : n13412;
  assign n13414 = pi11 ? n32 : n13413;
  assign n13415 = pi10 ? n32 : n13414;
  assign n13416 = pi19 ? n208 : ~n531;
  assign n13417 = pi18 ? n32 : n13416;
  assign n13418 = pi17 ? n32 : n13417;
  assign n13419 = pi16 ? n32 : n13418;
  assign n13420 = pi19 ? n244 : ~n531;
  assign n13421 = pi18 ? n32 : n13420;
  assign n13422 = pi17 ? n32 : n13421;
  assign n13423 = pi16 ? n32 : n13422;
  assign n13424 = pi15 ? n13419 : n13423;
  assign n13425 = pi14 ? n13424 : n13109;
  assign n13426 = pi21 ? n140 : n206;
  assign n13427 = pi20 ? n13426 : n321;
  assign n13428 = pi19 ? n2297 : ~n13427;
  assign n13429 = pi18 ? n32 : n13428;
  assign n13430 = pi17 ? n32 : n13429;
  assign n13431 = pi16 ? n32 : n13430;
  assign n13432 = pi19 ? n2297 : ~n1490;
  assign n13433 = pi18 ? n32 : n13432;
  assign n13434 = pi17 ? n32 : n13433;
  assign n13435 = pi16 ? n32 : n13434;
  assign n13436 = pi15 ? n13431 : n13435;
  assign n13437 = pi14 ? n13436 : n12835;
  assign n13438 = pi13 ? n13425 : n13437;
  assign n13439 = pi15 ? n12835 : n12565;
  assign n13440 = pi14 ? n12835 : n13439;
  assign n13441 = pi19 ? n2303 : ~n343;
  assign n13442 = pi18 ? n32 : n13441;
  assign n13443 = pi17 ? n32 : n13442;
  assign n13444 = pi16 ? n32 : n13443;
  assign n13445 = pi19 ? n2303 : ~n365;
  assign n13446 = pi18 ? n32 : n13445;
  assign n13447 = pi17 ? n32 : n13446;
  assign n13448 = pi16 ? n32 : n13447;
  assign n13449 = pi15 ? n13444 : n13448;
  assign n13450 = pi19 ? n2303 : ~n11250;
  assign n13451 = pi18 ? n32 : n13450;
  assign n13452 = pi17 ? n32 : n13451;
  assign n13453 = pi16 ? n32 : n13452;
  assign n13454 = pi15 ? n13140 : n13453;
  assign n13455 = pi14 ? n13449 : n13454;
  assign n13456 = pi13 ? n13440 : n13455;
  assign n13457 = pi12 ? n13438 : n13456;
  assign n13458 = pi19 ? n343 : n3692;
  assign n13459 = pi18 ? n32 : n13458;
  assign n13460 = pi17 ? n32 : n13459;
  assign n13461 = pi16 ? n32 : n13460;
  assign n13462 = pi19 ? n343 : ~n11250;
  assign n13463 = pi18 ? n32 : n13462;
  assign n13464 = pi17 ? n32 : n13463;
  assign n13465 = pi16 ? n32 : n13464;
  assign n13466 = pi15 ? n13461 : n13465;
  assign n13467 = pi19 ? n343 : ~n343;
  assign n13468 = pi18 ? n32 : n13467;
  assign n13469 = pi17 ? n32 : n13468;
  assign n13470 = pi16 ? n32 : n13469;
  assign n13471 = pi19 ? n343 : ~n11488;
  assign n13472 = pi18 ? n32 : n13471;
  assign n13473 = pi17 ? n32 : n13472;
  assign n13474 = pi16 ? n32 : n13473;
  assign n13475 = pi15 ? n13470 : n13474;
  assign n13476 = pi14 ? n13466 : n13475;
  assign n13477 = pi19 ? n343 : ~n422;
  assign n13478 = pi18 ? n32 : n13477;
  assign n13479 = pi17 ? n32 : n13478;
  assign n13480 = pi16 ? n32 : n13479;
  assign n13481 = pi19 ? n2317 : ~n11488;
  assign n13482 = pi18 ? n32 : n13481;
  assign n13483 = pi17 ? n32 : n13482;
  assign n13484 = pi16 ? n32 : n13483;
  assign n13485 = pi15 ? n13480 : n13484;
  assign n13486 = pi20 ? n428 : n1839;
  assign n13487 = pi19 ? n2317 : ~n13486;
  assign n13488 = pi18 ? n32 : n13487;
  assign n13489 = pi17 ? n32 : n13488;
  assign n13490 = pi16 ? n32 : n13489;
  assign n13491 = pi19 ? n589 : ~n11546;
  assign n13492 = pi18 ? n32 : n13491;
  assign n13493 = pi17 ? n32 : n13492;
  assign n13494 = pi16 ? n32 : n13493;
  assign n13495 = pi15 ? n13490 : n13494;
  assign n13496 = pi14 ? n13485 : n13495;
  assign n13497 = pi13 ? n13476 : n13496;
  assign n13498 = pi19 ? n2848 : ~n12416;
  assign n13499 = pi18 ? n32 : n13498;
  assign n13500 = pi17 ? n32 : n13499;
  assign n13501 = pi16 ? n32 : n13500;
  assign n13502 = pi20 ? n86 : n749;
  assign n13503 = pi19 ? n2848 : ~n13502;
  assign n13504 = pi18 ? n32 : n13503;
  assign n13505 = pi17 ? n32 : n13504;
  assign n13506 = pi16 ? n32 : n13505;
  assign n13507 = pi15 ? n13501 : n13506;
  assign n13508 = pi19 ? n2848 : ~n11504;
  assign n13509 = pi18 ? n32 : n13508;
  assign n13510 = pi17 ? n32 : n13509;
  assign n13511 = pi16 ? n32 : n13510;
  assign n13512 = pi20 ? n175 : n749;
  assign n13513 = pi19 ? n2848 : ~n13512;
  assign n13514 = pi18 ? n32 : n13513;
  assign n13515 = pi17 ? n32 : n13514;
  assign n13516 = pi16 ? n32 : n13515;
  assign n13517 = pi15 ? n13511 : n13516;
  assign n13518 = pi14 ? n13507 : n13517;
  assign n13519 = pi19 ? n2848 : ~n1265;
  assign n13520 = pi18 ? n32 : n13519;
  assign n13521 = pi17 ? n32 : n13520;
  assign n13522 = pi16 ? n32 : n13521;
  assign n13523 = pi20 ? n1839 : ~n1817;
  assign n13524 = pi19 ? n13523 : ~n12957;
  assign n13525 = pi18 ? n32 : n13524;
  assign n13526 = pi17 ? n32 : n13525;
  assign n13527 = pi16 ? n32 : n13526;
  assign n13528 = pi15 ? n13522 : n13527;
  assign n13529 = pi20 ? n321 : ~n1817;
  assign n13530 = pi19 ? n13529 : ~n340;
  assign n13531 = pi18 ? n32 : n13530;
  assign n13532 = pi17 ? n32 : n13531;
  assign n13533 = pi16 ? n32 : n13532;
  assign n13534 = pi19 ? n1812 : ~n12957;
  assign n13535 = pi18 ? n32 : n13534;
  assign n13536 = pi17 ? n32 : n13535;
  assign n13537 = pi16 ? n32 : n13536;
  assign n13538 = pi15 ? n13533 : n13537;
  assign n13539 = pi14 ? n13528 : n13538;
  assign n13540 = pi13 ? n13518 : n13539;
  assign n13541 = pi12 ? n13497 : n13540;
  assign n13542 = pi11 ? n13457 : n13541;
  assign n13543 = pi20 ? n3523 : n339;
  assign n13544 = pi19 ? n1812 : ~n13543;
  assign n13545 = pi18 ? n32 : n13544;
  assign n13546 = pi17 ? n32 : n13545;
  assign n13547 = pi16 ? n32 : n13546;
  assign n13548 = pi19 ? n1812 : ~n1265;
  assign n13549 = pi18 ? n32 : n13548;
  assign n13550 = pi17 ? n32 : n13549;
  assign n13551 = pi16 ? n32 : n13550;
  assign n13552 = pi15 ? n13547 : n13551;
  assign n13553 = pi19 ? n1812 : ~n2297;
  assign n13554 = pi18 ? n32 : n13553;
  assign n13555 = pi17 ? n32 : n13554;
  assign n13556 = pi16 ? n32 : n13555;
  assign n13557 = pi19 ? n1812 : ~n429;
  assign n13558 = pi18 ? n32 : n13557;
  assign n13559 = pi17 ? n32 : n13558;
  assign n13560 = pi16 ? n32 : n13559;
  assign n13561 = pi15 ? n13556 : n13560;
  assign n13562 = pi14 ? n13552 : n13561;
  assign n13563 = pi19 ? n1812 : ~n13263;
  assign n13564 = pi18 ? n32 : n13563;
  assign n13565 = pi17 ? n32 : n13564;
  assign n13566 = pi16 ? n32 : n13565;
  assign n13567 = pi15 ? n13566 : n13560;
  assign n13568 = pi19 ? n813 : ~n13270;
  assign n13569 = pi18 ? n32 : n13568;
  assign n13570 = pi17 ? n32 : n13569;
  assign n13571 = pi16 ? n32 : n13570;
  assign n13572 = pi19 ? n1941 : ~n589;
  assign n13573 = pi18 ? n32 : n13572;
  assign n13574 = pi17 ? n32 : n13573;
  assign n13575 = pi16 ? n32 : n13574;
  assign n13576 = pi15 ? n13571 : n13575;
  assign n13577 = pi14 ? n13567 : n13576;
  assign n13578 = pi13 ? n13562 : n13577;
  assign n13579 = pi19 ? n1941 : ~n10895;
  assign n13580 = pi18 ? n32 : n13579;
  assign n13581 = pi17 ? n32 : n13580;
  assign n13582 = pi16 ? n32 : n13581;
  assign n13583 = pi15 ? n13582 : n13575;
  assign n13584 = pi23 ? n33 : ~n33;
  assign n13585 = pi22 ? n173 : ~n13584;
  assign n13586 = pi21 ? n13585 : ~n32;
  assign n13587 = pi20 ? n13586 : ~n32;
  assign n13588 = pi19 ? n1941 : ~n13587;
  assign n13589 = pi18 ? n32 : n13588;
  assign n13590 = pi17 ? n32 : n13589;
  assign n13591 = pi16 ? n32 : n13590;
  assign n13592 = pi19 ? n1941 : ~n813;
  assign n13593 = pi18 ? n32 : n13592;
  assign n13594 = pi17 ? n32 : n13593;
  assign n13595 = pi16 ? n32 : n13594;
  assign n13596 = pi15 ? n13591 : n13595;
  assign n13597 = pi14 ? n13583 : n13596;
  assign n13598 = pi19 ? n1812 : ~n813;
  assign n13599 = pi18 ? n32 : n13598;
  assign n13600 = pi17 ? n32 : n13599;
  assign n13601 = pi16 ? n32 : n13600;
  assign n13602 = pi19 ? n1812 : ~n1941;
  assign n13603 = pi18 ? n32 : n13602;
  assign n13604 = pi17 ? n32 : n13603;
  assign n13605 = pi16 ? n32 : n13604;
  assign n13606 = pi15 ? n13601 : n13605;
  assign n13607 = pi19 ? n1812 : ~n617;
  assign n13608 = pi18 ? n32 : n13607;
  assign n13609 = pi17 ? n32 : n13608;
  assign n13610 = pi16 ? n32 : n13609;
  assign n13611 = pi14 ? n13606 : n13610;
  assign n13612 = pi13 ? n13597 : n13611;
  assign n13613 = pi12 ? n13578 : n13612;
  assign n13614 = pi19 ? n1812 : ~n1105;
  assign n13615 = pi18 ? n32 : n13614;
  assign n13616 = pi17 ? n32 : n13615;
  assign n13617 = pi16 ? n32 : n13616;
  assign n13618 = pi18 ? n32 : n6163;
  assign n13619 = pi17 ? n32 : n13618;
  assign n13620 = pi16 ? n32 : n13619;
  assign n13621 = pi15 ? n13617 : n13620;
  assign n13622 = pi20 ? n321 : ~n2140;
  assign n13623 = pi19 ? n13622 : n32;
  assign n13624 = pi18 ? n32 : n13623;
  assign n13625 = pi17 ? n32 : n13624;
  assign n13626 = pi16 ? n32 : n13625;
  assign n13627 = pi18 ? n32 : n5357;
  assign n13628 = pi17 ? n32 : n13627;
  assign n13629 = pi16 ? n32 : n13628;
  assign n13630 = pi15 ? n13626 : n13629;
  assign n13631 = pi14 ? n13621 : n13630;
  assign n13632 = pi20 ? n321 : ~n1319;
  assign n13633 = pi19 ? n13632 : n32;
  assign n13634 = pi18 ? n32 : n13633;
  assign n13635 = pi17 ? n32 : n13634;
  assign n13636 = pi16 ? n32 : n13635;
  assign n13637 = pi15 ? n13629 : n13636;
  assign n13638 = pi20 ? n518 : ~n518;
  assign n13639 = pi19 ? n13638 : n32;
  assign n13640 = pi18 ? n32 : n13639;
  assign n13641 = pi17 ? n32 : n13640;
  assign n13642 = pi16 ? n32 : n13641;
  assign n13643 = pi20 ? n518 : ~n1475;
  assign n13644 = pi19 ? n13643 : n32;
  assign n13645 = pi18 ? n32 : n13644;
  assign n13646 = pi17 ? n32 : n13645;
  assign n13647 = pi16 ? n32 : n13646;
  assign n13648 = pi15 ? n13642 : n13647;
  assign n13649 = pi14 ? n13637 : n13648;
  assign n13650 = pi13 ? n13631 : n13649;
  assign n13651 = pi20 ? n1319 : ~n1475;
  assign n13652 = pi19 ? n13651 : n32;
  assign n13653 = pi18 ? n32 : n13652;
  assign n13654 = pi17 ? n32 : n13653;
  assign n13655 = pi16 ? n32 : n13654;
  assign n13656 = pi20 ? n342 : ~n749;
  assign n13657 = pi19 ? n13656 : n32;
  assign n13658 = pi18 ? n32 : n13657;
  assign n13659 = pi17 ? n32 : n13658;
  assign n13660 = pi16 ? n32 : n13659;
  assign n13661 = pi15 ? n13655 : n13660;
  assign n13662 = pi20 ? n1319 : ~n207;
  assign n13663 = pi19 ? n13662 : n32;
  assign n13664 = pi18 ? n32 : n13663;
  assign n13665 = pi17 ? n32 : n13664;
  assign n13666 = pi16 ? n32 : n13665;
  assign n13667 = pi20 ? n342 : ~n339;
  assign n13668 = pi19 ? n13667 : n32;
  assign n13669 = pi18 ? n32 : n13668;
  assign n13670 = pi17 ? n32 : n13669;
  assign n13671 = pi16 ? n32 : n13670;
  assign n13672 = pi15 ? n13666 : n13671;
  assign n13673 = pi14 ? n13661 : n13672;
  assign n13674 = pi21 ? n32 : n11567;
  assign n13675 = pi20 ? n13674 : ~n141;
  assign n13676 = pi19 ? n13675 : n32;
  assign n13677 = pi18 ? n32 : n13676;
  assign n13678 = pi17 ? n32 : n13677;
  assign n13679 = pi16 ? n32 : n13678;
  assign n13680 = pi20 ? n428 : ~n141;
  assign n13681 = pi19 ? n13680 : n32;
  assign n13682 = pi18 ? n32 : n13681;
  assign n13683 = pi17 ? n32 : n13682;
  assign n13684 = pi16 ? n32 : n13683;
  assign n13685 = pi15 ? n13679 : n13684;
  assign n13686 = pi14 ? n13685 : n32;
  assign n13687 = pi13 ? n13673 : n13686;
  assign n13688 = pi12 ? n13650 : n13687;
  assign n13689 = pi11 ? n13613 : n13688;
  assign n13690 = pi10 ? n13542 : n13689;
  assign n13691 = pi09 ? n13415 : n13690;
  assign n13692 = pi19 ? n1476 : ~n343;
  assign n13693 = pi18 ? n32 : n13692;
  assign n13694 = pi17 ? n32 : n13693;
  assign n13695 = pi16 ? n32 : n13694;
  assign n13696 = pi15 ? n32 : n13695;
  assign n13697 = pi19 ? n1476 : ~n531;
  assign n13698 = pi18 ? n32 : n13697;
  assign n13699 = pi17 ? n32 : n13698;
  assign n13700 = pi16 ? n32 : n13699;
  assign n13701 = pi15 ? n13695 : n13700;
  assign n13702 = pi14 ? n13696 : n13701;
  assign n13703 = pi13 ? n32 : n13702;
  assign n13704 = pi12 ? n32 : n13703;
  assign n13705 = pi11 ? n32 : n13704;
  assign n13706 = pi10 ? n32 : n13705;
  assign n13707 = pi19 ? n750 : ~n531;
  assign n13708 = pi18 ? n32 : n13707;
  assign n13709 = pi17 ? n32 : n13708;
  assign n13710 = pi16 ? n32 : n13709;
  assign n13711 = pi15 ? n13710 : n13409;
  assign n13712 = pi15 ? n13409 : n13109;
  assign n13713 = pi14 ? n13711 : n13712;
  assign n13714 = pi20 ? n7939 : n321;
  assign n13715 = pi19 ? n365 : ~n13714;
  assign n13716 = pi18 ? n32 : n13715;
  assign n13717 = pi17 ? n32 : n13716;
  assign n13718 = pi16 ? n32 : n13717;
  assign n13719 = pi19 ? n365 : ~n1490;
  assign n13720 = pi18 ? n32 : n13719;
  assign n13721 = pi17 ? n32 : n13720;
  assign n13722 = pi16 ? n32 : n13721;
  assign n13723 = pi15 ? n13718 : n13722;
  assign n13724 = pi19 ? n365 : ~n531;
  assign n13725 = pi18 ? n32 : n13724;
  assign n13726 = pi17 ? n32 : n13725;
  assign n13727 = pi16 ? n32 : n13726;
  assign n13728 = pi14 ? n13723 : n13727;
  assign n13729 = pi13 ? n13713 : n13728;
  assign n13730 = pi19 ? n2297 : ~n343;
  assign n13731 = pi18 ? n32 : n13730;
  assign n13732 = pi17 ? n32 : n13731;
  assign n13733 = pi16 ? n32 : n13732;
  assign n13734 = pi15 ? n13733 : n12835;
  assign n13735 = pi19 ? n2297 : ~n11250;
  assign n13736 = pi18 ? n32 : n13735;
  assign n13737 = pi17 ? n32 : n13736;
  assign n13738 = pi16 ? n32 : n13737;
  assign n13739 = pi15 ? n12835 : n13738;
  assign n13740 = pi14 ? n13734 : n13739;
  assign n13741 = pi13 ? n12814 : n13740;
  assign n13742 = pi12 ? n13729 : n13741;
  assign n13743 = pi19 ? n2297 : n3692;
  assign n13744 = pi18 ? n32 : n13743;
  assign n13745 = pi17 ? n32 : n13744;
  assign n13746 = pi16 ? n32 : n13745;
  assign n13747 = pi20 ? n32 : ~n623;
  assign n13748 = pi19 ? n2297 : ~n13747;
  assign n13749 = pi18 ? n32 : n13748;
  assign n13750 = pi17 ? n32 : n13749;
  assign n13751 = pi16 ? n32 : n13750;
  assign n13752 = pi15 ? n13746 : n13751;
  assign n13753 = pi19 ? n429 : ~n11488;
  assign n13754 = pi18 ? n32 : n13753;
  assign n13755 = pi17 ? n32 : n13754;
  assign n13756 = pi16 ? n32 : n13755;
  assign n13757 = pi15 ? n13733 : n13756;
  assign n13758 = pi14 ? n13752 : n13757;
  assign n13759 = pi19 ? n429 : ~n422;
  assign n13760 = pi18 ? n32 : n13759;
  assign n13761 = pi17 ? n32 : n13760;
  assign n13762 = pi16 ? n32 : n13761;
  assign n13763 = pi19 ? n429 : ~n429;
  assign n13764 = pi18 ? n32 : n13763;
  assign n13765 = pi17 ? n32 : n13764;
  assign n13766 = pi16 ? n32 : n13765;
  assign n13767 = pi15 ? n13762 : n13766;
  assign n13768 = pi19 ? n429 : ~n1868;
  assign n13769 = pi18 ? n32 : n13768;
  assign n13770 = pi17 ? n32 : n13769;
  assign n13771 = pi16 ? n32 : n13770;
  assign n13772 = pi19 ? n429 : ~n6042;
  assign n13773 = pi18 ? n32 : n13772;
  assign n13774 = pi17 ? n32 : n13773;
  assign n13775 = pi16 ? n32 : n13774;
  assign n13776 = pi15 ? n13771 : n13775;
  assign n13777 = pi14 ? n13767 : n13776;
  assign n13778 = pi13 ? n13758 : n13777;
  assign n13779 = pi20 ? n1324 : ~n6229;
  assign n13780 = pi19 ? n2303 : ~n13779;
  assign n13781 = pi18 ? n32 : n13780;
  assign n13782 = pi17 ? n32 : n13781;
  assign n13783 = pi16 ? n32 : n13782;
  assign n13784 = pi22 ? n34 : ~n173;
  assign n13785 = pi21 ? n32 : n13784;
  assign n13786 = pi20 ? n13785 : n749;
  assign n13787 = pi19 ? n2303 : ~n13786;
  assign n13788 = pi18 ? n32 : n13787;
  assign n13789 = pi17 ? n32 : n13788;
  assign n13790 = pi16 ? n32 : n13789;
  assign n13791 = pi15 ? n13783 : n13790;
  assign n13792 = pi21 ? n32 : n7659;
  assign n13793 = pi20 ? n13792 : ~n32;
  assign n13794 = pi19 ? n2303 : ~n13793;
  assign n13795 = pi18 ? n32 : n13794;
  assign n13796 = pi17 ? n32 : n13795;
  assign n13797 = pi16 ? n32 : n13796;
  assign n13798 = pi20 ? n13785 : n339;
  assign n13799 = pi19 ? n2303 : ~n13798;
  assign n13800 = pi18 ? n32 : n13799;
  assign n13801 = pi17 ? n32 : n13800;
  assign n13802 = pi16 ? n32 : n13801;
  assign n13803 = pi15 ? n13797 : n13802;
  assign n13804 = pi14 ? n13791 : n13803;
  assign n13805 = pi19 ? n2303 : ~n1265;
  assign n13806 = pi18 ? n32 : n13805;
  assign n13807 = pi17 ? n32 : n13806;
  assign n13808 = pi16 ? n32 : n13807;
  assign n13809 = pi19 ? n10568 : ~n11541;
  assign n13810 = pi18 ? n32 : n13809;
  assign n13811 = pi17 ? n32 : n13810;
  assign n13812 = pi16 ? n32 : n13811;
  assign n13813 = pi15 ? n13808 : n13812;
  assign n13814 = pi19 ? n10568 : ~n340;
  assign n13815 = pi18 ? n32 : n13814;
  assign n13816 = pi17 ? n32 : n13815;
  assign n13817 = pi16 ? n32 : n13816;
  assign n13818 = pi19 ? n2317 : ~n11541;
  assign n13819 = pi18 ? n32 : n13818;
  assign n13820 = pi17 ? n32 : n13819;
  assign n13821 = pi16 ? n32 : n13820;
  assign n13822 = pi15 ? n13817 : n13821;
  assign n13823 = pi14 ? n13813 : n13822;
  assign n13824 = pi13 ? n13804 : n13823;
  assign n13825 = pi12 ? n13778 : n13824;
  assign n13826 = pi11 ? n13742 : n13825;
  assign n13827 = pi19 ? n2317 : ~n340;
  assign n13828 = pi18 ? n32 : n13827;
  assign n13829 = pi17 ? n32 : n13828;
  assign n13830 = pi16 ? n32 : n13829;
  assign n13831 = pi19 ? n2317 : ~n1265;
  assign n13832 = pi18 ? n32 : n13831;
  assign n13833 = pi17 ? n32 : n13832;
  assign n13834 = pi16 ? n32 : n13833;
  assign n13835 = pi15 ? n13830 : n13834;
  assign n13836 = pi19 ? n2317 : ~n2297;
  assign n13837 = pi18 ? n32 : n13836;
  assign n13838 = pi17 ? n32 : n13837;
  assign n13839 = pi16 ? n32 : n13838;
  assign n13840 = pi19 ? n2317 : ~n429;
  assign n13841 = pi18 ? n32 : n13840;
  assign n13842 = pi17 ? n32 : n13841;
  assign n13843 = pi16 ? n32 : n13842;
  assign n13844 = pi15 ? n13839 : n13843;
  assign n13845 = pi14 ? n13835 : n13844;
  assign n13846 = pi19 ? n2317 : ~n343;
  assign n13847 = pi18 ? n32 : n13846;
  assign n13848 = pi17 ? n32 : n13847;
  assign n13849 = pi16 ? n32 : n13848;
  assign n13850 = pi15 ? n13839 : n13849;
  assign n13851 = pi19 ? n589 : ~n589;
  assign n13852 = pi18 ? n32 : n13851;
  assign n13853 = pi17 ? n32 : n13852;
  assign n13854 = pi16 ? n32 : n13853;
  assign n13855 = pi19 ? n2848 : n10662;
  assign n13856 = pi18 ? n32 : n13855;
  assign n13857 = pi17 ? n32 : n13856;
  assign n13858 = pi16 ? n32 : n13857;
  assign n13859 = pi15 ? n13854 : n13858;
  assign n13860 = pi14 ? n13850 : n13859;
  assign n13861 = pi13 ? n13845 : n13860;
  assign n13862 = pi19 ? n2848 : ~n10895;
  assign n13863 = pi18 ? n32 : n13862;
  assign n13864 = pi17 ? n32 : n13863;
  assign n13865 = pi16 ? n32 : n13864;
  assign n13866 = pi19 ? n2848 : ~n589;
  assign n13867 = pi18 ? n32 : n13866;
  assign n13868 = pi17 ? n32 : n13867;
  assign n13869 = pi16 ? n32 : n13868;
  assign n13870 = pi15 ? n13865 : n13869;
  assign n13871 = pi19 ? n2848 : ~n1812;
  assign n13872 = pi18 ? n32 : n13871;
  assign n13873 = pi17 ? n32 : n13872;
  assign n13874 = pi16 ? n32 : n13873;
  assign n13875 = pi19 ? n2848 : ~n813;
  assign n13876 = pi18 ? n32 : n13875;
  assign n13877 = pi17 ? n32 : n13876;
  assign n13878 = pi16 ? n32 : n13877;
  assign n13879 = pi15 ? n13874 : n13878;
  assign n13880 = pi14 ? n13870 : n13879;
  assign n13881 = pi19 ? n2317 : ~n813;
  assign n13882 = pi18 ? n32 : n13881;
  assign n13883 = pi17 ? n32 : n13882;
  assign n13884 = pi16 ? n32 : n13883;
  assign n13885 = pi19 ? n2317 : ~n236;
  assign n13886 = pi18 ? n32 : n13885;
  assign n13887 = pi17 ? n32 : n13886;
  assign n13888 = pi16 ? n32 : n13887;
  assign n13889 = pi15 ? n13884 : n13888;
  assign n13890 = pi19 ? n2317 : ~n617;
  assign n13891 = pi18 ? n32 : n13890;
  assign n13892 = pi17 ? n32 : n13891;
  assign n13893 = pi16 ? n32 : n13892;
  assign n13894 = pi14 ? n13889 : n13893;
  assign n13895 = pi13 ? n13880 : n13894;
  assign n13896 = pi12 ? n13861 : n13895;
  assign n13897 = pi19 ? n2317 : ~n1105;
  assign n13898 = pi18 ? n32 : n13897;
  assign n13899 = pi17 ? n32 : n13898;
  assign n13900 = pi16 ? n32 : n13899;
  assign n13901 = pi19 ? n343 : n32;
  assign n13902 = pi18 ? n32 : n13901;
  assign n13903 = pi17 ? n32 : n13902;
  assign n13904 = pi16 ? n32 : n13903;
  assign n13905 = pi15 ? n13900 : n13904;
  assign n13906 = pi20 ? n342 : ~n2140;
  assign n13907 = pi19 ? n13906 : n32;
  assign n13908 = pi18 ? n32 : n13907;
  assign n13909 = pi17 ? n32 : n13908;
  assign n13910 = pi16 ? n32 : n13909;
  assign n13911 = pi18 ? n32 : n5742;
  assign n13912 = pi17 ? n32 : n13911;
  assign n13913 = pi16 ? n32 : n13912;
  assign n13914 = pi15 ? n13910 : n13913;
  assign n13915 = pi14 ? n13905 : n13914;
  assign n13916 = pi20 ? n342 : ~n518;
  assign n13917 = pi19 ? n13916 : n32;
  assign n13918 = pi18 ? n32 : n13917;
  assign n13919 = pi17 ? n32 : n13918;
  assign n13920 = pi16 ? n32 : n13919;
  assign n13921 = pi15 ? n13913 : n13920;
  assign n13922 = pi19 ? n9591 : n32;
  assign n13923 = pi18 ? n32 : n13922;
  assign n13924 = pi17 ? n32 : n13923;
  assign n13925 = pi16 ? n32 : n13924;
  assign n13926 = pi20 ? n428 : ~n1475;
  assign n13927 = pi19 ? n13926 : n32;
  assign n13928 = pi18 ? n32 : n13927;
  assign n13929 = pi17 ? n32 : n13928;
  assign n13930 = pi16 ? n32 : n13929;
  assign n13931 = pi15 ? n13925 : n13930;
  assign n13932 = pi14 ? n13921 : n13931;
  assign n13933 = pi13 ? n13915 : n13932;
  assign n13934 = pi20 ? n101 : ~n1475;
  assign n13935 = pi19 ? n13934 : n32;
  assign n13936 = pi18 ? n32 : n13935;
  assign n13937 = pi17 ? n32 : n13936;
  assign n13938 = pi16 ? n32 : n13937;
  assign n13939 = pi20 ? n32 : ~n749;
  assign n13940 = pi19 ? n13939 : n32;
  assign n13941 = pi18 ? n32 : n13940;
  assign n13942 = pi17 ? n32 : n13941;
  assign n13943 = pi16 ? n32 : n13942;
  assign n13944 = pi15 ? n13938 : n13943;
  assign n13945 = pi19 ? n9007 : n32;
  assign n13946 = pi18 ? n32 : n13945;
  assign n13947 = pi17 ? n32 : n13946;
  assign n13948 = pi16 ? n32 : n13947;
  assign n13949 = pi19 ? n8622 : n32;
  assign n13950 = pi18 ? n32 : n13949;
  assign n13951 = pi17 ? n32 : n13950;
  assign n13952 = pi16 ? n32 : n13951;
  assign n13953 = pi15 ? n13948 : n13952;
  assign n13954 = pi14 ? n13944 : n13953;
  assign n13955 = pi13 ? n13954 : n32;
  assign n13956 = pi12 ? n13933 : n13955;
  assign n13957 = pi11 ? n13896 : n13956;
  assign n13958 = pi10 ? n13826 : n13957;
  assign n13959 = pi09 ? n13706 : n13958;
  assign n13960 = pi08 ? n13691 : n13959;
  assign n13961 = pi07 ? n13400 : n13960;
  assign n13962 = pi06 ? n12800 : n13961;
  assign n13963 = pi05 ? n11873 : n13962;
  assign n13964 = pi04 ? n9997 : n13963;
  assign n13965 = pi19 ? n1840 : ~n531;
  assign n13966 = pi18 ? n32 : n13965;
  assign n13967 = pi17 ? n32 : n13966;
  assign n13968 = pi16 ? n32 : n13967;
  assign n13969 = pi15 ? n32 : n13968;
  assign n13970 = pi14 ? n13969 : n13968;
  assign n13971 = pi13 ? n32 : n13970;
  assign n13972 = pi12 ? n32 : n13971;
  assign n13973 = pi11 ? n32 : n13972;
  assign n13974 = pi10 ? n32 : n13973;
  assign n13975 = pi19 ? n322 : ~n531;
  assign n13976 = pi18 ? n32 : n13975;
  assign n13977 = pi17 ? n32 : n13976;
  assign n13978 = pi16 ? n32 : n13977;
  assign n13979 = pi15 ? n13978 : n13700;
  assign n13980 = pi15 ? n13700 : n13409;
  assign n13981 = pi14 ? n13979 : n13980;
  assign n13982 = pi19 ? n208 : ~n322;
  assign n13983 = pi18 ? n32 : n13982;
  assign n13984 = pi17 ? n32 : n13983;
  assign n13985 = pi16 ? n32 : n13984;
  assign n13986 = pi14 ? n13419 : n13985;
  assign n13987 = pi13 ? n13981 : n13986;
  assign n13988 = pi19 ? n244 : ~n322;
  assign n13989 = pi18 ? n32 : n13988;
  assign n13990 = pi17 ? n32 : n13989;
  assign n13991 = pi16 ? n32 : n13990;
  assign n13992 = pi19 ? n340 : ~n322;
  assign n13993 = pi18 ? n32 : n13992;
  assign n13994 = pi17 ? n32 : n13993;
  assign n13995 = pi16 ? n32 : n13994;
  assign n13996 = pi14 ? n13991 : n13995;
  assign n13997 = pi19 ? n365 : ~n11929;
  assign n13998 = pi18 ? n32 : n13997;
  assign n13999 = pi17 ? n32 : n13998;
  assign n14000 = pi16 ? n32 : n13999;
  assign n14001 = pi15 ? n13727 : n14000;
  assign n14002 = pi19 ? n365 : ~n343;
  assign n14003 = pi18 ? n32 : n14002;
  assign n14004 = pi17 ? n32 : n14003;
  assign n14005 = pi16 ? n32 : n14004;
  assign n14006 = pi19 ? n365 : ~n8546;
  assign n14007 = pi18 ? n32 : n14006;
  assign n14008 = pi17 ? n32 : n14007;
  assign n14009 = pi16 ? n32 : n14008;
  assign n14010 = pi15 ? n14005 : n14009;
  assign n14011 = pi14 ? n14001 : n14010;
  assign n14012 = pi13 ? n13996 : n14011;
  assign n14013 = pi12 ? n13987 : n14012;
  assign n14014 = pi18 ? n32 : n7042;
  assign n14015 = pi17 ? n32 : n14014;
  assign n14016 = pi16 ? n32 : n14015;
  assign n14017 = pi19 ? n531 : ~n11027;
  assign n14018 = pi18 ? n32 : n14017;
  assign n14019 = pi17 ? n32 : n14018;
  assign n14020 = pi16 ? n32 : n14019;
  assign n14021 = pi15 ? n14016 : n14020;
  assign n14022 = pi20 ? n32 : ~n915;
  assign n14023 = pi19 ? n531 : ~n14022;
  assign n14024 = pi18 ? n32 : n14023;
  assign n14025 = pi17 ? n32 : n14024;
  assign n14026 = pi16 ? n32 : n14025;
  assign n14027 = pi15 ? n14026 : n14020;
  assign n14028 = pi14 ? n14021 : n14027;
  assign n14029 = pi19 ? n531 : ~n10485;
  assign n14030 = pi18 ? n32 : n14029;
  assign n14031 = pi17 ? n32 : n14030;
  assign n14032 = pi16 ? n32 : n14031;
  assign n14033 = pi19 ? n531 : ~n1740;
  assign n14034 = pi18 ? n32 : n14033;
  assign n14035 = pi17 ? n32 : n14034;
  assign n14036 = pi16 ? n32 : n14035;
  assign n14037 = pi15 ? n12814 : n14036;
  assign n14038 = pi14 ? n14032 : n14037;
  assign n14039 = pi13 ? n14028 : n14038;
  assign n14040 = pi20 ? n86 : n11048;
  assign n14041 = pi19 ? n531 : ~n14040;
  assign n14042 = pi18 ? n32 : n14041;
  assign n14043 = pi17 ? n32 : n14042;
  assign n14044 = pi16 ? n32 : n14043;
  assign n14045 = pi19 ? n531 : ~n1053;
  assign n14046 = pi18 ? n32 : n14045;
  assign n14047 = pi17 ? n32 : n14046;
  assign n14048 = pi16 ? n32 : n14047;
  assign n14049 = pi15 ? n14044 : n14048;
  assign n14050 = pi20 ? n151 : n207;
  assign n14051 = pi19 ? n531 : ~n14050;
  assign n14052 = pi18 ? n32 : n14051;
  assign n14053 = pi17 ? n32 : n14052;
  assign n14054 = pi16 ? n32 : n14053;
  assign n14055 = pi19 ? n2297 : ~n1265;
  assign n14056 = pi18 ? n32 : n14055;
  assign n14057 = pi17 ? n32 : n14056;
  assign n14058 = pi16 ? n32 : n14057;
  assign n14059 = pi15 ? n14054 : n14058;
  assign n14060 = pi14 ? n14049 : n14059;
  assign n14061 = pi19 ? n2297 : ~n340;
  assign n14062 = pi18 ? n32 : n14061;
  assign n14063 = pi17 ? n32 : n14062;
  assign n14064 = pi16 ? n32 : n14063;
  assign n14065 = pi20 ? n175 : n243;
  assign n14066 = pi19 ? n2297 : ~n14065;
  assign n14067 = pi18 ? n32 : n14066;
  assign n14068 = pi17 ? n32 : n14067;
  assign n14069 = pi16 ? n32 : n14068;
  assign n14070 = pi15 ? n14064 : n14069;
  assign n14071 = pi19 ? n2297 : ~n12435;
  assign n14072 = pi18 ? n32 : n14071;
  assign n14073 = pi17 ? n32 : n14072;
  assign n14074 = pi16 ? n32 : n14073;
  assign n14075 = pi15 ? n14064 : n14074;
  assign n14076 = pi14 ? n14070 : n14075;
  assign n14077 = pi13 ? n14060 : n14076;
  assign n14078 = pi12 ? n14039 : n14077;
  assign n14079 = pi11 ? n14013 : n14078;
  assign n14080 = pi19 ? n2297 : ~n429;
  assign n14081 = pi18 ? n32 : n14080;
  assign n14082 = pi17 ? n32 : n14081;
  assign n14083 = pi16 ? n32 : n14082;
  assign n14084 = pi19 ? n2297 : ~n2297;
  assign n14085 = pi18 ? n32 : n14084;
  assign n14086 = pi17 ? n32 : n14085;
  assign n14087 = pi16 ? n32 : n14086;
  assign n14088 = pi14 ? n14083 : n14087;
  assign n14089 = pi19 ? n2297 : ~n2317;
  assign n14090 = pi18 ? n32 : n14089;
  assign n14091 = pi17 ? n32 : n14090;
  assign n14092 = pi16 ? n32 : n14091;
  assign n14093 = pi19 ? n429 : ~n2317;
  assign n14094 = pi18 ? n32 : n14093;
  assign n14095 = pi17 ? n32 : n14094;
  assign n14096 = pi16 ? n32 : n14095;
  assign n14097 = pi15 ? n14092 : n14096;
  assign n14098 = pi19 ? n429 : ~n589;
  assign n14099 = pi18 ? n32 : n14098;
  assign n14100 = pi17 ? n32 : n14099;
  assign n14101 = pi16 ? n32 : n14100;
  assign n14102 = pi19 ? n2303 : ~n589;
  assign n14103 = pi18 ? n32 : n14102;
  assign n14104 = pi17 ? n32 : n14103;
  assign n14105 = pi16 ? n32 : n14104;
  assign n14106 = pi15 ? n14101 : n14105;
  assign n14107 = pi14 ? n14097 : n14106;
  assign n14108 = pi13 ? n14088 : n14107;
  assign n14109 = pi19 ? n2303 : ~n1812;
  assign n14110 = pi18 ? n32 : n14109;
  assign n14111 = pi17 ? n32 : n14110;
  assign n14112 = pi16 ? n32 : n14111;
  assign n14113 = pi19 ? n2303 : ~n813;
  assign n14114 = pi18 ? n32 : n14113;
  assign n14115 = pi17 ? n32 : n14114;
  assign n14116 = pi16 ? n32 : n14115;
  assign n14117 = pi15 ? n14112 : n14116;
  assign n14118 = pi19 ? n2303 : ~n236;
  assign n14119 = pi18 ? n32 : n14118;
  assign n14120 = pi17 ? n32 : n14119;
  assign n14121 = pi16 ? n32 : n14120;
  assign n14122 = pi15 ? n14116 : n14121;
  assign n14123 = pi14 ? n14117 : n14122;
  assign n14124 = pi19 ? n2297 : ~n617;
  assign n14125 = pi18 ? n32 : n14124;
  assign n14126 = pi17 ? n32 : n14125;
  assign n14127 = pi16 ? n32 : n14126;
  assign n14128 = pi19 ? n531 : ~n1105;
  assign n14129 = pi18 ? n32 : n14128;
  assign n14130 = pi17 ? n32 : n14129;
  assign n14131 = pi16 ? n32 : n14130;
  assign n14132 = pi15 ? n14127 : n14131;
  assign n14133 = pi14 ? n14127 : n14132;
  assign n14134 = pi13 ? n14123 : n14133;
  assign n14135 = pi12 ? n14108 : n14134;
  assign n14136 = pi18 ? n32 : n5335;
  assign n14137 = pi17 ? n32 : n14136;
  assign n14138 = pi16 ? n32 : n14137;
  assign n14139 = pi20 ? n32 : ~n2140;
  assign n14140 = pi19 ? n14139 : n32;
  assign n14141 = pi18 ? n32 : n14140;
  assign n14142 = pi17 ? n32 : n14141;
  assign n14143 = pi16 ? n32 : n14142;
  assign n14144 = pi15 ? n14138 : n14143;
  assign n14145 = pi18 ? n32 : n4983;
  assign n14146 = pi17 ? n32 : n14145;
  assign n14147 = pi16 ? n32 : n14146;
  assign n14148 = pi15 ? n14143 : n14147;
  assign n14149 = pi14 ? n14144 : n14148;
  assign n14150 = pi18 ? n32 : n5731;
  assign n14151 = pi17 ? n32 : n14150;
  assign n14152 = pi16 ? n32 : n14151;
  assign n14153 = pi19 ? n5694 : n32;
  assign n14154 = pi18 ? n32 : n14153;
  assign n14155 = pi17 ? n32 : n14154;
  assign n14156 = pi16 ? n32 : n14155;
  assign n14157 = pi15 ? n14152 : n14156;
  assign n14158 = pi22 ? n173 : ~n34;
  assign n14159 = pi21 ? n14158 : n32;
  assign n14160 = pi20 ? n32 : n14159;
  assign n14161 = pi19 ? n14160 : n32;
  assign n14162 = pi18 ? n32 : n14161;
  assign n14163 = pi17 ? n32 : n14162;
  assign n14164 = pi16 ? n32 : n14163;
  assign n14165 = pi19 ? n572 : n32;
  assign n14166 = pi18 ? n32 : n14165;
  assign n14167 = pi17 ? n32 : n14166;
  assign n14168 = pi16 ? n32 : n14167;
  assign n14169 = pi15 ? n14164 : n14168;
  assign n14170 = pi14 ? n14157 : n14169;
  assign n14171 = pi13 ? n14149 : n14170;
  assign n14172 = pi12 ? n14171 : n32;
  assign n14173 = pi11 ? n14135 : n14172;
  assign n14174 = pi10 ? n14079 : n14173;
  assign n14175 = pi09 ? n13974 : n14174;
  assign n14176 = pi19 ? n519 : ~n531;
  assign n14177 = pi18 ? n32 : n14176;
  assign n14178 = pi17 ? n32 : n14177;
  assign n14179 = pi16 ? n32 : n14178;
  assign n14180 = pi15 ? n32 : n14179;
  assign n14181 = pi14 ? n14180 : n14179;
  assign n14182 = pi13 ? n32 : n14181;
  assign n14183 = pi12 ? n32 : n14182;
  assign n14184 = pi11 ? n32 : n14183;
  assign n14185 = pi10 ? n32 : n14184;
  assign n14186 = pi15 ? n14179 : n13968;
  assign n14187 = pi15 ? n13968 : n13700;
  assign n14188 = pi14 ? n14186 : n14187;
  assign n14189 = pi19 ? n750 : ~n322;
  assign n14190 = pi18 ? n32 : n14189;
  assign n14191 = pi17 ? n32 : n14190;
  assign n14192 = pi16 ? n32 : n14191;
  assign n14193 = pi14 ? n13710 : n14192;
  assign n14194 = pi13 ? n14188 : n14193;
  assign n14195 = pi19 ? n1969 : ~n322;
  assign n14196 = pi18 ? n32 : n14195;
  assign n14197 = pi17 ? n32 : n14196;
  assign n14198 = pi16 ? n32 : n14197;
  assign n14199 = pi19 ? n208 : ~n9001;
  assign n14200 = pi18 ? n32 : n14199;
  assign n14201 = pi17 ? n32 : n14200;
  assign n14202 = pi16 ? n32 : n14201;
  assign n14203 = pi15 ? n13419 : n14202;
  assign n14204 = pi19 ? n208 : ~n343;
  assign n14205 = pi18 ? n32 : n14204;
  assign n14206 = pi17 ? n32 : n14205;
  assign n14207 = pi16 ? n32 : n14206;
  assign n14208 = pi19 ? n208 : ~n8546;
  assign n14209 = pi18 ? n32 : n14208;
  assign n14210 = pi17 ? n32 : n14209;
  assign n14211 = pi16 ? n32 : n14210;
  assign n14212 = pi15 ? n14207 : n14211;
  assign n14213 = pi14 ? n14203 : n14212;
  assign n14214 = pi13 ? n14198 : n14213;
  assign n14215 = pi12 ? n14194 : n14214;
  assign n14216 = pi19 ? n244 : ~n343;
  assign n14217 = pi18 ? n32 : n14216;
  assign n14218 = pi17 ? n32 : n14217;
  assign n14219 = pi16 ? n32 : n14218;
  assign n14220 = pi19 ? n244 : ~n11027;
  assign n14221 = pi18 ? n32 : n14220;
  assign n14222 = pi17 ? n32 : n14221;
  assign n14223 = pi16 ? n32 : n14222;
  assign n14224 = pi15 ? n14219 : n14223;
  assign n14225 = pi19 ? n340 : ~n11027;
  assign n14226 = pi18 ? n32 : n14225;
  assign n14227 = pi17 ? n32 : n14226;
  assign n14228 = pi16 ? n32 : n14227;
  assign n14229 = pi15 ? n13995 : n14228;
  assign n14230 = pi14 ? n14224 : n14229;
  assign n14231 = pi19 ? n340 : ~n10485;
  assign n14232 = pi18 ? n32 : n14231;
  assign n14233 = pi17 ? n32 : n14232;
  assign n14234 = pi16 ? n32 : n14233;
  assign n14235 = pi19 ? n340 : ~n1490;
  assign n14236 = pi18 ? n32 : n14235;
  assign n14237 = pi17 ? n32 : n14236;
  assign n14238 = pi16 ? n32 : n14237;
  assign n14239 = pi15 ? n14234 : n14238;
  assign n14240 = pi19 ? n340 : ~n422;
  assign n14241 = pi18 ? n32 : n14240;
  assign n14242 = pi17 ? n32 : n14241;
  assign n14243 = pi16 ? n32 : n14242;
  assign n14244 = pi19 ? n340 : ~n1740;
  assign n14245 = pi18 ? n32 : n14244;
  assign n14246 = pi17 ? n32 : n14245;
  assign n14247 = pi16 ? n32 : n14246;
  assign n14248 = pi15 ? n14243 : n14247;
  assign n14249 = pi14 ? n14239 : n14248;
  assign n14250 = pi13 ? n14230 : n14249;
  assign n14251 = pi19 ? n365 : ~n11049;
  assign n14252 = pi18 ? n32 : n14251;
  assign n14253 = pi17 ? n32 : n14252;
  assign n14254 = pi16 ? n32 : n14253;
  assign n14255 = pi19 ? n365 : ~n1053;
  assign n14256 = pi18 ? n32 : n14255;
  assign n14257 = pi17 ? n32 : n14256;
  assign n14258 = pi16 ? n32 : n14257;
  assign n14259 = pi15 ? n14254 : n14258;
  assign n14260 = pi20 ? n3523 : n207;
  assign n14261 = pi19 ? n365 : ~n14260;
  assign n14262 = pi18 ? n32 : n14261;
  assign n14263 = pi17 ? n32 : n14262;
  assign n14264 = pi16 ? n32 : n14263;
  assign n14265 = pi19 ? n365 : ~n13793;
  assign n14266 = pi18 ? n32 : n14265;
  assign n14267 = pi17 ? n32 : n14266;
  assign n14268 = pi16 ? n32 : n14267;
  assign n14269 = pi15 ? n14264 : n14268;
  assign n14270 = pi14 ? n14259 : n14269;
  assign n14271 = pi19 ? n365 : ~n340;
  assign n14272 = pi18 ? n32 : n14271;
  assign n14273 = pi17 ? n32 : n14272;
  assign n14274 = pi16 ? n32 : n14273;
  assign n14275 = pi20 ? n13785 : n243;
  assign n14276 = pi19 ? n365 : ~n14275;
  assign n14277 = pi18 ? n32 : n14276;
  assign n14278 = pi17 ? n32 : n14277;
  assign n14279 = pi16 ? n32 : n14278;
  assign n14280 = pi15 ? n14274 : n14279;
  assign n14281 = pi20 ? n151 : n339;
  assign n14282 = pi19 ? n365 : ~n14281;
  assign n14283 = pi18 ? n32 : n14282;
  assign n14284 = pi17 ? n32 : n14283;
  assign n14285 = pi16 ? n32 : n14284;
  assign n14286 = pi21 ? n32 : n313;
  assign n14287 = pi20 ? n14286 : n339;
  assign n14288 = pi19 ? n340 : ~n14287;
  assign n14289 = pi18 ? n32 : n14288;
  assign n14290 = pi17 ? n32 : n14289;
  assign n14291 = pi16 ? n32 : n14290;
  assign n14292 = pi15 ? n14285 : n14291;
  assign n14293 = pi14 ? n14280 : n14292;
  assign n14294 = pi13 ? n14270 : n14293;
  assign n14295 = pi12 ? n14250 : n14294;
  assign n14296 = pi11 ? n14215 : n14295;
  assign n14297 = pi21 ? n32 : n34;
  assign n14298 = pi20 ? n14297 : ~n32;
  assign n14299 = pi19 ? n365 : ~n14298;
  assign n14300 = pi18 ? n32 : n14299;
  assign n14301 = pi17 ? n32 : n14300;
  assign n14302 = pi16 ? n32 : n14301;
  assign n14303 = pi19 ? n340 : ~n2297;
  assign n14304 = pi18 ? n32 : n14303;
  assign n14305 = pi17 ? n32 : n14304;
  assign n14306 = pi16 ? n32 : n14305;
  assign n14307 = pi15 ? n14302 : n14306;
  assign n14308 = pi19 ? n340 : ~n14298;
  assign n14309 = pi18 ? n32 : n14308;
  assign n14310 = pi17 ? n32 : n14309;
  assign n14311 = pi16 ? n32 : n14310;
  assign n14312 = pi19 ? n365 : ~n2297;
  assign n14313 = pi18 ? n32 : n14312;
  assign n14314 = pi17 ? n32 : n14313;
  assign n14315 = pi16 ? n32 : n14314;
  assign n14316 = pi15 ? n14311 : n14315;
  assign n14317 = pi14 ? n14307 : n14316;
  assign n14318 = pi21 ? n8275 : ~n32;
  assign n14319 = pi20 ? n32 : n14318;
  assign n14320 = pi19 ? n14319 : ~n2317;
  assign n14321 = pi18 ? n32 : n14320;
  assign n14322 = pi17 ? n32 : n14321;
  assign n14323 = pi16 ? n32 : n14322;
  assign n14324 = pi19 ? n365 : ~n2317;
  assign n14325 = pi18 ? n32 : n14324;
  assign n14326 = pi17 ? n32 : n14325;
  assign n14327 = pi16 ? n32 : n14326;
  assign n14328 = pi15 ? n14323 : n14327;
  assign n14329 = pi19 ? n531 : ~n2848;
  assign n14330 = pi18 ? n32 : n14329;
  assign n14331 = pi17 ? n32 : n14330;
  assign n14332 = pi16 ? n32 : n14331;
  assign n14333 = pi15 ? n14327 : n14332;
  assign n14334 = pi14 ? n14328 : n14333;
  assign n14335 = pi13 ? n14317 : n14334;
  assign n14336 = pi19 ? n531 : ~n1812;
  assign n14337 = pi18 ? n32 : n14336;
  assign n14338 = pi17 ? n32 : n14337;
  assign n14339 = pi16 ? n32 : n14338;
  assign n14340 = pi19 ? n365 : ~n813;
  assign n14341 = pi18 ? n32 : n14340;
  assign n14342 = pi17 ? n32 : n14341;
  assign n14343 = pi16 ? n32 : n14342;
  assign n14344 = pi15 ? n14339 : n14343;
  assign n14345 = pi19 ? n365 : ~n1941;
  assign n14346 = pi18 ? n32 : n14345;
  assign n14347 = pi17 ? n32 : n14346;
  assign n14348 = pi16 ? n32 : n14347;
  assign n14349 = pi15 ? n14343 : n14348;
  assign n14350 = pi14 ? n14344 : n14349;
  assign n14351 = pi19 ? n365 : ~n617;
  assign n14352 = pi18 ? n32 : n14351;
  assign n14353 = pi17 ? n32 : n14352;
  assign n14354 = pi16 ? n32 : n14353;
  assign n14355 = pi19 ? n340 : ~n617;
  assign n14356 = pi18 ? n32 : n14355;
  assign n14357 = pi17 ? n32 : n14356;
  assign n14358 = pi16 ? n32 : n14357;
  assign n14359 = pi15 ? n14354 : n14358;
  assign n14360 = pi19 ? n832 : n32;
  assign n14361 = pi18 ? n32 : n14360;
  assign n14362 = pi17 ? n32 : n14361;
  assign n14363 = pi16 ? n32 : n14362;
  assign n14364 = pi15 ? n14358 : n14363;
  assign n14365 = pi14 ? n14359 : n14364;
  assign n14366 = pi13 ? n14350 : n14365;
  assign n14367 = pi12 ? n14335 : n14366;
  assign n14368 = pi21 ? n242 : ~n405;
  assign n14369 = pi20 ? n32 : n14368;
  assign n14370 = pi19 ? n14369 : n32;
  assign n14371 = pi18 ? n32 : n14370;
  assign n14372 = pi17 ? n32 : n14371;
  assign n14373 = pi16 ? n32 : n14372;
  assign n14374 = pi21 ? n259 : ~n1939;
  assign n14375 = pi20 ? n32 : n14374;
  assign n14376 = pi19 ? n14375 : n32;
  assign n14377 = pi18 ? n32 : n14376;
  assign n14378 = pi17 ? n32 : n14377;
  assign n14379 = pi16 ? n32 : n14378;
  assign n14380 = pi15 ? n14373 : n14379;
  assign n14381 = pi21 ? n242 : ~n1939;
  assign n14382 = pi20 ? n32 : n14381;
  assign n14383 = pi19 ? n14382 : n32;
  assign n14384 = pi18 ? n32 : n14383;
  assign n14385 = pi17 ? n32 : n14384;
  assign n14386 = pi16 ? n32 : n14385;
  assign n14387 = pi18 ? n32 : n5502;
  assign n14388 = pi17 ? n32 : n14387;
  assign n14389 = pi16 ? n32 : n14388;
  assign n14390 = pi15 ? n14386 : n14389;
  assign n14391 = pi14 ? n14380 : n14390;
  assign n14392 = pi18 ? n32 : n5351;
  assign n14393 = pi17 ? n32 : n14392;
  assign n14394 = pi16 ? n32 : n14393;
  assign n14395 = pi18 ? n32 : n9012;
  assign n14396 = pi17 ? n32 : n14395;
  assign n14397 = pi16 ? n32 : n14396;
  assign n14398 = pi15 ? n14394 : n14397;
  assign n14399 = pi22 ? n32 : n13584;
  assign n14400 = pi21 ? n14399 : n32;
  assign n14401 = pi20 ? n32 : n14400;
  assign n14402 = pi19 ? n14401 : n32;
  assign n14403 = pi18 ? n32 : n14402;
  assign n14404 = pi17 ? n32 : n14403;
  assign n14405 = pi16 ? n32 : n14404;
  assign n14406 = pi14 ? n14398 : n14405;
  assign n14407 = pi13 ? n14391 : n14406;
  assign n14408 = pi12 ? n14407 : n32;
  assign n14409 = pi11 ? n14367 : n14408;
  assign n14410 = pi10 ? n14296 : n14409;
  assign n14411 = pi09 ? n14185 : n14410;
  assign n14412 = pi08 ? n14175 : n14411;
  assign n14413 = pi19 ? n507 : ~n531;
  assign n14414 = pi18 ? n32 : n14413;
  assign n14415 = pi17 ? n32 : n14414;
  assign n14416 = pi16 ? n32 : n14415;
  assign n14417 = pi15 ? n32 : n14416;
  assign n14418 = pi14 ? n14417 : n14416;
  assign n14419 = pi13 ? n32 : n14418;
  assign n14420 = pi12 ? n32 : n14419;
  assign n14421 = pi11 ? n32 : n14420;
  assign n14422 = pi10 ? n32 : n14421;
  assign n14423 = pi19 ? n1320 : ~n531;
  assign n14424 = pi18 ? n32 : n14423;
  assign n14425 = pi17 ? n32 : n14424;
  assign n14426 = pi16 ? n32 : n14425;
  assign n14427 = pi15 ? n14426 : n14179;
  assign n14428 = pi14 ? n14427 : n14186;
  assign n14429 = pi19 ? n322 : ~n322;
  assign n14430 = pi18 ? n32 : n14429;
  assign n14431 = pi17 ? n32 : n14430;
  assign n14432 = pi16 ? n32 : n14431;
  assign n14433 = pi14 ? n13978 : n14432;
  assign n14434 = pi13 ? n14428 : n14433;
  assign n14435 = pi19 ? n1476 : ~n322;
  assign n14436 = pi18 ? n32 : n14435;
  assign n14437 = pi17 ? n32 : n14436;
  assign n14438 = pi16 ? n32 : n14437;
  assign n14439 = pi19 ? n750 : ~n9001;
  assign n14440 = pi18 ? n32 : n14439;
  assign n14441 = pi17 ? n32 : n14440;
  assign n14442 = pi16 ? n32 : n14441;
  assign n14443 = pi15 ? n13710 : n14442;
  assign n14444 = pi19 ? n750 : ~n343;
  assign n14445 = pi18 ? n32 : n14444;
  assign n14446 = pi17 ? n32 : n14445;
  assign n14447 = pi16 ? n32 : n14446;
  assign n14448 = pi15 ? n14447 : n13710;
  assign n14449 = pi14 ? n14443 : n14448;
  assign n14450 = pi13 ? n14438 : n14449;
  assign n14451 = pi12 ? n14434 : n14450;
  assign n14452 = pi19 ? n1969 : ~n11027;
  assign n14453 = pi18 ? n32 : n14452;
  assign n14454 = pi17 ? n32 : n14453;
  assign n14455 = pi16 ? n32 : n14454;
  assign n14456 = pi15 ? n13404 : n14455;
  assign n14457 = pi15 ? n14198 : n13409;
  assign n14458 = pi14 ? n14456 : n14457;
  assign n14459 = pi19 ? n1969 : ~n1490;
  assign n14460 = pi18 ? n32 : n14459;
  assign n14461 = pi17 ? n32 : n14460;
  assign n14462 = pi16 ? n32 : n14461;
  assign n14463 = pi20 ? n1076 : n321;
  assign n14464 = pi19 ? n1969 : ~n14463;
  assign n14465 = pi18 ? n32 : n14464;
  assign n14466 = pi17 ? n32 : n14465;
  assign n14467 = pi16 ? n32 : n14466;
  assign n14468 = pi15 ? n14462 : n14467;
  assign n14469 = pi19 ? n1969 : ~n10593;
  assign n14470 = pi18 ? n32 : n14469;
  assign n14471 = pi17 ? n32 : n14470;
  assign n14472 = pi16 ? n32 : n14471;
  assign n14473 = pi19 ? n1969 : ~n750;
  assign n14474 = pi18 ? n32 : n14473;
  assign n14475 = pi17 ? n32 : n14474;
  assign n14476 = pi16 ? n32 : n14475;
  assign n14477 = pi15 ? n14472 : n14476;
  assign n14478 = pi14 ? n14468 : n14477;
  assign n14479 = pi13 ? n14458 : n14478;
  assign n14480 = pi20 ? n1319 : n749;
  assign n14481 = pi19 ? n208 : ~n14480;
  assign n14482 = pi18 ? n32 : n14481;
  assign n14483 = pi17 ? n32 : n14482;
  assign n14484 = pi16 ? n32 : n14483;
  assign n14485 = pi19 ? n208 : ~n2317;
  assign n14486 = pi18 ? n32 : n14485;
  assign n14487 = pi17 ? n32 : n14486;
  assign n14488 = pi16 ? n32 : n14487;
  assign n14489 = pi15 ? n14484 : n14488;
  assign n14490 = pi21 ? n32 : ~n85;
  assign n14491 = pi20 ? n14490 : n749;
  assign n14492 = pi19 ? n244 : ~n14491;
  assign n14493 = pi18 ? n32 : n14492;
  assign n14494 = pi17 ? n32 : n14493;
  assign n14495 = pi16 ? n32 : n14494;
  assign n14496 = pi20 ? n151 : n243;
  assign n14497 = pi19 ? n244 : ~n14496;
  assign n14498 = pi18 ? n32 : n14497;
  assign n14499 = pi17 ? n32 : n14498;
  assign n14500 = pi16 ? n32 : n14499;
  assign n14501 = pi15 ? n14495 : n14500;
  assign n14502 = pi14 ? n14489 : n14501;
  assign n14503 = pi19 ? n244 : ~n11546;
  assign n14504 = pi18 ? n32 : n14503;
  assign n14505 = pi17 ? n32 : n14504;
  assign n14506 = pi16 ? n32 : n14505;
  assign n14507 = pi20 ? n1319 : ~n481;
  assign n14508 = pi19 ? n244 : ~n14507;
  assign n14509 = pi18 ? n32 : n14508;
  assign n14510 = pi17 ? n32 : n14509;
  assign n14511 = pi16 ? n32 : n14510;
  assign n14512 = pi15 ? n14506 : n14511;
  assign n14513 = pi22 ? n84 : n173;
  assign n14514 = pi21 ? n32 : ~n14513;
  assign n14515 = pi20 ? n14514 : n339;
  assign n14516 = pi19 ? n244 : ~n14515;
  assign n14517 = pi18 ? n32 : n14516;
  assign n14518 = pi17 ? n32 : n14517;
  assign n14519 = pi16 ? n32 : n14518;
  assign n14520 = pi22 ? n84 : ~n173;
  assign n14521 = pi21 ? n32 : ~n14520;
  assign n14522 = pi20 ? n14521 : ~n32;
  assign n14523 = pi19 ? n244 : ~n14522;
  assign n14524 = pi18 ? n32 : n14523;
  assign n14525 = pi17 ? n32 : n14524;
  assign n14526 = pi16 ? n32 : n14525;
  assign n14527 = pi15 ? n14519 : n14526;
  assign n14528 = pi14 ? n14512 : n14527;
  assign n14529 = pi13 ? n14502 : n14528;
  assign n14530 = pi12 ? n14479 : n14529;
  assign n14531 = pi11 ? n14451 : n14530;
  assign n14532 = pi21 ? n32 : ~n84;
  assign n14533 = pi20 ? n14532 : ~n32;
  assign n14534 = pi19 ? n244 : ~n14533;
  assign n14535 = pi18 ? n32 : n14534;
  assign n14536 = pi17 ? n32 : n14535;
  assign n14537 = pi16 ? n32 : n14536;
  assign n14538 = pi19 ? n244 : ~n12020;
  assign n14539 = pi18 ? n32 : n14538;
  assign n14540 = pi17 ? n32 : n14539;
  assign n14541 = pi16 ? n32 : n14540;
  assign n14542 = pi15 ? n14537 : n14541;
  assign n14543 = pi22 ? n84 : ~n34;
  assign n14544 = pi21 ? n32 : ~n14543;
  assign n14545 = pi20 ? n14544 : ~n32;
  assign n14546 = pi19 ? n244 : ~n14545;
  assign n14547 = pi18 ? n32 : n14546;
  assign n14548 = pi17 ? n32 : n14547;
  assign n14549 = pi16 ? n32 : n14548;
  assign n14550 = pi15 ? n14549 : n14219;
  assign n14551 = pi14 ? n14542 : n14550;
  assign n14552 = pi20 ? n14490 : ~n32;
  assign n14553 = pi19 ? n208 : ~n14552;
  assign n14554 = pi18 ? n32 : n14553;
  assign n14555 = pi17 ? n32 : n14554;
  assign n14556 = pi16 ? n32 : n14555;
  assign n14557 = pi19 ? n340 : ~n813;
  assign n14558 = pi18 ? n32 : n14557;
  assign n14559 = pi17 ? n32 : n14558;
  assign n14560 = pi16 ? n32 : n14559;
  assign n14561 = pi14 ? n14556 : n14560;
  assign n14562 = pi13 ? n14551 : n14561;
  assign n14563 = pi19 ? n244 : ~n1812;
  assign n14564 = pi18 ? n32 : n14563;
  assign n14565 = pi17 ? n32 : n14564;
  assign n14566 = pi16 ? n32 : n14565;
  assign n14567 = pi19 ? n208 : ~n813;
  assign n14568 = pi18 ? n32 : n14567;
  assign n14569 = pi17 ? n32 : n14568;
  assign n14570 = pi16 ? n32 : n14569;
  assign n14571 = pi15 ? n14566 : n14570;
  assign n14572 = pi19 ? n208 : ~n1941;
  assign n14573 = pi18 ? n32 : n14572;
  assign n14574 = pi17 ? n32 : n14573;
  assign n14575 = pi16 ? n32 : n14574;
  assign n14576 = pi15 ? n14570 : n14575;
  assign n14577 = pi14 ? n14571 : n14576;
  assign n14578 = pi18 ? n32 : n6147;
  assign n14579 = pi17 ? n32 : n14578;
  assign n14580 = pi16 ? n32 : n14579;
  assign n14581 = pi19 ? n1969 : n32;
  assign n14582 = pi18 ? n32 : n14581;
  assign n14583 = pi17 ? n32 : n14582;
  assign n14584 = pi16 ? n32 : n14583;
  assign n14585 = pi15 ? n14580 : n14584;
  assign n14586 = pi14 ? n14580 : n14585;
  assign n14587 = pi13 ? n14577 : n14586;
  assign n14588 = pi12 ? n14562 : n14587;
  assign n14589 = pi20 ? n32 : n10644;
  assign n14590 = pi19 ? n14589 : n32;
  assign n14591 = pi18 ? n32 : n14590;
  assign n14592 = pi17 ? n32 : n14591;
  assign n14593 = pi16 ? n32 : n14592;
  assign n14594 = pi21 ? n1939 : ~n1939;
  assign n14595 = pi20 ? n32 : n14594;
  assign n14596 = pi19 ? n14595 : n32;
  assign n14597 = pi18 ? n32 : n14596;
  assign n14598 = pi17 ? n32 : n14597;
  assign n14599 = pi16 ? n32 : n14598;
  assign n14600 = pi15 ? n14593 : n14599;
  assign n14601 = pi21 ? n405 : ~n1939;
  assign n14602 = pi20 ? n32 : n14601;
  assign n14603 = pi19 ? n14602 : n32;
  assign n14604 = pi18 ? n32 : n14603;
  assign n14605 = pi17 ? n32 : n14604;
  assign n14606 = pi16 ? n32 : n14605;
  assign n14607 = pi15 ? n14606 : n658;
  assign n14608 = pi14 ? n14600 : n14607;
  assign n14609 = pi20 ? n32 : n6229;
  assign n14610 = pi19 ? n14609 : n32;
  assign n14611 = pi18 ? n32 : n14610;
  assign n14612 = pi17 ? n32 : n14611;
  assign n14613 = pi16 ? n32 : n14612;
  assign n14614 = pi14 ? n658 : n14613;
  assign n14615 = pi13 ? n14608 : n14614;
  assign n14616 = pi12 ? n14615 : n32;
  assign n14617 = pi11 ? n14588 : n14616;
  assign n14618 = pi10 ? n14531 : n14617;
  assign n14619 = pi09 ? n14422 : n14618;
  assign n14620 = pi19 ? n594 : ~n531;
  assign n14621 = pi18 ? n32 : n14620;
  assign n14622 = pi17 ? n32 : n14621;
  assign n14623 = pi16 ? n32 : n14622;
  assign n14624 = pi15 ? n32 : n14623;
  assign n14625 = pi14 ? n14624 : n14623;
  assign n14626 = pi13 ? n32 : n14625;
  assign n14627 = pi12 ? n32 : n14626;
  assign n14628 = pi11 ? n32 : n14627;
  assign n14629 = pi10 ? n32 : n14628;
  assign n14630 = pi19 ? n2141 : ~n531;
  assign n14631 = pi18 ? n32 : n14630;
  assign n14632 = pi17 ? n32 : n14631;
  assign n14633 = pi16 ? n32 : n14632;
  assign n14634 = pi15 ? n14633 : n14416;
  assign n14635 = pi15 ? n14416 : n14179;
  assign n14636 = pi14 ? n14634 : n14635;
  assign n14637 = pi19 ? n1840 : ~n322;
  assign n14638 = pi18 ? n32 : n14637;
  assign n14639 = pi17 ? n32 : n14638;
  assign n14640 = pi16 ? n32 : n14639;
  assign n14641 = pi14 ? n13968 : n14640;
  assign n14642 = pi13 ? n14636 : n14641;
  assign n14643 = pi19 ? n322 : ~n9001;
  assign n14644 = pi18 ? n32 : n14643;
  assign n14645 = pi17 ? n32 : n14644;
  assign n14646 = pi16 ? n32 : n14645;
  assign n14647 = pi15 ? n13978 : n14646;
  assign n14648 = pi19 ? n322 : ~n343;
  assign n14649 = pi18 ? n32 : n14648;
  assign n14650 = pi17 ? n32 : n14649;
  assign n14651 = pi16 ? n32 : n14650;
  assign n14652 = pi15 ? n14651 : n13978;
  assign n14653 = pi14 ? n14647 : n14652;
  assign n14654 = pi13 ? n14640 : n14653;
  assign n14655 = pi12 ? n14642 : n14654;
  assign n14656 = pi19 ? n1476 : ~n11027;
  assign n14657 = pi18 ? n32 : n14656;
  assign n14658 = pi17 ? n32 : n14657;
  assign n14659 = pi16 ? n32 : n14658;
  assign n14660 = pi15 ? n13695 : n14659;
  assign n14661 = pi20 ? n32 : ~n564;
  assign n14662 = pi19 ? n1476 : ~n14661;
  assign n14663 = pi18 ? n32 : n14662;
  assign n14664 = pi17 ? n32 : n14663;
  assign n14665 = pi16 ? n32 : n14664;
  assign n14666 = pi15 ? n14665 : n13700;
  assign n14667 = pi14 ? n14660 : n14666;
  assign n14668 = pi19 ? n1476 : ~n1490;
  assign n14669 = pi18 ? n32 : n14668;
  assign n14670 = pi17 ? n32 : n14669;
  assign n14671 = pi16 ? n32 : n14670;
  assign n14672 = pi19 ? n1476 : ~n321;
  assign n14673 = pi18 ? n32 : n14672;
  assign n14674 = pi17 ? n32 : n14673;
  assign n14675 = pi16 ? n32 : n14674;
  assign n14676 = pi15 ? n14671 : n14675;
  assign n14677 = pi19 ? n1476 : ~n10593;
  assign n14678 = pi18 ? n32 : n14677;
  assign n14679 = pi17 ? n32 : n14678;
  assign n14680 = pi16 ? n32 : n14679;
  assign n14681 = pi19 ? n1476 : ~n750;
  assign n14682 = pi18 ? n32 : n14681;
  assign n14683 = pi17 ? n32 : n14682;
  assign n14684 = pi16 ? n32 : n14683;
  assign n14685 = pi15 ? n14680 : n14684;
  assign n14686 = pi14 ? n14676 : n14685;
  assign n14687 = pi13 ? n14667 : n14686;
  assign n14688 = pi20 ? n321 : n749;
  assign n14689 = pi19 ? n750 : ~n14688;
  assign n14690 = pi18 ? n32 : n14689;
  assign n14691 = pi17 ? n32 : n14690;
  assign n14692 = pi16 ? n32 : n14691;
  assign n14693 = pi19 ? n750 : ~n589;
  assign n14694 = pi18 ? n32 : n14693;
  assign n14695 = pi17 ? n32 : n14694;
  assign n14696 = pi16 ? n32 : n14695;
  assign n14697 = pi15 ? n14692 : n14696;
  assign n14698 = pi20 ? n1076 : n749;
  assign n14699 = pi19 ? n750 : ~n14698;
  assign n14700 = pi18 ? n32 : n14699;
  assign n14701 = pi17 ? n32 : n14700;
  assign n14702 = pi16 ? n32 : n14701;
  assign n14703 = pi19 ? n750 : ~n14275;
  assign n14704 = pi18 ? n32 : n14703;
  assign n14705 = pi17 ? n32 : n14704;
  assign n14706 = pi16 ? n32 : n14705;
  assign n14707 = pi15 ? n14702 : n14706;
  assign n14708 = pi14 ? n14697 : n14707;
  assign n14709 = pi19 ? n750 : ~n14552;
  assign n14710 = pi18 ? n32 : n14709;
  assign n14711 = pi17 ? n32 : n14710;
  assign n14712 = pi16 ? n32 : n14711;
  assign n14713 = pi15 ? n14712 : n14696;
  assign n14714 = pi20 ? n14514 : n243;
  assign n14715 = pi19 ? n1969 : ~n14714;
  assign n14716 = pi18 ? n32 : n14715;
  assign n14717 = pi17 ? n32 : n14716;
  assign n14718 = pi16 ? n32 : n14717;
  assign n14719 = pi19 ? n750 : ~n6042;
  assign n14720 = pi18 ? n32 : n14719;
  assign n14721 = pi17 ? n32 : n14720;
  assign n14722 = pi16 ? n32 : n14721;
  assign n14723 = pi15 ? n14718 : n14722;
  assign n14724 = pi14 ? n14713 : n14723;
  assign n14725 = pi13 ? n14708 : n14724;
  assign n14726 = pi12 ? n14687 : n14725;
  assign n14727 = pi11 ? n14655 : n14726;
  assign n14728 = pi19 ? n1969 : ~n14533;
  assign n14729 = pi18 ? n32 : n14728;
  assign n14730 = pi17 ? n32 : n14729;
  assign n14731 = pi16 ? n32 : n14730;
  assign n14732 = pi19 ? n750 : ~n12020;
  assign n14733 = pi18 ? n32 : n14732;
  assign n14734 = pi17 ? n32 : n14733;
  assign n14735 = pi16 ? n32 : n14734;
  assign n14736 = pi15 ? n14731 : n14735;
  assign n14737 = pi19 ? n1969 : ~n14545;
  assign n14738 = pi18 ? n32 : n14737;
  assign n14739 = pi17 ? n32 : n14738;
  assign n14740 = pi16 ? n32 : n14739;
  assign n14741 = pi19 ? n1969 : ~n2317;
  assign n14742 = pi18 ? n32 : n14741;
  assign n14743 = pi17 ? n32 : n14742;
  assign n14744 = pi16 ? n32 : n14743;
  assign n14745 = pi15 ? n14740 : n14744;
  assign n14746 = pi14 ? n14736 : n14745;
  assign n14747 = pi19 ? n1969 : ~n349;
  assign n14748 = pi18 ? n32 : n14747;
  assign n14749 = pi17 ? n32 : n14748;
  assign n14750 = pi16 ? n32 : n14749;
  assign n14751 = pi19 ? n1969 : ~n813;
  assign n14752 = pi18 ? n32 : n14751;
  assign n14753 = pi17 ? n32 : n14752;
  assign n14754 = pi16 ? n32 : n14753;
  assign n14755 = pi19 ? n750 : ~n1812;
  assign n14756 = pi18 ? n32 : n14755;
  assign n14757 = pi17 ? n32 : n14756;
  assign n14758 = pi16 ? n32 : n14757;
  assign n14759 = pi15 ? n14754 : n14758;
  assign n14760 = pi14 ? n14750 : n14759;
  assign n14761 = pi13 ? n14746 : n14760;
  assign n14762 = pi19 ? n750 : ~n1941;
  assign n14763 = pi18 ? n32 : n14762;
  assign n14764 = pi17 ? n32 : n14763;
  assign n14765 = pi16 ? n32 : n14764;
  assign n14766 = pi19 ? n1476 : ~n617;
  assign n14767 = pi18 ? n32 : n14766;
  assign n14768 = pi17 ? n32 : n14767;
  assign n14769 = pi16 ? n32 : n14768;
  assign n14770 = pi15 ? n14765 : n14769;
  assign n14771 = pi14 ? n14759 : n14770;
  assign n14772 = pi19 ? n1476 : n32;
  assign n14773 = pi18 ? n32 : n14772;
  assign n14774 = pi17 ? n32 : n14773;
  assign n14775 = pi16 ? n32 : n14774;
  assign n14776 = pi15 ? n14769 : n14775;
  assign n14777 = pi14 ? n14769 : n14776;
  assign n14778 = pi13 ? n14771 : n14777;
  assign n14779 = pi12 ? n14761 : n14778;
  assign n14780 = pi21 ? n100 : ~n405;
  assign n14781 = pi20 ? n32 : n14780;
  assign n14782 = pi19 ? n14781 : n32;
  assign n14783 = pi18 ? n32 : n14782;
  assign n14784 = pi17 ? n32 : n14783;
  assign n14785 = pi16 ? n32 : n14784;
  assign n14786 = pi20 ? n32 : n7880;
  assign n14787 = pi19 ? n14786 : n32;
  assign n14788 = pi18 ? n32 : n14787;
  assign n14789 = pi17 ? n32 : n14788;
  assign n14790 = pi16 ? n32 : n14789;
  assign n14791 = pi15 ? n14785 : n14790;
  assign n14792 = pi22 ? n50 : ~n50;
  assign n14793 = pi21 ? n32 : n14792;
  assign n14794 = pi20 ? n32 : n14793;
  assign n14795 = pi19 ? n14794 : n32;
  assign n14796 = pi18 ? n32 : n14795;
  assign n14797 = pi17 ? n32 : n14796;
  assign n14798 = pi16 ? n32 : n14797;
  assign n14799 = pi15 ? n14798 : n32;
  assign n14800 = pi14 ? n14791 : n14799;
  assign n14801 = pi13 ? n14800 : n32;
  assign n14802 = pi12 ? n14801 : n32;
  assign n14803 = pi11 ? n14779 : n14802;
  assign n14804 = pi10 ? n14727 : n14803;
  assign n14805 = pi09 ? n14629 : n14804;
  assign n14806 = pi08 ? n14619 : n14805;
  assign n14807 = pi07 ? n14412 : n14806;
  assign n14808 = pi15 ? n14623 : n14633;
  assign n14809 = pi14 ? n14808 : n14416;
  assign n14810 = pi19 ? n1320 : ~n322;
  assign n14811 = pi18 ? n32 : n14810;
  assign n14812 = pi17 ? n32 : n14811;
  assign n14813 = pi16 ? n32 : n14812;
  assign n14814 = pi14 ? n14426 : n14813;
  assign n14815 = pi13 ? n14809 : n14814;
  assign n14816 = pi19 ? n519 : ~n1490;
  assign n14817 = pi18 ? n32 : n14816;
  assign n14818 = pi17 ? n32 : n14817;
  assign n14819 = pi16 ? n32 : n14818;
  assign n14820 = pi19 ? n519 : ~n322;
  assign n14821 = pi18 ? n32 : n14820;
  assign n14822 = pi17 ? n32 : n14821;
  assign n14823 = pi16 ? n32 : n14822;
  assign n14824 = pi15 ? n14819 : n14823;
  assign n14825 = pi14 ? n14824 : n14823;
  assign n14826 = pi20 ? n32 : ~n9013;
  assign n14827 = pi19 ? n1840 : ~n14826;
  assign n14828 = pi18 ? n32 : n14827;
  assign n14829 = pi17 ? n32 : n14828;
  assign n14830 = pi16 ? n32 : n14829;
  assign n14831 = pi15 ? n13968 : n14830;
  assign n14832 = pi19 ? n1840 : ~n365;
  assign n14833 = pi18 ? n32 : n14832;
  assign n14834 = pi17 ? n32 : n14833;
  assign n14835 = pi16 ? n32 : n14834;
  assign n14836 = pi15 ? n13968 : n14835;
  assign n14837 = pi14 ? n14831 : n14836;
  assign n14838 = pi13 ? n14825 : n14837;
  assign n14839 = pi12 ? n14815 : n14838;
  assign n14840 = pi19 ? n1840 : ~n12171;
  assign n14841 = pi18 ? n32 : n14840;
  assign n14842 = pi17 ? n32 : n14841;
  assign n14843 = pi16 ? n32 : n14842;
  assign n14844 = pi21 ? n1009 : ~n32;
  assign n14845 = pi20 ? n32 : n14844;
  assign n14846 = pi19 ? n1840 : ~n14845;
  assign n14847 = pi18 ? n32 : n14846;
  assign n14848 = pi17 ? n32 : n14847;
  assign n14849 = pi16 ? n32 : n14848;
  assign n14850 = pi15 ? n14843 : n14849;
  assign n14851 = pi19 ? n1840 : ~n11938;
  assign n14852 = pi18 ? n32 : n14851;
  assign n14853 = pi17 ? n32 : n14852;
  assign n14854 = pi16 ? n32 : n14853;
  assign n14855 = pi19 ? n1840 : ~n1490;
  assign n14856 = pi18 ? n32 : n14855;
  assign n14857 = pi17 ? n32 : n14856;
  assign n14858 = pi16 ? n32 : n14857;
  assign n14859 = pi15 ? n14854 : n14858;
  assign n14860 = pi14 ? n14850 : n14859;
  assign n14861 = pi20 ? n32 : ~n7487;
  assign n14862 = pi19 ? n1840 : ~n14861;
  assign n14863 = pi18 ? n32 : n14862;
  assign n14864 = pi17 ? n32 : n14863;
  assign n14865 = pi16 ? n32 : n14864;
  assign n14866 = pi19 ? n1840 : ~n750;
  assign n14867 = pi18 ? n32 : n14866;
  assign n14868 = pi17 ? n32 : n14867;
  assign n14869 = pi16 ? n32 : n14868;
  assign n14870 = pi15 ? n14865 : n14869;
  assign n14871 = pi14 ? n14640 : n14870;
  assign n14872 = pi13 ? n14860 : n14871;
  assign n14873 = pi19 ? n322 : ~n208;
  assign n14874 = pi18 ? n32 : n14873;
  assign n14875 = pi17 ? n32 : n14874;
  assign n14876 = pi16 ? n32 : n14875;
  assign n14877 = pi20 ? n342 : n749;
  assign n14878 = pi19 ? n322 : ~n14877;
  assign n14879 = pi18 ? n32 : n14878;
  assign n14880 = pi17 ? n32 : n14879;
  assign n14881 = pi16 ? n32 : n14880;
  assign n14882 = pi19 ? n322 : ~n14496;
  assign n14883 = pi18 ? n32 : n14882;
  assign n14884 = pi17 ? n32 : n14883;
  assign n14885 = pi16 ? n32 : n14884;
  assign n14886 = pi15 ? n14881 : n14885;
  assign n14887 = pi14 ? n14876 : n14886;
  assign n14888 = pi19 ? n322 : ~n11991;
  assign n14889 = pi18 ? n32 : n14888;
  assign n14890 = pi17 ? n32 : n14889;
  assign n14891 = pi16 ? n32 : n14890;
  assign n14892 = pi19 ? n322 : ~n429;
  assign n14893 = pi18 ? n32 : n14892;
  assign n14894 = pi17 ? n32 : n14893;
  assign n14895 = pi16 ? n32 : n14894;
  assign n14896 = pi15 ? n14891 : n14895;
  assign n14897 = pi19 ? n322 : ~n244;
  assign n14898 = pi18 ? n32 : n14897;
  assign n14899 = pi17 ? n32 : n14898;
  assign n14900 = pi16 ? n32 : n14899;
  assign n14901 = pi15 ? n14900 : n14895;
  assign n14902 = pi14 ? n14896 : n14901;
  assign n14903 = pi13 ? n14887 : n14902;
  assign n14904 = pi12 ? n14872 : n14903;
  assign n14905 = pi11 ? n14839 : n14904;
  assign n14906 = pi19 ? n322 : ~n2297;
  assign n14907 = pi18 ? n32 : n14906;
  assign n14908 = pi17 ? n32 : n14907;
  assign n14909 = pi16 ? n32 : n14908;
  assign n14910 = pi19 ? n322 : ~n12020;
  assign n14911 = pi18 ? n32 : n14910;
  assign n14912 = pi17 ? n32 : n14911;
  assign n14913 = pi16 ? n32 : n14912;
  assign n14914 = pi15 ? n14909 : n14913;
  assign n14915 = pi18 ? n32 : n6581;
  assign n14916 = pi17 ? n32 : n14915;
  assign n14917 = pi16 ? n32 : n14916;
  assign n14918 = pi15 ? n14895 : n14917;
  assign n14919 = pi14 ? n14914 : n14918;
  assign n14920 = pi19 ? n322 : ~n14552;
  assign n14921 = pi18 ? n32 : n14920;
  assign n14922 = pi17 ? n32 : n14921;
  assign n14923 = pi16 ? n32 : n14922;
  assign n14924 = pi15 ? n14651 : n14923;
  assign n14925 = pi19 ? n1476 : ~n589;
  assign n14926 = pi18 ? n32 : n14925;
  assign n14927 = pi17 ? n32 : n14926;
  assign n14928 = pi16 ? n32 : n14927;
  assign n14929 = pi19 ? n1476 : ~n1812;
  assign n14930 = pi18 ? n32 : n14929;
  assign n14931 = pi17 ? n32 : n14930;
  assign n14932 = pi16 ? n32 : n14931;
  assign n14933 = pi15 ? n14928 : n14932;
  assign n14934 = pi14 ? n14924 : n14933;
  assign n14935 = pi13 ? n14919 : n14934;
  assign n14936 = pi21 ? n32 : ~n66;
  assign n14937 = pi20 ? n32 : n14936;
  assign n14938 = pi19 ? n14937 : ~n1941;
  assign n14939 = pi18 ? n32 : n14938;
  assign n14940 = pi17 ? n32 : n14939;
  assign n14941 = pi16 ? n32 : n14940;
  assign n14942 = pi19 ? n1840 : ~n617;
  assign n14943 = pi18 ? n32 : n14942;
  assign n14944 = pi17 ? n32 : n14943;
  assign n14945 = pi16 ? n32 : n14944;
  assign n14946 = pi15 ? n14941 : n14945;
  assign n14947 = pi14 ? n14932 : n14946;
  assign n14948 = pi19 ? n519 : ~n617;
  assign n14949 = pi18 ? n32 : n14948;
  assign n14950 = pi17 ? n32 : n14949;
  assign n14951 = pi16 ? n32 : n14950;
  assign n14952 = pi15 ? n14945 : n14951;
  assign n14953 = pi21 ? n32 : n631;
  assign n14954 = pi20 ? n32 : n14953;
  assign n14955 = pi19 ? n14954 : n32;
  assign n14956 = pi18 ? n32 : n14955;
  assign n14957 = pi17 ? n32 : n14956;
  assign n14958 = pi16 ? n32 : n14957;
  assign n14959 = pi15 ? n14958 : n14798;
  assign n14960 = pi14 ? n14952 : n14959;
  assign n14961 = pi13 ? n14947 : n14960;
  assign n14962 = pi12 ? n14935 : n14961;
  assign n14963 = pi20 ? n32 : n14286;
  assign n14964 = pi19 ? n14963 : n32;
  assign n14965 = pi18 ? n32 : n14964;
  assign n14966 = pi17 ? n32 : n14965;
  assign n14967 = pi16 ? n32 : n14966;
  assign n14968 = pi21 ? n32 : n7500;
  assign n14969 = pi20 ? n32 : n14968;
  assign n14970 = pi19 ? n14969 : n32;
  assign n14971 = pi18 ? n32 : n14970;
  assign n14972 = pi17 ? n32 : n14971;
  assign n14973 = pi16 ? n32 : n14972;
  assign n14974 = pi15 ? n14967 : n14973;
  assign n14975 = pi15 ? n14973 : n32;
  assign n14976 = pi14 ? n14974 : n14975;
  assign n14977 = pi13 ? n14976 : n32;
  assign n14978 = pi12 ? n14977 : n32;
  assign n14979 = pi11 ? n14962 : n14978;
  assign n14980 = pi10 ? n14905 : n14979;
  assign n14981 = pi09 ? n14629 : n14980;
  assign n14982 = pi19 ? n32 : ~n531;
  assign n14983 = pi18 ? n32 : n14982;
  assign n14984 = pi17 ? n32 : n14983;
  assign n14985 = pi16 ? n32 : n14984;
  assign n14986 = pi15 ? n32 : n14985;
  assign n14987 = pi14 ? n14986 : n14985;
  assign n14988 = pi13 ? n32 : n14987;
  assign n14989 = pi12 ? n32 : n14988;
  assign n14990 = pi11 ? n32 : n14989;
  assign n14991 = pi10 ? n32 : n14990;
  assign n14992 = pi19 ? n1574 : ~n531;
  assign n14993 = pi18 ? n32 : n14992;
  assign n14994 = pi17 ? n32 : n14993;
  assign n14995 = pi16 ? n32 : n14994;
  assign n14996 = pi15 ? n14995 : n14623;
  assign n14997 = pi14 ? n14996 : n14633;
  assign n14998 = pi19 ? n2141 : ~n322;
  assign n14999 = pi18 ? n32 : n14998;
  assign n15000 = pi17 ? n32 : n14999;
  assign n15001 = pi16 ? n32 : n15000;
  assign n15002 = pi14 ? n14633 : n15001;
  assign n15003 = pi13 ? n14997 : n15002;
  assign n15004 = pi19 ? n507 : ~n1490;
  assign n15005 = pi18 ? n32 : n15004;
  assign n15006 = pi17 ? n32 : n15005;
  assign n15007 = pi16 ? n32 : n15006;
  assign n15008 = pi19 ? n507 : ~n322;
  assign n15009 = pi18 ? n32 : n15008;
  assign n15010 = pi17 ? n32 : n15009;
  assign n15011 = pi16 ? n32 : n15010;
  assign n15012 = pi15 ? n15007 : n15011;
  assign n15013 = pi14 ? n15012 : n15011;
  assign n15014 = pi19 ? n1320 : ~n365;
  assign n15015 = pi18 ? n32 : n15014;
  assign n15016 = pi17 ? n32 : n15015;
  assign n15017 = pi16 ? n32 : n15016;
  assign n15018 = pi14 ? n14426 : n15017;
  assign n15019 = pi13 ? n15013 : n15018;
  assign n15020 = pi12 ? n15003 : n15019;
  assign n15021 = pi19 ? n519 : ~n12171;
  assign n15022 = pi18 ? n32 : n15021;
  assign n15023 = pi17 ? n32 : n15022;
  assign n15024 = pi16 ? n32 : n15023;
  assign n15025 = pi19 ? n519 : ~n14845;
  assign n15026 = pi18 ? n32 : n15025;
  assign n15027 = pi17 ? n32 : n15026;
  assign n15028 = pi16 ? n32 : n15027;
  assign n15029 = pi15 ? n15024 : n15028;
  assign n15030 = pi15 ? n14179 : n14819;
  assign n15031 = pi14 ? n15029 : n15030;
  assign n15032 = pi19 ? n519 : ~n14861;
  assign n15033 = pi18 ? n32 : n15032;
  assign n15034 = pi17 ? n32 : n15033;
  assign n15035 = pi16 ? n32 : n15034;
  assign n15036 = pi19 ? n519 : ~n750;
  assign n15037 = pi18 ? n32 : n15036;
  assign n15038 = pi17 ? n32 : n15037;
  assign n15039 = pi16 ? n32 : n15038;
  assign n15040 = pi15 ? n15035 : n15039;
  assign n15041 = pi14 ? n14823 : n15040;
  assign n15042 = pi13 ? n15031 : n15041;
  assign n15043 = pi19 ? n519 : ~n208;
  assign n15044 = pi18 ? n32 : n15043;
  assign n15045 = pi17 ? n32 : n15044;
  assign n15046 = pi16 ? n32 : n15045;
  assign n15047 = pi19 ? n519 : ~n1740;
  assign n15048 = pi18 ? n32 : n15047;
  assign n15049 = pi17 ? n32 : n15048;
  assign n15050 = pi16 ? n32 : n15049;
  assign n15051 = pi20 ? n3523 : n243;
  assign n15052 = pi19 ? n1840 : ~n15051;
  assign n15053 = pi18 ? n32 : n15052;
  assign n15054 = pi17 ? n32 : n15053;
  assign n15055 = pi16 ? n32 : n15054;
  assign n15056 = pi15 ? n15050 : n15055;
  assign n15057 = pi14 ? n15046 : n15056;
  assign n15058 = pi19 ? n519 : ~n12957;
  assign n15059 = pi18 ? n32 : n15058;
  assign n15060 = pi17 ? n32 : n15059;
  assign n15061 = pi16 ? n32 : n15060;
  assign n15062 = pi15 ? n14179 : n15061;
  assign n15063 = pi19 ? n519 : ~n429;
  assign n15064 = pi18 ? n32 : n15063;
  assign n15065 = pi17 ? n32 : n15064;
  assign n15066 = pi16 ? n32 : n15065;
  assign n15067 = pi15 ? n14179 : n15066;
  assign n15068 = pi14 ? n15062 : n15067;
  assign n15069 = pi13 ? n15057 : n15068;
  assign n15070 = pi12 ? n15042 : n15069;
  assign n15071 = pi11 ? n15020 : n15070;
  assign n15072 = pi19 ? n519 : ~n343;
  assign n15073 = pi18 ? n32 : n15072;
  assign n15074 = pi17 ? n32 : n15073;
  assign n15075 = pi16 ? n32 : n15074;
  assign n15076 = pi15 ? n15066 : n15075;
  assign n15077 = pi19 ? n519 : ~n349;
  assign n15078 = pi18 ? n32 : n15077;
  assign n15079 = pi17 ? n32 : n15078;
  assign n15080 = pi16 ? n32 : n15079;
  assign n15081 = pi15 ? n15075 : n15080;
  assign n15082 = pi14 ? n15076 : n15081;
  assign n15083 = pi19 ? n1840 : ~n349;
  assign n15084 = pi18 ? n32 : n15083;
  assign n15085 = pi17 ? n32 : n15084;
  assign n15086 = pi16 ? n32 : n15085;
  assign n15087 = pi19 ? n519 : ~n1812;
  assign n15088 = pi18 ? n32 : n15087;
  assign n15089 = pi17 ? n32 : n15088;
  assign n15090 = pi16 ? n32 : n15089;
  assign n15091 = pi15 ? n15086 : n15090;
  assign n15092 = pi14 ? n15081 : n15091;
  assign n15093 = pi13 ? n15082 : n15092;
  assign n15094 = pi22 ? n50 : ~n65;
  assign n15095 = pi21 ? n32 : n15094;
  assign n15096 = pi20 ? n32 : n15095;
  assign n15097 = pi19 ? n15096 : ~n1812;
  assign n15098 = pi18 ? n32 : n15097;
  assign n15099 = pi17 ? n32 : n15098;
  assign n15100 = pi16 ? n32 : n15099;
  assign n15101 = pi15 ? n15100 : n15090;
  assign n15102 = pi19 ? n519 : ~n1941;
  assign n15103 = pi18 ? n32 : n15102;
  assign n15104 = pi17 ? n32 : n15103;
  assign n15105 = pi16 ? n32 : n15104;
  assign n15106 = pi19 ? n519 : ~n2614;
  assign n15107 = pi18 ? n32 : n15106;
  assign n15108 = pi17 ? n32 : n15107;
  assign n15109 = pi16 ? n32 : n15108;
  assign n15110 = pi15 ? n15105 : n15109;
  assign n15111 = pi14 ? n15101 : n15110;
  assign n15112 = pi19 ? n1320 : ~n617;
  assign n15113 = pi18 ? n32 : n15112;
  assign n15114 = pi17 ? n32 : n15113;
  assign n15115 = pi16 ? n32 : n15114;
  assign n15116 = pi19 ? n507 : ~n617;
  assign n15117 = pi18 ? n32 : n15116;
  assign n15118 = pi17 ? n32 : n15117;
  assign n15119 = pi16 ? n32 : n15118;
  assign n15120 = pi15 ? n15115 : n15119;
  assign n15121 = pi18 ? n32 : n8106;
  assign n15122 = pi17 ? n32 : n15121;
  assign n15123 = pi16 ? n32 : n15122;
  assign n15124 = pi14 ? n15120 : n15123;
  assign n15125 = pi13 ? n15111 : n15124;
  assign n15126 = pi12 ? n15093 : n15125;
  assign n15127 = pi15 ? n15123 : n32;
  assign n15128 = pi14 ? n15127 : n32;
  assign n15129 = pi13 ? n15128 : n32;
  assign n15130 = pi12 ? n15129 : n32;
  assign n15131 = pi11 ? n15126 : n15130;
  assign n15132 = pi10 ? n15071 : n15131;
  assign n15133 = pi09 ? n14991 : n15132;
  assign n15134 = pi08 ? n14981 : n15133;
  assign n15135 = pi20 ? n339 : n32;
  assign n15136 = pi19 ? n32 : n15135;
  assign n15137 = pi18 ? n32 : n15136;
  assign n15138 = pi17 ? n32 : n15137;
  assign n15139 = pi16 ? n32 : n15138;
  assign n15140 = pi15 ? n32 : n15139;
  assign n15141 = pi14 ? n15140 : n15139;
  assign n15142 = pi13 ? n32 : n15141;
  assign n15143 = pi12 ? n32 : n15142;
  assign n15144 = pi11 ? n32 : n15143;
  assign n15145 = pi10 ? n32 : n15144;
  assign n15146 = pi20 ? n141 : n32;
  assign n15147 = pi19 ? n32 : n15146;
  assign n15148 = pi18 ? n32 : n15147;
  assign n15149 = pi17 ? n32 : n15148;
  assign n15150 = pi16 ? n32 : n15149;
  assign n15151 = pi15 ? n15150 : n14985;
  assign n15152 = pi14 ? n15151 : n14623;
  assign n15153 = pi13 ? n15152 : n15002;
  assign n15154 = pi19 ? n2141 : ~n1490;
  assign n15155 = pi18 ? n32 : n15154;
  assign n15156 = pi17 ? n32 : n15155;
  assign n15157 = pi16 ? n32 : n15156;
  assign n15158 = pi15 ? n15157 : n15001;
  assign n15159 = pi14 ? n15158 : n15001;
  assign n15160 = pi19 ? n2141 : ~n365;
  assign n15161 = pi18 ? n32 : n15160;
  assign n15162 = pi17 ? n32 : n15161;
  assign n15163 = pi16 ? n32 : n15162;
  assign n15164 = pi15 ? n15163 : n14633;
  assign n15165 = pi14 ? n14633 : n15164;
  assign n15166 = pi13 ? n15159 : n15165;
  assign n15167 = pi12 ? n15153 : n15166;
  assign n15168 = pi19 ? n507 : ~n11250;
  assign n15169 = pi18 ? n32 : n15168;
  assign n15170 = pi17 ? n32 : n15169;
  assign n15171 = pi16 ? n32 : n15170;
  assign n15172 = pi19 ? n507 : ~n14022;
  assign n15173 = pi18 ? n32 : n15172;
  assign n15174 = pi17 ? n32 : n15173;
  assign n15175 = pi16 ? n32 : n15174;
  assign n15176 = pi15 ? n15171 : n15175;
  assign n15177 = pi15 ? n14416 : n15007;
  assign n15178 = pi14 ? n15176 : n15177;
  assign n15179 = pi19 ? n507 : ~n519;
  assign n15180 = pi18 ? n32 : n15179;
  assign n15181 = pi17 ? n32 : n15180;
  assign n15182 = pi16 ? n32 : n15181;
  assign n15183 = pi19 ? n507 : ~n1840;
  assign n15184 = pi18 ? n32 : n15183;
  assign n15185 = pi17 ? n32 : n15184;
  assign n15186 = pi16 ? n32 : n15185;
  assign n15187 = pi15 ? n15182 : n15186;
  assign n15188 = pi19 ? n507 : ~n1476;
  assign n15189 = pi18 ? n32 : n15188;
  assign n15190 = pi17 ? n32 : n15189;
  assign n15191 = pi16 ? n32 : n15190;
  assign n15192 = pi15 ? n14416 : n15191;
  assign n15193 = pi14 ? n15187 : n15192;
  assign n15194 = pi13 ? n15178 : n15193;
  assign n15195 = pi19 ? n1320 : ~n1476;
  assign n15196 = pi18 ? n32 : n15195;
  assign n15197 = pi17 ? n32 : n15196;
  assign n15198 = pi16 ? n32 : n15197;
  assign n15199 = pi19 ? n1320 : ~n1740;
  assign n15200 = pi18 ? n32 : n15199;
  assign n15201 = pi17 ? n32 : n15200;
  assign n15202 = pi16 ? n32 : n15201;
  assign n15203 = pi19 ? n1320 : ~n244;
  assign n15204 = pi18 ? n32 : n15203;
  assign n15205 = pi17 ? n32 : n15204;
  assign n15206 = pi16 ? n32 : n15205;
  assign n15207 = pi15 ? n15202 : n15206;
  assign n15208 = pi14 ? n15198 : n15207;
  assign n15209 = pi19 ? n1320 : ~n343;
  assign n15210 = pi18 ? n32 : n15209;
  assign n15211 = pi17 ? n32 : n15210;
  assign n15212 = pi16 ? n32 : n15211;
  assign n15213 = pi15 ? n15212 : n14426;
  assign n15214 = pi14 ? n15206 : n15213;
  assign n15215 = pi13 ? n15208 : n15214;
  assign n15216 = pi12 ? n15194 : n15215;
  assign n15217 = pi11 ? n15167 : n15216;
  assign n15218 = pi19 ? n1320 : ~n2297;
  assign n15219 = pi18 ? n32 : n15218;
  assign n15220 = pi17 ? n32 : n15219;
  assign n15221 = pi16 ? n32 : n15220;
  assign n15222 = pi19 ? n507 : ~n1265;
  assign n15223 = pi18 ? n32 : n15222;
  assign n15224 = pi17 ? n32 : n15223;
  assign n15225 = pi16 ? n32 : n15224;
  assign n15226 = pi15 ? n15221 : n15225;
  assign n15227 = pi19 ? n507 : ~n343;
  assign n15228 = pi18 ? n32 : n15227;
  assign n15229 = pi17 ? n32 : n15228;
  assign n15230 = pi16 ? n32 : n15229;
  assign n15231 = pi14 ? n15226 : n15230;
  assign n15232 = pi19 ? n2141 : ~n343;
  assign n15233 = pi18 ? n32 : n15232;
  assign n15234 = pi17 ? n32 : n15233;
  assign n15235 = pi16 ? n32 : n15234;
  assign n15236 = pi19 ? n2141 : ~n589;
  assign n15237 = pi18 ? n32 : n15236;
  assign n15238 = pi17 ? n32 : n15237;
  assign n15239 = pi16 ? n32 : n15238;
  assign n15240 = pi15 ? n15235 : n15239;
  assign n15241 = pi19 ? n507 : ~n349;
  assign n15242 = pi18 ? n32 : n15241;
  assign n15243 = pi17 ? n32 : n15242;
  assign n15244 = pi16 ? n32 : n15243;
  assign n15245 = pi19 ? n507 : ~n1812;
  assign n15246 = pi18 ? n32 : n15245;
  assign n15247 = pi17 ? n32 : n15246;
  assign n15248 = pi16 ? n32 : n15247;
  assign n15249 = pi15 ? n15244 : n15248;
  assign n15250 = pi14 ? n15240 : n15249;
  assign n15251 = pi13 ? n15231 : n15250;
  assign n15252 = pi19 ? n507 : ~n2614;
  assign n15253 = pi18 ? n32 : n15252;
  assign n15254 = pi17 ? n32 : n15253;
  assign n15255 = pi16 ? n32 : n15254;
  assign n15256 = pi15 ? n15248 : n15255;
  assign n15257 = pi19 ? n2141 : ~n2614;
  assign n15258 = pi18 ? n32 : n15257;
  assign n15259 = pi17 ? n32 : n15258;
  assign n15260 = pi16 ? n32 : n15259;
  assign n15261 = pi15 ? n15260 : n15255;
  assign n15262 = pi14 ? n15256 : n15261;
  assign n15263 = pi16 ? n32 : n1788;
  assign n15264 = pi14 ? n15119 : n15263;
  assign n15265 = pi13 ? n15262 : n15264;
  assign n15266 = pi12 ? n15251 : n15265;
  assign n15267 = pi15 ? n15263 : n32;
  assign n15268 = pi14 ? n15267 : n32;
  assign n15269 = pi13 ? n15268 : n32;
  assign n15270 = pi12 ? n15269 : n32;
  assign n15271 = pi11 ? n15266 : n15270;
  assign n15272 = pi10 ? n15217 : n15271;
  assign n15273 = pi09 ? n15145 : n15272;
  assign n15274 = pi14 ? n15139 : n14985;
  assign n15275 = pi19 ? n1574 : ~n322;
  assign n15276 = pi18 ? n32 : n15275;
  assign n15277 = pi17 ? n32 : n15276;
  assign n15278 = pi16 ? n32 : n15277;
  assign n15279 = pi14 ? n14995 : n15278;
  assign n15280 = pi13 ? n15274 : n15279;
  assign n15281 = pi19 ? n594 : ~n1490;
  assign n15282 = pi18 ? n32 : n15281;
  assign n15283 = pi17 ? n32 : n15282;
  assign n15284 = pi16 ? n32 : n15283;
  assign n15285 = pi19 ? n594 : ~n322;
  assign n15286 = pi18 ? n32 : n15285;
  assign n15287 = pi17 ? n32 : n15286;
  assign n15288 = pi16 ? n32 : n15287;
  assign n15289 = pi15 ? n15284 : n15288;
  assign n15290 = pi14 ? n15289 : n15288;
  assign n15291 = pi13 ? n15290 : n14633;
  assign n15292 = pi12 ? n15280 : n15291;
  assign n15293 = pi19 ? n2141 : ~n507;
  assign n15294 = pi18 ? n32 : n15293;
  assign n15295 = pi17 ? n32 : n15294;
  assign n15296 = pi16 ? n32 : n15295;
  assign n15297 = pi19 ? n2141 : ~n14661;
  assign n15298 = pi18 ? n32 : n15297;
  assign n15299 = pi17 ? n32 : n15298;
  assign n15300 = pi16 ? n32 : n15299;
  assign n15301 = pi15 ? n15296 : n15300;
  assign n15302 = pi15 ? n15163 : n15157;
  assign n15303 = pi14 ? n15301 : n15302;
  assign n15304 = pi19 ? n2141 : ~n519;
  assign n15305 = pi18 ? n32 : n15304;
  assign n15306 = pi17 ? n32 : n15305;
  assign n15307 = pi16 ? n32 : n15306;
  assign n15308 = pi19 ? n2141 : ~n1840;
  assign n15309 = pi18 ? n32 : n15308;
  assign n15310 = pi17 ? n32 : n15309;
  assign n15311 = pi16 ? n32 : n15310;
  assign n15312 = pi15 ? n15307 : n15311;
  assign n15313 = pi19 ? n594 : ~n1476;
  assign n15314 = pi18 ? n32 : n15313;
  assign n15315 = pi17 ? n32 : n15314;
  assign n15316 = pi16 ? n32 : n15315;
  assign n15317 = pi15 ? n14623 : n15316;
  assign n15318 = pi14 ? n15312 : n15317;
  assign n15319 = pi13 ? n15303 : n15318;
  assign n15320 = pi19 ? n2141 : ~n1476;
  assign n15321 = pi18 ? n32 : n15320;
  assign n15322 = pi17 ? n32 : n15321;
  assign n15323 = pi16 ? n32 : n15322;
  assign n15324 = pi19 ? n2141 : ~n1740;
  assign n15325 = pi18 ? n32 : n15324;
  assign n15326 = pi17 ? n32 : n15325;
  assign n15327 = pi16 ? n32 : n15326;
  assign n15328 = pi19 ? n2141 : ~n244;
  assign n15329 = pi18 ? n32 : n15328;
  assign n15330 = pi17 ? n32 : n15329;
  assign n15331 = pi16 ? n32 : n15330;
  assign n15332 = pi15 ? n15327 : n15331;
  assign n15333 = pi14 ? n15323 : n15332;
  assign n15334 = pi19 ? n2141 : ~n340;
  assign n15335 = pi18 ? n32 : n15334;
  assign n15336 = pi17 ? n32 : n15335;
  assign n15337 = pi16 ? n32 : n15336;
  assign n15338 = pi15 ? n15331 : n15337;
  assign n15339 = pi15 ? n15235 : n14633;
  assign n15340 = pi14 ? n15338 : n15339;
  assign n15341 = pi13 ? n15333 : n15340;
  assign n15342 = pi12 ? n15319 : n15341;
  assign n15343 = pi11 ? n15292 : n15342;
  assign n15344 = pi19 ? n2141 : ~n2297;
  assign n15345 = pi18 ? n32 : n15344;
  assign n15346 = pi17 ? n32 : n15345;
  assign n15347 = pi16 ? n32 : n15346;
  assign n15348 = pi19 ? n2141 : ~n1265;
  assign n15349 = pi18 ? n32 : n15348;
  assign n15350 = pi17 ? n32 : n15349;
  assign n15351 = pi16 ? n32 : n15350;
  assign n15352 = pi15 ? n15347 : n15351;
  assign n15353 = pi14 ? n15352 : n15235;
  assign n15354 = pi19 ? n594 : ~n589;
  assign n15355 = pi18 ? n32 : n15354;
  assign n15356 = pi17 ? n32 : n15355;
  assign n15357 = pi16 ? n32 : n15356;
  assign n15358 = pi15 ? n15235 : n15357;
  assign n15359 = pi19 ? n594 : ~n349;
  assign n15360 = pi18 ? n32 : n15359;
  assign n15361 = pi17 ? n32 : n15360;
  assign n15362 = pi16 ? n32 : n15361;
  assign n15363 = pi19 ? n2141 : ~n1812;
  assign n15364 = pi18 ? n32 : n15363;
  assign n15365 = pi17 ? n32 : n15364;
  assign n15366 = pi16 ? n32 : n15365;
  assign n15367 = pi15 ? n15362 : n15366;
  assign n15368 = pi14 ? n15358 : n15367;
  assign n15369 = pi13 ? n15353 : n15368;
  assign n15370 = pi19 ? n11404 : ~n1812;
  assign n15371 = pi18 ? n32 : n15370;
  assign n15372 = pi17 ? n32 : n15371;
  assign n15373 = pi16 ? n32 : n15372;
  assign n15374 = pi19 ? n11404 : ~n2614;
  assign n15375 = pi18 ? n32 : n15374;
  assign n15376 = pi17 ? n32 : n15375;
  assign n15377 = pi16 ? n32 : n15376;
  assign n15378 = pi15 ? n15373 : n15377;
  assign n15379 = pi19 ? n1574 : ~n2614;
  assign n15380 = pi18 ? n32 : n15379;
  assign n15381 = pi17 ? n32 : n15380;
  assign n15382 = pi16 ? n32 : n15381;
  assign n15383 = pi19 ? n594 : ~n2614;
  assign n15384 = pi18 ? n32 : n15383;
  assign n15385 = pi17 ? n32 : n15384;
  assign n15386 = pi16 ? n32 : n15385;
  assign n15387 = pi15 ? n15382 : n15386;
  assign n15388 = pi14 ? n15378 : n15387;
  assign n15389 = pi16 ? n32 : n2081;
  assign n15390 = pi15 ? n15389 : n32;
  assign n15391 = pi14 ? n15390 : n32;
  assign n15392 = pi13 ? n15388 : n15391;
  assign n15393 = pi12 ? n15369 : n15392;
  assign n15394 = pi11 ? n15393 : n32;
  assign n15395 = pi10 ? n15343 : n15394;
  assign n15396 = pi09 ? n15145 : n15395;
  assign n15397 = pi08 ? n15273 : n15396;
  assign n15398 = pi07 ? n15134 : n15397;
  assign n15399 = pi06 ? n14807 : n15398;
  assign n15400 = pi19 ? n32 : n5707;
  assign n15401 = pi18 ? n32 : n15400;
  assign n15402 = pi17 ? n32 : n15401;
  assign n15403 = pi16 ? n32 : n15402;
  assign n15404 = pi15 ? n32 : n15403;
  assign n15405 = pi20 ? n207 : ~n321;
  assign n15406 = pi19 ? n32 : n15405;
  assign n15407 = pi18 ? n32 : n15406;
  assign n15408 = pi17 ? n32 : n15407;
  assign n15409 = pi16 ? n32 : n15408;
  assign n15410 = pi20 ? n243 : ~n321;
  assign n15411 = pi19 ? n32 : n15410;
  assign n15412 = pi18 ? n32 : n15411;
  assign n15413 = pi17 ? n32 : n15412;
  assign n15414 = pi16 ? n32 : n15413;
  assign n15415 = pi15 ? n15409 : n15414;
  assign n15416 = pi14 ? n15404 : n15415;
  assign n15417 = pi13 ? n32 : n15416;
  assign n15418 = pi12 ? n32 : n15417;
  assign n15419 = pi11 ? n32 : n15418;
  assign n15420 = pi10 ? n32 : n15419;
  assign n15421 = pi19 ? n32 : n6800;
  assign n15422 = pi18 ? n32 : n15421;
  assign n15423 = pi17 ? n32 : n15422;
  assign n15424 = pi16 ? n32 : n15423;
  assign n15425 = pi15 ? n15414 : n15424;
  assign n15426 = pi14 ? n15425 : n15139;
  assign n15427 = pi13 ? n15426 : n15150;
  assign n15428 = pi19 ? n1574 : ~n365;
  assign n15429 = pi18 ? n32 : n15428;
  assign n15430 = pi17 ? n32 : n15429;
  assign n15431 = pi16 ? n32 : n15430;
  assign n15432 = pi15 ? n14995 : n15431;
  assign n15433 = pi19 ? n1574 : ~n1508;
  assign n15434 = pi18 ? n32 : n15433;
  assign n15435 = pi17 ? n32 : n15434;
  assign n15436 = pi16 ? n32 : n15435;
  assign n15437 = pi15 ? n15436 : n15431;
  assign n15438 = pi14 ? n15432 : n15437;
  assign n15439 = pi13 ? n14985 : n15438;
  assign n15440 = pi12 ? n15427 : n15439;
  assign n15441 = pi19 ? n594 : ~n507;
  assign n15442 = pi18 ? n32 : n15441;
  assign n15443 = pi17 ? n32 : n15442;
  assign n15444 = pi16 ? n32 : n15443;
  assign n15445 = pi15 ? n15444 : n14623;
  assign n15446 = pi19 ? n594 : ~n14845;
  assign n15447 = pi18 ? n32 : n15446;
  assign n15448 = pi17 ? n32 : n15447;
  assign n15449 = pi16 ? n32 : n15448;
  assign n15450 = pi19 ? n594 : ~n365;
  assign n15451 = pi18 ? n32 : n15450;
  assign n15452 = pi17 ? n32 : n15451;
  assign n15453 = pi16 ? n32 : n15452;
  assign n15454 = pi15 ? n15449 : n15453;
  assign n15455 = pi14 ? n15445 : n15454;
  assign n15456 = pi19 ? n594 : ~n519;
  assign n15457 = pi18 ? n32 : n15456;
  assign n15458 = pi17 ? n32 : n15457;
  assign n15459 = pi16 ? n32 : n15458;
  assign n15460 = pi20 ? n32 : ~n6229;
  assign n15461 = pi19 ? n594 : ~n15460;
  assign n15462 = pi18 ? n32 : n15461;
  assign n15463 = pi17 ? n32 : n15462;
  assign n15464 = pi16 ? n32 : n15463;
  assign n15465 = pi15 ? n15459 : n15464;
  assign n15466 = pi19 ? n594 : ~n11972;
  assign n15467 = pi18 ? n32 : n15466;
  assign n15468 = pi17 ? n32 : n15467;
  assign n15469 = pi16 ? n32 : n15468;
  assign n15470 = pi15 ? n15469 : n15464;
  assign n15471 = pi14 ? n15465 : n15470;
  assign n15472 = pi13 ? n15455 : n15471;
  assign n15473 = pi19 ? n594 : ~n208;
  assign n15474 = pi18 ? n32 : n15473;
  assign n15475 = pi17 ? n32 : n15474;
  assign n15476 = pi16 ? n32 : n15475;
  assign n15477 = pi15 ? n15316 : n15476;
  assign n15478 = pi19 ? n594 : ~n11991;
  assign n15479 = pi18 ? n32 : n15478;
  assign n15480 = pi17 ? n32 : n15479;
  assign n15481 = pi16 ? n32 : n15480;
  assign n15482 = pi15 ? n14623 : n15481;
  assign n15483 = pi14 ? n15477 : n15482;
  assign n15484 = pi19 ? n594 : ~n340;
  assign n15485 = pi18 ? n32 : n15484;
  assign n15486 = pi17 ? n32 : n15485;
  assign n15487 = pi16 ? n32 : n15486;
  assign n15488 = pi15 ? n15487 : n14995;
  assign n15489 = pi15 ? n14623 : n14995;
  assign n15490 = pi14 ? n15488 : n15489;
  assign n15491 = pi13 ? n15483 : n15490;
  assign n15492 = pi12 ? n15472 : n15491;
  assign n15493 = pi11 ? n15440 : n15492;
  assign n15494 = pi19 ? n1574 : ~n429;
  assign n15495 = pi18 ? n32 : n15494;
  assign n15496 = pi17 ? n32 : n15495;
  assign n15497 = pi16 ? n32 : n15496;
  assign n15498 = pi19 ? n1574 : ~n343;
  assign n15499 = pi18 ? n32 : n15498;
  assign n15500 = pi17 ? n32 : n15499;
  assign n15501 = pi16 ? n32 : n15500;
  assign n15502 = pi15 ? n15497 : n15501;
  assign n15503 = pi14 ? n15502 : n15501;
  assign n15504 = pi19 ? n1574 : ~n349;
  assign n15505 = pi18 ? n32 : n15504;
  assign n15506 = pi17 ? n32 : n15505;
  assign n15507 = pi16 ? n32 : n15506;
  assign n15508 = pi19 ? n1574 : ~n1812;
  assign n15509 = pi18 ? n32 : n15508;
  assign n15510 = pi17 ? n32 : n15509;
  assign n15511 = pi16 ? n32 : n15510;
  assign n15512 = pi15 ? n15507 : n15511;
  assign n15513 = pi14 ? n15507 : n15512;
  assign n15514 = pi13 ? n15503 : n15513;
  assign n15515 = pi19 ? n32 : ~n2614;
  assign n15516 = pi18 ? n32 : n15515;
  assign n15517 = pi17 ? n32 : n15516;
  assign n15518 = pi16 ? n32 : n15517;
  assign n15519 = pi15 ? n15511 : n15518;
  assign n15520 = pi15 ? n15518 : n15382;
  assign n15521 = pi14 ? n15519 : n15520;
  assign n15522 = pi13 ? n15521 : n32;
  assign n15523 = pi12 ? n15514 : n15522;
  assign n15524 = pi11 ? n15523 : n32;
  assign n15525 = pi10 ? n15493 : n15524;
  assign n15526 = pi09 ? n15420 : n15525;
  assign n15527 = pi20 ? n749 : n32;
  assign n15528 = pi19 ? n32 : n15527;
  assign n15529 = pi18 ? n32 : n15528;
  assign n15530 = pi17 ? n32 : n15529;
  assign n15531 = pi16 ? n32 : n15530;
  assign n15532 = pi15 ? n32 : n15531;
  assign n15533 = pi20 ? n749 : ~n321;
  assign n15534 = pi19 ? n32 : n15533;
  assign n15535 = pi18 ? n32 : n15534;
  assign n15536 = pi17 ? n32 : n15535;
  assign n15537 = pi16 ? n32 : n15536;
  assign n15538 = pi14 ? n15532 : n15537;
  assign n15539 = pi13 ? n32 : n15538;
  assign n15540 = pi12 ? n32 : n15539;
  assign n15541 = pi11 ? n32 : n15540;
  assign n15542 = pi10 ? n32 : n15541;
  assign n15543 = pi15 ? n15537 : n15424;
  assign n15544 = pi21 ? n14158 : ~n32;
  assign n15545 = pi20 ? n15544 : n32;
  assign n15546 = pi19 ? n32 : n15545;
  assign n15547 = pi18 ? n32 : n15546;
  assign n15548 = pi17 ? n32 : n15547;
  assign n15549 = pi16 ? n32 : n15548;
  assign n15550 = pi15 ? n15139 : n15549;
  assign n15551 = pi14 ? n15543 : n15550;
  assign n15552 = pi13 ? n15551 : n15150;
  assign n15553 = pi15 ? n15150 : n15139;
  assign n15554 = pi14 ? n15150 : n15553;
  assign n15555 = pi20 ? n141 : ~n141;
  assign n15556 = pi19 ? n32 : n15555;
  assign n15557 = pi18 ? n32 : n15556;
  assign n15558 = pi17 ? n32 : n15557;
  assign n15559 = pi16 ? n32 : n15558;
  assign n15560 = pi15 ? n15150 : n15559;
  assign n15561 = pi20 ? n141 : n220;
  assign n15562 = pi19 ? n32 : n15561;
  assign n15563 = pi18 ? n32 : n15562;
  assign n15564 = pi17 ? n32 : n15563;
  assign n15565 = pi16 ? n32 : n15564;
  assign n15566 = pi15 ? n15565 : n15559;
  assign n15567 = pi14 ? n15560 : n15566;
  assign n15568 = pi13 ? n15554 : n15567;
  assign n15569 = pi12 ? n15552 : n15568;
  assign n15570 = pi19 ? n32 : ~n507;
  assign n15571 = pi18 ? n32 : n15570;
  assign n15572 = pi17 ? n32 : n15571;
  assign n15573 = pi16 ? n32 : n15572;
  assign n15574 = pi19 ? n32 : ~n365;
  assign n15575 = pi18 ? n32 : n15574;
  assign n15576 = pi17 ? n32 : n15575;
  assign n15577 = pi16 ? n32 : n15576;
  assign n15578 = pi15 ? n15573 : n15577;
  assign n15579 = pi19 ? n32 : ~n1248;
  assign n15580 = pi18 ? n32 : n15579;
  assign n15581 = pi17 ? n32 : n15580;
  assign n15582 = pi16 ? n32 : n15581;
  assign n15583 = pi15 ? n15582 : n14985;
  assign n15584 = pi14 ? n15578 : n15583;
  assign n15585 = pi19 ? n32 : ~n519;
  assign n15586 = pi18 ? n32 : n15585;
  assign n15587 = pi17 ? n32 : n15586;
  assign n15588 = pi16 ? n32 : n15587;
  assign n15589 = pi15 ? n15588 : n14985;
  assign n15590 = pi19 ? n32 : ~n11972;
  assign n15591 = pi18 ? n32 : n15590;
  assign n15592 = pi17 ? n32 : n15591;
  assign n15593 = pi16 ? n32 : n15592;
  assign n15594 = pi19 ? n32 : ~n15460;
  assign n15595 = pi18 ? n32 : n15594;
  assign n15596 = pi17 ? n32 : n15595;
  assign n15597 = pi16 ? n32 : n15596;
  assign n15598 = pi15 ? n15593 : n15597;
  assign n15599 = pi14 ? n15589 : n15598;
  assign n15600 = pi13 ? n15584 : n15599;
  assign n15601 = pi19 ? n1574 : ~n1476;
  assign n15602 = pi18 ? n32 : n15601;
  assign n15603 = pi17 ? n32 : n15602;
  assign n15604 = pi16 ? n32 : n15603;
  assign n15605 = pi19 ? n1574 : ~n208;
  assign n15606 = pi18 ? n32 : n15605;
  assign n15607 = pi17 ? n32 : n15606;
  assign n15608 = pi16 ? n32 : n15607;
  assign n15609 = pi15 ? n15604 : n15608;
  assign n15610 = pi20 ? n1817 : ~n481;
  assign n15611 = pi19 ? n1574 : ~n15610;
  assign n15612 = pi18 ? n32 : n15611;
  assign n15613 = pi17 ? n32 : n15612;
  assign n15614 = pi16 ? n32 : n15613;
  assign n15615 = pi15 ? n14995 : n15614;
  assign n15616 = pi14 ? n15609 : n15615;
  assign n15617 = pi19 ? n1574 : ~n340;
  assign n15618 = pi18 ? n32 : n15617;
  assign n15619 = pi17 ? n32 : n15618;
  assign n15620 = pi16 ? n32 : n15619;
  assign n15621 = pi19 ? n1574 : ~n11531;
  assign n15622 = pi18 ? n32 : n15621;
  assign n15623 = pi17 ? n32 : n15622;
  assign n15624 = pi16 ? n32 : n15623;
  assign n15625 = pi15 ? n15620 : n15624;
  assign n15626 = pi14 ? n15625 : n15624;
  assign n15627 = pi13 ? n15616 : n15626;
  assign n15628 = pi12 ? n15600 : n15627;
  assign n15629 = pi11 ? n15569 : n15628;
  assign n15630 = pi19 ? n32 : ~n11546;
  assign n15631 = pi18 ? n32 : n15630;
  assign n15632 = pi17 ? n32 : n15631;
  assign n15633 = pi16 ? n32 : n15632;
  assign n15634 = pi19 ? n32 : ~n1077;
  assign n15635 = pi18 ? n32 : n15634;
  assign n15636 = pi17 ? n32 : n15635;
  assign n15637 = pi16 ? n32 : n15636;
  assign n15638 = pi15 ? n15633 : n15637;
  assign n15639 = pi20 ? n726 : n32;
  assign n15640 = pi19 ? n32 : n15639;
  assign n15641 = pi18 ? n32 : n15640;
  assign n15642 = pi17 ? n32 : n15641;
  assign n15643 = pi16 ? n32 : n15642;
  assign n15644 = pi15 ? n15637 : n15643;
  assign n15645 = pi14 ? n15638 : n15644;
  assign n15646 = pi20 ? n564 : n32;
  assign n15647 = pi19 ? n32 : n15646;
  assign n15648 = pi18 ? n32 : n15647;
  assign n15649 = pi17 ? n32 : n15648;
  assign n15650 = pi16 ? n32 : n15649;
  assign n15651 = pi20 ? n1010 : n32;
  assign n15652 = pi19 ? n32 : n15651;
  assign n15653 = pi18 ? n32 : n15652;
  assign n15654 = pi17 ? n32 : n15653;
  assign n15655 = pi16 ? n32 : n15654;
  assign n15656 = pi15 ? n15650 : n15655;
  assign n15657 = pi14 ? n15650 : n15656;
  assign n15658 = pi13 ? n15645 : n15657;
  assign n15659 = pi22 ? n13584 : n32;
  assign n15660 = pi21 ? n15659 : n32;
  assign n15661 = pi20 ? n15660 : n32;
  assign n15662 = pi19 ? n32 : n15661;
  assign n15663 = pi18 ? n32 : n15662;
  assign n15664 = pi17 ? n32 : n15663;
  assign n15665 = pi16 ? n32 : n15664;
  assign n15666 = pi15 ? n15665 : n15518;
  assign n15667 = pi14 ? n15665 : n15666;
  assign n15668 = pi13 ? n15667 : n32;
  assign n15669 = pi12 ? n15658 : n15668;
  assign n15670 = pi11 ? n15669 : n32;
  assign n15671 = pi10 ? n15629 : n15670;
  assign n15672 = pi09 ? n15542 : n15671;
  assign n15673 = pi08 ? n15526 : n15672;
  assign n15674 = pi20 ? n1475 : n32;
  assign n15675 = pi19 ? n32 : n15674;
  assign n15676 = pi18 ? n32 : n15675;
  assign n15677 = pi17 ? n32 : n15676;
  assign n15678 = pi16 ? n32 : n15677;
  assign n15679 = pi15 ? n32 : n15678;
  assign n15680 = pi14 ? n15679 : n15537;
  assign n15681 = pi13 ? n32 : n15680;
  assign n15682 = pi12 ? n32 : n15681;
  assign n15683 = pi11 ? n32 : n15682;
  assign n15684 = pi10 ? n32 : n15683;
  assign n15685 = pi20 ? n1940 : ~n321;
  assign n15686 = pi19 ? n32 : n15685;
  assign n15687 = pi18 ? n32 : n15686;
  assign n15688 = pi17 ? n32 : n15687;
  assign n15689 = pi16 ? n32 : n15688;
  assign n15690 = pi15 ? n15537 : n15689;
  assign n15691 = pi20 ? n12244 : n32;
  assign n15692 = pi19 ? n32 : n15691;
  assign n15693 = pi18 ? n32 : n15692;
  assign n15694 = pi17 ? n32 : n15693;
  assign n15695 = pi16 ? n32 : n15694;
  assign n15696 = pi20 ? n11086 : n32;
  assign n15697 = pi19 ? n32 : n15696;
  assign n15698 = pi18 ? n32 : n15697;
  assign n15699 = pi17 ? n32 : n15698;
  assign n15700 = pi16 ? n32 : n15699;
  assign n15701 = pi15 ? n15695 : n15700;
  assign n15702 = pi14 ? n15690 : n15701;
  assign n15703 = pi20 ? n243 : n32;
  assign n15704 = pi19 ? n32 : n15703;
  assign n15705 = pi18 ? n32 : n15704;
  assign n15706 = pi17 ? n32 : n15705;
  assign n15707 = pi16 ? n32 : n15706;
  assign n15708 = pi15 ? n15403 : n15707;
  assign n15709 = pi15 ? n15707 : n15139;
  assign n15710 = pi14 ? n15708 : n15709;
  assign n15711 = pi13 ? n15702 : n15710;
  assign n15712 = pi14 ? n15139 : n15550;
  assign n15713 = pi20 ? n141 : n9000;
  assign n15714 = pi19 ? n32 : n15713;
  assign n15715 = pi18 ? n32 : n15714;
  assign n15716 = pi17 ? n32 : n15715;
  assign n15717 = pi16 ? n32 : n15716;
  assign n15718 = pi20 ? n141 : n111;
  assign n15719 = pi19 ? n32 : n15718;
  assign n15720 = pi18 ? n32 : n15719;
  assign n15721 = pi17 ? n32 : n15720;
  assign n15722 = pi16 ? n32 : n15721;
  assign n15723 = pi15 ? n15717 : n15722;
  assign n15724 = pi14 ? n15150 : n15723;
  assign n15725 = pi13 ? n15712 : n15724;
  assign n15726 = pi12 ? n15711 : n15725;
  assign n15727 = pi20 ? n141 : n726;
  assign n15728 = pi19 ? n32 : n15727;
  assign n15729 = pi18 ? n32 : n15728;
  assign n15730 = pi17 ? n32 : n15729;
  assign n15731 = pi16 ? n32 : n15730;
  assign n15732 = pi21 ? n140 : n259;
  assign n15733 = pi20 ? n141 : ~n15732;
  assign n15734 = pi19 ? n32 : n15733;
  assign n15735 = pi18 ? n32 : n15734;
  assign n15736 = pi17 ? n32 : n15735;
  assign n15737 = pi16 ? n32 : n15736;
  assign n15738 = pi15 ? n15731 : n15737;
  assign n15739 = pi20 ? n141 : n1445;
  assign n15740 = pi19 ? n32 : n15739;
  assign n15741 = pi18 ? n32 : n15740;
  assign n15742 = pi17 ? n32 : n15741;
  assign n15743 = pi16 ? n32 : n15742;
  assign n15744 = pi20 ? n141 : n1817;
  assign n15745 = pi19 ? n32 : n15744;
  assign n15746 = pi18 ? n32 : n15745;
  assign n15747 = pi17 ? n32 : n15746;
  assign n15748 = pi16 ? n32 : n15747;
  assign n15749 = pi15 ? n15743 : n15748;
  assign n15750 = pi14 ? n15738 : n15749;
  assign n15751 = pi20 ? n339 : ~n518;
  assign n15752 = pi19 ? n32 : n15751;
  assign n15753 = pi18 ? n32 : n15752;
  assign n15754 = pi17 ? n32 : n15753;
  assign n15755 = pi16 ? n32 : n15754;
  assign n15756 = pi20 ? n339 : n6229;
  assign n15757 = pi19 ? n32 : n15756;
  assign n15758 = pi18 ? n32 : n15757;
  assign n15759 = pi17 ? n32 : n15758;
  assign n15760 = pi16 ? n32 : n15759;
  assign n15761 = pi15 ? n15755 : n15760;
  assign n15762 = pi20 ? n339 : ~n749;
  assign n15763 = pi19 ? n32 : n15762;
  assign n15764 = pi18 ? n32 : n15763;
  assign n15765 = pi17 ? n32 : n15764;
  assign n15766 = pi16 ? n32 : n15765;
  assign n15767 = pi15 ? n15766 : n15760;
  assign n15768 = pi14 ? n15761 : n15767;
  assign n15769 = pi13 ? n15750 : n15768;
  assign n15770 = pi20 ? n141 : ~n749;
  assign n15771 = pi19 ? n32 : n15770;
  assign n15772 = pi18 ? n32 : n15771;
  assign n15773 = pi17 ? n32 : n15772;
  assign n15774 = pi16 ? n32 : n15773;
  assign n15775 = pi20 ? n141 : ~n207;
  assign n15776 = pi19 ? n32 : n15775;
  assign n15777 = pi18 ? n32 : n15776;
  assign n15778 = pi17 ? n32 : n15777;
  assign n15779 = pi16 ? n32 : n15778;
  assign n15780 = pi15 ? n15774 : n15779;
  assign n15781 = pi21 ? n631 : ~n32;
  assign n15782 = pi20 ? n15781 : n32;
  assign n15783 = pi19 ? n32 : n15782;
  assign n15784 = pi18 ? n32 : n15783;
  assign n15785 = pi17 ? n32 : n15784;
  assign n15786 = pi16 ? n32 : n15785;
  assign n15787 = pi20 ? n141 : n481;
  assign n15788 = pi19 ? n32 : n15787;
  assign n15789 = pi18 ? n32 : n15788;
  assign n15790 = pi17 ? n32 : n15789;
  assign n15791 = pi16 ? n32 : n15790;
  assign n15792 = pi15 ? n15786 : n15791;
  assign n15793 = pi14 ? n15780 : n15792;
  assign n15794 = pi20 ? n15781 : ~n339;
  assign n15795 = pi19 ? n32 : n15794;
  assign n15796 = pi18 ? n32 : n15795;
  assign n15797 = pi17 ? n32 : n15796;
  assign n15798 = pi16 ? n32 : n15797;
  assign n15799 = pi21 ? n50 : ~n32;
  assign n15800 = pi20 ? n15799 : n32;
  assign n15801 = pi19 ? n32 : n15800;
  assign n15802 = pi18 ? n32 : n15801;
  assign n15803 = pi17 ? n32 : n15802;
  assign n15804 = pi16 ? n32 : n15803;
  assign n15805 = pi15 ? n15798 : n15804;
  assign n15806 = pi20 ? n1188 : n32;
  assign n15807 = pi19 ? n32 : n15806;
  assign n15808 = pi18 ? n32 : n15807;
  assign n15809 = pi17 ? n32 : n15808;
  assign n15810 = pi16 ? n32 : n15809;
  assign n15811 = pi15 ? n15810 : n15150;
  assign n15812 = pi14 ? n15805 : n15811;
  assign n15813 = pi13 ? n15793 : n15812;
  assign n15814 = pi12 ? n15769 : n15813;
  assign n15815 = pi11 ? n15726 : n15814;
  assign n15816 = pi22 ? n50 : n65;
  assign n15817 = pi21 ? n15816 : ~n206;
  assign n15818 = pi20 ? n15817 : n32;
  assign n15819 = pi19 ? n32 : n15818;
  assign n15820 = pi18 ? n32 : n15819;
  assign n15821 = pi17 ? n32 : n15820;
  assign n15822 = pi16 ? n32 : n15821;
  assign n15823 = pi15 ? n15810 : n15822;
  assign n15824 = pi21 ? n50 : ~n206;
  assign n15825 = pi20 ? n15824 : n32;
  assign n15826 = pi19 ? n32 : n15825;
  assign n15827 = pi18 ? n32 : n15826;
  assign n15828 = pi17 ? n32 : n15827;
  assign n15829 = pi16 ? n32 : n15828;
  assign n15830 = pi14 ? n15823 : n15829;
  assign n15831 = pi19 ? n32 : n1885;
  assign n15832 = pi18 ? n32 : n15831;
  assign n15833 = pi17 ? n32 : n15832;
  assign n15834 = pi16 ? n32 : n15833;
  assign n15835 = pi15 ? n15834 : n15650;
  assign n15836 = pi16 ? n32 : n2055;
  assign n15837 = pi15 ? n15834 : n15836;
  assign n15838 = pi14 ? n15835 : n15837;
  assign n15839 = pi13 ? n15830 : n15838;
  assign n15840 = pi12 ? n15839 : n32;
  assign n15841 = pi11 ? n15840 : n32;
  assign n15842 = pi10 ? n15815 : n15841;
  assign n15843 = pi09 ? n15684 : n15842;
  assign n15844 = pi19 ? n32 : n4342;
  assign n15845 = pi18 ? n32 : n15844;
  assign n15846 = pi17 ? n32 : n15845;
  assign n15847 = pi16 ? n32 : n15846;
  assign n15848 = pi15 ? n32 : n15847;
  assign n15849 = pi19 ? n32 : n4964;
  assign n15850 = pi18 ? n32 : n15849;
  assign n15851 = pi17 ? n32 : n15850;
  assign n15852 = pi16 ? n32 : n15851;
  assign n15853 = pi14 ? n15848 : n15852;
  assign n15854 = pi13 ? n32 : n15853;
  assign n15855 = pi12 ? n32 : n15854;
  assign n15856 = pi11 ? n32 : n15855;
  assign n15857 = pi10 ? n32 : n15856;
  assign n15858 = pi15 ? n15852 : n15689;
  assign n15859 = pi20 ? n1940 : n32;
  assign n15860 = pi19 ? n32 : n15859;
  assign n15861 = pi18 ? n32 : n15860;
  assign n15862 = pi17 ? n32 : n15861;
  assign n15863 = pi16 ? n32 : n15862;
  assign n15864 = pi19 ? n32 : n7435;
  assign n15865 = pi18 ? n32 : n15864;
  assign n15866 = pi17 ? n32 : n15865;
  assign n15867 = pi16 ? n32 : n15866;
  assign n15868 = pi15 ? n15863 : n15867;
  assign n15869 = pi14 ? n15858 : n15868;
  assign n15870 = pi15 ? n15403 : n15863;
  assign n15871 = pi14 ? n15870 : n15863;
  assign n15872 = pi13 ? n15869 : n15871;
  assign n15873 = pi20 ? n243 : n9000;
  assign n15874 = pi19 ? n32 : n15873;
  assign n15875 = pi18 ? n32 : n15874;
  assign n15876 = pi17 ? n32 : n15875;
  assign n15877 = pi16 ? n32 : n15876;
  assign n15878 = pi20 ? n339 : n111;
  assign n15879 = pi19 ? n32 : n15878;
  assign n15880 = pi18 ? n32 : n15879;
  assign n15881 = pi17 ? n32 : n15880;
  assign n15882 = pi16 ? n32 : n15881;
  assign n15883 = pi15 ? n15877 : n15882;
  assign n15884 = pi14 ? n15708 : n15883;
  assign n15885 = pi13 ? n15863 : n15884;
  assign n15886 = pi12 ? n15872 : n15885;
  assign n15887 = pi20 ? n339 : n623;
  assign n15888 = pi19 ? n32 : n15887;
  assign n15889 = pi18 ? n32 : n15888;
  assign n15890 = pi17 ? n32 : n15889;
  assign n15891 = pi16 ? n32 : n15890;
  assign n15892 = pi20 ? n339 : ~n15732;
  assign n15893 = pi19 ? n32 : n15892;
  assign n15894 = pi18 ? n32 : n15893;
  assign n15895 = pi17 ? n32 : n15894;
  assign n15896 = pi16 ? n32 : n15895;
  assign n15897 = pi15 ? n15891 : n15896;
  assign n15898 = pi20 ? n339 : n1445;
  assign n15899 = pi19 ? n32 : n15898;
  assign n15900 = pi18 ? n32 : n15899;
  assign n15901 = pi17 ? n32 : n15900;
  assign n15902 = pi16 ? n32 : n15901;
  assign n15903 = pi20 ? n339 : n1817;
  assign n15904 = pi19 ? n32 : n15903;
  assign n15905 = pi18 ? n32 : n15904;
  assign n15906 = pi17 ? n32 : n15905;
  assign n15907 = pi16 ? n32 : n15906;
  assign n15908 = pi15 ? n15902 : n15907;
  assign n15909 = pi14 ? n15897 : n15908;
  assign n15910 = pi15 ? n15766 : n15139;
  assign n15911 = pi14 ? n15767 : n15910;
  assign n15912 = pi13 ? n15909 : n15911;
  assign n15913 = pi19 ? n32 : n6120;
  assign n15914 = pi18 ? n32 : n15913;
  assign n15915 = pi17 ? n32 : n15914;
  assign n15916 = pi16 ? n32 : n15915;
  assign n15917 = pi20 ? n10446 : ~n207;
  assign n15918 = pi19 ? n32 : n15917;
  assign n15919 = pi18 ? n32 : n15918;
  assign n15920 = pi17 ? n32 : n15919;
  assign n15921 = pi16 ? n32 : n15920;
  assign n15922 = pi15 ? n15916 : n15921;
  assign n15923 = pi20 ? n2358 : n32;
  assign n15924 = pi19 ? n32 : n15923;
  assign n15925 = pi18 ? n32 : n15924;
  assign n15926 = pi17 ? n32 : n15925;
  assign n15927 = pi16 ? n32 : n15926;
  assign n15928 = pi15 ? n15927 : n15139;
  assign n15929 = pi14 ? n15922 : n15928;
  assign n15930 = pi21 ? n35 : ~n32;
  assign n15931 = pi20 ? n15930 : n32;
  assign n15932 = pi19 ? n32 : n15931;
  assign n15933 = pi18 ? n32 : n15932;
  assign n15934 = pi17 ? n32 : n15933;
  assign n15935 = pi16 ? n32 : n15934;
  assign n15936 = pi15 ? n15935 : n15707;
  assign n15937 = pi20 ? n14368 : n32;
  assign n15938 = pi19 ? n32 : n15937;
  assign n15939 = pi18 ? n32 : n15938;
  assign n15940 = pi17 ? n32 : n15939;
  assign n15941 = pi16 ? n32 : n15940;
  assign n15942 = pi21 ? n242 : ~n206;
  assign n15943 = pi20 ? n15942 : n32;
  assign n15944 = pi19 ? n32 : n15943;
  assign n15945 = pi18 ? n32 : n15944;
  assign n15946 = pi17 ? n32 : n15945;
  assign n15947 = pi16 ? n32 : n15946;
  assign n15948 = pi15 ? n15941 : n15947;
  assign n15949 = pi14 ? n15936 : n15948;
  assign n15950 = pi13 ? n15929 : n15949;
  assign n15951 = pi12 ? n15912 : n15950;
  assign n15952 = pi11 ? n15886 : n15951;
  assign n15953 = pi22 ? n34 : ~n65;
  assign n15954 = pi21 ? n15953 : ~n206;
  assign n15955 = pi20 ? n15954 : n32;
  assign n15956 = pi19 ? n32 : n15955;
  assign n15957 = pi18 ? n32 : n15956;
  assign n15958 = pi17 ? n32 : n15957;
  assign n15959 = pi16 ? n32 : n15958;
  assign n15960 = pi15 ? n15947 : n15959;
  assign n15961 = pi21 ? n242 : n32;
  assign n15962 = pi20 ? n15961 : n32;
  assign n15963 = pi19 ? n32 : n15962;
  assign n15964 = pi18 ? n32 : n15963;
  assign n15965 = pi17 ? n32 : n15964;
  assign n15966 = pi16 ? n32 : n15965;
  assign n15967 = pi14 ? n15960 : n15966;
  assign n15968 = pi15 ? n15966 : n15836;
  assign n15969 = pi14 ? n15966 : n15968;
  assign n15970 = pi13 ? n15967 : n15969;
  assign n15971 = pi12 ? n15970 : n32;
  assign n15972 = pi11 ? n15971 : n32;
  assign n15973 = pi10 ? n15952 : n15972;
  assign n15974 = pi09 ? n15857 : n15973;
  assign n15975 = pi08 ? n15843 : n15974;
  assign n15976 = pi07 ? n15673 : n15975;
  assign n15977 = pi20 ? n1839 : ~n321;
  assign n15978 = pi19 ? n32 : n15977;
  assign n15979 = pi18 ? n32 : n15978;
  assign n15980 = pi17 ? n32 : n15979;
  assign n15981 = pi16 ? n32 : n15980;
  assign n15982 = pi15 ? n32 : n15981;
  assign n15983 = pi20 ? n518 : ~n321;
  assign n15984 = pi19 ? n32 : n15983;
  assign n15985 = pi18 ? n32 : n15984;
  assign n15986 = pi17 ? n32 : n15985;
  assign n15987 = pi16 ? n32 : n15986;
  assign n15988 = pi14 ? n15982 : n15987;
  assign n15989 = pi13 ? n32 : n15988;
  assign n15990 = pi12 ? n32 : n15989;
  assign n15991 = pi11 ? n32 : n15990;
  assign n15992 = pi10 ? n32 : n15991;
  assign n15993 = pi20 ? n1475 : ~n321;
  assign n15994 = pi19 ? n32 : n15993;
  assign n15995 = pi18 ? n32 : n15994;
  assign n15996 = pi17 ? n32 : n15995;
  assign n15997 = pi16 ? n32 : n15996;
  assign n15998 = pi15 ? n15987 : n15997;
  assign n15999 = pi14 ? n15998 : n15531;
  assign n16000 = pi14 ? n15531 : n15863;
  assign n16001 = pi13 ? n15999 : n16000;
  assign n16002 = pi20 ? n207 : n220;
  assign n16003 = pi19 ? n32 : n16002;
  assign n16004 = pi18 ? n32 : n16003;
  assign n16005 = pi17 ? n32 : n16004;
  assign n16006 = pi16 ? n32 : n16005;
  assign n16007 = pi15 ? n16006 : n15403;
  assign n16008 = pi21 ? n206 : ~n51;
  assign n16009 = pi20 ? n207 : ~n16008;
  assign n16010 = pi19 ? n32 : n16009;
  assign n16011 = pi18 ? n32 : n16010;
  assign n16012 = pi17 ? n32 : n16011;
  assign n16013 = pi16 ? n32 : n16012;
  assign n16014 = pi20 ? n11048 : n111;
  assign n16015 = pi19 ? n32 : n16014;
  assign n16016 = pi18 ? n32 : n16015;
  assign n16017 = pi17 ? n32 : n16016;
  assign n16018 = pi16 ? n32 : n16017;
  assign n16019 = pi15 ? n16013 : n16018;
  assign n16020 = pi14 ? n16007 : n16019;
  assign n16021 = pi13 ? n15863 : n16020;
  assign n16022 = pi12 ? n16001 : n16021;
  assign n16023 = pi20 ? n1940 : n266;
  assign n16024 = pi19 ? n32 : n16023;
  assign n16025 = pi18 ? n32 : n16024;
  assign n16026 = pi17 ? n32 : n16025;
  assign n16027 = pi16 ? n32 : n16026;
  assign n16028 = pi20 ? n1940 : n1817;
  assign n16029 = pi19 ? n32 : n16028;
  assign n16030 = pi18 ? n32 : n16029;
  assign n16031 = pi17 ? n32 : n16030;
  assign n16032 = pi16 ? n32 : n16031;
  assign n16033 = pi15 ? n16027 : n16032;
  assign n16034 = pi20 ? n207 : n1010;
  assign n16035 = pi19 ? n32 : n16034;
  assign n16036 = pi18 ? n32 : n16035;
  assign n16037 = pi17 ? n32 : n16036;
  assign n16038 = pi16 ? n32 : n16037;
  assign n16039 = pi15 ? n16038 : n16032;
  assign n16040 = pi14 ? n16033 : n16039;
  assign n16041 = pi19 ? n32 : n13069;
  assign n16042 = pi18 ? n32 : n16041;
  assign n16043 = pi17 ? n32 : n16042;
  assign n16044 = pi16 ? n32 : n16043;
  assign n16045 = pi20 ? n1940 : ~n11048;
  assign n16046 = pi19 ? n32 : n16045;
  assign n16047 = pi18 ? n32 : n16046;
  assign n16048 = pi17 ? n32 : n16047;
  assign n16049 = pi16 ? n32 : n16048;
  assign n16050 = pi15 ? n16044 : n16049;
  assign n16051 = pi20 ? n207 : n274;
  assign n16052 = pi19 ? n32 : n16051;
  assign n16053 = pi18 ? n32 : n16052;
  assign n16054 = pi17 ? n32 : n16053;
  assign n16055 = pi16 ? n32 : n16054;
  assign n16056 = pi15 ? n16055 : n16044;
  assign n16057 = pi14 ? n16050 : n16056;
  assign n16058 = pi13 ? n16040 : n16057;
  assign n16059 = pi22 ? n34 : ~n13584;
  assign n16060 = pi21 ? n16059 : ~n32;
  assign n16061 = pi20 ? n16060 : ~n207;
  assign n16062 = pi19 ? n32 : n16061;
  assign n16063 = pi18 ? n32 : n16062;
  assign n16064 = pi17 ? n32 : n16063;
  assign n16065 = pi16 ? n32 : n16064;
  assign n16066 = pi20 ? n243 : ~n339;
  assign n16067 = pi19 ? n32 : n16066;
  assign n16068 = pi18 ? n32 : n16067;
  assign n16069 = pi17 ? n32 : n16068;
  assign n16070 = pi16 ? n32 : n16069;
  assign n16071 = pi15 ? n16065 : n16070;
  assign n16072 = pi14 ? n15707 : n16071;
  assign n16073 = pi21 ? n15953 : ~n32;
  assign n16074 = pi20 ? n16073 : n32;
  assign n16075 = pi19 ? n32 : n16074;
  assign n16076 = pi18 ? n32 : n16075;
  assign n16077 = pi17 ? n32 : n16076;
  assign n16078 = pi16 ? n32 : n16077;
  assign n16079 = pi21 ? n242 : n206;
  assign n16080 = pi20 ? n16079 : n32;
  assign n16081 = pi19 ? n32 : n16080;
  assign n16082 = pi18 ? n32 : n16081;
  assign n16083 = pi17 ? n32 : n16082;
  assign n16084 = pi16 ? n32 : n16083;
  assign n16085 = pi15 ? n16078 : n16084;
  assign n16086 = pi15 ? n15707 : n15947;
  assign n16087 = pi14 ? n16085 : n16086;
  assign n16088 = pi13 ? n16072 : n16087;
  assign n16089 = pi12 ? n16058 : n16088;
  assign n16090 = pi11 ? n16022 : n16089;
  assign n16091 = pi22 ? n34 : ~n84;
  assign n16092 = pi21 ? n16091 : ~n206;
  assign n16093 = pi20 ? n16092 : n32;
  assign n16094 = pi19 ? n32 : n16093;
  assign n16095 = pi18 ? n32 : n16094;
  assign n16096 = pi17 ? n32 : n16095;
  assign n16097 = pi16 ? n32 : n16096;
  assign n16098 = pi19 ? n32 : n3692;
  assign n16099 = pi18 ? n32 : n16098;
  assign n16100 = pi17 ? n32 : n16099;
  assign n16101 = pi16 ? n32 : n16100;
  assign n16102 = pi15 ? n16097 : n16101;
  assign n16103 = pi18 ? n32 : n5657;
  assign n16104 = pi17 ? n32 : n16103;
  assign n16105 = pi16 ? n32 : n16104;
  assign n16106 = pi15 ? n15700 : n16105;
  assign n16107 = pi14 ? n16102 : n16106;
  assign n16108 = pi16 ? n32 : n1528;
  assign n16109 = pi15 ? n16105 : n16108;
  assign n16110 = pi15 ? n16108 : n32;
  assign n16111 = pi14 ? n16109 : n16110;
  assign n16112 = pi13 ? n16107 : n16111;
  assign n16113 = pi12 ? n16112 : n32;
  assign n16114 = pi11 ? n16113 : n32;
  assign n16115 = pi10 ? n16090 : n16114;
  assign n16116 = pi09 ? n15992 : n16115;
  assign n16117 = pi14 ? n15982 : n15981;
  assign n16118 = pi13 ? n32 : n16117;
  assign n16119 = pi12 ? n32 : n16118;
  assign n16120 = pi11 ? n32 : n16119;
  assign n16121 = pi10 ? n32 : n16120;
  assign n16122 = pi15 ? n15981 : n15852;
  assign n16123 = pi14 ? n16122 : n15678;
  assign n16124 = pi13 ? n16123 : n15678;
  assign n16125 = pi15 ? n15678 : n15531;
  assign n16126 = pi14 ? n15678 : n16125;
  assign n16127 = pi20 ? n749 : n220;
  assign n16128 = pi19 ? n32 : n16127;
  assign n16129 = pi18 ? n32 : n16128;
  assign n16130 = pi17 ? n32 : n16129;
  assign n16131 = pi16 ? n32 : n16130;
  assign n16132 = pi15 ? n16131 : n15531;
  assign n16133 = pi20 ? n749 : n8760;
  assign n16134 = pi19 ? n32 : n16133;
  assign n16135 = pi18 ? n32 : n16134;
  assign n16136 = pi17 ? n32 : n16135;
  assign n16137 = pi16 ? n32 : n16136;
  assign n16138 = pi20 ? n1940 : n111;
  assign n16139 = pi19 ? n32 : n16138;
  assign n16140 = pi18 ? n32 : n16139;
  assign n16141 = pi17 ? n32 : n16140;
  assign n16142 = pi16 ? n32 : n16141;
  assign n16143 = pi15 ? n16137 : n16142;
  assign n16144 = pi14 ? n16132 : n16143;
  assign n16145 = pi13 ? n16126 : n16144;
  assign n16146 = pi12 ? n16124 : n16145;
  assign n16147 = pi20 ? n1940 : n1010;
  assign n16148 = pi19 ? n32 : n16147;
  assign n16149 = pi18 ? n32 : n16148;
  assign n16150 = pi17 ? n32 : n16149;
  assign n16151 = pi16 ? n32 : n16150;
  assign n16152 = pi15 ? n16151 : n15863;
  assign n16153 = pi14 ? n16033 : n16152;
  assign n16154 = pi20 ? n1940 : ~n207;
  assign n16155 = pi19 ? n32 : n16154;
  assign n16156 = pi18 ? n32 : n16155;
  assign n16157 = pi17 ? n32 : n16156;
  assign n16158 = pi16 ? n32 : n16157;
  assign n16159 = pi15 ? n16158 : n16049;
  assign n16160 = pi20 ? n1940 : n274;
  assign n16161 = pi19 ? n32 : n16160;
  assign n16162 = pi18 ? n32 : n16161;
  assign n16163 = pi17 ? n32 : n16162;
  assign n16164 = pi16 ? n32 : n16163;
  assign n16165 = pi15 ? n16164 : n16158;
  assign n16166 = pi14 ? n16159 : n16165;
  assign n16167 = pi13 ? n16153 : n16166;
  assign n16168 = pi21 ? n2076 : ~n32;
  assign n16169 = pi20 ? n16168 : n32;
  assign n16170 = pi19 ? n32 : n16169;
  assign n16171 = pi18 ? n32 : n16170;
  assign n16172 = pi17 ? n32 : n16171;
  assign n16173 = pi16 ? n32 : n16172;
  assign n16174 = pi15 ? n15531 : n16173;
  assign n16175 = pi22 ? n32 : ~n13584;
  assign n16176 = pi21 ? n16175 : ~n32;
  assign n16177 = pi20 ? n16176 : ~n207;
  assign n16178 = pi19 ? n32 : n16177;
  assign n16179 = pi18 ? n32 : n16178;
  assign n16180 = pi17 ? n32 : n16179;
  assign n16181 = pi16 ? n32 : n16180;
  assign n16182 = pi20 ? n12244 : ~n339;
  assign n16183 = pi19 ? n32 : n16182;
  assign n16184 = pi18 ? n32 : n16183;
  assign n16185 = pi17 ? n32 : n16184;
  assign n16186 = pi16 ? n32 : n16185;
  assign n16187 = pi15 ? n16181 : n16186;
  assign n16188 = pi14 ? n16174 : n16187;
  assign n16189 = pi20 ? n785 : n32;
  assign n16190 = pi19 ? n32 : n16189;
  assign n16191 = pi18 ? n32 : n16190;
  assign n16192 = pi17 ? n32 : n16191;
  assign n16193 = pi16 ? n32 : n16192;
  assign n16194 = pi15 ? n15403 : n16193;
  assign n16195 = pi21 ? n11567 : ~n32;
  assign n16196 = pi20 ? n16195 : n32;
  assign n16197 = pi19 ? n32 : n16196;
  assign n16198 = pi18 ? n32 : n16197;
  assign n16199 = pi17 ? n32 : n16198;
  assign n16200 = pi16 ? n32 : n16199;
  assign n16201 = pi19 ? n32 : n10863;
  assign n16202 = pi18 ? n32 : n16201;
  assign n16203 = pi17 ? n32 : n16202;
  assign n16204 = pi16 ? n32 : n16203;
  assign n16205 = pi15 ? n16200 : n16204;
  assign n16206 = pi14 ? n16194 : n16205;
  assign n16207 = pi13 ? n16188 : n16206;
  assign n16208 = pi12 ? n16167 : n16207;
  assign n16209 = pi11 ? n16146 : n16208;
  assign n16210 = pi21 ? n1939 : ~n140;
  assign n16211 = pi20 ? n16210 : n32;
  assign n16212 = pi19 ? n32 : n16211;
  assign n16213 = pi18 ? n32 : n16212;
  assign n16214 = pi17 ? n32 : n16213;
  assign n16215 = pi16 ? n32 : n16214;
  assign n16216 = pi15 ? n16215 : n15700;
  assign n16217 = pi14 ? n16204 : n16216;
  assign n16218 = pi15 ? n15700 : n32;
  assign n16219 = pi14 ? n16218 : n32;
  assign n16220 = pi13 ? n16217 : n16219;
  assign n16221 = pi12 ? n16220 : n32;
  assign n16222 = pi11 ? n16221 : n32;
  assign n16223 = pi10 ? n16209 : n16222;
  assign n16224 = pi09 ? n16121 : n16223;
  assign n16225 = pi08 ? n16116 : n16224;
  assign n16226 = pi15 ? n32 : n15987;
  assign n16227 = pi14 ? n16226 : n15987;
  assign n16228 = pi13 ? n32 : n16227;
  assign n16229 = pi12 ? n32 : n16228;
  assign n16230 = pi11 ? n32 : n16229;
  assign n16231 = pi10 ? n32 : n16230;
  assign n16232 = pi15 ? n15847 : n15678;
  assign n16233 = pi14 ? n16122 : n16232;
  assign n16234 = pi19 ? n32 : n5004;
  assign n16235 = pi18 ? n32 : n16234;
  assign n16236 = pi17 ? n32 : n16235;
  assign n16237 = pi16 ? n32 : n16236;
  assign n16238 = pi15 ? n15847 : n16237;
  assign n16239 = pi14 ? n15678 : n16238;
  assign n16240 = pi13 ? n16233 : n16239;
  assign n16241 = pi14 ? n15847 : n16232;
  assign n16242 = pi20 ? n1475 : ~n2140;
  assign n16243 = pi19 ? n32 : n16242;
  assign n16244 = pi18 ? n32 : n16243;
  assign n16245 = pi17 ? n32 : n16244;
  assign n16246 = pi16 ? n32 : n16245;
  assign n16247 = pi20 ? n1475 : ~n141;
  assign n16248 = pi19 ? n32 : n16247;
  assign n16249 = pi18 ? n32 : n16248;
  assign n16250 = pi17 ? n32 : n16249;
  assign n16251 = pi16 ? n32 : n16250;
  assign n16252 = pi15 ? n16246 : n16251;
  assign n16253 = pi21 ? n140 : ~n51;
  assign n16254 = pi20 ? n749 : ~n16253;
  assign n16255 = pi19 ? n32 : n16254;
  assign n16256 = pi18 ? n32 : n16255;
  assign n16257 = pi17 ? n32 : n16256;
  assign n16258 = pi16 ? n32 : n16257;
  assign n16259 = pi15 ? n15678 : n16258;
  assign n16260 = pi14 ? n16252 : n16259;
  assign n16261 = pi13 ? n16241 : n16260;
  assign n16262 = pi12 ? n16240 : n16261;
  assign n16263 = pi20 ? n1475 : n564;
  assign n16264 = pi19 ? n32 : n16263;
  assign n16265 = pi18 ? n32 : n16264;
  assign n16266 = pi17 ? n32 : n16265;
  assign n16267 = pi16 ? n32 : n16266;
  assign n16268 = pi15 ? n16267 : n15678;
  assign n16269 = pi14 ? n16268 : n15678;
  assign n16270 = pi20 ? n749 : ~n749;
  assign n16271 = pi19 ? n32 : n16270;
  assign n16272 = pi18 ? n32 : n16271;
  assign n16273 = pi17 ? n32 : n16272;
  assign n16274 = pi16 ? n32 : n16273;
  assign n16275 = pi19 ? n32 : n13362;
  assign n16276 = pi18 ? n32 : n16275;
  assign n16277 = pi17 ? n32 : n16276;
  assign n16278 = pi16 ? n32 : n16277;
  assign n16279 = pi15 ? n15531 : n16278;
  assign n16280 = pi14 ? n16274 : n16279;
  assign n16281 = pi13 ? n16269 : n16280;
  assign n16282 = pi20 ? n749 : ~n207;
  assign n16283 = pi19 ? n32 : n16282;
  assign n16284 = pi18 ? n32 : n16283;
  assign n16285 = pi17 ? n32 : n16284;
  assign n16286 = pi16 ? n32 : n16285;
  assign n16287 = pi15 ? n16286 : n15531;
  assign n16288 = pi14 ? n15531 : n16287;
  assign n16289 = pi20 ? n9897 : n32;
  assign n16290 = pi19 ? n32 : n16289;
  assign n16291 = pi18 ? n32 : n16290;
  assign n16292 = pi17 ? n32 : n16291;
  assign n16293 = pi16 ? n32 : n16292;
  assign n16294 = pi20 ? n7839 : n32;
  assign n16295 = pi19 ? n32 : n16294;
  assign n16296 = pi18 ? n32 : n16295;
  assign n16297 = pi17 ? n32 : n16296;
  assign n16298 = pi16 ? n32 : n16297;
  assign n16299 = pi15 ? n16293 : n16298;
  assign n16300 = pi14 ? n15531 : n16299;
  assign n16301 = pi13 ? n16288 : n16300;
  assign n16302 = pi12 ? n16281 : n16301;
  assign n16303 = pi11 ? n16262 : n16302;
  assign n16304 = pi20 ? n9863 : n32;
  assign n16305 = pi19 ? n32 : n16304;
  assign n16306 = pi18 ? n32 : n16305;
  assign n16307 = pi17 ? n32 : n16306;
  assign n16308 = pi16 ? n32 : n16307;
  assign n16309 = pi21 ? n405 : ~n140;
  assign n16310 = pi20 ? n16309 : n32;
  assign n16311 = pi19 ? n32 : n16310;
  assign n16312 = pi18 ? n32 : n16311;
  assign n16313 = pi17 ? n32 : n16312;
  assign n16314 = pi16 ? n32 : n16313;
  assign n16315 = pi15 ? n16308 : n16314;
  assign n16316 = pi19 ? n32 : n1844;
  assign n16317 = pi18 ? n32 : n16316;
  assign n16318 = pi17 ? n32 : n16317;
  assign n16319 = pi16 ? n32 : n16318;
  assign n16320 = pi14 ? n16315 : n16319;
  assign n16321 = pi15 ? n16319 : n32;
  assign n16322 = pi14 ? n16321 : n32;
  assign n16323 = pi13 ? n16320 : n16322;
  assign n16324 = pi12 ? n16323 : n32;
  assign n16325 = pi11 ? n16324 : n32;
  assign n16326 = pi10 ? n16303 : n16325;
  assign n16327 = pi09 ? n16231 : n16326;
  assign n16328 = pi15 ? n15987 : n15981;
  assign n16329 = pi20 ? n1839 : n32;
  assign n16330 = pi19 ? n32 : n16329;
  assign n16331 = pi18 ? n32 : n16330;
  assign n16332 = pi17 ? n32 : n16331;
  assign n16333 = pi16 ? n32 : n16332;
  assign n16334 = pi15 ? n16333 : n15847;
  assign n16335 = pi14 ? n16328 : n16334;
  assign n16336 = pi14 ? n15847 : n16238;
  assign n16337 = pi13 ? n16335 : n16336;
  assign n16338 = pi20 ? n1475 : ~n16253;
  assign n16339 = pi19 ? n32 : n16338;
  assign n16340 = pi18 ? n32 : n16339;
  assign n16341 = pi17 ? n32 : n16340;
  assign n16342 = pi16 ? n32 : n16341;
  assign n16343 = pi15 ? n15678 : n16342;
  assign n16344 = pi14 ? n16252 : n16343;
  assign n16345 = pi13 ? n15847 : n16344;
  assign n16346 = pi12 ? n16337 : n16345;
  assign n16347 = pi15 ? n16267 : n15847;
  assign n16348 = pi14 ? n16347 : n15847;
  assign n16349 = pi19 ? n32 : n5163;
  assign n16350 = pi18 ? n32 : n16349;
  assign n16351 = pi17 ? n32 : n16350;
  assign n16352 = pi16 ? n32 : n16351;
  assign n16353 = pi15 ? n15678 : n16352;
  assign n16354 = pi14 ? n16278 : n16353;
  assign n16355 = pi13 ? n16348 : n16354;
  assign n16356 = pi15 ? n16286 : n15847;
  assign n16357 = pi14 ? n15678 : n16356;
  assign n16358 = pi21 ? n100 : ~n1392;
  assign n16359 = pi20 ? n16358 : n32;
  assign n16360 = pi19 ? n32 : n16359;
  assign n16361 = pi18 ? n32 : n16360;
  assign n16362 = pi17 ? n32 : n16361;
  assign n16363 = pi16 ? n32 : n16362;
  assign n16364 = pi15 ? n16363 : n16293;
  assign n16365 = pi14 ? n16232 : n16364;
  assign n16366 = pi13 ? n16357 : n16365;
  assign n16367 = pi12 ? n16355 : n16366;
  assign n16368 = pi11 ? n16346 : n16367;
  assign n16369 = pi21 ? n100 : ~n259;
  assign n16370 = pi20 ? n16369 : n32;
  assign n16371 = pi19 ? n32 : n16370;
  assign n16372 = pi18 ? n32 : n16371;
  assign n16373 = pi17 ? n32 : n16372;
  assign n16374 = pi16 ? n32 : n16373;
  assign n16375 = pi15 ? n16374 : n32;
  assign n16376 = pi17 ? n32 : n3243;
  assign n16377 = pi16 ? n32 : n16376;
  assign n16378 = pi15 ? n16377 : n32;
  assign n16379 = pi14 ? n16375 : n16378;
  assign n16380 = pi13 ? n16379 : n32;
  assign n16381 = pi12 ? n16380 : n32;
  assign n16382 = pi11 ? n16381 : n32;
  assign n16383 = pi10 ? n16368 : n16382;
  assign n16384 = pi09 ? n16231 : n16383;
  assign n16385 = pi08 ? n16327 : n16384;
  assign n16386 = pi07 ? n16225 : n16385;
  assign n16387 = pi06 ? n15976 : n16386;
  assign n16388 = pi05 ? n15399 : n16387;
  assign n16389 = pi19 ? n32 : n4670;
  assign n16390 = pi18 ? n32 : n16389;
  assign n16391 = pi17 ? n32 : n16390;
  assign n16392 = pi16 ? n32 : n16391;
  assign n16393 = pi15 ? n32 : n16392;
  assign n16394 = pi19 ? n32 : n6988;
  assign n16395 = pi18 ? n32 : n16394;
  assign n16396 = pi17 ? n32 : n16395;
  assign n16397 = pi16 ? n32 : n16396;
  assign n16398 = pi20 ? n1319 : ~n321;
  assign n16399 = pi19 ? n32 : n16398;
  assign n16400 = pi18 ? n32 : n16399;
  assign n16401 = pi17 ? n32 : n16400;
  assign n16402 = pi16 ? n32 : n16401;
  assign n16403 = pi15 ? n16397 : n16402;
  assign n16404 = pi14 ? n16393 : n16403;
  assign n16405 = pi13 ? n32 : n16404;
  assign n16406 = pi12 ? n32 : n16405;
  assign n16407 = pi11 ? n32 : n16406;
  assign n16408 = pi10 ? n32 : n16407;
  assign n16409 = pi20 ? n1839 : ~n207;
  assign n16410 = pi19 ? n32 : n16409;
  assign n16411 = pi18 ? n32 : n16410;
  assign n16412 = pi17 ? n32 : n16411;
  assign n16413 = pi16 ? n32 : n16412;
  assign n16414 = pi15 ? n16413 : n16333;
  assign n16415 = pi14 ? n15981 : n16414;
  assign n16416 = pi13 ? n15981 : n16415;
  assign n16417 = pi20 ? n321 : n8760;
  assign n16418 = pi19 ? n32 : n16417;
  assign n16419 = pi18 ? n32 : n16418;
  assign n16420 = pi17 ? n32 : n16419;
  assign n16421 = pi16 ? n32 : n16420;
  assign n16422 = pi15 ? n16421 : n15847;
  assign n16423 = pi19 ? n32 : n6173;
  assign n16424 = pi18 ? n32 : n16423;
  assign n16425 = pi17 ? n32 : n16424;
  assign n16426 = pi16 ? n32 : n16425;
  assign n16427 = pi15 ? n15847 : n16426;
  assign n16428 = pi14 ? n16422 : n16427;
  assign n16429 = pi13 ? n15981 : n16428;
  assign n16430 = pi12 ? n16416 : n16429;
  assign n16431 = pi20 ? n321 : n266;
  assign n16432 = pi19 ? n32 : n16431;
  assign n16433 = pi18 ? n32 : n16432;
  assign n16434 = pi17 ? n32 : n16433;
  assign n16435 = pi16 ? n32 : n16434;
  assign n16436 = pi15 ? n16237 : n16435;
  assign n16437 = pi20 ? n321 : ~n14844;
  assign n16438 = pi19 ? n32 : n16437;
  assign n16439 = pi18 ? n32 : n16438;
  assign n16440 = pi17 ? n32 : n16439;
  assign n16441 = pi16 ? n32 : n16440;
  assign n16442 = pi14 ? n16436 : n16441;
  assign n16443 = pi15 ? n16352 : n16237;
  assign n16444 = pi15 ? n16237 : n16352;
  assign n16445 = pi14 ? n16443 : n16444;
  assign n16446 = pi13 ? n16442 : n16445;
  assign n16447 = pi15 ? n16237 : n16413;
  assign n16448 = pi14 ? n16447 : n16414;
  assign n16449 = pi19 ? n32 : n247;
  assign n16450 = pi18 ? n32 : n16449;
  assign n16451 = pi17 ? n32 : n16450;
  assign n16452 = pi16 ? n32 : n16451;
  assign n16453 = pi14 ? n16334 : n16452;
  assign n16454 = pi13 ? n16448 : n16453;
  assign n16455 = pi12 ? n16446 : n16454;
  assign n16456 = pi11 ? n16430 : n16455;
  assign n16457 = pi15 ? n16452 : n16377;
  assign n16458 = pi14 ? n16457 : n32;
  assign n16459 = pi13 ? n16458 : n32;
  assign n16460 = pi12 ? n16459 : n32;
  assign n16461 = pi11 ? n16460 : n32;
  assign n16462 = pi10 ? n16456 : n16461;
  assign n16463 = pi09 ? n16408 : n16462;
  assign n16464 = pi19 ? n32 : n13382;
  assign n16465 = pi18 ? n32 : n16464;
  assign n16466 = pi17 ? n32 : n16465;
  assign n16467 = pi16 ? n32 : n16466;
  assign n16468 = pi15 ? n32 : n16467;
  assign n16469 = pi14 ? n16468 : n16402;
  assign n16470 = pi13 ? n32 : n16469;
  assign n16471 = pi12 ? n32 : n16470;
  assign n16472 = pi11 ? n32 : n16471;
  assign n16473 = pi10 ? n32 : n16472;
  assign n16474 = pi14 ? n15987 : n16328;
  assign n16475 = pi13 ? n16474 : n16415;
  assign n16476 = pi20 ? n1839 : ~n16008;
  assign n16477 = pi19 ? n32 : n16476;
  assign n16478 = pi18 ? n32 : n16477;
  assign n16479 = pi17 ? n32 : n16478;
  assign n16480 = pi16 ? n32 : n16479;
  assign n16481 = pi15 ? n16480 : n16333;
  assign n16482 = pi19 ? n32 : n13376;
  assign n16483 = pi18 ? n32 : n16482;
  assign n16484 = pi17 ? n32 : n16483;
  assign n16485 = pi16 ? n32 : n16484;
  assign n16486 = pi20 ? n1839 : ~n10066;
  assign n16487 = pi19 ? n32 : n16486;
  assign n16488 = pi18 ? n32 : n16487;
  assign n16489 = pi17 ? n32 : n16488;
  assign n16490 = pi16 ? n32 : n16489;
  assign n16491 = pi15 ? n16485 : n16490;
  assign n16492 = pi14 ? n16481 : n16491;
  assign n16493 = pi13 ? n15981 : n16492;
  assign n16494 = pi12 ? n16475 : n16493;
  assign n16495 = pi20 ? n1839 : ~n14844;
  assign n16496 = pi19 ? n32 : n16495;
  assign n16497 = pi18 ? n32 : n16496;
  assign n16498 = pi17 ? n32 : n16497;
  assign n16499 = pi16 ? n32 : n16498;
  assign n16500 = pi15 ? n16413 : n16499;
  assign n16501 = pi14 ? n16500 : n16499;
  assign n16502 = pi20 ? n1839 : ~n749;
  assign n16503 = pi19 ? n32 : n16502;
  assign n16504 = pi18 ? n32 : n16503;
  assign n16505 = pi17 ? n32 : n16504;
  assign n16506 = pi16 ? n32 : n16505;
  assign n16507 = pi15 ? n16506 : n16413;
  assign n16508 = pi14 ? n16507 : n16413;
  assign n16509 = pi13 ? n16501 : n16508;
  assign n16510 = pi14 ? n16413 : n16333;
  assign n16511 = pi20 ? n7377 : n32;
  assign n16512 = pi19 ? n32 : n16511;
  assign n16513 = pi18 ? n32 : n16512;
  assign n16514 = pi17 ? n32 : n16513;
  assign n16515 = pi16 ? n32 : n16514;
  assign n16516 = pi15 ? n16333 : n16515;
  assign n16517 = pi19 ? n32 : n7881;
  assign n16518 = pi18 ? n32 : n16517;
  assign n16519 = pi17 ? n32 : n16518;
  assign n16520 = pi16 ? n32 : n16519;
  assign n16521 = pi21 ? n32 : ~n1392;
  assign n16522 = pi20 ? n16521 : n32;
  assign n16523 = pi19 ? n32 : n16522;
  assign n16524 = pi18 ? n32 : n16523;
  assign n16525 = pi17 ? n32 : n16524;
  assign n16526 = pi16 ? n32 : n16525;
  assign n16527 = pi15 ? n16520 : n16526;
  assign n16528 = pi14 ? n16516 : n16527;
  assign n16529 = pi13 ? n16510 : n16528;
  assign n16530 = pi12 ? n16509 : n16529;
  assign n16531 = pi11 ? n16494 : n16530;
  assign n16532 = pi10 ? n16531 : n32;
  assign n16533 = pi09 ? n16473 : n16532;
  assign n16534 = pi08 ? n16463 : n16533;
  assign n16535 = pi14 ? n16393 : n16397;
  assign n16536 = pi13 ? n32 : n16535;
  assign n16537 = pi12 ? n32 : n16536;
  assign n16538 = pi11 ? n32 : n16537;
  assign n16539 = pi10 ? n32 : n16538;
  assign n16540 = pi15 ? n16402 : n15987;
  assign n16541 = pi14 ? n16402 : n16540;
  assign n16542 = pi20 ? n518 : n32;
  assign n16543 = pi19 ? n32 : n16542;
  assign n16544 = pi18 ? n32 : n16543;
  assign n16545 = pi17 ? n32 : n16544;
  assign n16546 = pi16 ? n32 : n16545;
  assign n16547 = pi14 ? n15987 : n16546;
  assign n16548 = pi13 ? n16541 : n16547;
  assign n16549 = pi20 ? n1839 : ~n141;
  assign n16550 = pi19 ? n32 : n16549;
  assign n16551 = pi18 ? n32 : n16550;
  assign n16552 = pi17 ? n32 : n16551;
  assign n16553 = pi16 ? n32 : n16552;
  assign n16554 = pi15 ? n16553 : n16333;
  assign n16555 = pi20 ? n1839 : ~n342;
  assign n16556 = pi19 ? n32 : n16555;
  assign n16557 = pi18 ? n32 : n16556;
  assign n16558 = pi17 ? n32 : n16557;
  assign n16559 = pi16 ? n32 : n16558;
  assign n16560 = pi15 ? n16553 : n16559;
  assign n16561 = pi14 ? n16554 : n16560;
  assign n16562 = pi13 ? n15987 : n16561;
  assign n16563 = pi12 ? n16548 : n16562;
  assign n16564 = pi15 ? n16333 : n15981;
  assign n16565 = pi20 ? n1839 : n1445;
  assign n16566 = pi19 ? n32 : n16565;
  assign n16567 = pi18 ? n32 : n16566;
  assign n16568 = pi17 ? n32 : n16567;
  assign n16569 = pi16 ? n32 : n16568;
  assign n16570 = pi21 ? n140 : ~n140;
  assign n16571 = pi20 ? n1839 : n16570;
  assign n16572 = pi19 ? n32 : n16571;
  assign n16573 = pi18 ? n32 : n16572;
  assign n16574 = pi17 ? n32 : n16573;
  assign n16575 = pi16 ? n32 : n16574;
  assign n16576 = pi15 ? n16569 : n16575;
  assign n16577 = pi14 ? n16564 : n16576;
  assign n16578 = pi20 ? n1839 : ~n1475;
  assign n16579 = pi19 ? n32 : n16578;
  assign n16580 = pi18 ? n32 : n16579;
  assign n16581 = pi17 ? n32 : n16580;
  assign n16582 = pi16 ? n32 : n16581;
  assign n16583 = pi20 ? n14286 : ~n207;
  assign n16584 = pi19 ? n32 : n16583;
  assign n16585 = pi18 ? n32 : n16584;
  assign n16586 = pi17 ? n32 : n16585;
  assign n16587 = pi16 ? n32 : n16586;
  assign n16588 = pi15 ? n16582 : n16587;
  assign n16589 = pi14 ? n16582 : n16588;
  assign n16590 = pi13 ? n16577 : n16589;
  assign n16591 = pi20 ? n518 : ~n207;
  assign n16592 = pi19 ? n32 : n16591;
  assign n16593 = pi18 ? n32 : n16592;
  assign n16594 = pi17 ? n32 : n16593;
  assign n16595 = pi16 ? n32 : n16594;
  assign n16596 = pi14 ? n16595 : n16546;
  assign n16597 = pi20 ? n14968 : n32;
  assign n16598 = pi19 ? n32 : n16597;
  assign n16599 = pi18 ? n32 : n16598;
  assign n16600 = pi17 ? n32 : n16599;
  assign n16601 = pi16 ? n32 : n16600;
  assign n16602 = pi15 ? n16546 : n16601;
  assign n16603 = pi19 ? n32 : n9169;
  assign n16604 = pi18 ? n32 : n16603;
  assign n16605 = pi17 ? n32 : n16604;
  assign n16606 = pi16 ? n32 : n16605;
  assign n16607 = pi15 ? n16601 : n16606;
  assign n16608 = pi14 ? n16602 : n16607;
  assign n16609 = pi13 ? n16596 : n16608;
  assign n16610 = pi12 ? n16590 : n16609;
  assign n16611 = pi11 ? n16563 : n16610;
  assign n16612 = pi10 ? n16611 : n32;
  assign n16613 = pi09 ? n16539 : n16612;
  assign n16614 = pi15 ? n15987 : n16402;
  assign n16615 = pi14 ? n15987 : n16614;
  assign n16616 = pi20 ? n518 : n726;
  assign n16617 = pi19 ? n32 : n16616;
  assign n16618 = pi18 ? n32 : n16617;
  assign n16619 = pi17 ? n32 : n16618;
  assign n16620 = pi16 ? n32 : n16619;
  assign n16621 = pi15 ? n16546 : n16620;
  assign n16622 = pi14 ? n16546 : n16621;
  assign n16623 = pi13 ? n16615 : n16622;
  assign n16624 = pi12 ? n16548 : n16623;
  assign n16625 = pi20 ? n518 : ~n141;
  assign n16626 = pi19 ? n32 : n16625;
  assign n16627 = pi18 ? n32 : n16626;
  assign n16628 = pi17 ? n32 : n16627;
  assign n16629 = pi16 ? n32 : n16628;
  assign n16630 = pi15 ? n16629 : n15987;
  assign n16631 = pi19 ? n32 : n13638;
  assign n16632 = pi18 ? n32 : n16631;
  assign n16633 = pi17 ? n32 : n16632;
  assign n16634 = pi16 ? n32 : n16633;
  assign n16635 = pi20 ? n518 : n16570;
  assign n16636 = pi19 ? n32 : n16635;
  assign n16637 = pi18 ? n32 : n16636;
  assign n16638 = pi17 ? n32 : n16637;
  assign n16639 = pi16 ? n32 : n16638;
  assign n16640 = pi15 ? n16634 : n16639;
  assign n16641 = pi14 ? n16630 : n16640;
  assign n16642 = pi19 ? n32 : n13643;
  assign n16643 = pi18 ? n32 : n16642;
  assign n16644 = pi17 ? n32 : n16643;
  assign n16645 = pi16 ? n32 : n16644;
  assign n16646 = pi15 ? n16645 : n16587;
  assign n16647 = pi14 ? n16645 : n16646;
  assign n16648 = pi13 ? n16641 : n16647;
  assign n16649 = pi22 ? n34 : ~n50;
  assign n16650 = pi21 ? n32 : n16649;
  assign n16651 = pi20 ? n16650 : n32;
  assign n16652 = pi19 ? n32 : n16651;
  assign n16653 = pi18 ? n32 : n16652;
  assign n16654 = pi17 ? n32 : n16653;
  assign n16655 = pi16 ? n32 : n16654;
  assign n16656 = pi15 ? n16655 : n32;
  assign n16657 = pi14 ? n16602 : n16656;
  assign n16658 = pi13 ? n16596 : n16657;
  assign n16659 = pi12 ? n16648 : n16658;
  assign n16660 = pi11 ? n16624 : n16659;
  assign n16661 = pi10 ? n16660 : n32;
  assign n16662 = pi09 ? n16539 : n16661;
  assign n16663 = pi08 ? n16613 : n16662;
  assign n16664 = pi07 ? n16534 : n16663;
  assign n16665 = pi20 ? n2140 : ~n321;
  assign n16666 = pi19 ? n32 : n16665;
  assign n16667 = pi18 ? n32 : n16666;
  assign n16668 = pi17 ? n32 : n16667;
  assign n16669 = pi16 ? n32 : n16668;
  assign n16670 = pi15 ? n32 : n16669;
  assign n16671 = pi14 ? n16670 : n16669;
  assign n16672 = pi13 ? n32 : n16671;
  assign n16673 = pi12 ? n32 : n16672;
  assign n16674 = pi11 ? n32 : n16673;
  assign n16675 = pi10 ? n32 : n16674;
  assign n16676 = pi14 ? n16397 : n16403;
  assign n16677 = pi15 ? n16467 : n16402;
  assign n16678 = pi14 ? n16402 : n16677;
  assign n16679 = pi13 ? n16676 : n16678;
  assign n16680 = pi20 ? n518 : ~n10066;
  assign n16681 = pi19 ? n32 : n16680;
  assign n16682 = pi18 ? n32 : n16681;
  assign n16683 = pi17 ? n32 : n16682;
  assign n16684 = pi16 ? n32 : n16683;
  assign n16685 = pi15 ? n16629 : n16684;
  assign n16686 = pi15 ? n16629 : n16620;
  assign n16687 = pi14 ? n16685 : n16686;
  assign n16688 = pi13 ? n16402 : n16687;
  assign n16689 = pi12 ? n16679 : n16688;
  assign n16690 = pi20 ? n518 : ~n14844;
  assign n16691 = pi19 ? n32 : n16690;
  assign n16692 = pi18 ? n32 : n16691;
  assign n16693 = pi17 ? n32 : n16692;
  assign n16694 = pi16 ? n32 : n16693;
  assign n16695 = pi20 ? n14286 : ~n141;
  assign n16696 = pi19 ? n32 : n16695;
  assign n16697 = pi18 ? n32 : n16696;
  assign n16698 = pi17 ? n32 : n16697;
  assign n16699 = pi16 ? n32 : n16698;
  assign n16700 = pi15 ? n16694 : n16699;
  assign n16701 = pi15 ? n16634 : n16595;
  assign n16702 = pi14 ? n16700 : n16701;
  assign n16703 = pi19 ? n32 : n13651;
  assign n16704 = pi18 ? n32 : n16703;
  assign n16705 = pi17 ? n32 : n16704;
  assign n16706 = pi16 ? n32 : n16705;
  assign n16707 = pi15 ? n16546 : n16706;
  assign n16708 = pi19 ? n32 : n13662;
  assign n16709 = pi18 ? n32 : n16708;
  assign n16710 = pi17 ? n32 : n16709;
  assign n16711 = pi16 ? n32 : n16710;
  assign n16712 = pi14 ? n16707 : n16711;
  assign n16713 = pi13 ? n16702 : n16712;
  assign n16714 = pi20 ? n13785 : ~n207;
  assign n16715 = pi19 ? n32 : n16714;
  assign n16716 = pi18 ? n32 : n16715;
  assign n16717 = pi17 ? n32 : n16716;
  assign n16718 = pi16 ? n32 : n16717;
  assign n16719 = pi15 ? n16718 : n16467;
  assign n16720 = pi20 ? n1319 : ~n141;
  assign n16721 = pi19 ? n32 : n16720;
  assign n16722 = pi18 ? n32 : n16721;
  assign n16723 = pi17 ? n32 : n16722;
  assign n16724 = pi16 ? n32 : n16723;
  assign n16725 = pi15 ? n16724 : n16467;
  assign n16726 = pi14 ? n16719 : n16725;
  assign n16727 = pi14 ? n16655 : n32;
  assign n16728 = pi13 ? n16726 : n16727;
  assign n16729 = pi12 ? n16713 : n16728;
  assign n16730 = pi11 ? n16689 : n16729;
  assign n16731 = pi10 ? n16730 : n32;
  assign n16732 = pi09 ? n16675 : n16731;
  assign n16733 = pi19 ? n32 : n9591;
  assign n16734 = pi18 ? n32 : n16733;
  assign n16735 = pi17 ? n32 : n16734;
  assign n16736 = pi16 ? n32 : n16735;
  assign n16737 = pi15 ? n32 : n16736;
  assign n16738 = pi15 ? n16736 : n16669;
  assign n16739 = pi14 ? n16737 : n16738;
  assign n16740 = pi13 ? n32 : n16739;
  assign n16741 = pi12 ? n32 : n16740;
  assign n16742 = pi11 ? n32 : n16741;
  assign n16743 = pi10 ? n32 : n16742;
  assign n16744 = pi14 ? n16402 : n16397;
  assign n16745 = pi20 ? n1319 : ~n10066;
  assign n16746 = pi19 ? n32 : n16745;
  assign n16747 = pi18 ? n32 : n16746;
  assign n16748 = pi17 ? n32 : n16747;
  assign n16749 = pi16 ? n32 : n16748;
  assign n16750 = pi15 ? n16724 : n16749;
  assign n16751 = pi20 ? n1319 : n726;
  assign n16752 = pi19 ? n32 : n16751;
  assign n16753 = pi18 ? n32 : n16752;
  assign n16754 = pi17 ? n32 : n16753;
  assign n16755 = pi16 ? n32 : n16754;
  assign n16756 = pi15 ? n16724 : n16755;
  assign n16757 = pi14 ? n16750 : n16756;
  assign n16758 = pi13 ? n16744 : n16757;
  assign n16759 = pi12 ? n16679 : n16758;
  assign n16760 = pi20 ? n1319 : n266;
  assign n16761 = pi19 ? n32 : n16760;
  assign n16762 = pi18 ? n32 : n16761;
  assign n16763 = pi17 ? n32 : n16762;
  assign n16764 = pi16 ? n32 : n16763;
  assign n16765 = pi20 ? n13785 : ~n141;
  assign n16766 = pi19 ? n32 : n16765;
  assign n16767 = pi18 ? n32 : n16766;
  assign n16768 = pi17 ? n32 : n16767;
  assign n16769 = pi16 ? n32 : n16768;
  assign n16770 = pi15 ? n16764 : n16769;
  assign n16771 = pi20 ? n1319 : n1445;
  assign n16772 = pi19 ? n32 : n16771;
  assign n16773 = pi18 ? n32 : n16772;
  assign n16774 = pi17 ? n32 : n16773;
  assign n16775 = pi16 ? n32 : n16774;
  assign n16776 = pi15 ? n16775 : n16711;
  assign n16777 = pi14 ? n16770 : n16776;
  assign n16778 = pi15 ? n16467 : n16706;
  assign n16779 = pi14 ? n16778 : n16711;
  assign n16780 = pi13 ? n16777 : n16779;
  assign n16781 = pi15 ? n16718 : n16724;
  assign n16782 = pi14 ? n16781 : n16725;
  assign n16783 = pi19 ? n32 : n112;
  assign n16784 = pi18 ? n32 : n16783;
  assign n16785 = pi17 ? n32 : n16784;
  assign n16786 = pi16 ? n32 : n16785;
  assign n16787 = pi14 ? n16786 : n32;
  assign n16788 = pi13 ? n16782 : n16787;
  assign n16789 = pi12 ? n16780 : n16788;
  assign n16790 = pi11 ? n16759 : n16789;
  assign n16791 = pi10 ? n16790 : n32;
  assign n16792 = pi09 ? n16743 : n16791;
  assign n16793 = pi08 ? n16732 : n16792;
  assign n16794 = pi14 ? n16737 : n16736;
  assign n16795 = pi13 ? n32 : n16794;
  assign n16796 = pi12 ? n32 : n16795;
  assign n16797 = pi11 ? n32 : n16796;
  assign n16798 = pi10 ? n32 : n16797;
  assign n16799 = pi15 ? n16669 : n16397;
  assign n16800 = pi14 ? n16669 : n16799;
  assign n16801 = pi19 ? n32 : n5748;
  assign n16802 = pi18 ? n32 : n16801;
  assign n16803 = pi17 ? n32 : n16802;
  assign n16804 = pi16 ? n32 : n16803;
  assign n16805 = pi15 ? n16804 : n16397;
  assign n16806 = pi14 ? n16397 : n16805;
  assign n16807 = pi13 ? n16800 : n16806;
  assign n16808 = pi20 ? n1319 : ~n2140;
  assign n16809 = pi19 ? n32 : n16808;
  assign n16810 = pi18 ? n32 : n16809;
  assign n16811 = pi17 ? n32 : n16810;
  assign n16812 = pi16 ? n32 : n16811;
  assign n16813 = pi15 ? n16467 : n16812;
  assign n16814 = pi14 ? n16813 : n16756;
  assign n16815 = pi13 ? n16397 : n16814;
  assign n16816 = pi12 ? n16807 : n16815;
  assign n16817 = pi15 ? n16775 : n16724;
  assign n16818 = pi15 ? n16775 : n16706;
  assign n16819 = pi14 ? n16817 : n16818;
  assign n16820 = pi20 ? n342 : ~n1475;
  assign n16821 = pi19 ? n32 : n16820;
  assign n16822 = pi18 ? n32 : n16821;
  assign n16823 = pi17 ? n32 : n16822;
  assign n16824 = pi16 ? n32 : n16823;
  assign n16825 = pi15 ? n16392 : n16824;
  assign n16826 = pi14 ? n16825 : n16804;
  assign n16827 = pi13 ? n16819 : n16826;
  assign n16828 = pi20 ? n342 : ~n141;
  assign n16829 = pi19 ? n32 : n16828;
  assign n16830 = pi18 ? n32 : n16829;
  assign n16831 = pi17 ? n32 : n16830;
  assign n16832 = pi16 ? n32 : n16831;
  assign n16833 = pi15 ? n16804 : n16832;
  assign n16834 = pi19 ? n32 : n176;
  assign n16835 = pi18 ? n32 : n16834;
  assign n16836 = pi17 ? n32 : n16835;
  assign n16837 = pi16 ? n32 : n16836;
  assign n16838 = pi15 ? n16832 : n16837;
  assign n16839 = pi14 ? n16833 : n16838;
  assign n16840 = pi15 ? n16786 : n32;
  assign n16841 = pi14 ? n16840 : n32;
  assign n16842 = pi13 ? n16839 : n16841;
  assign n16843 = pi12 ? n16827 : n16842;
  assign n16844 = pi11 ? n16816 : n16843;
  assign n16845 = pi10 ? n16844 : n32;
  assign n16846 = pi09 ? n16798 : n16845;
  assign n16847 = pi19 ? n32 : n5694;
  assign n16848 = pi18 ? n32 : n16847;
  assign n16849 = pi17 ? n32 : n16848;
  assign n16850 = pi16 ? n32 : n16849;
  assign n16851 = pi15 ? n32 : n16850;
  assign n16852 = pi15 ? n16850 : n16736;
  assign n16853 = pi14 ? n16851 : n16852;
  assign n16854 = pi13 ? n32 : n16853;
  assign n16855 = pi12 ? n32 : n16854;
  assign n16856 = pi11 ? n32 : n16855;
  assign n16857 = pi10 ? n32 : n16856;
  assign n16858 = pi20 ? n2140 : ~n207;
  assign n16859 = pi19 ? n32 : n16858;
  assign n16860 = pi18 ? n32 : n16859;
  assign n16861 = pi17 ? n32 : n16860;
  assign n16862 = pi16 ? n32 : n16861;
  assign n16863 = pi15 ? n16862 : n16669;
  assign n16864 = pi14 ? n16799 : n16863;
  assign n16865 = pi13 ? n16800 : n16864;
  assign n16866 = pi19 ? n32 : n13906;
  assign n16867 = pi18 ? n32 : n16866;
  assign n16868 = pi17 ? n32 : n16867;
  assign n16869 = pi16 ? n32 : n16868;
  assign n16870 = pi15 ? n16392 : n16869;
  assign n16871 = pi20 ? n342 : n623;
  assign n16872 = pi19 ? n32 : n16871;
  assign n16873 = pi18 ? n32 : n16872;
  assign n16874 = pi17 ? n32 : n16873;
  assign n16875 = pi16 ? n32 : n16874;
  assign n16876 = pi15 ? n16832 : n16875;
  assign n16877 = pi14 ? n16870 : n16876;
  assign n16878 = pi13 ? n16669 : n16877;
  assign n16879 = pi12 ? n16865 : n16878;
  assign n16880 = pi20 ? n342 : n1445;
  assign n16881 = pi19 ? n32 : n16880;
  assign n16882 = pi18 ? n32 : n16881;
  assign n16883 = pi17 ? n32 : n16882;
  assign n16884 = pi16 ? n32 : n16883;
  assign n16885 = pi15 ? n16884 : n16832;
  assign n16886 = pi20 ? n342 : n439;
  assign n16887 = pi19 ? n32 : n16886;
  assign n16888 = pi18 ? n32 : n16887;
  assign n16889 = pi17 ? n32 : n16888;
  assign n16890 = pi16 ? n32 : n16889;
  assign n16891 = pi15 ? n16890 : n16824;
  assign n16892 = pi14 ? n16885 : n16891;
  assign n16893 = pi15 ? n16392 : n16804;
  assign n16894 = pi14 ? n16893 : n16804;
  assign n16895 = pi13 ? n16892 : n16894;
  assign n16896 = pi19 ? n32 : n13388;
  assign n16897 = pi18 ? n32 : n16896;
  assign n16898 = pi17 ? n32 : n16897;
  assign n16899 = pi16 ? n32 : n16898;
  assign n16900 = pi15 ? n16899 : n32;
  assign n16901 = pi14 ? n16832 : n16900;
  assign n16902 = pi13 ? n16901 : n32;
  assign n16903 = pi12 ? n16895 : n16902;
  assign n16904 = pi11 ? n16879 : n16903;
  assign n16905 = pi10 ? n16904 : n32;
  assign n16906 = pi09 ? n16857 : n16905;
  assign n16907 = pi08 ? n16846 : n16906;
  assign n16908 = pi07 ? n16793 : n16907;
  assign n16909 = pi06 ? n16664 : n16908;
  assign n16910 = pi19 ? n32 : n102;
  assign n16911 = pi18 ? n32 : n16910;
  assign n16912 = pi17 ? n32 : n16911;
  assign n16913 = pi16 ? n32 : n16912;
  assign n16914 = pi15 ? n32 : n16913;
  assign n16915 = pi20 ? n101 : ~n321;
  assign n16916 = pi19 ? n32 : n16915;
  assign n16917 = pi18 ? n32 : n16916;
  assign n16918 = pi17 ? n32 : n16917;
  assign n16919 = pi16 ? n32 : n16918;
  assign n16920 = pi14 ? n16914 : n16919;
  assign n16921 = pi13 ? n32 : n16920;
  assign n16922 = pi12 ? n32 : n16921;
  assign n16923 = pi11 ? n32 : n16922;
  assign n16924 = pi10 ? n32 : n16923;
  assign n16925 = pi14 ? n16736 : n16738;
  assign n16926 = pi20 ? n67 : ~n321;
  assign n16927 = pi19 ? n32 : n16926;
  assign n16928 = pi18 ? n32 : n16927;
  assign n16929 = pi17 ? n32 : n16928;
  assign n16930 = pi16 ? n32 : n16929;
  assign n16931 = pi15 ? n16669 : n16930;
  assign n16932 = pi14 ? n16931 : n16669;
  assign n16933 = pi13 ? n16925 : n16932;
  assign n16934 = pi20 ? n342 : n8760;
  assign n16935 = pi19 ? n32 : n16934;
  assign n16936 = pi18 ? n32 : n16935;
  assign n16937 = pi17 ? n32 : n16936;
  assign n16938 = pi16 ? n32 : n16937;
  assign n16939 = pi15 ? n16392 : n16938;
  assign n16940 = pi15 ? n16392 : n16832;
  assign n16941 = pi14 ? n16939 : n16940;
  assign n16942 = pi13 ? n16669 : n16941;
  assign n16943 = pi12 ? n16933 : n16942;
  assign n16944 = pi20 ? n2140 : ~n287;
  assign n16945 = pi19 ? n32 : n16944;
  assign n16946 = pi18 ? n32 : n16945;
  assign n16947 = pi17 ? n32 : n16946;
  assign n16948 = pi16 ? n32 : n16947;
  assign n16949 = pi20 ? n2140 : ~n141;
  assign n16950 = pi19 ? n32 : n16949;
  assign n16951 = pi18 ? n32 : n16950;
  assign n16952 = pi17 ? n32 : n16951;
  assign n16953 = pi16 ? n32 : n16952;
  assign n16954 = pi15 ? n16948 : n16953;
  assign n16955 = pi20 ? n2140 : ~n1475;
  assign n16956 = pi19 ? n32 : n16955;
  assign n16957 = pi18 ? n32 : n16956;
  assign n16958 = pi17 ? n32 : n16957;
  assign n16959 = pi16 ? n32 : n16958;
  assign n16960 = pi15 ? n16953 : n16959;
  assign n16961 = pi14 ? n16954 : n16960;
  assign n16962 = pi19 ? n32 : n6324;
  assign n16963 = pi18 ? n32 : n16962;
  assign n16964 = pi17 ? n32 : n16963;
  assign n16965 = pi16 ? n32 : n16964;
  assign n16966 = pi15 ? n16862 : n16965;
  assign n16967 = pi14 ? n16966 : n16862;
  assign n16968 = pi13 ? n16961 : n16967;
  assign n16969 = pi20 ? n2077 : n32;
  assign n16970 = pi19 ? n32 : n16969;
  assign n16971 = pi18 ? n32 : n16970;
  assign n16972 = pi17 ? n32 : n16971;
  assign n16973 = pi16 ? n32 : n16972;
  assign n16974 = pi15 ? n16973 : n32;
  assign n16975 = pi14 ? n16953 : n16974;
  assign n16976 = pi13 ? n16975 : n32;
  assign n16977 = pi12 ? n16968 : n16976;
  assign n16978 = pi11 ? n16943 : n16977;
  assign n16979 = pi10 ? n16978 : n32;
  assign n16980 = pi09 ? n16924 : n16979;
  assign n16981 = pi19 ? n32 : n8622;
  assign n16982 = pi18 ? n32 : n16981;
  assign n16983 = pi17 ? n32 : n16982;
  assign n16984 = pi16 ? n32 : n16983;
  assign n16985 = pi15 ? n32 : n16984;
  assign n16986 = pi14 ? n16985 : n16919;
  assign n16987 = pi13 ? n32 : n16986;
  assign n16988 = pi12 ? n32 : n16987;
  assign n16989 = pi11 ? n32 : n16988;
  assign n16990 = pi10 ? n32 : n16989;
  assign n16991 = pi20 ? n2140 : ~n16008;
  assign n16992 = pi19 ? n32 : n16991;
  assign n16993 = pi18 ? n32 : n16992;
  assign n16994 = pi17 ? n32 : n16993;
  assign n16995 = pi16 ? n32 : n16994;
  assign n16996 = pi15 ? n16953 : n16995;
  assign n16997 = pi21 ? n32 : n14399;
  assign n16998 = pi20 ? n16997 : n32;
  assign n16999 = pi19 ? n32 : n16998;
  assign n17000 = pi18 ? n32 : n16999;
  assign n17001 = pi17 ? n32 : n17000;
  assign n17002 = pi16 ? n32 : n17001;
  assign n17003 = pi15 ? n17002 : n16953;
  assign n17004 = pi14 ? n16996 : n17003;
  assign n17005 = pi13 ? n16736 : n17004;
  assign n17006 = pi12 ? n16736 : n17005;
  assign n17007 = pi15 ? n16948 : n16965;
  assign n17008 = pi14 ? n17007 : n16960;
  assign n17009 = pi20 ? n2140 : ~n339;
  assign n17010 = pi19 ? n32 : n17009;
  assign n17011 = pi18 ? n32 : n17010;
  assign n17012 = pi17 ? n32 : n17011;
  assign n17013 = pi16 ? n32 : n17012;
  assign n17014 = pi15 ? n16862 : n17013;
  assign n17015 = pi14 ? n16966 : n17014;
  assign n17016 = pi13 ? n17008 : n17015;
  assign n17017 = pi15 ? n16953 : n16973;
  assign n17018 = pi14 ? n17017 : n32;
  assign n17019 = pi13 ? n17018 : n32;
  assign n17020 = pi12 ? n17016 : n17019;
  assign n17021 = pi11 ? n17006 : n17020;
  assign n17022 = pi10 ? n17021 : n32;
  assign n17023 = pi09 ? n16990 : n17022;
  assign n17024 = pi08 ? n16980 : n17023;
  assign n17025 = pi14 ? n16985 : n16850;
  assign n17026 = pi13 ? n32 : n17025;
  assign n17027 = pi12 ? n32 : n17026;
  assign n17028 = pi11 ? n32 : n17027;
  assign n17029 = pi10 ? n32 : n17028;
  assign n17030 = pi15 ? n16919 : n16736;
  assign n17031 = pi14 ? n17030 : n16736;
  assign n17032 = pi13 ? n16919 : n17031;
  assign n17033 = pi19 ? n32 : n13680;
  assign n17034 = pi18 ? n32 : n17033;
  assign n17035 = pi17 ? n32 : n17034;
  assign n17036 = pi16 ? n32 : n17035;
  assign n17037 = pi18 ? n32 : n6071;
  assign n17038 = pi17 ? n32 : n17037;
  assign n17039 = pi16 ? n32 : n17038;
  assign n17040 = pi14 ? n17036 : n17039;
  assign n17041 = pi13 ? n16736 : n17040;
  assign n17042 = pi12 ? n17032 : n17041;
  assign n17043 = pi15 ? n17036 : n17039;
  assign n17044 = pi22 ? n50 : ~n34;
  assign n17045 = pi21 ? n17044 : n32;
  assign n17046 = pi20 ? n428 : n17045;
  assign n17047 = pi19 ? n32 : n17046;
  assign n17048 = pi18 ? n32 : n17047;
  assign n17049 = pi17 ? n32 : n17048;
  assign n17050 = pi16 ? n32 : n17049;
  assign n17051 = pi15 ? n17050 : n16953;
  assign n17052 = pi14 ? n17043 : n17051;
  assign n17053 = pi19 ? n32 : n13926;
  assign n17054 = pi18 ? n32 : n17053;
  assign n17055 = pi17 ? n32 : n17054;
  assign n17056 = pi16 ? n32 : n17055;
  assign n17057 = pi15 ? n17056 : n17039;
  assign n17058 = pi19 ? n32 : n7349;
  assign n17059 = pi18 ? n32 : n17058;
  assign n17060 = pi17 ? n32 : n17059;
  assign n17061 = pi16 ? n32 : n17060;
  assign n17062 = pi20 ? n428 : ~n339;
  assign n17063 = pi19 ? n32 : n17062;
  assign n17064 = pi18 ? n32 : n17063;
  assign n17065 = pi17 ? n32 : n17064;
  assign n17066 = pi16 ? n32 : n17065;
  assign n17067 = pi15 ? n17061 : n17066;
  assign n17068 = pi14 ? n17057 : n17067;
  assign n17069 = pi13 ? n17052 : n17068;
  assign n17070 = pi15 ? n17036 : n32;
  assign n17071 = pi14 ? n17070 : n32;
  assign n17072 = pi13 ? n17071 : n32;
  assign n17073 = pi12 ? n17069 : n17072;
  assign n17074 = pi11 ? n17042 : n17073;
  assign n17075 = pi10 ? n17074 : n32;
  assign n17076 = pi09 ? n17029 : n17075;
  assign n17077 = pi14 ? n32 : n16850;
  assign n17078 = pi13 ? n32 : n17077;
  assign n17079 = pi12 ? n32 : n17078;
  assign n17080 = pi11 ? n32 : n17079;
  assign n17081 = pi10 ? n32 : n17080;
  assign n17082 = pi14 ? n16919 : n16850;
  assign n17083 = pi15 ? n16850 : n16919;
  assign n17084 = pi14 ? n17083 : n16852;
  assign n17085 = pi13 ? n17082 : n17084;
  assign n17086 = pi20 ? n101 : ~n141;
  assign n17087 = pi19 ? n32 : n17086;
  assign n17088 = pi18 ? n32 : n17087;
  assign n17089 = pi17 ? n32 : n17088;
  assign n17090 = pi16 ? n32 : n17089;
  assign n17091 = pi15 ? n17090 : n17036;
  assign n17092 = pi14 ? n17090 : n17091;
  assign n17093 = pi13 ? n16919 : n17092;
  assign n17094 = pi12 ? n17085 : n17093;
  assign n17095 = pi15 ? n17056 : n17036;
  assign n17096 = pi14 ? n17036 : n17095;
  assign n17097 = pi15 ? n17061 : n16984;
  assign n17098 = pi14 ? n17057 : n17097;
  assign n17099 = pi13 ? n17096 : n17098;
  assign n17100 = pi15 ? n17090 : n32;
  assign n17101 = pi14 ? n17100 : n32;
  assign n17102 = pi13 ? n17101 : n32;
  assign n17103 = pi12 ? n17099 : n17102;
  assign n17104 = pi11 ? n17094 : n17103;
  assign n17105 = pi10 ? n17104 : n32;
  assign n17106 = pi09 ? n17081 : n17105;
  assign n17107 = pi08 ? n17076 : n17106;
  assign n17108 = pi07 ? n17024 : n17107;
  assign n17109 = pi18 ? n32 : n127;
  assign n17110 = pi17 ? n32 : n17109;
  assign n17111 = pi16 ? n32 : n17110;
  assign n17112 = pi15 ? n32 : n17111;
  assign n17113 = pi14 ? n17112 : n32;
  assign n17114 = pi13 ? n32 : n17113;
  assign n17115 = pi12 ? n32 : n17114;
  assign n17116 = pi11 ? n32 : n17115;
  assign n17117 = pi10 ? n32 : n17116;
  assign n17118 = pi19 ? n32 : n9007;
  assign n17119 = pi18 ? n32 : n17118;
  assign n17120 = pi17 ? n32 : n17119;
  assign n17121 = pi16 ? n32 : n17120;
  assign n17122 = pi15 ? n17121 : n16984;
  assign n17123 = pi14 ? n17121 : n17122;
  assign n17124 = pi20 ? n101 : ~n207;
  assign n17125 = pi19 ? n32 : n17124;
  assign n17126 = pi18 ? n32 : n17125;
  assign n17127 = pi17 ? n32 : n17126;
  assign n17128 = pi16 ? n32 : n17127;
  assign n17129 = pi15 ? n17128 : n16919;
  assign n17130 = pi14 ? n17122 : n17129;
  assign n17131 = pi13 ? n17123 : n17130;
  assign n17132 = pi14 ? n17128 : n17129;
  assign n17133 = pi15 ? n17090 : n16913;
  assign n17134 = pi21 ? n124 : n206;
  assign n17135 = pi20 ? n32 : ~n17134;
  assign n17136 = pi19 ? n32 : n17135;
  assign n17137 = pi18 ? n32 : n17136;
  assign n17138 = pi17 ? n32 : n17137;
  assign n17139 = pi16 ? n32 : n17138;
  assign n17140 = pi21 ? n1392 : n259;
  assign n17141 = pi20 ? n101 : ~n17140;
  assign n17142 = pi19 ? n32 : n17141;
  assign n17143 = pi18 ? n32 : n17142;
  assign n17144 = pi17 ? n32 : n17143;
  assign n17145 = pi16 ? n32 : n17144;
  assign n17146 = pi15 ? n17139 : n17145;
  assign n17147 = pi14 ? n17133 : n17146;
  assign n17148 = pi13 ? n17132 : n17147;
  assign n17149 = pi12 ? n17131 : n17148;
  assign n17150 = pi18 ? n32 : n625;
  assign n17151 = pi17 ? n32 : n17150;
  assign n17152 = pi16 ? n32 : n17151;
  assign n17153 = pi20 ? n428 : ~n13269;
  assign n17154 = pi19 ? n32 : n17153;
  assign n17155 = pi18 ? n32 : n17154;
  assign n17156 = pi17 ? n32 : n17155;
  assign n17157 = pi16 ? n32 : n17156;
  assign n17158 = pi15 ? n17152 : n17157;
  assign n17159 = pi21 ? n10182 : ~n32;
  assign n17160 = pi20 ? n428 : ~n17159;
  assign n17161 = pi19 ? n32 : n17160;
  assign n17162 = pi18 ? n32 : n17161;
  assign n17163 = pi17 ? n32 : n17162;
  assign n17164 = pi16 ? n32 : n17163;
  assign n17165 = pi14 ? n17158 : n17164;
  assign n17166 = pi20 ? n101 : ~n339;
  assign n17167 = pi19 ? n32 : n17166;
  assign n17168 = pi18 ? n32 : n17167;
  assign n17169 = pi17 ? n32 : n17168;
  assign n17170 = pi16 ? n32 : n17169;
  assign n17171 = pi15 ? n17170 : n32;
  assign n17172 = pi14 ? n17128 : n17171;
  assign n17173 = pi13 ? n17165 : n17172;
  assign n17174 = pi12 ? n17173 : n32;
  assign n17175 = pi11 ? n17149 : n17174;
  assign n17176 = pi10 ? n17175 : n32;
  assign n17177 = pi09 ? n17117 : n17176;
  assign n17178 = pi15 ? n17121 : n32;
  assign n17179 = pi14 ? n17121 : n17178;
  assign n17180 = pi14 ? n17178 : n17129;
  assign n17181 = pi13 ? n17179 : n17180;
  assign n17182 = pi15 ? n17128 : n17121;
  assign n17183 = pi15 ? n17121 : n16850;
  assign n17184 = pi14 ? n17182 : n17183;
  assign n17185 = pi19 ? n32 : n142;
  assign n17186 = pi18 ? n32 : n17185;
  assign n17187 = pi17 ? n32 : n17186;
  assign n17188 = pi16 ? n32 : n17187;
  assign n17189 = pi15 ? n17188 : n32;
  assign n17190 = pi19 ? n32 : n14139;
  assign n17191 = pi18 ? n32 : n17190;
  assign n17192 = pi17 ? n32 : n17191;
  assign n17193 = pi16 ? n32 : n17192;
  assign n17194 = pi20 ? n32 : ~n287;
  assign n17195 = pi19 ? n32 : n17194;
  assign n17196 = pi18 ? n32 : n17195;
  assign n17197 = pi17 ? n32 : n17196;
  assign n17198 = pi16 ? n32 : n17197;
  assign n17199 = pi15 ? n17193 : n17198;
  assign n17200 = pi14 ? n17189 : n17199;
  assign n17201 = pi13 ? n17184 : n17200;
  assign n17202 = pi12 ? n17181 : n17201;
  assign n17203 = pi18 ? n32 : n1447;
  assign n17204 = pi17 ? n32 : n17203;
  assign n17205 = pi16 ? n32 : n17204;
  assign n17206 = pi20 ? n101 : n1445;
  assign n17207 = pi19 ? n32 : n17206;
  assign n17208 = pi18 ? n32 : n17207;
  assign n17209 = pi17 ? n32 : n17208;
  assign n17210 = pi16 ? n32 : n17209;
  assign n17211 = pi15 ? n17205 : n17210;
  assign n17212 = pi20 ? n32 : ~n1475;
  assign n17213 = pi19 ? n32 : n17212;
  assign n17214 = pi18 ? n32 : n17213;
  assign n17215 = pi17 ? n32 : n17214;
  assign n17216 = pi16 ? n32 : n17215;
  assign n17217 = pi20 ? n101 : n17045;
  assign n17218 = pi19 ? n32 : n17217;
  assign n17219 = pi18 ? n32 : n17218;
  assign n17220 = pi17 ? n32 : n17219;
  assign n17221 = pi16 ? n32 : n17220;
  assign n17222 = pi15 ? n17216 : n17221;
  assign n17223 = pi14 ? n17211 : n17222;
  assign n17224 = pi20 ? n101 : ~n1940;
  assign n17225 = pi19 ? n32 : n17224;
  assign n17226 = pi18 ? n32 : n17225;
  assign n17227 = pi17 ? n32 : n17226;
  assign n17228 = pi16 ? n32 : n17227;
  assign n17229 = pi15 ? n17228 : n17121;
  assign n17230 = pi15 ? n16984 : n17090;
  assign n17231 = pi14 ? n17229 : n17230;
  assign n17232 = pi13 ? n17223 : n17231;
  assign n17233 = pi12 ? n17232 : n32;
  assign n17234 = pi11 ? n17202 : n17233;
  assign n17235 = pi10 ? n17234 : n32;
  assign n17236 = pi09 ? n17117 : n17235;
  assign n17237 = pi08 ? n17177 : n17236;
  assign n17238 = pi15 ? n16984 : n16850;
  assign n17239 = pi14 ? n32 : n17238;
  assign n17240 = pi13 ? n32 : n17239;
  assign n17241 = pi15 ? n16984 : n17121;
  assign n17242 = pi14 ? n17241 : n17183;
  assign n17243 = pi15 ? n17193 : n17111;
  assign n17244 = pi14 ? n17188 : n17243;
  assign n17245 = pi13 ? n17242 : n17244;
  assign n17246 = pi12 ? n17240 : n17245;
  assign n17247 = pi20 ? n101 : ~n518;
  assign n17248 = pi19 ? n32 : n17247;
  assign n17249 = pi18 ? n32 : n17248;
  assign n17250 = pi17 ? n32 : n17249;
  assign n17251 = pi16 ? n32 : n17250;
  assign n17252 = pi19 ? n32 : n13934;
  assign n17253 = pi18 ? n32 : n17252;
  assign n17254 = pi17 ? n32 : n17253;
  assign n17255 = pi16 ? n32 : n17254;
  assign n17256 = pi14 ? n17251 : n17255;
  assign n17257 = pi20 ? n32 : ~n1940;
  assign n17258 = pi19 ? n32 : n17257;
  assign n17259 = pi18 ? n32 : n17258;
  assign n17260 = pi17 ? n32 : n17259;
  assign n17261 = pi16 ? n32 : n17260;
  assign n17262 = pi15 ? n17261 : n17121;
  assign n17263 = pi14 ? n17262 : n17230;
  assign n17264 = pi13 ? n17256 : n17263;
  assign n17265 = pi12 ? n17264 : n32;
  assign n17266 = pi11 ? n17246 : n17265;
  assign n17267 = pi10 ? n17266 : n32;
  assign n17268 = pi09 ? n32 : n17267;
  assign n17269 = pi14 ? n32 : n16851;
  assign n17270 = pi13 ? n32 : n17269;
  assign n17271 = pi15 ? n32 : n17121;
  assign n17272 = pi14 ? n17271 : n17183;
  assign n17273 = pi15 ? n32 : n17188;
  assign n17274 = pi20 ? n32 : n9000;
  assign n17275 = pi19 ? n32 : n17274;
  assign n17276 = pi18 ? n32 : n17275;
  assign n17277 = pi17 ? n32 : n17276;
  assign n17278 = pi16 ? n32 : n17277;
  assign n17279 = pi15 ? n17278 : n32;
  assign n17280 = pi14 ? n17273 : n17279;
  assign n17281 = pi13 ? n17272 : n17280;
  assign n17282 = pi12 ? n17270 : n17281;
  assign n17283 = pi19 ? n32 : n5730;
  assign n17284 = pi18 ? n32 : n17283;
  assign n17285 = pi17 ? n32 : n17284;
  assign n17286 = pi16 ? n32 : n17285;
  assign n17287 = pi21 ? n124 : ~n32;
  assign n17288 = pi20 ? n32 : ~n17287;
  assign n17289 = pi19 ? n32 : n17288;
  assign n17290 = pi18 ? n32 : n17289;
  assign n17291 = pi17 ? n32 : n17290;
  assign n17292 = pi16 ? n32 : n17291;
  assign n17293 = pi15 ? n17286 : n17292;
  assign n17294 = pi20 ? n32 : n7501;
  assign n17295 = pi19 ? n32 : n17294;
  assign n17296 = pi18 ? n32 : n17295;
  assign n17297 = pi17 ? n32 : n17296;
  assign n17298 = pi16 ? n32 : n17297;
  assign n17299 = pi15 ? n17255 : n17298;
  assign n17300 = pi14 ? n17293 : n17299;
  assign n17301 = pi14 ? n17122 : n17189;
  assign n17302 = pi13 ? n17300 : n17301;
  assign n17303 = pi12 ? n17302 : n32;
  assign n17304 = pi11 ? n17282 : n17303;
  assign n17305 = pi10 ? n17304 : n32;
  assign n17306 = pi09 ? n32 : n17305;
  assign n17307 = pi08 ? n17268 : n17306;
  assign n17308 = pi07 ? n17237 : n17307;
  assign n17309 = pi06 ? n17108 : n17308;
  assign n17310 = pi05 ? n16909 : n17309;
  assign n17311 = pi04 ? n16388 : n17310;
  assign n17312 = pi03 ? n13964 : n17311;
  assign n17313 = pi14 ? n32 : n16985;
  assign n17314 = pi18 ? n32 : n262;
  assign n17315 = pi17 ? n32 : n17314;
  assign n17316 = pi16 ? n32 : n17315;
  assign n17317 = pi15 ? n17316 : n32;
  assign n17318 = pi14 ? n17317 : n17279;
  assign n17319 = pi13 ? n17313 : n17318;
  assign n17320 = pi12 ? n32 : n17319;
  assign n17321 = pi20 ? n32 : ~n14844;
  assign n17322 = pi19 ? n32 : n17321;
  assign n17323 = pi18 ? n32 : n17322;
  assign n17324 = pi17 ? n32 : n17323;
  assign n17325 = pi16 ? n32 : n17324;
  assign n17326 = pi15 ? n17205 : n17325;
  assign n17327 = pi20 ? n32 : n17045;
  assign n17328 = pi19 ? n32 : n17327;
  assign n17329 = pi18 ? n32 : n17328;
  assign n17330 = pi17 ? n32 : n17329;
  assign n17331 = pi16 ? n32 : n17330;
  assign n17332 = pi20 ? n32 : n52;
  assign n17333 = pi19 ? n32 : n17332;
  assign n17334 = pi18 ? n32 : n17333;
  assign n17335 = pi17 ? n32 : n17334;
  assign n17336 = pi16 ? n32 : n17335;
  assign n17337 = pi15 ? n17331 : n17336;
  assign n17338 = pi14 ? n17326 : n17337;
  assign n17339 = pi13 ? n17338 : n17301;
  assign n17340 = pi12 ? n17339 : n32;
  assign n17341 = pi11 ? n17320 : n17340;
  assign n17342 = pi10 ? n17341 : n32;
  assign n17343 = pi09 ? n32 : n17342;
  assign n17344 = pi13 ? n32 : n17279;
  assign n17345 = pi12 ? n32 : n17344;
  assign n17346 = pi18 ? n32 : n268;
  assign n17347 = pi17 ? n32 : n17346;
  assign n17348 = pi16 ? n32 : n17347;
  assign n17349 = pi15 ? n17205 : n17348;
  assign n17350 = pi14 ? n17349 : n17337;
  assign n17351 = pi13 ? n17350 : n17301;
  assign n17352 = pi12 ? n17351 : n32;
  assign n17353 = pi11 ? n17345 : n17352;
  assign n17354 = pi10 ? n17353 : n32;
  assign n17355 = pi09 ? n32 : n17354;
  assign n17356 = pi08 ? n17343 : n17355;
  assign n17357 = pi15 ? n17205 : n32;
  assign n17358 = pi14 ? n17279 : n17357;
  assign n17359 = pi13 ? n32 : n17358;
  assign n17360 = pi12 ? n32 : n17359;
  assign n17361 = pi18 ? n32 : n566;
  assign n17362 = pi17 ? n32 : n17361;
  assign n17363 = pi16 ? n32 : n17362;
  assign n17364 = pi15 ? n17363 : n32;
  assign n17365 = pi18 ? n32 : n1012;
  assign n17366 = pi17 ? n32 : n17365;
  assign n17367 = pi16 ? n32 : n17366;
  assign n17368 = pi15 ? n17367 : n32;
  assign n17369 = pi14 ? n17364 : n17368;
  assign n17370 = pi13 ? n17369 : n32;
  assign n17371 = pi12 ? n17370 : n32;
  assign n17372 = pi11 ? n17360 : n17371;
  assign n17373 = pi10 ? n17372 : n32;
  assign n17374 = pi09 ? n32 : n17373;
  assign n17375 = pi14 ? n17273 : n32;
  assign n17376 = pi13 ? n17369 : n17375;
  assign n17377 = pi12 ? n17376 : n32;
  assign n17378 = pi11 ? n17360 : n17377;
  assign n17379 = pi10 ? n17378 : n32;
  assign n17380 = pi09 ? n32 : n17379;
  assign n17381 = pi08 ? n17374 : n17380;
  assign n17382 = pi07 ? n17356 : n17381;
  assign n17383 = pi20 ? n32 : n8760;
  assign n17384 = pi19 ? n32 : n17383;
  assign n17385 = pi18 ? n32 : n17384;
  assign n17386 = pi17 ? n32 : n17385;
  assign n17387 = pi16 ? n32 : n17386;
  assign n17388 = pi15 ? n17387 : n32;
  assign n17389 = pi21 ? n1009 : ~n259;
  assign n17390 = pi20 ? n32 : n17389;
  assign n17391 = pi19 ? n32 : n17390;
  assign n17392 = pi18 ? n32 : n17391;
  assign n17393 = pi17 ? n32 : n17392;
  assign n17394 = pi16 ? n32 : n17393;
  assign n17395 = pi15 ? n17394 : n32;
  assign n17396 = pi14 ? n17388 : n17395;
  assign n17397 = pi13 ? n32 : n17396;
  assign n17398 = pi12 ? n32 : n17397;
  assign n17399 = pi14 ? n17368 : n17178;
  assign n17400 = pi13 ? n17399 : n17375;
  assign n17401 = pi12 ? n17400 : n32;
  assign n17402 = pi11 ? n17398 : n17401;
  assign n17403 = pi10 ? n17402 : n32;
  assign n17404 = pi09 ? n32 : n17403;
  assign n17405 = pi13 ? n17399 : n32;
  assign n17406 = pi12 ? n17405 : n32;
  assign n17407 = pi11 ? n17398 : n17406;
  assign n17408 = pi10 ? n17407 : n32;
  assign n17409 = pi09 ? n32 : n17408;
  assign n17410 = pi08 ? n17404 : n17409;
  assign n17411 = pi14 ? n32 : n17271;
  assign n17412 = pi15 ? n16984 : n32;
  assign n17413 = pi14 ? n17412 : n32;
  assign n17414 = pi13 ? n17411 : n17413;
  assign n17415 = pi12 ? n17414 : n32;
  assign n17416 = pi11 ? n32 : n17415;
  assign n17417 = pi10 ? n17416 : n32;
  assign n17418 = pi09 ? n32 : n17417;
  assign n17419 = pi07 ? n17410 : n17418;
  assign n17420 = pi06 ? n17382 : n17419;
  assign n17421 = pi15 ? n32 : n17316;
  assign n17422 = pi15 ? n32 : n17152;
  assign n17423 = pi14 ? n17421 : n17422;
  assign n17424 = pi13 ? n32 : n17423;
  assign n17425 = pi12 ? n32 : n17424;
  assign n17426 = pi18 ? n32 : n917;
  assign n17427 = pi17 ? n32 : n17426;
  assign n17428 = pi16 ? n32 : n17427;
  assign n17429 = pi18 ? n32 : n573;
  assign n17430 = pi17 ? n32 : n17429;
  assign n17431 = pi16 ? n32 : n17430;
  assign n17432 = pi15 ? n17428 : n17431;
  assign n17433 = pi18 ? n32 : n463;
  assign n17434 = pi17 ? n32 : n17433;
  assign n17435 = pi16 ? n32 : n17434;
  assign n17436 = pi15 ? n17435 : n16984;
  assign n17437 = pi14 ? n17432 : n17436;
  assign n17438 = pi13 ? n17437 : n32;
  assign n17439 = pi12 ? n17438 : n32;
  assign n17440 = pi11 ? n17425 : n17439;
  assign n17441 = pi10 ? n17440 : n32;
  assign n17442 = pi09 ? n32 : n17441;
  assign n17443 = pi15 ? n32 : n17278;
  assign n17444 = pi15 ? n32 : n17205;
  assign n17445 = pi14 ? n17443 : n17444;
  assign n17446 = pi13 ? n32 : n17445;
  assign n17447 = pi12 ? n32 : n17446;
  assign n17448 = pi15 ? n17363 : n17331;
  assign n17449 = pi21 ? n14792 : n32;
  assign n17450 = pi20 ? n32 : n17449;
  assign n17451 = pi19 ? n32 : n17450;
  assign n17452 = pi18 ? n32 : n17451;
  assign n17453 = pi17 ? n32 : n17452;
  assign n17454 = pi16 ? n32 : n17453;
  assign n17455 = pi15 ? n17454 : n16984;
  assign n17456 = pi14 ? n17448 : n17455;
  assign n17457 = pi13 ? n17456 : n32;
  assign n17458 = pi12 ? n17457 : n32;
  assign n17459 = pi11 ? n17447 : n17458;
  assign n17460 = pi10 ? n17459 : n32;
  assign n17461 = pi09 ? n32 : n17460;
  assign n17462 = pi08 ? n17442 : n17461;
  assign n17463 = pi18 ? n32 : n222;
  assign n17464 = pi17 ? n32 : n17463;
  assign n17465 = pi16 ? n32 : n17464;
  assign n17466 = pi15 ? n32 : n17465;
  assign n17467 = pi14 ? n17466 : n17444;
  assign n17468 = pi13 ? n32 : n17467;
  assign n17469 = pi12 ? n32 : n17468;
  assign n17470 = pi15 ? n17454 : n17188;
  assign n17471 = pi14 ? n17448 : n17470;
  assign n17472 = pi13 ? n17471 : n32;
  assign n17473 = pi12 ? n17472 : n32;
  assign n17474 = pi11 ? n17469 : n17473;
  assign n17475 = pi10 ? n17474 : n32;
  assign n17476 = pi09 ? n32 : n17475;
  assign n17477 = pi15 ? n17363 : n17454;
  assign n17478 = pi14 ? n17477 : n32;
  assign n17479 = pi13 ? n17478 : n32;
  assign n17480 = pi12 ? n17479 : n32;
  assign n17481 = pi11 ? n17469 : n17480;
  assign n17482 = pi10 ? n17481 : n32;
  assign n17483 = pi09 ? n32 : n17482;
  assign n17484 = pi08 ? n17476 : n17483;
  assign n17485 = pi07 ? n17462 : n17484;
  assign n17486 = pi17 ? n32 : n4261;
  assign n17487 = pi16 ? n32 : n17486;
  assign n17488 = pi15 ? n32 : n17487;
  assign n17489 = pi14 ? n17488 : n32;
  assign n17490 = pi13 ? n32 : n17489;
  assign n17491 = pi12 ? n32 : n17490;
  assign n17492 = pi11 ? n32 : n17491;
  assign n17493 = pi10 ? n32 : n17492;
  assign n17494 = pi15 ? n17278 : n17205;
  assign n17495 = pi14 ? n32 : n17494;
  assign n17496 = pi13 ? n32 : n17495;
  assign n17497 = pi12 ? n32 : n17496;
  assign n17498 = pi11 ? n17497 : n17480;
  assign n17499 = pi10 ? n17498 : n32;
  assign n17500 = pi09 ? n17493 : n17499;
  assign n17501 = pi15 ? n17363 : n17367;
  assign n17502 = pi14 ? n17501 : n32;
  assign n17503 = pi13 ? n17502 : n32;
  assign n17504 = pi12 ? n17503 : n32;
  assign n17505 = pi11 ? n17497 : n17504;
  assign n17506 = pi10 ? n17505 : n32;
  assign n17507 = pi09 ? n17493 : n17506;
  assign n17508 = pi08 ? n17500 : n17507;
  assign n17509 = pi21 ? n206 : n85;
  assign n17510 = pi20 ? n32 : n17509;
  assign n17511 = pi19 ? n32 : n17510;
  assign n17512 = pi18 ? n32 : n17511;
  assign n17513 = pi17 ? n32 : n17512;
  assign n17514 = pi16 ? n32 : n17513;
  assign n17515 = pi15 ? n17514 : n17348;
  assign n17516 = pi14 ? n32 : n17515;
  assign n17517 = pi13 ? n32 : n17516;
  assign n17518 = pi12 ? n32 : n17517;
  assign n17519 = pi14 ? n17368 : n32;
  assign n17520 = pi13 ? n17519 : n32;
  assign n17521 = pi12 ? n17520 : n32;
  assign n17522 = pi11 ? n17518 : n17521;
  assign n17523 = pi10 ? n17522 : n32;
  assign n17524 = pi09 ? n17493 : n17523;
  assign n17525 = pi07 ? n17508 : n17524;
  assign n17526 = pi06 ? n17485 : n17525;
  assign n17527 = pi05 ? n17420 : n17526;
  assign n17528 = pi19 ? n32 : n2092;
  assign n17529 = pi18 ? n32 : n17528;
  assign n17530 = pi17 ? n32 : n17529;
  assign n17531 = pi16 ? n32 : n17530;
  assign n17532 = pi15 ? n17531 : n17431;
  assign n17533 = pi14 ? n32 : n17532;
  assign n17534 = pi13 ? n32 : n17533;
  assign n17535 = pi12 ? n32 : n17534;
  assign n17536 = pi11 ? n17535 : n32;
  assign n17537 = pi10 ? n17536 : n32;
  assign n17538 = pi09 ? n32 : n17537;
  assign n17539 = pi15 ? n17531 : n17331;
  assign n17540 = pi14 ? n32 : n17539;
  assign n17541 = pi13 ? n32 : n17540;
  assign n17542 = pi12 ? n32 : n17541;
  assign n17543 = pi11 ? n17542 : n32;
  assign n17544 = pi10 ? n17543 : n32;
  assign n17545 = pi09 ? n32 : n17544;
  assign n17546 = pi08 ? n17538 : n17545;
  assign n17547 = pi08 ? n17545 : n32;
  assign n17548 = pi07 ? n17546 : n17547;
  assign n17549 = pi14 ? n17443 : n17357;
  assign n17550 = pi13 ? n32 : n17549;
  assign n17551 = pi12 ? n32 : n17550;
  assign n17552 = pi11 ? n17551 : n32;
  assign n17553 = pi10 ? n17552 : n32;
  assign n17554 = pi09 ? n32 : n17553;
  assign n17555 = pi14 ? n17443 : n32;
  assign n17556 = pi13 ? n32 : n17555;
  assign n17557 = pi12 ? n32 : n17556;
  assign n17558 = pi11 ? n17557 : n32;
  assign n17559 = pi10 ? n17558 : n32;
  assign n17560 = pi09 ? n32 : n17559;
  assign n17561 = pi07 ? n17554 : n17560;
  assign n17562 = pi06 ? n17548 : n17561;
  assign n17563 = pi08 ? n17560 : n32;
  assign n17564 = pi07 ? n17563 : n32;
  assign n17565 = pi06 ? n17564 : n32;
  assign n17566 = pi05 ? n17562 : n17565;
  assign n17567 = pi04 ? n17527 : n17566;
  assign n17568 = pi09 ? n17493 : n32;
  assign n17569 = pi07 ? n17568 : n32;
  assign n17570 = pi06 ? n32 : n17569;
  assign n17571 = pi05 ? n17570 : n32;
  assign n17572 = pi06 ? n17569 : n32;
  assign n17573 = pi05 ? n32 : n17572;
  assign n17574 = pi04 ? n17571 : n17573;
  assign n17575 = pi03 ? n17567 : n17574;
  assign n17576 = pi02 ? n17312 : n17575;
  assign n17577 = pi05 ? n32 : n17570;
  assign n17578 = pi15 ? n32 : n17435;
  assign n17579 = pi14 ? n17578 : n32;
  assign n17580 = pi13 ? n32 : n17579;
  assign n17581 = pi12 ? n32 : n17580;
  assign n17582 = pi11 ? n32 : n17581;
  assign n17583 = pi10 ? n32 : n17582;
  assign n17584 = pi09 ? n17583 : n32;
  assign n17585 = pi07 ? n17584 : n32;
  assign n17586 = pi07 ? n32 : n17568;
  assign n17587 = pi06 ? n17585 : n17586;
  assign n17588 = pi05 ? n32 : n17587;
  assign n17589 = pi04 ? n17577 : n17588;
  assign n17590 = pi14 ? n17466 : n32;
  assign n17591 = pi13 ? n32 : n17590;
  assign n17592 = pi12 ? n32 : n17591;
  assign n17593 = pi11 ? n32 : n17592;
  assign n17594 = pi10 ? n32 : n17593;
  assign n17595 = pi09 ? n17594 : n32;
  assign n17596 = pi14 ? n17421 : n32;
  assign n17597 = pi13 ? n32 : n17596;
  assign n17598 = pi12 ? n32 : n17597;
  assign n17599 = pi11 ? n32 : n17598;
  assign n17600 = pi10 ? n32 : n17599;
  assign n17601 = pi09 ? n17600 : n32;
  assign n17602 = pi07 ? n17595 : n17601;
  assign n17603 = pi06 ? n17602 : n32;
  assign n17604 = pi05 ? n17572 : n17603;
  assign n17605 = pi18 ? n32 : n833;
  assign n17606 = pi17 ? n32 : n17605;
  assign n17607 = pi16 ? n32 : n17606;
  assign n17608 = pi15 ? n32 : n17607;
  assign n17609 = pi14 ? n17608 : n32;
  assign n17610 = pi13 ? n32 : n17609;
  assign n17611 = pi12 ? n32 : n17610;
  assign n17612 = pi11 ? n32 : n17611;
  assign n17613 = pi10 ? n32 : n17612;
  assign n17614 = pi09 ? n17613 : n32;
  assign n17615 = pi19 ? n32 : n14375;
  assign n17616 = pi18 ? n32 : n17615;
  assign n17617 = pi17 ? n32 : n17616;
  assign n17618 = pi16 ? n32 : n17617;
  assign n17619 = pi15 ? n32 : n17618;
  assign n17620 = pi14 ? n17619 : n32;
  assign n17621 = pi13 ? n32 : n17620;
  assign n17622 = pi12 ? n32 : n17621;
  assign n17623 = pi11 ? n32 : n17622;
  assign n17624 = pi10 ? n32 : n17623;
  assign n17625 = pi09 ? n17624 : n32;
  assign n17626 = pi08 ? n17614 : n17625;
  assign n17627 = pi07 ? n17626 : n32;
  assign n17628 = pi06 ? n17568 : n17627;
  assign n17629 = pi05 ? n17628 : n32;
  assign n17630 = pi04 ? n17604 : n17629;
  assign n17631 = pi03 ? n17589 : n17630;
  assign n17632 = pi02 ? n17631 : n32;
  assign n17633 = pi01 ? n17576 : n17632;
  assign n17634 = pi00 ? n6528 : n17633;
  assign n17635 = pi18 ? n858 : n32;
  assign n17636 = pi17 ? n32 : n17635;
  assign n17637 = pi16 ? n32 : n17636;
  assign n17638 = pi15 ? n32 : n17637;
  assign n17639 = pi14 ? n17638 : n17637;
  assign n17640 = pi13 ? n32 : n17639;
  assign n17641 = pi20 ? n342 : n274;
  assign n17642 = pi19 ? n17641 : n32;
  assign n17643 = pi18 ? n32 : n17642;
  assign n17644 = pi20 ? n1076 : n5854;
  assign n17645 = pi19 ? n17644 : ~n9536;
  assign n17646 = pi18 ? n17645 : n32;
  assign n17647 = pi17 ? n17643 : n17646;
  assign n17648 = pi16 ? n32 : n17647;
  assign n17649 = pi20 ? n342 : n357;
  assign n17650 = pi19 ? n17649 : n32;
  assign n17651 = pi18 ? n32 : n17650;
  assign n17652 = pi21 ? n174 : ~n174;
  assign n17653 = pi20 ? n321 : n17652;
  assign n17654 = pi21 ? n32 : ~n100;
  assign n17655 = pi20 ? n32 : n17654;
  assign n17656 = pi19 ? n17653 : n17655;
  assign n17657 = pi18 ? n17656 : n32;
  assign n17658 = pi17 ? n17651 : n17657;
  assign n17659 = pi16 ? n32 : n17658;
  assign n17660 = pi15 ? n17648 : n17659;
  assign n17661 = pi18 ? n858 : n177;
  assign n17662 = pi17 ? n32 : n17661;
  assign n17663 = pi20 ? n1368 : n175;
  assign n17664 = pi19 ? n32 : n17663;
  assign n17665 = pi21 ? n309 : ~n259;
  assign n17666 = pi20 ? n1611 : n17665;
  assign n17667 = pi19 ? n17666 : n11145;
  assign n17668 = pi18 ? n17664 : n17667;
  assign n17669 = pi21 ? n309 : ~n174;
  assign n17670 = pi20 ? n333 : ~n17669;
  assign n17671 = pi21 ? n174 : n405;
  assign n17672 = pi21 ? n174 : ~n9326;
  assign n17673 = pi20 ? n17671 : n17672;
  assign n17674 = pi19 ? n17670 : ~n17673;
  assign n17675 = pi18 ? n17674 : ~n32;
  assign n17676 = pi17 ? n17668 : ~n17675;
  assign n17677 = pi16 ? n17662 : n17676;
  assign n17678 = pi20 ? n2385 : n17669;
  assign n17679 = pi19 ? n17678 : n17655;
  assign n17680 = pi18 ? n17679 : n32;
  assign n17681 = pi17 ? n17651 : n17680;
  assign n17682 = pi16 ? n32 : n17681;
  assign n17683 = pi15 ? n17677 : n17682;
  assign n17684 = pi14 ? n17660 : n17683;
  assign n17685 = pi20 ? n32 : n13387;
  assign n17686 = pi19 ? n507 : n17685;
  assign n17687 = pi18 ? n17686 : n32;
  assign n17688 = pi17 ? n13946 : n17687;
  assign n17689 = pi16 ? n32 : n17688;
  assign n17690 = pi15 ? n17689 : n32;
  assign n17691 = pi14 ? n17690 : n32;
  assign n17692 = pi13 ? n17684 : n17691;
  assign n17693 = pi12 ? n17640 : n17692;
  assign n17694 = pi11 ? n32 : n17693;
  assign n17695 = pi19 ? n32 : n14969;
  assign n17696 = pi18 ? n17695 : n32;
  assign n17697 = pi17 ? n32 : n17696;
  assign n17698 = pi16 ? n32 : n17697;
  assign n17699 = pi19 ? n32 : n14786;
  assign n17700 = pi18 ? n17699 : n32;
  assign n17701 = pi17 ? n32 : n17700;
  assign n17702 = pi16 ? n32 : n17701;
  assign n17703 = pi15 ? n17698 : n17702;
  assign n17704 = pi14 ? n32 : n17703;
  assign n17705 = pi18 ? n1819 : n32;
  assign n17706 = pi17 ? n32 : n17705;
  assign n17707 = pi16 ? n32 : n17706;
  assign n17708 = pi15 ? n17707 : n32;
  assign n17709 = pi14 ? n17698 : n17708;
  assign n17710 = pi13 ? n17704 : n17709;
  assign n17711 = pi12 ? n32 : n17710;
  assign n17712 = pi21 ? n32 : ~n242;
  assign n17713 = pi20 ? n32 : n17712;
  assign n17714 = pi19 ? n32 : n17713;
  assign n17715 = pi18 ? n17714 : n32;
  assign n17716 = pi17 ? n32 : n17715;
  assign n17717 = pi16 ? n32 : n17716;
  assign n17718 = pi20 ? n32 : n7467;
  assign n17719 = pi19 ? n32 : n17718;
  assign n17720 = pi18 ? n17719 : n32;
  assign n17721 = pi17 ? n32 : n17720;
  assign n17722 = pi16 ? n32 : n17721;
  assign n17723 = pi15 ? n17717 : n17722;
  assign n17724 = pi21 ? n32 : n15659;
  assign n17725 = pi20 ? n32 : n17724;
  assign n17726 = pi19 ? n32 : n17725;
  assign n17727 = pi18 ? n17726 : n32;
  assign n17728 = pi17 ? n32 : n17727;
  assign n17729 = pi16 ? n32 : n17728;
  assign n17730 = pi14 ? n17723 : n17729;
  assign n17731 = pi14 ? n17729 : n17717;
  assign n17732 = pi13 ? n17730 : n17731;
  assign n17733 = pi19 ? n32 : n5350;
  assign n17734 = pi18 ? n17733 : n32;
  assign n17735 = pi17 ? n32 : n17734;
  assign n17736 = pi16 ? n32 : n17735;
  assign n17737 = pi20 ? n175 : n1817;
  assign n17738 = pi19 ? n32 : n17737;
  assign n17739 = pi18 ? n17738 : n32;
  assign n17740 = pi17 ? n32 : n17739;
  assign n17741 = pi16 ? n32 : n17740;
  assign n17742 = pi15 ? n17736 : n17741;
  assign n17743 = pi18 ? n16432 : n32;
  assign n17744 = pi18 ? n17283 : n32;
  assign n17745 = pi17 ? n17743 : n17744;
  assign n17746 = pi16 ? n32 : n17745;
  assign n17747 = pi15 ? n17736 : n17746;
  assign n17748 = pi14 ? n17742 : n17747;
  assign n17749 = pi20 ? n206 : ~n220;
  assign n17750 = pi19 ? n17749 : ~n32;
  assign n17751 = pi18 ? n496 : ~n17750;
  assign n17752 = pi20 ? n246 : ~n1839;
  assign n17753 = pi19 ? n221 : n17752;
  assign n17754 = pi18 ? n17753 : n32;
  assign n17755 = pi17 ? n17751 : n17754;
  assign n17756 = pi16 ? n32 : n17755;
  assign n17757 = pi20 ? n266 : n206;
  assign n17758 = pi19 ? n32 : ~n17757;
  assign n17759 = pi18 ? n17758 : ~n5372;
  assign n17760 = pi20 ? n266 : n7388;
  assign n17761 = pi19 ? n221 : n17760;
  assign n17762 = pi18 ? n17761 : n32;
  assign n17763 = pi17 ? n17759 : n17762;
  assign n17764 = pi16 ? n32 : n17763;
  assign n17765 = pi15 ? n17756 : n17764;
  assign n17766 = pi20 ? n246 : ~n207;
  assign n17767 = pi19 ? n32 : n17766;
  assign n17768 = pi18 ? n17767 : n32;
  assign n17769 = pi20 ? n266 : n1331;
  assign n17770 = pi19 ? n267 : n17769;
  assign n17771 = pi18 ? n17770 : n32;
  assign n17772 = pi17 ? n17768 : n17771;
  assign n17773 = pi16 ? n32 : n17772;
  assign n17774 = pi17 ? n17768 : n269;
  assign n17775 = pi16 ? n32 : n17774;
  assign n17776 = pi15 ? n17773 : n17775;
  assign n17777 = pi14 ? n17765 : n17776;
  assign n17778 = pi13 ? n17748 : n17777;
  assign n17779 = pi12 ? n17732 : n17778;
  assign n17780 = pi11 ? n17711 : n17779;
  assign n17781 = pi10 ? n17694 : n17780;
  assign n17782 = pi09 ? n32 : n17781;
  assign n17783 = pi14 ? n32 : n17638;
  assign n17784 = pi13 ? n32 : n17783;
  assign n17785 = pi20 ? n339 : ~n13387;
  assign n17786 = pi19 ? n17644 : ~n17785;
  assign n17787 = pi18 ? n17786 : n32;
  assign n17788 = pi17 ? n17643 : n17787;
  assign n17789 = pi16 ? n32 : n17788;
  assign n17790 = pi19 ? n17653 : n4518;
  assign n17791 = pi18 ? n17790 : n32;
  assign n17792 = pi17 ? n17651 : n17791;
  assign n17793 = pi16 ? n32 : n17792;
  assign n17794 = pi15 ? n17789 : n17793;
  assign n17795 = pi21 ? n174 : ~n11567;
  assign n17796 = pi20 ? n17671 : n17795;
  assign n17797 = pi19 ? n17670 : ~n17796;
  assign n17798 = pi18 ? n17797 : ~n32;
  assign n17799 = pi17 ? n17668 : ~n17798;
  assign n17800 = pi16 ? n17662 : n17799;
  assign n17801 = pi19 ? n17678 : n4518;
  assign n17802 = pi18 ? n17801 : n32;
  assign n17803 = pi17 ? n17651 : n17802;
  assign n17804 = pi16 ? n32 : n17803;
  assign n17805 = pi15 ? n17800 : n17804;
  assign n17806 = pi14 ? n17794 : n17805;
  assign n17807 = pi18 ? n507 : n32;
  assign n17808 = pi17 ? n13946 : n17807;
  assign n17809 = pi16 ? n32 : n17808;
  assign n17810 = pi19 ? n32 : n2078;
  assign n17811 = pi18 ? n17810 : n32;
  assign n17812 = pi17 ? n32 : n17811;
  assign n17813 = pi16 ? n32 : n17812;
  assign n17814 = pi15 ? n17809 : n17813;
  assign n17815 = pi14 ? n17814 : n32;
  assign n17816 = pi13 ? n17806 : n17815;
  assign n17817 = pi12 ? n17784 : n17816;
  assign n17818 = pi11 ? n32 : n17817;
  assign n17819 = pi19 ? n32 : n14963;
  assign n17820 = pi18 ? n17819 : n32;
  assign n17821 = pi17 ? n32 : n17820;
  assign n17822 = pi16 ? n32 : n17821;
  assign n17823 = pi18 ? n4519 : n32;
  assign n17824 = pi17 ? n32 : n17823;
  assign n17825 = pi16 ? n32 : n17824;
  assign n17826 = pi15 ? n17822 : n17825;
  assign n17827 = pi14 ? n17638 : n17826;
  assign n17828 = pi21 ? n32 : ~n10445;
  assign n17829 = pi20 ? n32 : n17828;
  assign n17830 = pi19 ? n32 : n17829;
  assign n17831 = pi18 ? n17830 : n32;
  assign n17832 = pi17 ? n32 : n17831;
  assign n17833 = pi16 ? n32 : n17832;
  assign n17834 = pi19 ? n32 : n644;
  assign n17835 = pi18 ? n17834 : n32;
  assign n17836 = pi17 ? n32 : n17835;
  assign n17837 = pi16 ? n32 : n17836;
  assign n17838 = pi15 ? n17833 : n17837;
  assign n17839 = pi14 ? n17822 : n17838;
  assign n17840 = pi13 ? n17827 : n17839;
  assign n17841 = pi12 ? n32 : n17840;
  assign n17842 = pi20 ? n32 : n7442;
  assign n17843 = pi19 ? n32 : n17842;
  assign n17844 = pi18 ? n17843 : n32;
  assign n17845 = pi17 ? n32 : n17844;
  assign n17846 = pi16 ? n32 : n17845;
  assign n17847 = pi15 ? n17702 : n17846;
  assign n17848 = pi19 ? n32 : n6398;
  assign n17849 = pi18 ? n17848 : n32;
  assign n17850 = pi17 ? n32 : n17849;
  assign n17851 = pi16 ? n32 : n17850;
  assign n17852 = pi15 ? n17851 : n32;
  assign n17853 = pi14 ? n17847 : n17852;
  assign n17854 = pi18 ? n17528 : n32;
  assign n17855 = pi17 ? n32 : n17854;
  assign n17856 = pi16 ? n32 : n17855;
  assign n17857 = pi14 ? n17856 : n17717;
  assign n17858 = pi13 ? n17853 : n17857;
  assign n17859 = pi20 ? n32 : n11086;
  assign n17860 = pi19 ? n32 : n17859;
  assign n17861 = pi18 ? n17860 : n32;
  assign n17862 = pi17 ? n17768 : n17861;
  assign n17863 = pi16 ? n32 : n17862;
  assign n17864 = pi15 ? n17773 : n17863;
  assign n17865 = pi14 ? n17765 : n17864;
  assign n17866 = pi13 ? n17748 : n17865;
  assign n17867 = pi12 ? n17858 : n17866;
  assign n17868 = pi11 ? n17841 : n17867;
  assign n17869 = pi10 ? n17818 : n17868;
  assign n17870 = pi09 ? n32 : n17869;
  assign n17871 = pi08 ? n17782 : n17870;
  assign n17872 = pi07 ? n32 : n17871;
  assign n17873 = pi06 ? n32 : n17872;
  assign n17874 = pi18 ? n1575 : n32;
  assign n17875 = pi17 ? n32 : n17874;
  assign n17876 = pi16 ? n32 : n17875;
  assign n17877 = pi15 ? n17876 : n32;
  assign n17878 = pi14 ? n32 : n17877;
  assign n17879 = pi19 ? n857 : n594;
  assign n17880 = pi18 ? n17879 : n32;
  assign n17881 = pi17 ? n32 : n17880;
  assign n17882 = pi16 ? n32 : n17881;
  assign n17883 = pi18 ? n936 : n32;
  assign n17884 = pi17 ? n32 : n17883;
  assign n17885 = pi16 ? n32 : n17884;
  assign n17886 = pi15 ? n17882 : n17885;
  assign n17887 = pi14 ? n17886 : n32;
  assign n17888 = pi13 ? n17878 : n17887;
  assign n17889 = pi18 ? n863 : ~n1676;
  assign n17890 = pi17 ? n32 : n17889;
  assign n17891 = pi16 ? n32 : n17890;
  assign n17892 = pi18 ? n32 : ~n1676;
  assign n17893 = pi17 ? n32 : n17892;
  assign n17894 = pi16 ? n32 : n17893;
  assign n17895 = pi15 ? n17891 : n17894;
  assign n17896 = pi14 ? n17895 : n17894;
  assign n17897 = pi14 ? n17876 : n32;
  assign n17898 = pi13 ? n17896 : n17897;
  assign n17899 = pi12 ? n17888 : n17898;
  assign n17900 = pi11 ? n32 : n17899;
  assign n17901 = pi18 ? n863 : n32;
  assign n17902 = pi17 ? n32 : n17901;
  assign n17903 = pi16 ? n32 : n17902;
  assign n17904 = pi15 ? n17903 : n17876;
  assign n17905 = pi14 ? n32 : n17904;
  assign n17906 = pi13 ? n32 : n17905;
  assign n17907 = pi19 ? n32 : n17685;
  assign n17908 = pi18 ? n17907 : n32;
  assign n17909 = pi17 ? n32 : n17908;
  assign n17910 = pi16 ? n32 : n17909;
  assign n17911 = pi15 ? n32 : n17910;
  assign n17912 = pi19 ? n32 : n17655;
  assign n17913 = pi18 ? n17912 : n32;
  assign n17914 = pi17 ? n32 : n17913;
  assign n17915 = pi16 ? n32 : n17914;
  assign n17916 = pi15 ? n17910 : n17915;
  assign n17917 = pi14 ? n17911 : n17916;
  assign n17918 = pi20 ? n32 : ~n428;
  assign n17919 = pi19 ? n32 : n17918;
  assign n17920 = pi18 ? n17919 : n32;
  assign n17921 = pi17 ? n32 : n17920;
  assign n17922 = pi16 ? n32 : n17921;
  assign n17923 = pi15 ? n17825 : n17922;
  assign n17924 = pi14 ? n17916 : n17923;
  assign n17925 = pi13 ? n17917 : n17924;
  assign n17926 = pi12 ? n17906 : n17925;
  assign n17927 = pi19 ? n32 : n14589;
  assign n17928 = pi18 ? n17927 : n32;
  assign n17929 = pi17 ? n32 : n17928;
  assign n17930 = pi16 ? n32 : n17929;
  assign n17931 = pi15 ? n17930 : n17825;
  assign n17932 = pi15 ? n17698 : n17851;
  assign n17933 = pi14 ? n17931 : n17932;
  assign n17934 = pi18 ? n312 : n32;
  assign n17935 = pi17 ? n32 : n17934;
  assign n17936 = pi16 ? n32 : n17935;
  assign n17937 = pi16 ? n32 : n264;
  assign n17938 = pi15 ? n17936 : n17937;
  assign n17939 = pi14 ? n17851 : n17938;
  assign n17940 = pi13 ? n17933 : n17939;
  assign n17941 = pi20 ? n32 : ~n1319;
  assign n17942 = pi19 ? n32 : n17941;
  assign n17943 = pi18 ? n17942 : n32;
  assign n17944 = pi17 ? n32 : n17943;
  assign n17945 = pi16 ? n32 : n17944;
  assign n17946 = pi19 ? n32 : n13632;
  assign n17947 = pi18 ? n17946 : n32;
  assign n17948 = pi17 ? n32 : n17947;
  assign n17949 = pi16 ? n32 : n17948;
  assign n17950 = pi15 ? n17945 : n17949;
  assign n17951 = pi18 ? n6071 : n32;
  assign n17952 = pi17 ? n17951 : n17947;
  assign n17953 = pi16 ? n32 : n17952;
  assign n17954 = pi20 ? n207 : n7467;
  assign n17955 = pi19 ? n322 : n17954;
  assign n17956 = pi18 ? n17955 : n32;
  assign n17957 = pi17 ? n17951 : n17956;
  assign n17958 = pi16 ? n32 : n17957;
  assign n17959 = pi15 ? n17953 : n17958;
  assign n17960 = pi14 ? n17950 : n17959;
  assign n17961 = pi20 ? n2385 : n1331;
  assign n17962 = pi19 ? n32 : n17961;
  assign n17963 = pi18 ? n17962 : n32;
  assign n17964 = pi20 ? n321 : ~n1685;
  assign n17965 = pi19 ? n322 : ~n17964;
  assign n17966 = pi18 ? n17965 : n32;
  assign n17967 = pi17 ? n17963 : n17966;
  assign n17968 = pi16 ? n32 : n17967;
  assign n17969 = pi19 ? n208 : ~n17964;
  assign n17970 = pi18 ? n17969 : n32;
  assign n17971 = pi17 ? n32 : n17970;
  assign n17972 = pi16 ? n32 : n17971;
  assign n17973 = pi15 ? n17968 : n17972;
  assign n17974 = pi20 ? n174 : n32;
  assign n17975 = pi19 ? n32 : n17974;
  assign n17976 = pi18 ? n17975 : n32;
  assign n17977 = pi20 ? n915 : n7388;
  assign n17978 = pi19 ? n786 : n17977;
  assign n17979 = pi18 ? n17978 : n32;
  assign n17980 = pi17 ? n17976 : n17979;
  assign n17981 = pi16 ? n32 : n17980;
  assign n17982 = pi20 ? n32 : n7388;
  assign n17983 = pi19 ? n1818 : n17982;
  assign n17984 = pi18 ? n17983 : n32;
  assign n17985 = pi17 ? n32 : n17984;
  assign n17986 = pi16 ? n32 : n17985;
  assign n17987 = pi15 ? n17981 : n17986;
  assign n17988 = pi14 ? n17973 : n17987;
  assign n17989 = pi13 ? n17960 : n17988;
  assign n17990 = pi12 ? n17940 : n17989;
  assign n17991 = pi11 ? n17926 : n17990;
  assign n17992 = pi10 ? n17900 : n17991;
  assign n17993 = pi09 ? n32 : n17992;
  assign n17994 = pi19 ? n5635 : n32;
  assign n17995 = pi18 ? n32 : n17994;
  assign n17996 = pi17 ? n32 : n17995;
  assign n17997 = pi16 ? n32 : n17996;
  assign n17998 = pi14 ? n32 : n17997;
  assign n17999 = pi18 ? n8106 : n32;
  assign n18000 = pi17 ? n32 : n17999;
  assign n18001 = pi16 ? n32 : n18000;
  assign n18002 = pi15 ? n18001 : n32;
  assign n18003 = pi14 ? n18002 : n32;
  assign n18004 = pi13 ? n17998 : n18003;
  assign n18005 = pi15 ? n17903 : n32;
  assign n18006 = pi18 ? n32 : ~n618;
  assign n18007 = pi17 ? n32 : n18006;
  assign n18008 = pi16 ? n32 : n18007;
  assign n18009 = pi14 ? n18005 : n18008;
  assign n18010 = pi14 ? n18008 : n32;
  assign n18011 = pi13 ? n18009 : n18010;
  assign n18012 = pi12 ? n18004 : n18011;
  assign n18013 = pi11 ? n32 : n18012;
  assign n18014 = pi14 ? n32 : n17895;
  assign n18015 = pi13 ? n32 : n18014;
  assign n18016 = pi15 ? n32 : n17903;
  assign n18017 = pi18 ? n940 : n32;
  assign n18018 = pi17 ? n32 : n18017;
  assign n18019 = pi16 ? n32 : n18018;
  assign n18020 = pi15 ? n17903 : n18019;
  assign n18021 = pi14 ? n18016 : n18020;
  assign n18022 = pi20 ? n32 : ~n101;
  assign n18023 = pi19 ? n32 : n18022;
  assign n18024 = pi18 ? n18023 : n32;
  assign n18025 = pi17 ? n32 : n18024;
  assign n18026 = pi16 ? n32 : n18025;
  assign n18027 = pi15 ? n17915 : n18026;
  assign n18028 = pi14 ? n18020 : n18027;
  assign n18029 = pi13 ? n18021 : n18028;
  assign n18030 = pi12 ? n18015 : n18029;
  assign n18031 = pi20 ? n32 : n13084;
  assign n18032 = pi19 ? n32 : n18031;
  assign n18033 = pi18 ? n18032 : n32;
  assign n18034 = pi17 ? n32 : n18033;
  assign n18035 = pi16 ? n32 : n18034;
  assign n18036 = pi15 ? n18035 : n17825;
  assign n18037 = pi14 ? n18036 : n17932;
  assign n18038 = pi13 ? n18037 : n17939;
  assign n18039 = pi17 ? n32 : n17744;
  assign n18040 = pi16 ? n32 : n18039;
  assign n18041 = pi20 ? n321 : ~n518;
  assign n18042 = pi19 ? n594 : n18041;
  assign n18043 = pi18 ? n18042 : n32;
  assign n18044 = pi17 ? n32 : n18043;
  assign n18045 = pi16 ? n32 : n18044;
  assign n18046 = pi15 ? n18040 : n18045;
  assign n18047 = pi17 ? n32 : n17956;
  assign n18048 = pi16 ? n32 : n18047;
  assign n18049 = pi15 ? n17949 : n18048;
  assign n18050 = pi14 ? n18046 : n18049;
  assign n18051 = pi17 ? n32 : n17966;
  assign n18052 = pi16 ? n32 : n18051;
  assign n18053 = pi15 ? n18052 : n17972;
  assign n18054 = pi19 ? n4126 : n17977;
  assign n18055 = pi18 ? n18054 : n32;
  assign n18056 = pi17 ? n32 : n18055;
  assign n18057 = pi16 ? n32 : n18056;
  assign n18058 = pi19 ? n32 : n17982;
  assign n18059 = pi18 ? n18058 : n32;
  assign n18060 = pi17 ? n32 : n18059;
  assign n18061 = pi16 ? n32 : n18060;
  assign n18062 = pi15 ? n18057 : n18061;
  assign n18063 = pi14 ? n18053 : n18062;
  assign n18064 = pi13 ? n18050 : n18063;
  assign n18065 = pi12 ? n18038 : n18064;
  assign n18066 = pi11 ? n18030 : n18065;
  assign n18067 = pi10 ? n18013 : n18066;
  assign n18068 = pi09 ? n32 : n18067;
  assign n18069 = pi08 ? n17993 : n18068;
  assign n18070 = pi20 ? n32 : ~n820;
  assign n18071 = pi19 ? n18070 : n32;
  assign n18072 = pi18 ? n32 : n18071;
  assign n18073 = pi21 ? n309 : ~n313;
  assign n18074 = pi20 ? n246 : ~n18073;
  assign n18075 = pi19 ? n18074 : ~n617;
  assign n18076 = pi19 ? n5626 : n32;
  assign n18077 = pi18 ? n18075 : n18076;
  assign n18078 = pi17 ? n18072 : n18077;
  assign n18079 = pi16 ? n32 : n18078;
  assign n18080 = pi15 ? n18079 : n32;
  assign n18081 = pi14 ? n32 : n18080;
  assign n18082 = pi18 ? n32 : n4492;
  assign n18083 = pi17 ? n32 : n18082;
  assign n18084 = pi20 ? n274 : n246;
  assign n18085 = pi19 ? n32 : n18084;
  assign n18086 = pi19 ? n247 : n428;
  assign n18087 = pi18 ? n18085 : n18086;
  assign n18088 = pi19 ? n8044 : n175;
  assign n18089 = pi18 ? n18088 : n32;
  assign n18090 = pi17 ? n18087 : n18089;
  assign n18091 = pi16 ? n18083 : n18090;
  assign n18092 = pi15 ? n32 : n18091;
  assign n18093 = pi14 ? n32 : n18092;
  assign n18094 = pi13 ? n18081 : n18093;
  assign n18095 = pi20 ? n1331 : ~n785;
  assign n18096 = pi19 ? n220 : ~n18095;
  assign n18097 = pi18 ? n863 : ~n18096;
  assign n18098 = pi17 ? n32 : n18097;
  assign n18099 = pi20 ? n11107 : n246;
  assign n18100 = pi19 ? n18099 : n12801;
  assign n18101 = pi18 ? n18100 : ~n32;
  assign n18102 = pi19 ? n32 : n246;
  assign n18103 = pi18 ? n18102 : n237;
  assign n18104 = pi17 ? n18101 : ~n18103;
  assign n18105 = pi16 ? n18098 : n18104;
  assign n18106 = pi20 ? n785 : ~n11107;
  assign n18107 = pi19 ? n17961 : ~n18106;
  assign n18108 = pi18 ? n863 : n18107;
  assign n18109 = pi17 ? n32 : n18108;
  assign n18110 = pi20 ? n246 : n1611;
  assign n18111 = pi20 ? n342 : n1331;
  assign n18112 = pi19 ? n18110 : n18111;
  assign n18113 = pi20 ? n1331 : n342;
  assign n18114 = pi19 ? n18113 : n1331;
  assign n18115 = pi18 ? n18112 : n18114;
  assign n18116 = pi20 ? n2385 : n32;
  assign n18117 = pi19 ? n18116 : n246;
  assign n18118 = pi18 ? n18117 : ~n237;
  assign n18119 = pi17 ? n18115 : n18118;
  assign n18120 = pi16 ? n18109 : n18119;
  assign n18121 = pi15 ? n18105 : n18120;
  assign n18122 = pi20 ? n749 : n1331;
  assign n18123 = pi19 ? n18122 : ~n18106;
  assign n18124 = pi18 ? n863 : n18123;
  assign n18125 = pi17 ? n32 : n18124;
  assign n18126 = pi20 ? n1611 : n2385;
  assign n18127 = pi19 ? n18110 : n18126;
  assign n18128 = pi20 ? n2385 : n1611;
  assign n18129 = pi21 ? n405 : n174;
  assign n18130 = pi20 ? n18129 : ~n17652;
  assign n18131 = pi19 ? n18128 : n18130;
  assign n18132 = pi18 ? n18127 : n18131;
  assign n18133 = pi20 ? n5854 : ~n17669;
  assign n18134 = pi19 ? n18133 : ~n1324;
  assign n18135 = pi18 ? n18134 : n237;
  assign n18136 = pi17 ? n18132 : ~n18135;
  assign n18137 = pi16 ? n18125 : n18136;
  assign n18138 = pi15 ? n18137 : n32;
  assign n18139 = pi14 ? n18121 : n18138;
  assign n18140 = pi18 ? n32 : n18076;
  assign n18141 = pi17 ? n32 : n18140;
  assign n18142 = pi16 ? n32 : n18141;
  assign n18143 = pi15 ? n32 : n18008;
  assign n18144 = pi14 ? n18142 : n18143;
  assign n18145 = pi13 ? n18139 : n18144;
  assign n18146 = pi12 ? n18094 : n18145;
  assign n18147 = pi11 ? n32 : n18146;
  assign n18148 = pi15 ? n17997 : n32;
  assign n18149 = pi14 ? n18008 : n18148;
  assign n18150 = pi14 ? n32 : n17894;
  assign n18151 = pi13 ? n18149 : n18150;
  assign n18152 = pi15 ? n17903 : n17891;
  assign n18153 = pi14 ? n18152 : n18020;
  assign n18154 = pi18 ? n751 : n32;
  assign n18155 = pi17 ? n32 : n18154;
  assign n18156 = pi16 ? n32 : n18155;
  assign n18157 = pi15 ? n17903 : n18156;
  assign n18158 = pi21 ? n32 : n14158;
  assign n18159 = pi20 ? n32 : n18158;
  assign n18160 = pi19 ? n32 : n18159;
  assign n18161 = pi18 ? n18160 : n32;
  assign n18162 = pi17 ? n32 : n18161;
  assign n18163 = pi16 ? n32 : n18162;
  assign n18164 = pi15 ? n18163 : n17910;
  assign n18165 = pi14 ? n18157 : n18164;
  assign n18166 = pi13 ? n18153 : n18165;
  assign n18167 = pi12 ? n18151 : n18166;
  assign n18168 = pi15 ? n17825 : n17702;
  assign n18169 = pi14 ? n18163 : n18168;
  assign n18170 = pi15 ? n17702 : n17698;
  assign n18171 = pi14 ? n18170 : n17846;
  assign n18172 = pi13 ? n18169 : n18171;
  assign n18173 = pi21 ? n259 : ~n309;
  assign n18174 = pi20 ? n18173 : n342;
  assign n18175 = pi19 ? n32 : ~n18174;
  assign n18176 = pi18 ? n18175 : n32;
  assign n18177 = pi17 ? n32 : n18176;
  assign n18178 = pi16 ? n32 : n18177;
  assign n18179 = pi18 ? n15570 : n32;
  assign n18180 = pi17 ? n32 : n18179;
  assign n18181 = pi16 ? n32 : n18180;
  assign n18182 = pi15 ? n18178 : n18181;
  assign n18183 = pi19 ? n32 : n5356;
  assign n18184 = pi18 ? n18183 : n32;
  assign n18185 = pi17 ? n32 : n18184;
  assign n18186 = pi16 ? n32 : n18185;
  assign n18187 = pi19 ? n322 : n16002;
  assign n18188 = pi18 ? n18187 : n32;
  assign n18189 = pi17 ? n32 : n18188;
  assign n18190 = pi16 ? n32 : n18189;
  assign n18191 = pi15 ? n18186 : n18190;
  assign n18192 = pi14 ? n18182 : n18191;
  assign n18193 = pi19 ? n322 : ~n9028;
  assign n18194 = pi18 ? n18193 : n32;
  assign n18195 = pi17 ? n32 : n18194;
  assign n18196 = pi16 ? n32 : n18195;
  assign n18197 = pi21 ? n1392 : n206;
  assign n18198 = pi20 ? n32 : n18197;
  assign n18199 = pi19 ? n32 : n18198;
  assign n18200 = pi20 ? n266 : n10644;
  assign n18201 = pi19 ? n18200 : n5004;
  assign n18202 = pi18 ? n18199 : ~n18201;
  assign n18203 = pi17 ? n32 : n18202;
  assign n18204 = pi20 ? n518 : n1319;
  assign n18205 = pi19 ? n32 : n18204;
  assign n18206 = pi18 ? n18205 : ~n32;
  assign n18207 = pi17 ? n1028 : ~n18206;
  assign n18208 = pi16 ? n18203 : n18207;
  assign n18209 = pi15 ? n18196 : n18208;
  assign n18210 = pi19 ? n208 : ~n507;
  assign n18211 = pi20 ? n220 : ~n321;
  assign n18212 = pi19 ? n15405 : n18211;
  assign n18213 = pi18 ? n18210 : n18212;
  assign n18214 = pi19 ? n236 : ~n17964;
  assign n18215 = pi18 ? n18214 : n32;
  assign n18216 = pi17 ? n18213 : n18215;
  assign n18217 = pi16 ? n17902 : n18216;
  assign n18218 = pi20 ? n32 : n16309;
  assign n18219 = pi19 ? n32 : n18218;
  assign n18220 = pi18 ? n18219 : n32;
  assign n18221 = pi17 ? n32 : n18220;
  assign n18222 = pi16 ? n32 : n18221;
  assign n18223 = pi15 ? n18217 : n18222;
  assign n18224 = pi14 ? n18209 : n18223;
  assign n18225 = pi13 ? n18192 : n18224;
  assign n18226 = pi12 ? n18172 : n18225;
  assign n18227 = pi11 ? n18167 : n18226;
  assign n18228 = pi10 ? n18147 : n18227;
  assign n18229 = pi09 ? n32 : n18228;
  assign n18230 = pi18 ? n18075 : n32;
  assign n18231 = pi17 ? n18072 : n18230;
  assign n18232 = pi16 ? n32 : n18231;
  assign n18233 = pi15 ? n18232 : n32;
  assign n18234 = pi14 ? n32 : n18233;
  assign n18235 = pi18 ? n18088 : n359;
  assign n18236 = pi17 ? n18087 : n18235;
  assign n18237 = pi16 ? n18083 : n18236;
  assign n18238 = pi15 ? n32 : n18237;
  assign n18239 = pi14 ? n32 : n18238;
  assign n18240 = pi13 ? n18234 : n18239;
  assign n18241 = pi20 ? n9194 : n18129;
  assign n18242 = pi19 ? n6303 : n18241;
  assign n18243 = pi18 ? n2387 : ~n18242;
  assign n18244 = pi17 ? n32 : n18243;
  assign n18245 = pi21 ? n173 : ~n405;
  assign n18246 = pi20 ? n18173 : n18245;
  assign n18247 = pi19 ? n18246 : ~n247;
  assign n18248 = pi18 ? n18247 : ~n32;
  assign n18249 = pi19 ? n32 : n3523;
  assign n18250 = pi18 ? n18249 : n1942;
  assign n18251 = pi17 ? n18248 : ~n18250;
  assign n18252 = pi16 ? n18244 : n18251;
  assign n18253 = pi21 ? n313 : ~n309;
  assign n18254 = pi20 ? n1091 : n18253;
  assign n18255 = pi21 ? n405 : ~n173;
  assign n18256 = pi21 ? n206 : ~n313;
  assign n18257 = pi20 ? n18255 : ~n18256;
  assign n18258 = pi19 ? n18254 : n18257;
  assign n18259 = pi18 ? n863 : ~n18258;
  assign n18260 = pi17 ? n32 : n18259;
  assign n18261 = pi21 ? n173 : n206;
  assign n18262 = pi20 ? n3695 : n18261;
  assign n18263 = pi20 ? n260 : n314;
  assign n18264 = pi19 ? n18262 : ~n18263;
  assign n18265 = pi20 ? n314 : ~n2385;
  assign n18266 = pi20 ? n18253 : ~n3843;
  assign n18267 = pi19 ? n18265 : n18266;
  assign n18268 = pi18 ? n18264 : ~n18267;
  assign n18269 = pi19 ? n18116 : n12884;
  assign n18270 = pi18 ? n18269 : ~n1942;
  assign n18271 = pi17 ? n18268 : n18270;
  assign n18272 = pi16 ? n18260 : n18271;
  assign n18273 = pi15 ? n18252 : n18272;
  assign n18274 = pi20 ? n439 : n18253;
  assign n18275 = pi19 ? n18274 : n18257;
  assign n18276 = pi18 ? n2387 : ~n18275;
  assign n18277 = pi17 ? n32 : n18276;
  assign n18278 = pi20 ? n5854 : n13171;
  assign n18279 = pi19 ? n18262 : ~n18278;
  assign n18280 = pi20 ? n13171 : ~n18261;
  assign n18281 = pi21 ? n313 : ~n313;
  assign n18282 = pi21 ? n174 : ~n313;
  assign n18283 = pi20 ? n18281 : n18282;
  assign n18284 = pi19 ? n18280 : n18283;
  assign n18285 = pi18 ? n18279 : ~n18284;
  assign n18286 = pi19 ? n18133 : ~n17669;
  assign n18287 = pi18 ? n18286 : n1942;
  assign n18288 = pi17 ? n18285 : ~n18287;
  assign n18289 = pi16 ? n18277 : n18288;
  assign n18290 = pi15 ? n18289 : n32;
  assign n18291 = pi14 ? n18273 : n18290;
  assign n18292 = pi18 ? n32 : n359;
  assign n18293 = pi17 ? n32 : n18292;
  assign n18294 = pi16 ? n32 : n18293;
  assign n18295 = pi18 ? n32 : ~n3350;
  assign n18296 = pi17 ? n32 : n18295;
  assign n18297 = pi16 ? n32 : n18296;
  assign n18298 = pi15 ? n32 : n18297;
  assign n18299 = pi14 ? n18294 : n18298;
  assign n18300 = pi13 ? n18291 : n18299;
  assign n18301 = pi12 ? n18240 : n18300;
  assign n18302 = pi11 ? n32 : n18301;
  assign n18303 = pi15 ? n18297 : n18142;
  assign n18304 = pi15 ? n18142 : n32;
  assign n18305 = pi14 ? n18303 : n18304;
  assign n18306 = pi13 ? n18305 : n17998;
  assign n18307 = pi18 ? n940 : ~n1676;
  assign n18308 = pi17 ? n32 : n18307;
  assign n18309 = pi16 ? n32 : n18308;
  assign n18310 = pi15 ? n17891 : n18309;
  assign n18311 = pi14 ? n17891 : n18310;
  assign n18312 = pi18 ? n751 : ~n1676;
  assign n18313 = pi17 ? n32 : n18312;
  assign n18314 = pi16 ? n32 : n18313;
  assign n18315 = pi15 ? n17891 : n18314;
  assign n18316 = pi18 ? n1592 : n32;
  assign n18317 = pi17 ? n32 : n18316;
  assign n18318 = pi16 ? n32 : n18317;
  assign n18319 = pi15 ? n18318 : n17903;
  assign n18320 = pi14 ? n18315 : n18319;
  assign n18321 = pi13 ? n18311 : n18320;
  assign n18322 = pi12 ? n18306 : n18321;
  assign n18323 = pi15 ? n18318 : n18163;
  assign n18324 = pi18 ? n4380 : n32;
  assign n18325 = pi17 ? n32 : n18324;
  assign n18326 = pi16 ? n32 : n18325;
  assign n18327 = pi15 ? n17825 : n18326;
  assign n18328 = pi14 ? n18323 : n18327;
  assign n18329 = pi13 ? n18328 : n18171;
  assign n18330 = pi20 ? n32 : n17671;
  assign n18331 = pi19 ? n32 : n18330;
  assign n18332 = pi20 ? n18173 : n339;
  assign n18333 = pi20 ? n314 : ~n18129;
  assign n18334 = pi19 ? n18332 : n18333;
  assign n18335 = pi18 ? n18331 : ~n18334;
  assign n18336 = pi17 ? n32 : n18335;
  assign n18337 = pi21 ? n174 : n313;
  assign n18338 = pi20 ? n9641 : n18337;
  assign n18339 = pi20 ? n313 : n12884;
  assign n18340 = pi19 ? n18338 : n18339;
  assign n18341 = pi20 ? n313 : ~n6621;
  assign n18342 = pi20 ? n18073 : n6621;
  assign n18343 = pi19 ? n18341 : ~n18342;
  assign n18344 = pi18 ? n18340 : ~n18343;
  assign n18345 = pi20 ? n12884 : ~n266;
  assign n18346 = pi19 ? n18345 : n16002;
  assign n18347 = pi18 ? n18346 : n32;
  assign n18348 = pi17 ? n18344 : n18347;
  assign n18349 = pi16 ? n18336 : n18348;
  assign n18350 = pi15 ? n18186 : n18349;
  assign n18351 = pi14 ? n18182 : n18350;
  assign n18352 = pi19 ? n18345 : ~n9028;
  assign n18353 = pi18 ? n18352 : n32;
  assign n18354 = pi17 ? n18344 : n18353;
  assign n18355 = pi16 ? n18336 : n18354;
  assign n18356 = pi18 ? n4127 : ~n18201;
  assign n18357 = pi17 ? n32 : n18356;
  assign n18358 = pi16 ? n18357 : n18207;
  assign n18359 = pi15 ? n18355 : n18358;
  assign n18360 = pi19 ? n32 : n9864;
  assign n18361 = pi18 ? n18360 : n32;
  assign n18362 = pi17 ? n32 : n18361;
  assign n18363 = pi16 ? n32 : n18362;
  assign n18364 = pi15 ? n18217 : n18363;
  assign n18365 = pi14 ? n18359 : n18364;
  assign n18366 = pi13 ? n18351 : n18365;
  assign n18367 = pi12 ? n18329 : n18366;
  assign n18368 = pi11 ? n18322 : n18367;
  assign n18369 = pi10 ? n18302 : n18368;
  assign n18370 = pi09 ? n32 : n18369;
  assign n18371 = pi08 ? n18229 : n18370;
  assign n18372 = pi07 ? n18069 : n18371;
  assign n18373 = pi19 ? n18099 : n8946;
  assign n18374 = pi20 ? n339 : ~n266;
  assign n18375 = pi19 ? n18374 : ~n275;
  assign n18376 = pi18 ? n18373 : n18375;
  assign n18377 = pi20 ? n206 : n11107;
  assign n18378 = pi19 ? n5614 : ~n18377;
  assign n18379 = pi18 ? n18378 : n237;
  assign n18380 = pi17 ? n18376 : ~n18379;
  assign n18381 = pi16 ? n18098 : n18380;
  assign n18382 = pi15 ? n32 : n18381;
  assign n18383 = pi14 ? n32 : n18382;
  assign n18384 = pi13 ? n32 : n18383;
  assign n18385 = pi19 ? n18110 : n14877;
  assign n18386 = pi20 ? n749 : ~n220;
  assign n18387 = pi20 ? n2385 : ~n5854;
  assign n18388 = pi19 ? n18386 : n18387;
  assign n18389 = pi18 ? n18385 : n18388;
  assign n18390 = pi20 ? n321 : n246;
  assign n18391 = pi19 ? n5614 : ~n18390;
  assign n18392 = pi18 ? n18391 : n237;
  assign n18393 = pi17 ? n18389 : ~n18392;
  assign n18394 = pi16 ? n18109 : n18393;
  assign n18395 = pi18 ? n32 : n4671;
  assign n18396 = pi20 ? n342 : n246;
  assign n18397 = pi19 ? n18396 : n246;
  assign n18398 = pi18 ? n18397 : ~n237;
  assign n18399 = pi17 ? n18395 : n18398;
  assign n18400 = pi16 ? n32 : n18399;
  assign n18401 = pi15 ? n18394 : n18400;
  assign n18402 = pi19 ? n32 : n1325;
  assign n18403 = pi20 ? n18073 : n9194;
  assign n18404 = pi20 ? n9488 : ~n18253;
  assign n18405 = pi19 ? n18403 : n18404;
  assign n18406 = pi18 ? n18402 : n18405;
  assign n18407 = pi17 ? n32 : n18406;
  assign n18408 = pi21 ? n173 : ~n173;
  assign n18409 = pi20 ? n18408 : ~n18282;
  assign n18410 = pi20 ? n17669 : n9491;
  assign n18411 = pi19 ? n18409 : ~n18410;
  assign n18412 = pi20 ? n9491 : n18281;
  assign n18413 = pi19 ? n18412 : n9194;
  assign n18414 = pi18 ? n18411 : ~n18413;
  assign n18415 = pi21 ? n313 : ~n174;
  assign n18416 = pi20 ? n17669 : n18415;
  assign n18417 = pi19 ? n18416 : ~n18408;
  assign n18418 = pi18 ? n18417 : ~n237;
  assign n18419 = pi17 ? n18414 : ~n18418;
  assign n18420 = pi16 ? n18407 : ~n18419;
  assign n18421 = pi15 ? n18420 : n32;
  assign n18422 = pi14 ? n18401 : n18421;
  assign n18423 = pi21 ? n16649 : n32;
  assign n18424 = pi20 ? n18423 : n32;
  assign n18425 = pi19 ? n18424 : n32;
  assign n18426 = pi18 ? n32 : n18425;
  assign n18427 = pi17 ? n32 : n18426;
  assign n18428 = pi16 ? n32 : n18427;
  assign n18429 = pi15 ? n57 : n18428;
  assign n18430 = pi15 ? n41 : n18294;
  assign n18431 = pi14 ? n18429 : n18430;
  assign n18432 = pi13 ? n18422 : n18431;
  assign n18433 = pi12 ? n18384 : n18432;
  assign n18434 = pi11 ? n32 : n18433;
  assign n18435 = pi15 ? n18294 : n18142;
  assign n18436 = pi14 ? n18435 : n18304;
  assign n18437 = pi18 ? n863 : ~n618;
  assign n18438 = pi17 ? n32 : n18437;
  assign n18439 = pi16 ? n32 : n18438;
  assign n18440 = pi15 ? n18008 : n18439;
  assign n18441 = pi14 ? n32 : n18440;
  assign n18442 = pi13 ? n18436 : n18441;
  assign n18443 = pi15 ? n17894 : n17891;
  assign n18444 = pi14 ? n18143 : n18443;
  assign n18445 = pi18 ? n209 : ~n1676;
  assign n18446 = pi17 ? n32 : n18445;
  assign n18447 = pi16 ? n32 : n18446;
  assign n18448 = pi15 ? n18309 : n18447;
  assign n18449 = pi15 ? n18019 : n17903;
  assign n18450 = pi14 ? n18448 : n18449;
  assign n18451 = pi13 ? n18444 : n18450;
  assign n18452 = pi12 ? n18442 : n18451;
  assign n18453 = pi15 ? n17825 : n17637;
  assign n18454 = pi14 ? n18020 : n18453;
  assign n18455 = pi15 ? n17637 : n17825;
  assign n18456 = pi20 ? n1331 : ~n428;
  assign n18457 = pi19 ? n32 : n18456;
  assign n18458 = pi18 ? n18457 : n32;
  assign n18459 = pi17 ? n32 : n18458;
  assign n18460 = pi16 ? n32 : n18459;
  assign n18461 = pi15 ? n17922 : n18460;
  assign n18462 = pi14 ? n18455 : n18461;
  assign n18463 = pi13 ? n18454 : n18462;
  assign n18464 = pi20 ? n266 : n2140;
  assign n18465 = pi19 ? n32 : ~n18464;
  assign n18466 = pi18 ? n18465 : n32;
  assign n18467 = pi17 ? n32 : n18466;
  assign n18468 = pi16 ? n32 : n18467;
  assign n18469 = pi19 ? n594 : ~n2141;
  assign n18470 = pi18 ? n18469 : n32;
  assign n18471 = pi17 ? n32 : n18470;
  assign n18472 = pi16 ? n32 : n18471;
  assign n18473 = pi15 ? n18468 : n18472;
  assign n18474 = pi19 ? n594 : ~n236;
  assign n18475 = pi18 ? n209 : ~n18474;
  assign n18476 = pi17 ? n32 : n18475;
  assign n18477 = pi16 ? n18476 : ~n2144;
  assign n18478 = pi20 ? n207 : n321;
  assign n18479 = pi19 ? n9037 : ~n18478;
  assign n18480 = pi18 ? n222 : ~n18479;
  assign n18481 = pi17 ? n32 : n18480;
  assign n18482 = pi18 ? n6059 : n32;
  assign n18483 = pi17 ? n18482 : n2143;
  assign n18484 = pi16 ? n18481 : ~n18483;
  assign n18485 = pi15 ? n18477 : n18484;
  assign n18486 = pi14 ? n18473 : n18485;
  assign n18487 = pi18 ? n32 : ~n350;
  assign n18488 = pi17 ? n32 : n18487;
  assign n18489 = pi20 ? n266 : n342;
  assign n18490 = pi19 ? n18489 : ~n18390;
  assign n18491 = pi18 ? n508 : ~n18490;
  assign n18492 = pi19 ? n349 : ~n2141;
  assign n18493 = pi18 ? n18492 : n32;
  assign n18494 = pi17 ? n18491 : n18493;
  assign n18495 = pi16 ? n18488 : n18494;
  assign n18496 = pi20 ? n246 : ~n266;
  assign n18497 = pi20 ? n220 : n246;
  assign n18498 = pi19 ? n18496 : ~n18497;
  assign n18499 = pi18 ? n222 : ~n18498;
  assign n18500 = pi17 ? n32 : n18499;
  assign n18501 = pi19 ? n1757 : n1464;
  assign n18502 = pi20 ? n207 : ~n266;
  assign n18503 = pi19 ? n18502 : ~n267;
  assign n18504 = pi18 ? n18501 : ~n18503;
  assign n18505 = pi20 ? n206 : n1319;
  assign n18506 = pi19 ? n32 : n18505;
  assign n18507 = pi18 ? n18506 : ~n32;
  assign n18508 = pi17 ? n18504 : n18507;
  assign n18509 = pi16 ? n18500 : ~n18508;
  assign n18510 = pi15 ? n18495 : n18509;
  assign n18511 = pi14 ? n18510 : n17707;
  assign n18512 = pi13 ? n18486 : n18511;
  assign n18513 = pi12 ? n18463 : n18512;
  assign n18514 = pi11 ? n18452 : n18513;
  assign n18515 = pi10 ? n18434 : n18514;
  assign n18516 = pi09 ? n32 : n18515;
  assign n18517 = pi19 ? n176 : n8622;
  assign n18518 = pi18 ? n858 : n18517;
  assign n18519 = pi20 ? n354 : ~n357;
  assign n18520 = pi19 ? n18519 : ~n4491;
  assign n18521 = pi19 ? n7488 : n32;
  assign n18522 = pi18 ? n18520 : ~n18521;
  assign n18523 = pi17 ? n18518 : ~n18522;
  assign n18524 = pi16 ? n32 : n18523;
  assign n18525 = pi15 ? n18524 : n32;
  assign n18526 = pi14 ? n32 : n18525;
  assign n18527 = pi13 ? n32 : n18526;
  assign n18528 = pi12 ? n32 : n18527;
  assign n18529 = pi18 ? n32 : n18521;
  assign n18530 = pi17 ? n32 : n18529;
  assign n18531 = pi16 ? n32 : n18530;
  assign n18532 = pi19 ? n5614 : n32;
  assign n18533 = pi18 ? n32 : n18532;
  assign n18534 = pi17 ? n32 : n18533;
  assign n18535 = pi16 ? n32 : n18534;
  assign n18536 = pi15 ? n18535 : n32;
  assign n18537 = pi14 ? n18531 : n18536;
  assign n18538 = pi19 ? n18246 : ~n5855;
  assign n18539 = pi18 ? n18538 : ~n275;
  assign n18540 = pi21 ? n259 : ~n313;
  assign n18541 = pi20 ? n18173 : n18540;
  assign n18542 = pi19 ? n5614 : ~n18541;
  assign n18543 = pi18 ? n18542 : n814;
  assign n18544 = pi17 ? n18539 : ~n18543;
  assign n18545 = pi16 ? n18244 : n18544;
  assign n18546 = pi15 ? n32 : n18545;
  assign n18547 = pi14 ? n32 : n18546;
  assign n18548 = pi13 ? n18537 : n18547;
  assign n18549 = pi20 ? n260 : n439;
  assign n18550 = pi19 ? n18262 : ~n18549;
  assign n18551 = pi20 ? n439 : n5854;
  assign n18552 = pi20 ? n1091 : n6303;
  assign n18553 = pi19 ? n18551 : n18552;
  assign n18554 = pi18 ? n18550 : ~n18553;
  assign n18555 = pi20 ? n2358 : n12884;
  assign n18556 = pi19 ? n5614 : ~n18555;
  assign n18557 = pi18 ? n18556 : n814;
  assign n18558 = pi17 ? n18554 : ~n18557;
  assign n18559 = pi16 ? n18260 : n18558;
  assign n18560 = pi18 ? n32 : n9170;
  assign n18561 = pi17 ? n32 : n18560;
  assign n18562 = pi18 ? n18397 : ~n814;
  assign n18563 = pi17 ? n18395 : n18562;
  assign n18564 = pi16 ? n18561 : n18563;
  assign n18565 = pi15 ? n18559 : n18564;
  assign n18566 = pi20 ? n9641 : n1817;
  assign n18567 = pi20 ? n6085 : n1331;
  assign n18568 = pi19 ? n18566 : n18567;
  assign n18569 = pi18 ? n18402 : n18568;
  assign n18570 = pi17 ? n32 : n18569;
  assign n18571 = pi20 ? n18173 : ~n17671;
  assign n18572 = pi20 ? n1324 : n9641;
  assign n18573 = pi19 ? n18571 : ~n18572;
  assign n18574 = pi20 ? n9641 : n17671;
  assign n18575 = pi20 ? n1817 : n17665;
  assign n18576 = pi19 ? n18574 : n18575;
  assign n18577 = pi18 ? n18573 : ~n18576;
  assign n18578 = pi20 ? n17669 : n333;
  assign n18579 = pi19 ? n18578 : ~n18173;
  assign n18580 = pi18 ? n18579 : ~n618;
  assign n18581 = pi17 ? n18577 : ~n18580;
  assign n18582 = pi16 ? n18570 : ~n18581;
  assign n18583 = pi15 ? n18582 : n32;
  assign n18584 = pi14 ? n18565 : n18583;
  assign n18585 = pi15 ? n32 : n18294;
  assign n18586 = pi14 ? n57 : n18585;
  assign n18587 = pi13 ? n18584 : n18586;
  assign n18588 = pi12 ? n18548 : n18587;
  assign n18589 = pi11 ? n18528 : n18588;
  assign n18590 = pi15 ? n18294 : n32;
  assign n18591 = pi14 ? n41 : n18590;
  assign n18592 = pi18 ? n863 : ~n3350;
  assign n18593 = pi17 ? n32 : n18592;
  assign n18594 = pi16 ? n32 : n18593;
  assign n18595 = pi15 ? n18297 : n18594;
  assign n18596 = pi14 ? n32 : n18595;
  assign n18597 = pi13 ? n18591 : n18596;
  assign n18598 = pi14 ? n18008 : n18440;
  assign n18599 = pi18 ? n940 : ~n618;
  assign n18600 = pi17 ? n32 : n18599;
  assign n18601 = pi16 ? n32 : n18600;
  assign n18602 = pi18 ? n209 : ~n618;
  assign n18603 = pi17 ? n32 : n18602;
  assign n18604 = pi16 ? n32 : n18603;
  assign n18605 = pi15 ? n18601 : n18604;
  assign n18606 = pi15 ? n18309 : n17891;
  assign n18607 = pi14 ? n18605 : n18606;
  assign n18608 = pi13 ? n18598 : n18607;
  assign n18609 = pi12 ? n18597 : n18608;
  assign n18610 = pi21 ? n32 : n10445;
  assign n18611 = pi20 ? n266 : n18610;
  assign n18612 = pi19 ? n32 : ~n18611;
  assign n18613 = pi18 ? n18612 : n32;
  assign n18614 = pi17 ? n32 : n18613;
  assign n18615 = pi16 ? n32 : n18614;
  assign n18616 = pi20 ? n17669 : n6822;
  assign n18617 = pi20 ? n8644 : n9491;
  assign n18618 = pi19 ? n18616 : ~n18617;
  assign n18619 = pi18 ? n335 : ~n18618;
  assign n18620 = pi17 ? n32 : n18619;
  assign n18621 = pi20 ? n18281 : n333;
  assign n18622 = pi20 ? n405 : n6621;
  assign n18623 = pi19 ? n18621 : ~n18622;
  assign n18624 = pi21 ? n206 : n313;
  assign n18625 = pi20 ? n333 : ~n18624;
  assign n18626 = pi20 ? n18073 : ~n18073;
  assign n18627 = pi19 ? n18625 : ~n18626;
  assign n18628 = pi18 ? n18623 : ~n18627;
  assign n18629 = pi20 ? n18073 : ~n313;
  assign n18630 = pi19 ? n18629 : ~n2141;
  assign n18631 = pi18 ? n18630 : n32;
  assign n18632 = pi17 ? n18628 : n18631;
  assign n18633 = pi16 ? n18620 : n18632;
  assign n18634 = pi15 ? n18615 : n18633;
  assign n18635 = pi14 ? n18634 : n18485;
  assign n18636 = pi15 ? n17717 : n17707;
  assign n18637 = pi14 ? n18510 : n18636;
  assign n18638 = pi13 ? n18635 : n18637;
  assign n18639 = pi12 ? n18463 : n18638;
  assign n18640 = pi11 ? n18609 : n18639;
  assign n18641 = pi10 ? n18589 : n18640;
  assign n18642 = pi09 ? n32 : n18641;
  assign n18643 = pi08 ? n18516 : n18642;
  assign n18644 = pi20 ? n357 : n17665;
  assign n18645 = pi19 ? n18644 : n1464;
  assign n18646 = pi18 ? n6071 : n18645;
  assign n18647 = pi19 ? n18572 : n274;
  assign n18648 = pi18 ? n18647 : n6059;
  assign n18649 = pi17 ? n18646 : n18648;
  assign n18650 = pi16 ? n32 : n18649;
  assign n18651 = pi15 ? n18650 : n32;
  assign n18652 = pi14 ? n32 : n18651;
  assign n18653 = pi13 ? n32 : n18652;
  assign n18654 = pi12 ? n32 : n18653;
  assign n18655 = pi18 ? n32 : n6867;
  assign n18656 = pi17 ? n32 : n18655;
  assign n18657 = pi16 ? n32 : n18656;
  assign n18658 = pi19 ? n6230 : n32;
  assign n18659 = pi18 ? n32 : n18658;
  assign n18660 = pi17 ? n32 : n18659;
  assign n18661 = pi16 ? n32 : n18660;
  assign n18662 = pi15 ? n18657 : n18661;
  assign n18663 = pi15 ? n18661 : n32;
  assign n18664 = pi14 ? n18662 : n18663;
  assign n18665 = pi20 ? n357 : n246;
  assign n18666 = pi19 ? n18665 : n32;
  assign n18667 = pi18 ? n32 : n18666;
  assign n18668 = pi19 ? n32 : n266;
  assign n18669 = pi18 ? n18668 : n18532;
  assign n18670 = pi17 ? n18667 : n18669;
  assign n18671 = pi16 ? n32 : n18670;
  assign n18672 = pi16 ? n1705 : ~n2137;
  assign n18673 = pi15 ? n18671 : n18672;
  assign n18674 = pi14 ? n32 : n18673;
  assign n18675 = pi13 ? n18664 : n18674;
  assign n18676 = pi16 ? n1471 : ~n2137;
  assign n18677 = pi20 ? n2358 : ~n266;
  assign n18678 = pi20 ? n246 : n342;
  assign n18679 = pi19 ? n18677 : ~n18678;
  assign n18680 = pi18 ? n1862 : n18679;
  assign n18681 = pi17 ? n32 : n18680;
  assign n18682 = pi16 ? n18681 : ~n2137;
  assign n18683 = pi15 ? n18676 : n18682;
  assign n18684 = pi14 ? n18683 : n32;
  assign n18685 = pi19 ? n7502 : n32;
  assign n18686 = pi18 ? n32 : n18685;
  assign n18687 = pi17 ? n32 : n18686;
  assign n18688 = pi16 ? n32 : n18687;
  assign n18689 = pi15 ? n57 : n18688;
  assign n18690 = pi14 ? n18535 : n18689;
  assign n18691 = pi13 ? n18684 : n18690;
  assign n18692 = pi12 ? n18675 : n18691;
  assign n18693 = pi11 ? n18654 : n18692;
  assign n18694 = pi15 ? n18688 : n18294;
  assign n18695 = pi15 ? n41 : n32;
  assign n18696 = pi14 ? n18694 : n18695;
  assign n18697 = pi15 ? n18142 : n18594;
  assign n18698 = pi14 ? n32 : n18697;
  assign n18699 = pi13 ? n18696 : n18698;
  assign n18700 = pi12 ? n18699 : n18608;
  assign n18701 = pi14 ? n18309 : n17910;
  assign n18702 = pi20 ? n274 : ~n101;
  assign n18703 = pi19 ? n32 : n18702;
  assign n18704 = pi18 ? n18703 : n32;
  assign n18705 = pi17 ? n32 : n18704;
  assign n18706 = pi16 ? n32 : n18705;
  assign n18707 = pi15 ? n18026 : n18706;
  assign n18708 = pi14 ? n17916 : n18707;
  assign n18709 = pi13 ? n18701 : n18708;
  assign n18710 = pi19 ? n32 : n2359;
  assign n18711 = pi18 ? n18710 : ~n3496;
  assign n18712 = pi17 ? n32 : n18711;
  assign n18713 = pi16 ? n18712 : ~n1834;
  assign n18714 = pi20 ? n1685 : n207;
  assign n18715 = pi19 ? n11879 : n18714;
  assign n18716 = pi18 ? n863 : ~n18715;
  assign n18717 = pi17 ? n32 : n18716;
  assign n18718 = pi18 ? n4671 : n32;
  assign n18719 = pi17 ? n18718 : n1833;
  assign n18720 = pi16 ? n18717 : ~n18719;
  assign n18721 = pi15 ? n18713 : n18720;
  assign n18722 = pi20 ? n266 : ~n220;
  assign n18723 = pi19 ? n18722 : ~n15983;
  assign n18724 = pi18 ? n863 : ~n18723;
  assign n18725 = pi17 ? n32 : n18724;
  assign n18726 = pi16 ? n18725 : ~n18719;
  assign n18727 = pi19 ? n267 : ~n206;
  assign n18728 = pi20 ? n246 : n266;
  assign n18729 = pi19 ? n267 : n18728;
  assign n18730 = pi18 ? n18727 : n18729;
  assign n18731 = pi19 ? n5435 : ~n594;
  assign n18732 = pi18 ? n18731 : n32;
  assign n18733 = pi17 ? n18730 : n18732;
  assign n18734 = pi16 ? n32 : n18733;
  assign n18735 = pi15 ? n18726 : n18734;
  assign n18736 = pi14 ? n18721 : n18735;
  assign n18737 = pi19 ? n208 : ~n594;
  assign n18738 = pi18 ? n18737 : n32;
  assign n18739 = pi17 ? n32 : n18738;
  assign n18740 = pi16 ? n32 : n18739;
  assign n18741 = pi20 ? n32 : n9641;
  assign n18742 = pi19 ? n18741 : n334;
  assign n18743 = pi18 ? n18742 : n32;
  assign n18744 = pi17 ? n32 : n18743;
  assign n18745 = pi16 ? n32 : n18744;
  assign n18746 = pi15 ? n18740 : n18745;
  assign n18747 = pi14 ? n18746 : n17717;
  assign n18748 = pi13 ? n18736 : n18747;
  assign n18749 = pi12 ? n18709 : n18748;
  assign n18750 = pi11 ? n18700 : n18749;
  assign n18751 = pi10 ? n18693 : n18750;
  assign n18752 = pi09 ? n32 : n18751;
  assign n18753 = pi19 ? n339 : ~n32;
  assign n18754 = pi18 ? n32 : ~n18753;
  assign n18755 = pi17 ? n32 : n18754;
  assign n18756 = pi20 ? n18129 : ~n18281;
  assign n18757 = pi19 ? n32 : n18756;
  assign n18758 = pi20 ? n18281 : n18415;
  assign n18759 = pi19 ? n18758 : n18253;
  assign n18760 = pi18 ? n18757 : ~n18759;
  assign n18761 = pi20 ? n18281 : n17652;
  assign n18762 = pi21 ? n309 : n405;
  assign n18763 = pi20 ? n1611 : n18762;
  assign n18764 = pi19 ? n18761 : ~n18763;
  assign n18765 = pi18 ? n18764 : ~n359;
  assign n18766 = pi17 ? n18760 : ~n18765;
  assign n18767 = pi16 ? n18755 : n18766;
  assign n18768 = pi15 ? n32 : n18767;
  assign n18769 = pi18 ? n6071 : n4380;
  assign n18770 = pi19 ? n6171 : n32;
  assign n18771 = pi18 ? n18770 : n6867;
  assign n18772 = pi17 ? n18769 : n18771;
  assign n18773 = pi16 ? n32 : n18772;
  assign n18774 = pi15 ? n18773 : n18657;
  assign n18775 = pi14 ? n18768 : n18774;
  assign n18776 = pi13 ? n32 : n18775;
  assign n18777 = pi12 ? n32 : n18776;
  assign n18778 = pi20 ? n18253 : n18408;
  assign n18779 = pi19 ? n9488 : ~n18778;
  assign n18780 = pi18 ? n858 : n18779;
  assign n18781 = pi17 ? n32 : n18780;
  assign n18782 = pi20 ? n18282 : n9194;
  assign n18783 = pi20 ? n6085 : n448;
  assign n18784 = pi19 ? n18782 : n18783;
  assign n18785 = pi20 ? n448 : n1385;
  assign n18786 = pi20 ? n9488 : n18129;
  assign n18787 = pi19 ? n18785 : n18786;
  assign n18788 = pi18 ? n18784 : n18787;
  assign n18789 = pi20 ? n18129 : n32;
  assign n18790 = pi19 ? n18789 : n1685;
  assign n18791 = pi18 ? n18790 : n18532;
  assign n18792 = pi17 ? n18788 : n18791;
  assign n18793 = pi16 ? n18781 : n18792;
  assign n18794 = pi16 ? n1705 : ~n1815;
  assign n18795 = pi15 ? n18793 : n18794;
  assign n18796 = pi14 ? n32 : n18795;
  assign n18797 = pi13 ? n18664 : n18796;
  assign n18798 = pi16 ? n1471 : ~n1815;
  assign n18799 = pi16 ? n18681 : ~n1815;
  assign n18800 = pi15 ? n18798 : n18799;
  assign n18801 = pi14 ? n18800 : n32;
  assign n18802 = pi19 ? n1630 : n32;
  assign n18803 = pi18 ? n32 : n18802;
  assign n18804 = pi17 ? n32 : n18803;
  assign n18805 = pi16 ? n32 : n18804;
  assign n18806 = pi15 ? n32 : n18688;
  assign n18807 = pi14 ? n18805 : n18806;
  assign n18808 = pi13 ? n18801 : n18807;
  assign n18809 = pi12 ? n18797 : n18808;
  assign n18810 = pi11 ? n18777 : n18809;
  assign n18811 = pi14 ? n18688 : n32;
  assign n18812 = pi18 ? n863 : ~n237;
  assign n18813 = pi17 ? n32 : n18812;
  assign n18814 = pi16 ? n32 : n18813;
  assign n18815 = pi15 ? n18294 : n18814;
  assign n18816 = pi14 ? n32 : n18815;
  assign n18817 = pi13 ? n18811 : n18816;
  assign n18818 = pi14 ? n18297 : n18595;
  assign n18819 = pi18 ? n940 : ~n3350;
  assign n18820 = pi17 ? n32 : n18819;
  assign n18821 = pi16 ? n32 : n18820;
  assign n18822 = pi15 ? n18821 : n18604;
  assign n18823 = pi15 ? n18601 : n17891;
  assign n18824 = pi14 ? n18822 : n18823;
  assign n18825 = pi13 ? n18818 : n18824;
  assign n18826 = pi12 ? n18817 : n18825;
  assign n18827 = pi15 ? n18309 : n18019;
  assign n18828 = pi14 ? n18827 : n17910;
  assign n18829 = pi21 ? n10182 : n309;
  assign n18830 = pi20 ? n32 : n18829;
  assign n18831 = pi19 ? n32 : n18830;
  assign n18832 = pi21 ? n173 : ~n309;
  assign n18833 = pi20 ? n18281 : ~n18832;
  assign n18834 = pi21 ? n313 : n206;
  assign n18835 = pi20 ? n18834 : n18281;
  assign n18836 = pi19 ? n18833 : ~n18835;
  assign n18837 = pi18 ? n18831 : ~n18836;
  assign n18838 = pi17 ? n32 : n18837;
  assign n18839 = pi20 ? n18415 : n333;
  assign n18840 = pi21 ? n313 : n174;
  assign n18841 = pi20 ? n18840 : n18337;
  assign n18842 = pi19 ? n18839 : ~n18841;
  assign n18843 = pi20 ? n309 : ~n313;
  assign n18844 = pi20 ? n18624 : ~n18624;
  assign n18845 = pi19 ? n18843 : n18844;
  assign n18846 = pi18 ? n18842 : ~n18845;
  assign n18847 = pi20 ? n18624 : ~n6621;
  assign n18848 = pi20 ? n1685 : ~n428;
  assign n18849 = pi19 ? n18847 : ~n18848;
  assign n18850 = pi18 ? n18849 : ~n32;
  assign n18851 = pi17 ? n18846 : ~n18850;
  assign n18852 = pi16 ? n18838 : n18851;
  assign n18853 = pi15 ? n18026 : n18852;
  assign n18854 = pi14 ? n17916 : n18853;
  assign n18855 = pi13 ? n18828 : n18854;
  assign n18856 = pi19 ? n208 : ~n2141;
  assign n18857 = pi18 ? n18856 : n32;
  assign n18858 = pi17 ? n32 : n18857;
  assign n18859 = pi16 ? n32 : n18858;
  assign n18860 = pi19 ? n1818 : n6398;
  assign n18861 = pi18 ? n18860 : n32;
  assign n18862 = pi17 ? n32 : n18861;
  assign n18863 = pi16 ? n32 : n18862;
  assign n18864 = pi15 ? n18859 : n18863;
  assign n18865 = pi20 ? n32 : n7377;
  assign n18866 = pi19 ? n32 : n18865;
  assign n18867 = pi18 ? n18866 : n32;
  assign n18868 = pi17 ? n32 : n18867;
  assign n18869 = pi16 ? n32 : n18868;
  assign n18870 = pi15 ? n18869 : n17729;
  assign n18871 = pi14 ? n18864 : n18870;
  assign n18872 = pi13 ? n18736 : n18871;
  assign n18873 = pi12 ? n18855 : n18872;
  assign n18874 = pi11 ? n18826 : n18873;
  assign n18875 = pi10 ? n18810 : n18874;
  assign n18876 = pi09 ? n32 : n18875;
  assign n18877 = pi08 ? n18752 : n18876;
  assign n18878 = pi07 ? n18643 : n18877;
  assign n18879 = pi06 ? n18372 : n18878;
  assign n18880 = pi05 ? n17873 : n18879;
  assign n18881 = pi04 ? n32 : n18880;
  assign n18882 = pi19 ? n6350 : n32;
  assign n18883 = pi18 ? n32 : ~n18882;
  assign n18884 = pi17 ? n32 : n18883;
  assign n18885 = pi16 ? n18884 : ~n3338;
  assign n18886 = pi15 ? n32 : n18885;
  assign n18887 = pi19 ? n5446 : n32;
  assign n18888 = pi18 ? n32 : n18887;
  assign n18889 = pi17 ? n32 : n18888;
  assign n18890 = pi16 ? n32 : n18889;
  assign n18891 = pi19 ? n207 : ~n32;
  assign n18892 = pi18 ? n32 : ~n18891;
  assign n18893 = pi19 ? n1508 : n4670;
  assign n18894 = pi19 ? n16310 : n32;
  assign n18895 = pi18 ? n18893 : n18894;
  assign n18896 = pi17 ? n18892 : n18895;
  assign n18897 = pi16 ? n32 : n18896;
  assign n18898 = pi15 ? n18890 : n18897;
  assign n18899 = pi14 ? n18886 : n18898;
  assign n18900 = pi13 ? n32 : n18899;
  assign n18901 = pi12 ? n32 : n18900;
  assign n18902 = pi18 ? n32 : n18894;
  assign n18903 = pi17 ? n32 : n18902;
  assign n18904 = pi16 ? n32 : n18903;
  assign n18905 = pi15 ? n18904 : n18657;
  assign n18906 = pi15 ? n18657 : n32;
  assign n18907 = pi14 ? n18905 : n18906;
  assign n18908 = pi19 ? n32 : n18741;
  assign n18909 = pi20 ? n18282 : n17652;
  assign n18910 = pi20 ? n18253 : ~n333;
  assign n18911 = pi19 ? n18909 : n18910;
  assign n18912 = pi18 ? n18908 : n18911;
  assign n18913 = pi17 ? n32 : n18912;
  assign n18914 = pi19 ? n32 : n18130;
  assign n18915 = pi20 ? n2180 : n18253;
  assign n18916 = pi19 ? n17652 : n18915;
  assign n18917 = pi18 ? n18914 : ~n18916;
  assign n18918 = pi20 ? n18415 : ~n9491;
  assign n18919 = pi20 ? n9641 : n428;
  assign n18920 = pi19 ? n18918 : ~n18919;
  assign n18921 = pi18 ? n18920 : ~n618;
  assign n18922 = pi17 ? n18917 : ~n18921;
  assign n18923 = pi16 ? n18913 : ~n18922;
  assign n18924 = pi20 ? n17652 : n32;
  assign n18925 = pi19 ? n857 : ~n18924;
  assign n18926 = pi18 ? n32 : n18925;
  assign n18927 = pi17 ? n32 : n18926;
  assign n18928 = pi19 ? n1757 : n266;
  assign n18929 = pi18 ? n268 : n18928;
  assign n18930 = pi18 ? n6059 : n1813;
  assign n18931 = pi17 ? n18929 : n18930;
  assign n18932 = pi16 ? n18927 : ~n18931;
  assign n18933 = pi15 ? n18923 : n18932;
  assign n18934 = pi14 ? n32 : n18933;
  assign n18935 = pi13 ? n18907 : n18934;
  assign n18936 = pi19 ? n32 : n18404;
  assign n18937 = pi18 ? n32 : n18936;
  assign n18938 = pi17 ? n32 : n18937;
  assign n18939 = pi19 ? n358 : n267;
  assign n18940 = pi18 ? n18939 : n18928;
  assign n18941 = pi19 ? n266 : n32;
  assign n18942 = pi18 ? n18941 : n1813;
  assign n18943 = pi17 ? n18940 : n18942;
  assign n18944 = pi16 ? n18938 : ~n18943;
  assign n18945 = pi15 ? n18944 : n32;
  assign n18946 = pi14 ? n18945 : n32;
  assign n18947 = pi15 ? n18661 : n18531;
  assign n18948 = pi15 ? n18805 : n18535;
  assign n18949 = pi14 ? n18947 : n18948;
  assign n18950 = pi13 ? n18946 : n18949;
  assign n18951 = pi12 ? n18935 : n18950;
  assign n18952 = pi11 ? n18901 : n18951;
  assign n18953 = pi14 ? n57 : n32;
  assign n18954 = pi15 ? n18814 : n18294;
  assign n18955 = pi14 ? n32 : n18954;
  assign n18956 = pi13 ? n18953 : n18955;
  assign n18957 = pi18 ? n863 : n18076;
  assign n18958 = pi17 ? n32 : n18957;
  assign n18959 = pi16 ? n32 : n18958;
  assign n18960 = pi15 ? n18142 : n18959;
  assign n18961 = pi14 ? n18142 : n18960;
  assign n18962 = pi15 ? n18821 : n18601;
  assign n18963 = pi18 ? n1139 : ~n618;
  assign n18964 = pi17 ? n32 : n18963;
  assign n18965 = pi16 ? n32 : n18964;
  assign n18966 = pi15 ? n18965 : n18439;
  assign n18967 = pi14 ? n18962 : n18966;
  assign n18968 = pi13 ? n18961 : n18967;
  assign n18969 = pi12 ? n18956 : n18968;
  assign n18970 = pi18 ? n936 : ~n1676;
  assign n18971 = pi17 ? n32 : n18970;
  assign n18972 = pi16 ? n32 : n18971;
  assign n18973 = pi15 ? n18601 : n18972;
  assign n18974 = pi14 ? n18973 : n17885;
  assign n18975 = pi18 ? n2043 : n32;
  assign n18976 = pi17 ? n32 : n18975;
  assign n18977 = pi16 ? n32 : n18976;
  assign n18978 = pi15 ? n17903 : n18977;
  assign n18979 = pi16 ? n1135 : ~n1683;
  assign n18980 = pi18 ? n341 : ~n16389;
  assign n18981 = pi17 ? n32 : n18980;
  assign n18982 = pi20 ? n32 : n12019;
  assign n18983 = pi19 ? n32 : n18982;
  assign n18984 = pi18 ? n18983 : ~n32;
  assign n18985 = pi17 ? n32 : n18984;
  assign n18986 = pi16 ? n18981 : ~n18985;
  assign n18987 = pi15 ? n18979 : n18986;
  assign n18988 = pi14 ? n18978 : n18987;
  assign n18989 = pi13 ? n18974 : n18988;
  assign n18990 = pi18 ? n341 : ~n15844;
  assign n18991 = pi17 ? n32 : n18990;
  assign n18992 = pi16 ? n18991 : ~n18985;
  assign n18993 = pi18 ? n940 : ~n15849;
  assign n18994 = pi17 ? n32 : n18993;
  assign n18995 = pi16 ? n18994 : ~n1577;
  assign n18996 = pi15 ? n18992 : n18995;
  assign n18997 = pi19 ? n507 : ~n1574;
  assign n18998 = pi18 ? n18997 : n32;
  assign n18999 = pi17 ? n32 : n18998;
  assign n19000 = pi16 ? n32 : n18999;
  assign n19001 = pi19 ? n32 : n12578;
  assign n19002 = pi18 ? n19001 : n32;
  assign n19003 = pi17 ? n32 : n19002;
  assign n19004 = pi16 ? n32 : n19003;
  assign n19005 = pi15 ? n19000 : n19004;
  assign n19006 = pi14 ? n18996 : n19005;
  assign n19007 = pi19 ? n32 : n12572;
  assign n19008 = pi18 ? n19007 : n32;
  assign n19009 = pi17 ? n32 : n19008;
  assign n19010 = pi16 ? n32 : n19009;
  assign n19011 = pi15 ? n19010 : n18326;
  assign n19012 = pi15 ? n17851 : n18326;
  assign n19013 = pi14 ? n19011 : n19012;
  assign n19014 = pi13 ? n19006 : n19013;
  assign n19015 = pi12 ? n18989 : n19014;
  assign n19016 = pi11 ? n18969 : n19015;
  assign n19017 = pi10 ? n18952 : n19016;
  assign n19018 = pi09 ? n32 : n19017;
  assign n19019 = pi20 ? n2102 : n32;
  assign n19020 = pi19 ? n19019 : n32;
  assign n19021 = pi18 ? n18893 : n19020;
  assign n19022 = pi17 ? n18892 : n19021;
  assign n19023 = pi16 ? n32 : n19022;
  assign n19024 = pi15 ? n165 : n19023;
  assign n19025 = pi14 ? n18886 : n19024;
  assign n19026 = pi13 ? n32 : n19025;
  assign n19027 = pi12 ? n32 : n19026;
  assign n19028 = pi18 ? n32 : n19020;
  assign n19029 = pi17 ? n32 : n19028;
  assign n19030 = pi16 ? n32 : n19029;
  assign n19031 = pi15 ? n19030 : n18890;
  assign n19032 = pi15 ? n18890 : n32;
  assign n19033 = pi14 ? n19031 : n19032;
  assign n19034 = pi20 ? n6085 : ~n5854;
  assign n19035 = pi19 ? n32 : n19034;
  assign n19036 = pi18 ? n32 : n19035;
  assign n19037 = pi17 ? n32 : n19036;
  assign n19038 = pi16 ? n19037 : ~n18922;
  assign n19039 = pi18 ? n6059 : n814;
  assign n19040 = pi17 ? n18929 : n19039;
  assign n19041 = pi16 ? n18927 : ~n19040;
  assign n19042 = pi15 ? n19038 : n19041;
  assign n19043 = pi14 ? n32 : n19042;
  assign n19044 = pi13 ? n19033 : n19043;
  assign n19045 = pi20 ? n32 : ~n18173;
  assign n19046 = pi19 ? n32 : n19045;
  assign n19047 = pi18 ? n32 : n19046;
  assign n19048 = pi17 ? n32 : n19047;
  assign n19049 = pi18 ? n18941 : n814;
  assign n19050 = pi17 ? n18940 : n19049;
  assign n19051 = pi16 ? n19048 : ~n19050;
  assign n19052 = pi15 ? n19051 : n32;
  assign n19053 = pi14 ? n19052 : n32;
  assign n19054 = pi14 ? n18947 : n18535;
  assign n19055 = pi13 ? n19053 : n19054;
  assign n19056 = pi12 ? n19044 : n19055;
  assign n19057 = pi11 ? n19027 : n19056;
  assign n19058 = pi14 ? n18805 : n32;
  assign n19059 = pi18 ? n863 : ~n1942;
  assign n19060 = pi17 ? n32 : n19059;
  assign n19061 = pi16 ? n32 : n19060;
  assign n19062 = pi15 ? n19061 : n18688;
  assign n19063 = pi14 ? n32 : n19062;
  assign n19064 = pi13 ? n19058 : n19063;
  assign n19065 = pi19 ? n15651 : n32;
  assign n19066 = pi18 ? n863 : n19065;
  assign n19067 = pi17 ? n32 : n19066;
  assign n19068 = pi16 ? n32 : n19067;
  assign n19069 = pi15 ? n18294 : n19068;
  assign n19070 = pi14 ? n18294 : n19069;
  assign n19071 = pi18 ? n940 : ~n237;
  assign n19072 = pi17 ? n32 : n19071;
  assign n19073 = pi16 ? n32 : n19072;
  assign n19074 = pi18 ? n751 : ~n3350;
  assign n19075 = pi17 ? n32 : n19074;
  assign n19076 = pi16 ? n32 : n19075;
  assign n19077 = pi15 ? n19073 : n19076;
  assign n19078 = pi15 ? n18821 : n18439;
  assign n19079 = pi14 ? n19077 : n19078;
  assign n19080 = pi13 ? n19070 : n19079;
  assign n19081 = pi12 ? n19064 : n19080;
  assign n19082 = pi19 ? n32 : n6057;
  assign n19083 = pi20 ? n1331 : n18762;
  assign n19084 = pi19 ? n19083 : n333;
  assign n19085 = pi18 ? n19082 : n19084;
  assign n19086 = pi17 ? n32 : n19085;
  assign n19087 = pi20 ? n3523 : ~n18173;
  assign n19088 = pi20 ? n13171 : n313;
  assign n19089 = pi19 ? n19087 : ~n19088;
  assign n19090 = pi20 ? n206 : n333;
  assign n19091 = pi20 ? n18624 : ~n18337;
  assign n19092 = pi19 ? n19090 : ~n19091;
  assign n19093 = pi18 ? n19089 : n19092;
  assign n19094 = pi20 ? n18073 : n18337;
  assign n19095 = pi19 ? n19094 : n4558;
  assign n19096 = pi18 ? n19095 : n32;
  assign n19097 = pi17 ? n19093 : n19096;
  assign n19098 = pi16 ? n19086 : n19097;
  assign n19099 = pi15 ? n17903 : n19098;
  assign n19100 = pi16 ? n1233 : ~n1683;
  assign n19101 = pi16 ? n18981 : ~n1581;
  assign n19102 = pi15 ? n19100 : n19101;
  assign n19103 = pi14 ? n19099 : n19102;
  assign n19104 = pi13 ? n18974 : n19103;
  assign n19105 = pi15 ? n19010 : n17702;
  assign n19106 = pi14 ? n19105 : n19012;
  assign n19107 = pi13 ? n19006 : n19106;
  assign n19108 = pi12 ? n19104 : n19107;
  assign n19109 = pi11 ? n19081 : n19108;
  assign n19110 = pi10 ? n19057 : n19109;
  assign n19111 = pi09 ? n32 : n19110;
  assign n19112 = pi08 ? n19018 : n19111;
  assign n19113 = pi20 ? n2385 : n175;
  assign n19114 = pi19 ? n32 : n19113;
  assign n19115 = pi20 ? n6050 : n501;
  assign n19116 = pi20 ? n32 : ~n2358;
  assign n19117 = pi19 ? n19115 : ~n19116;
  assign n19118 = pi18 ? n19114 : ~n19117;
  assign n19119 = pi20 ? n12884 : n333;
  assign n19120 = pi19 ? n19119 : ~n1611;
  assign n19121 = pi19 ? n10662 : n32;
  assign n19122 = pi18 ? n19120 : ~n19121;
  assign n19123 = pi17 ? n19118 : ~n19122;
  assign n19124 = pi16 ? n32 : n19123;
  assign n19125 = pi15 ? n165 : n19124;
  assign n19126 = pi14 ? n166 : n19125;
  assign n19127 = pi13 ? n32 : n19126;
  assign n19128 = pi12 ? n32 : n19127;
  assign n19129 = pi20 ? n18129 : n175;
  assign n19130 = pi19 ? n32 : n19129;
  assign n19131 = pi20 ? n354 : n501;
  assign n19132 = pi19 ? n19131 : ~n19116;
  assign n19133 = pi18 ? n19130 : ~n19132;
  assign n19134 = pi20 ? n17669 : ~n18832;
  assign n19135 = pi19 ? n19134 : ~n18762;
  assign n19136 = pi20 ? n2019 : n32;
  assign n19137 = pi19 ? n19136 : n32;
  assign n19138 = pi18 ? n19135 : ~n19137;
  assign n19139 = pi17 ? n19133 : ~n19138;
  assign n19140 = pi16 ? n32 : n19139;
  assign n19141 = pi20 ? n32 : n18129;
  assign n19142 = pi19 ? n19141 : n357;
  assign n19143 = pi18 ? n19142 : n18894;
  assign n19144 = pi17 ? n13950 : n19143;
  assign n19145 = pi16 ? n32 : n19144;
  assign n19146 = pi15 ? n19140 : n19145;
  assign n19147 = pi15 ? n18904 : n32;
  assign n19148 = pi14 ? n19146 : n19147;
  assign n19149 = pi19 ? n507 : n342;
  assign n19150 = pi18 ? n19149 : n342;
  assign n19151 = pi20 ? n206 : n342;
  assign n19152 = pi19 ? n18396 : ~n19151;
  assign n19153 = pi18 ? n19152 : n6059;
  assign n19154 = pi17 ? n19150 : n19153;
  assign n19155 = pi16 ? n32 : n19154;
  assign n19156 = pi15 ? n18657 : n19155;
  assign n19157 = pi14 ? n32 : n19156;
  assign n19158 = pi13 ? n19148 : n19157;
  assign n19159 = pi14 ? n18657 : n18531;
  assign n19160 = pi13 ? n32 : n19159;
  assign n19161 = pi12 ? n19158 : n19160;
  assign n19162 = pi11 ? n19128 : n19161;
  assign n19163 = pi14 ? n18535 : n32;
  assign n19164 = pi18 ? n32 : ~n1942;
  assign n19165 = pi17 ? n32 : n19164;
  assign n19166 = pi16 ? n32 : n19165;
  assign n19167 = pi15 ? n19166 : n18688;
  assign n19168 = pi14 ? n32 : n19167;
  assign n19169 = pi13 ? n19163 : n19168;
  assign n19170 = pi18 ? n32 : ~n237;
  assign n19171 = pi17 ? n32 : n19170;
  assign n19172 = pi16 ? n32 : n19171;
  assign n19173 = pi15 ? n18294 : n19172;
  assign n19174 = pi15 ? n19172 : n18814;
  assign n19175 = pi14 ? n19173 : n19174;
  assign n19176 = pi15 ? n19073 : n18821;
  assign n19177 = pi15 ? n18821 : n18594;
  assign n19178 = pi14 ? n19176 : n19177;
  assign n19179 = pi13 ? n19175 : n19178;
  assign n19180 = pi12 ? n19169 : n19179;
  assign n19181 = pi15 ? n18594 : n18439;
  assign n19182 = pi18 ? n1575 : ~n1676;
  assign n19183 = pi17 ? n32 : n19182;
  assign n19184 = pi16 ? n32 : n19183;
  assign n19185 = pi15 ? n17891 : n19184;
  assign n19186 = pi14 ? n19181 : n19185;
  assign n19187 = pi20 ? n175 : n1685;
  assign n19188 = pi19 ? n19187 : n18497;
  assign n19189 = pi18 ? n858 : n19188;
  assign n19190 = pi17 ? n32 : n19189;
  assign n19191 = pi20 ? n339 : n321;
  assign n19192 = pi19 ? n19191 : n247;
  assign n19193 = pi18 ? n19192 : n17118;
  assign n19194 = pi19 ? n11879 : n32;
  assign n19195 = pi18 ? n19194 : n1676;
  assign n19196 = pi17 ? n19193 : n19195;
  assign n19197 = pi16 ? n19190 : ~n19196;
  assign n19198 = pi15 ? n17891 : n19197;
  assign n19199 = pi18 ? n341 : ~n17118;
  assign n19200 = pi17 ? n32 : n19199;
  assign n19201 = pi16 ? n19200 : ~n1678;
  assign n19202 = pi19 ? n32 : n13939;
  assign n19203 = pi18 ? n209 : ~n19202;
  assign n19204 = pi17 ? n32 : n19203;
  assign n19205 = pi16 ? n19204 : ~n1683;
  assign n19206 = pi15 ? n19201 : n19205;
  assign n19207 = pi14 ? n19198 : n19206;
  assign n19208 = pi13 ? n19186 : n19207;
  assign n19209 = pi19 ? n32 : n13656;
  assign n19210 = pi18 ? n209 : ~n19209;
  assign n19211 = pi17 ? n32 : n19210;
  assign n19212 = pi16 ? n19211 : ~n1683;
  assign n19213 = pi16 ? n18994 : ~n1683;
  assign n19214 = pi15 ? n19212 : n19213;
  assign n19215 = pi18 ? n880 : n32;
  assign n19216 = pi17 ? n32 : n19215;
  assign n19217 = pi16 ? n32 : n19216;
  assign n19218 = pi20 ? n206 : ~n101;
  assign n19219 = pi19 ? n32 : n19218;
  assign n19220 = pi18 ? n19219 : n32;
  assign n19221 = pi17 ? n32 : n19220;
  assign n19222 = pi16 ? n32 : n19221;
  assign n19223 = pi15 ? n19217 : n19222;
  assign n19224 = pi14 ? n19214 : n19223;
  assign n19225 = pi15 ? n17637 : n17698;
  assign n19226 = pi14 ? n19225 : n17698;
  assign n19227 = pi13 ? n19224 : n19226;
  assign n19228 = pi12 ? n19208 : n19227;
  assign n19229 = pi11 ? n19180 : n19228;
  assign n19230 = pi10 ? n19162 : n19229;
  assign n19231 = pi09 ? n32 : n19230;
  assign n19232 = pi19 ? n3495 : n32;
  assign n19233 = pi18 ? n32 : n19232;
  assign n19234 = pi17 ? n32 : n19233;
  assign n19235 = pi16 ? n32 : n19234;
  assign n19236 = pi15 ? n32 : n19235;
  assign n19237 = pi19 ? n5597 : n32;
  assign n19238 = pi18 ? n32 : n19237;
  assign n19239 = pi17 ? n32 : n19238;
  assign n19240 = pi16 ? n32 : n19239;
  assign n19241 = pi15 ? n19240 : n19124;
  assign n19242 = pi14 ? n19236 : n19241;
  assign n19243 = pi13 ? n32 : n19242;
  assign n19244 = pi12 ? n32 : n19243;
  assign n19245 = pi19 ? n32 : n18789;
  assign n19246 = pi20 ? n339 : n314;
  assign n19247 = pi19 ? n19246 : ~n19116;
  assign n19248 = pi18 ? n19245 : ~n19247;
  assign n19249 = pi20 ? n17669 : ~n18129;
  assign n19250 = pi19 ? n19249 : ~n357;
  assign n19251 = pi18 ? n19250 : ~n19137;
  assign n19252 = pi17 ? n19248 : ~n19251;
  assign n19253 = pi16 ? n32 : n19252;
  assign n19254 = pi15 ? n19253 : n19145;
  assign n19255 = pi14 ? n19254 : n19147;
  assign n19256 = pi13 ? n19255 : n19157;
  assign n19257 = pi14 ? n18890 : n18531;
  assign n19258 = pi13 ? n32 : n19257;
  assign n19259 = pi12 ? n19256 : n19258;
  assign n19260 = pi11 ? n19244 : n19259;
  assign n19261 = pi14 ? n18661 : n32;
  assign n19262 = pi18 ? n32 : ~n814;
  assign n19263 = pi17 ? n32 : n19262;
  assign n19264 = pi16 ? n32 : n19263;
  assign n19265 = pi18 ? n32 : n441;
  assign n19266 = pi17 ? n32 : n19265;
  assign n19267 = pi16 ? n32 : n19266;
  assign n19268 = pi15 ? n19264 : n19267;
  assign n19269 = pi14 ? n32 : n19268;
  assign n19270 = pi13 ? n19261 : n19269;
  assign n19271 = pi15 ? n18688 : n19166;
  assign n19272 = pi15 ? n19166 : n19061;
  assign n19273 = pi14 ? n19271 : n19272;
  assign n19274 = pi15 ? n19073 : n18594;
  assign n19275 = pi14 ? n19073 : n19274;
  assign n19276 = pi13 ? n19273 : n19275;
  assign n19277 = pi12 ? n19270 : n19276;
  assign n19278 = pi15 ? n17903 : n17894;
  assign n19279 = pi14 ? n19181 : n19278;
  assign n19280 = pi20 ? n220 : ~n7939;
  assign n19281 = pi19 ? n19187 : n19280;
  assign n19282 = pi18 ? n858 : n19281;
  assign n19283 = pi17 ? n32 : n19282;
  assign n19284 = pi16 ? n19283 : ~n19196;
  assign n19285 = pi15 ? n17891 : n19284;
  assign n19286 = pi18 ? n341 : ~n463;
  assign n19287 = pi17 ? n32 : n19286;
  assign n19288 = pi16 ? n19287 : ~n1678;
  assign n19289 = pi15 ? n19288 : n19205;
  assign n19290 = pi14 ? n19285 : n19289;
  assign n19291 = pi13 ? n19279 : n19290;
  assign n19292 = pi18 ? n4407 : n32;
  assign n19293 = pi17 ? n32 : n19292;
  assign n19294 = pi16 ? n32 : n19293;
  assign n19295 = pi15 ? n19217 : n19294;
  assign n19296 = pi14 ? n19214 : n19295;
  assign n19297 = pi15 ? n17910 : n17822;
  assign n19298 = pi14 ? n19297 : n17698;
  assign n19299 = pi13 ? n19296 : n19298;
  assign n19300 = pi12 ? n19291 : n19299;
  assign n19301 = pi11 ? n19277 : n19300;
  assign n19302 = pi10 ? n19260 : n19301;
  assign n19303 = pi09 ? n32 : n19302;
  assign n19304 = pi08 ? n19231 : n19303;
  assign n19305 = pi07 ? n19112 : n19304;
  assign n19306 = pi20 ? n357 : ~n207;
  assign n19307 = pi19 ? n311 : ~n19306;
  assign n19308 = pi18 ? n32 : n19307;
  assign n19309 = pi17 ? n32 : n19308;
  assign n19310 = pi17 ? n18482 : n2319;
  assign n19311 = pi16 ? n19309 : ~n19310;
  assign n19312 = pi15 ? n19235 : n19311;
  assign n19313 = pi14 ? n19236 : n19312;
  assign n19314 = pi13 ? n32 : n19313;
  assign n19315 = pi12 ? n32 : n19314;
  assign n19316 = pi19 ? n6622 : ~n207;
  assign n19317 = pi20 ? n17712 : n32;
  assign n19318 = pi19 ? n19317 : n32;
  assign n19319 = pi18 ? n19316 : n19318;
  assign n19320 = pi17 ? n13950 : n19319;
  assign n19321 = pi16 ? n32 : n19320;
  assign n19322 = pi18 ? n19316 : n19232;
  assign n19323 = pi17 ? n13950 : n19322;
  assign n19324 = pi16 ? n32 : n19323;
  assign n19325 = pi15 ? n19321 : n19324;
  assign n19326 = pi15 ? n19235 : n32;
  assign n19327 = pi14 ? n19325 : n19326;
  assign n19328 = pi13 ? n19327 : n32;
  assign n19329 = pi14 ? n18904 : n18657;
  assign n19330 = pi13 ? n32 : n19329;
  assign n19331 = pi12 ? n19328 : n19330;
  assign n19332 = pi11 ? n19315 : n19331;
  assign n19333 = pi15 ? n32 : n18535;
  assign n19334 = pi15 ? n18535 : n19264;
  assign n19335 = pi14 ? n19333 : n19334;
  assign n19336 = pi13 ? n19261 : n19335;
  assign n19337 = pi14 ? n18689 : n19166;
  assign n19338 = pi15 ? n19073 : n18814;
  assign n19339 = pi15 ? n18814 : n19172;
  assign n19340 = pi14 ? n19338 : n19339;
  assign n19341 = pi13 ? n19337 : n19340;
  assign n19342 = pi12 ? n19336 : n19341;
  assign n19343 = pi15 ? n19172 : n18297;
  assign n19344 = pi14 ? n19343 : n18440;
  assign n19345 = pi18 ? n341 : ~n4380;
  assign n19346 = pi17 ? n32 : n19345;
  assign n19347 = pi16 ? n19346 : ~n3356;
  assign n19348 = pi15 ? n18439 : n19347;
  assign n19349 = pi16 ? n1135 : ~n3356;
  assign n19350 = pi19 ? n32 : n9220;
  assign n19351 = pi18 ? n341 : ~n19350;
  assign n19352 = pi17 ? n32 : n19351;
  assign n19353 = pi16 ? n19352 : ~n1678;
  assign n19354 = pi15 ? n19349 : n19353;
  assign n19355 = pi14 ? n19348 : n19354;
  assign n19356 = pi13 ? n19344 : n19355;
  assign n19357 = pi18 ? n18710 : ~n222;
  assign n19358 = pi17 ? n32 : n19357;
  assign n19359 = pi16 ? n19358 : ~n1678;
  assign n19360 = pi17 ? n1500 : ~n1677;
  assign n19361 = pi16 ? n11695 : n19360;
  assign n19362 = pi15 ? n19359 : n19361;
  assign n19363 = pi20 ? n3523 : ~n623;
  assign n19364 = pi19 ? n32 : n19363;
  assign n19365 = pi18 ? n19364 : n32;
  assign n19366 = pi17 ? n32 : n19365;
  assign n19367 = pi16 ? n32 : n19366;
  assign n19368 = pi15 ? n18309 : n19367;
  assign n19369 = pi14 ? n19362 : n19368;
  assign n19370 = pi20 ? n32 : n16997;
  assign n19371 = pi19 ? n32 : n19370;
  assign n19372 = pi18 ? n19371 : n32;
  assign n19373 = pi17 ? n32 : n19372;
  assign n19374 = pi16 ? n32 : n19373;
  assign n19375 = pi15 ? n19374 : n17637;
  assign n19376 = pi14 ? n19375 : n17637;
  assign n19377 = pi13 ? n19369 : n19376;
  assign n19378 = pi12 ? n19356 : n19377;
  assign n19379 = pi11 ? n19342 : n19378;
  assign n19380 = pi10 ? n19332 : n19379;
  assign n19381 = pi09 ? n32 : n19380;
  assign n19382 = pi18 ? n32 : n19318;
  assign n19383 = pi17 ? n32 : n19382;
  assign n19384 = pi16 ? n32 : n19383;
  assign n19385 = pi15 ? n32 : n19384;
  assign n19386 = pi15 ? n19384 : n19311;
  assign n19387 = pi14 ? n19385 : n19386;
  assign n19388 = pi13 ? n32 : n19387;
  assign n19389 = pi12 ? n32 : n19388;
  assign n19390 = pi14 ? n165 : n18657;
  assign n19391 = pi13 ? n32 : n19390;
  assign n19392 = pi12 ? n19328 : n19391;
  assign n19393 = pi11 ? n19389 : n19392;
  assign n19394 = pi14 ? n18657 : n32;
  assign n19395 = pi15 ? n32 : n18531;
  assign n19396 = pi18 ? n32 : ~n1813;
  assign n19397 = pi17 ? n32 : n19396;
  assign n19398 = pi16 ? n32 : n19397;
  assign n19399 = pi15 ? n18531 : n19398;
  assign n19400 = pi14 ? n19395 : n19399;
  assign n19401 = pi13 ? n19394 : n19400;
  assign n19402 = pi14 ? n18535 : n19264;
  assign n19403 = pi18 ? n940 : ~n1942;
  assign n19404 = pi17 ? n32 : n19403;
  assign n19405 = pi16 ? n32 : n19404;
  assign n19406 = pi15 ? n19405 : n19061;
  assign n19407 = pi15 ? n19061 : n19172;
  assign n19408 = pi14 ? n19406 : n19407;
  assign n19409 = pi13 ? n19402 : n19408;
  assign n19410 = pi12 ? n19401 : n19409;
  assign n19411 = pi20 ? n3523 : n342;
  assign n19412 = pi19 ? n32 : n19411;
  assign n19413 = pi18 ? n19412 : n32;
  assign n19414 = pi17 ? n32 : n19413;
  assign n19415 = pi16 ? n32 : n19414;
  assign n19416 = pi15 ? n18309 : n19415;
  assign n19417 = pi14 ? n19362 : n19416;
  assign n19418 = pi15 ? n17903 : n17910;
  assign n19419 = pi14 ? n19418 : n17637;
  assign n19420 = pi13 ? n19417 : n19419;
  assign n19421 = pi12 ? n19356 : n19420;
  assign n19422 = pi11 ? n19410 : n19421;
  assign n19423 = pi10 ? n19393 : n19422;
  assign n19424 = pi09 ? n32 : n19423;
  assign n19425 = pi08 ? n19381 : n19424;
  assign n19426 = pi20 ? n501 : n314;
  assign n19427 = pi19 ? n975 : n19426;
  assign n19428 = pi18 ? n32 : n19427;
  assign n19429 = pi17 ? n32 : n19428;
  assign n19430 = pi16 ? n19429 : ~n1934;
  assign n19431 = pi17 ? n32 : n3296;
  assign n19432 = pi18 ? n18532 : n32;
  assign n19433 = pi17 ? n19432 : n1933;
  assign n19434 = pi16 ? n19431 : ~n19433;
  assign n19435 = pi15 ? n19430 : n19434;
  assign n19436 = pi14 ? n92 : n19435;
  assign n19437 = pi13 ? n32 : n19436;
  assign n19438 = pi12 ? n32 : n19437;
  assign n19439 = pi19 ? n334 : ~n339;
  assign n19440 = pi18 ? n19439 : n248;
  assign n19441 = pi17 ? n18082 : n19440;
  assign n19442 = pi16 ? n32 : n19441;
  assign n19443 = pi18 ? n19439 : n19318;
  assign n19444 = pi17 ? n18082 : n19443;
  assign n19445 = pi16 ? n32 : n19444;
  assign n19446 = pi15 ? n19442 : n19445;
  assign n19447 = pi15 ? n91 : n32;
  assign n19448 = pi14 ? n19446 : n19447;
  assign n19449 = pi13 ? n19448 : n32;
  assign n19450 = pi14 ? n19235 : n19030;
  assign n19451 = pi13 ? n32 : n19450;
  assign n19452 = pi12 ? n19449 : n19451;
  assign n19453 = pi11 ? n19438 : n19452;
  assign n19454 = pi14 ? n18890 : n32;
  assign n19455 = pi14 ? n18535 : n18531;
  assign n19456 = pi13 ? n19454 : n19455;
  assign n19457 = pi18 ? n940 : ~n814;
  assign n19458 = pi17 ? n32 : n19457;
  assign n19459 = pi16 ? n32 : n19458;
  assign n19460 = pi15 ? n19459 : n19061;
  assign n19461 = pi15 ? n19061 : n19166;
  assign n19462 = pi14 ? n19460 : n19461;
  assign n19463 = pi13 ? n19402 : n19462;
  assign n19464 = pi12 ? n19456 : n19463;
  assign n19465 = pi15 ? n19166 : n19172;
  assign n19466 = pi18 ? n1575 : ~n3350;
  assign n19467 = pi17 ? n32 : n19466;
  assign n19468 = pi16 ? n32 : n19467;
  assign n19469 = pi15 ? n19468 : n18594;
  assign n19470 = pi14 ? n19465 : n19469;
  assign n19471 = pi18 ? n209 : ~n936;
  assign n19472 = pi17 ? n32 : n19471;
  assign n19473 = pi17 ? n2008 : ~n3351;
  assign n19474 = pi16 ? n19472 : n19473;
  assign n19475 = pi15 ? n18594 : n19474;
  assign n19476 = pi16 ? n1135 : ~n3352;
  assign n19477 = pi18 ? n209 : ~n863;
  assign n19478 = pi17 ? n32 : n19477;
  assign n19479 = pi17 ? n2008 : ~n2123;
  assign n19480 = pi16 ? n19478 : n19479;
  assign n19481 = pi15 ? n19476 : n19480;
  assign n19482 = pi14 ? n19475 : n19481;
  assign n19483 = pi13 ? n19470 : n19482;
  assign n19484 = pi18 ? n940 : ~n209;
  assign n19485 = pi17 ? n32 : n19484;
  assign n19486 = pi16 ? n19485 : n5310;
  assign n19487 = pi17 ? n1500 : ~n2123;
  assign n19488 = pi16 ? n11695 : n19487;
  assign n19489 = pi15 ? n19486 : n19488;
  assign n19490 = pi18 ? n1249 : ~n618;
  assign n19491 = pi17 ? n32 : n19490;
  assign n19492 = pi16 ? n32 : n19491;
  assign n19493 = pi15 ? n19492 : n17891;
  assign n19494 = pi14 ? n19489 : n19493;
  assign n19495 = pi15 ? n17885 : n17910;
  assign n19496 = pi15 ? n17910 : n17637;
  assign n19497 = pi14 ? n19495 : n19496;
  assign n19498 = pi13 ? n19494 : n19497;
  assign n19499 = pi12 ? n19483 : n19498;
  assign n19500 = pi11 ? n19464 : n19499;
  assign n19501 = pi10 ? n19453 : n19500;
  assign n19502 = pi09 ? n32 : n19501;
  assign n19503 = pi16 ? n32 : n18561;
  assign n19504 = pi15 ? n32 : n19503;
  assign n19505 = pi20 ? n1076 : n2358;
  assign n19506 = pi19 ? n594 : n19505;
  assign n19507 = pi18 ? n32 : n19506;
  assign n19508 = pi17 ? n32 : n19507;
  assign n19509 = pi16 ? n19508 : ~n1934;
  assign n19510 = pi15 ? n19509 : n19434;
  assign n19511 = pi14 ? n19504 : n19510;
  assign n19512 = pi13 ? n32 : n19511;
  assign n19513 = pi12 ? n32 : n19512;
  assign n19514 = pi18 ? n19439 : n9170;
  assign n19515 = pi17 ? n18082 : n19514;
  assign n19516 = pi16 ? n32 : n19515;
  assign n19517 = pi18 ? n19439 : n88;
  assign n19518 = pi17 ? n18082 : n19517;
  assign n19519 = pi16 ? n32 : n19518;
  assign n19520 = pi15 ? n19516 : n19519;
  assign n19521 = pi14 ? n19520 : n19447;
  assign n19522 = pi13 ? n19521 : n32;
  assign n19523 = pi15 ? n165 : n19235;
  assign n19524 = pi14 ? n19326 : n19523;
  assign n19525 = pi13 ? n32 : n19524;
  assign n19526 = pi12 ? n19522 : n19525;
  assign n19527 = pi11 ? n19513 : n19526;
  assign n19528 = pi14 ? n165 : n32;
  assign n19529 = pi18 ? n32 : n6059;
  assign n19530 = pi17 ? n32 : n19529;
  assign n19531 = pi16 ? n32 : n19530;
  assign n19532 = pi13 ? n19528 : n19531;
  assign n19533 = pi14 ? n18531 : n19398;
  assign n19534 = pi18 ? n863 : ~n814;
  assign n19535 = pi17 ? n32 : n19534;
  assign n19536 = pi16 ? n32 : n19535;
  assign n19537 = pi15 ? n19459 : n19536;
  assign n19538 = pi15 ? n19536 : n19166;
  assign n19539 = pi14 ? n19537 : n19538;
  assign n19540 = pi13 ? n19533 : n19539;
  assign n19541 = pi12 ? n19532 : n19540;
  assign n19542 = pi18 ? n936 : ~n3350;
  assign n19543 = pi17 ? n32 : n19542;
  assign n19544 = pi16 ? n32 : n19543;
  assign n19545 = pi15 ? n19544 : n18594;
  assign n19546 = pi14 ? n19465 : n19545;
  assign n19547 = pi20 ? n274 : ~n18415;
  assign n19548 = pi19 ? n1817 : n19547;
  assign n19549 = pi18 ? n1819 : n19548;
  assign n19550 = pi17 ? n32 : n19549;
  assign n19551 = pi20 ? n6085 : n18073;
  assign n19552 = pi19 ? n19129 : n19551;
  assign n19553 = pi20 ? n206 : n313;
  assign n19554 = pi21 ? n313 : n309;
  assign n19555 = pi20 ? n18415 : ~n19554;
  assign n19556 = pi19 ? n19553 : n19555;
  assign n19557 = pi18 ? n19552 : ~n19556;
  assign n19558 = pi20 ? n13171 : ~n333;
  assign n19559 = pi20 ? n13171 : ~n2385;
  assign n19560 = pi19 ? n19558 : n19559;
  assign n19561 = pi18 ? n19560 : n3350;
  assign n19562 = pi17 ? n19557 : ~n19561;
  assign n19563 = pi16 ? n19550 : n19562;
  assign n19564 = pi15 ? n19563 : n19474;
  assign n19565 = pi14 ? n19564 : n19481;
  assign n19566 = pi13 ? n19546 : n19565;
  assign n19567 = pi15 ? n18972 : n17910;
  assign n19568 = pi14 ? n19567 : n19496;
  assign n19569 = pi13 ? n19494 : n19568;
  assign n19570 = pi12 ? n19566 : n19569;
  assign n19571 = pi11 ? n19541 : n19570;
  assign n19572 = pi10 ? n19527 : n19571;
  assign n19573 = pi09 ? n32 : n19572;
  assign n19574 = pi08 ? n19502 : n19573;
  assign n19575 = pi07 ? n19425 : n19574;
  assign n19576 = pi06 ? n19305 : n19575;
  assign n19577 = pi20 ? n3523 : ~n357;
  assign n19578 = pi19 ? n19577 : ~n32;
  assign n19579 = pi18 ? n19578 : ~n32;
  assign n19580 = pi17 ? n19579 : ~n2305;
  assign n19581 = pi16 ? n32 : n19580;
  assign n19582 = pi20 ? n32 : n17652;
  assign n19583 = pi20 ? n501 : n207;
  assign n19584 = pi19 ? n19582 : n19583;
  assign n19585 = pi20 ? n32 : ~n4279;
  assign n19586 = pi19 ? n19585 : ~n236;
  assign n19587 = pi18 ? n19584 : ~n19586;
  assign n19588 = pi19 ? n32 : n357;
  assign n19589 = pi18 ? n19588 : n2304;
  assign n19590 = pi17 ? n19587 : ~n19589;
  assign n19591 = pi16 ? n32 : n19590;
  assign n19592 = pi15 ? n19581 : n19591;
  assign n19593 = pi14 ? n19504 : n19592;
  assign n19594 = pi13 ? n32 : n19593;
  assign n19595 = pi12 ? n32 : n19594;
  assign n19596 = pi20 ? n1817 : n1076;
  assign n19597 = pi19 ? n32 : n19596;
  assign n19598 = pi20 ? n342 : n1611;
  assign n19599 = pi19 ? n6350 : n19598;
  assign n19600 = pi18 ? n19597 : n19599;
  assign n19601 = pi20 ? n2358 : n5854;
  assign n19602 = pi20 ? n7939 : n9491;
  assign n19603 = pi19 ? n19601 : ~n19602;
  assign n19604 = pi21 ? n32 : ~n7500;
  assign n19605 = pi20 ? n19604 : ~n32;
  assign n19606 = pi19 ? n19605 : ~n32;
  assign n19607 = pi18 ? n19603 : ~n19606;
  assign n19608 = pi17 ? n19600 : n19607;
  assign n19609 = pi16 ? n32 : n19608;
  assign n19610 = pi20 ? n9491 : n32;
  assign n19611 = pi19 ? n19610 : n6398;
  assign n19612 = pi20 ? n9491 : ~n32;
  assign n19613 = pi19 ? n19612 : ~n32;
  assign n19614 = pi18 ? n19611 : ~n19613;
  assign n19615 = pi17 ? n32 : n19614;
  assign n19616 = pi16 ? n32 : n19615;
  assign n19617 = pi15 ? n19609 : n19616;
  assign n19618 = pi15 ? n19503 : n32;
  assign n19619 = pi14 ? n19617 : n19618;
  assign n19620 = pi13 ? n19619 : n32;
  assign n19621 = pi15 ? n19384 : n19235;
  assign n19622 = pi14 ? n19621 : n19235;
  assign n19623 = pi13 ? n32 : n19622;
  assign n19624 = pi12 ? n19620 : n19623;
  assign n19625 = pi11 ? n19595 : n19624;
  assign n19626 = pi15 ? n32 : n19531;
  assign n19627 = pi14 ? n165 : n19626;
  assign n19628 = pi16 ? n32 : n18488;
  assign n19629 = pi19 ? n15962 : n32;
  assign n19630 = pi18 ? n32 : n19629;
  assign n19631 = pi17 ? n32 : n19630;
  assign n19632 = pi16 ? n32 : n19631;
  assign n19633 = pi15 ? n19628 : n19632;
  assign n19634 = pi14 ? n19531 : n19633;
  assign n19635 = pi13 ? n19627 : n19634;
  assign n19636 = pi18 ? n209 : ~n1813;
  assign n19637 = pi17 ? n32 : n19636;
  assign n19638 = pi16 ? n32 : n19637;
  assign n19639 = pi15 ? n19398 : n19638;
  assign n19640 = pi14 ? n19399 : n19639;
  assign n19641 = pi18 ? n684 : ~n1813;
  assign n19642 = pi17 ? n32 : n19641;
  assign n19643 = pi16 ? n32 : n19642;
  assign n19644 = pi15 ? n19643 : n19536;
  assign n19645 = pi14 ? n19644 : n19264;
  assign n19646 = pi13 ? n19640 : n19645;
  assign n19647 = pi12 ? n19635 : n19646;
  assign n19648 = pi14 ? n19166 : n19172;
  assign n19649 = pi17 ? n18482 : n2325;
  assign n19650 = pi16 ? n1214 : ~n19649;
  assign n19651 = pi18 ? n1395 : ~n32;
  assign n19652 = pi17 ? n32 : n19651;
  assign n19653 = pi16 ? n19652 : ~n2326;
  assign n19654 = pi19 ? n1885 : n32;
  assign n19655 = pi18 ? n19654 : n32;
  assign n19656 = pi17 ? n19655 : n3351;
  assign n19657 = pi16 ? n1214 : ~n19656;
  assign n19658 = pi15 ? n19653 : n19657;
  assign n19659 = pi14 ? n19650 : n19658;
  assign n19660 = pi13 ? n19648 : n19659;
  assign n19661 = pi18 ? n880 : ~n3350;
  assign n19662 = pi17 ? n32 : n19661;
  assign n19663 = pi16 ? n32 : n19662;
  assign n19664 = pi18 ? n209 : ~n3350;
  assign n19665 = pi17 ? n32 : n19664;
  assign n19666 = pi16 ? n32 : n19665;
  assign n19667 = pi15 ? n19663 : n19666;
  assign n19668 = pi15 ? n18008 : n18972;
  assign n19669 = pi14 ? n19667 : n19668;
  assign n19670 = pi15 ? n18972 : n17885;
  assign n19671 = pi15 ? n17885 : n17813;
  assign n19672 = pi14 ? n19670 : n19671;
  assign n19673 = pi13 ? n19669 : n19672;
  assign n19674 = pi12 ? n19660 : n19673;
  assign n19675 = pi11 ? n19647 : n19674;
  assign n19676 = pi10 ? n19625 : n19675;
  assign n19677 = pi09 ? n32 : n19676;
  assign n19678 = pi14 ? n117 : n19592;
  assign n19679 = pi13 ? n32 : n19678;
  assign n19680 = pi12 ? n32 : n19679;
  assign n19681 = pi15 ? n91 : n19384;
  assign n19682 = pi15 ? n19235 : n19384;
  assign n19683 = pi14 ? n19681 : n19682;
  assign n19684 = pi13 ? n32 : n19683;
  assign n19685 = pi12 ? n19620 : n19684;
  assign n19686 = pi11 ? n19680 : n19685;
  assign n19687 = pi14 ? n19235 : n19626;
  assign n19688 = pi19 ? n7693 : n32;
  assign n19689 = pi18 ? n32 : n19688;
  assign n19690 = pi17 ? n32 : n19689;
  assign n19691 = pi16 ? n32 : n19690;
  assign n19692 = pi18 ? n32 : ~n3336;
  assign n19693 = pi17 ? n32 : n19692;
  assign n19694 = pi16 ? n32 : n19693;
  assign n19695 = pi15 ? n19694 : n18904;
  assign n19696 = pi14 ? n19691 : n19695;
  assign n19697 = pi13 ? n19687 : n19696;
  assign n19698 = pi15 ? n19531 : n19628;
  assign n19699 = pi18 ? n209 : ~n350;
  assign n19700 = pi17 ? n32 : n19699;
  assign n19701 = pi16 ? n32 : n19700;
  assign n19702 = pi15 ? n19628 : n19701;
  assign n19703 = pi14 ? n19698 : n19702;
  assign n19704 = pi18 ? n863 : ~n1813;
  assign n19705 = pi17 ? n32 : n19704;
  assign n19706 = pi16 ? n32 : n19705;
  assign n19707 = pi15 ? n19643 : n19706;
  assign n19708 = pi14 ? n19707 : n19264;
  assign n19709 = pi13 ? n19703 : n19708;
  assign n19710 = pi12 ? n19697 : n19709;
  assign n19711 = pi16 ? n1214 : ~n2326;
  assign n19712 = pi15 ? n19711 : n19657;
  assign n19713 = pi14 ? n19650 : n19712;
  assign n19714 = pi13 ? n19648 : n19713;
  assign n19715 = pi18 ? n936 : ~n618;
  assign n19716 = pi17 ? n32 : n19715;
  assign n19717 = pi16 ? n32 : n19716;
  assign n19718 = pi15 ? n18008 : n19717;
  assign n19719 = pi14 ? n19667 : n19718;
  assign n19720 = pi15 ? n19717 : n17885;
  assign n19721 = pi14 ? n19720 : n19671;
  assign n19722 = pi13 ? n19719 : n19721;
  assign n19723 = pi12 ? n19714 : n19722;
  assign n19724 = pi11 ? n19710 : n19723;
  assign n19725 = pi10 ? n19686 : n19724;
  assign n19726 = pi09 ? n32 : n19725;
  assign n19727 = pi08 ? n19677 : n19726;
  assign n19728 = pi20 ? n207 : n6050;
  assign n19729 = pi19 ? n1265 : n19728;
  assign n19730 = pi18 ? n6356 : ~n19729;
  assign n19731 = pi21 ? n405 : n313;
  assign n19732 = pi20 ? n32 : n19731;
  assign n19733 = pi20 ? n6050 : n1324;
  assign n19734 = pi19 ? n19732 : ~n19733;
  assign n19735 = pi18 ? n19734 : n430;
  assign n19736 = pi17 ? n19730 : ~n19735;
  assign n19737 = pi16 ? n32 : n19736;
  assign n19738 = pi20 ? n310 : ~n439;
  assign n19739 = pi19 ? n19738 : ~n594;
  assign n19740 = pi19 ? n10394 : ~n32;
  assign n19741 = pi18 ? n19739 : n19740;
  assign n19742 = pi17 ? n19170 : ~n19741;
  assign n19743 = pi16 ? n32 : n19742;
  assign n19744 = pi15 ? n19737 : n19743;
  assign n19745 = pi14 ? n117 : n19744;
  assign n19746 = pi13 ? n32 : n19745;
  assign n19747 = pi12 ? n32 : n19746;
  assign n19748 = pi19 ? n462 : n594;
  assign n19749 = pi20 ? n1385 : n32;
  assign n19750 = pi19 ? n19749 : n32;
  assign n19751 = pi18 ? n19748 : n19750;
  assign n19752 = pi17 ? n32 : n19751;
  assign n19753 = pi16 ? n32 : n19752;
  assign n19754 = pi15 ? n19753 : n180;
  assign n19755 = pi15 ? n116 : n32;
  assign n19756 = pi14 ? n19754 : n19755;
  assign n19757 = pi13 ? n19756 : n32;
  assign n19758 = pi15 ? n19503 : n91;
  assign n19759 = pi14 ? n19758 : n19384;
  assign n19760 = pi13 ? n32 : n19759;
  assign n19761 = pi12 ? n19757 : n19760;
  assign n19762 = pi11 ? n19747 : n19761;
  assign n19763 = pi15 ? n32 : n19691;
  assign n19764 = pi14 ? n19240 : n19763;
  assign n19765 = pi13 ? n19764 : n19691;
  assign n19766 = pi15 ? n19531 : n19701;
  assign n19767 = pi14 ? n19698 : n19766;
  assign n19768 = pi15 ? n19643 : n19398;
  assign n19769 = pi14 ? n19768 : n19398;
  assign n19770 = pi13 ? n19767 : n19769;
  assign n19771 = pi12 ? n19765 : n19770;
  assign n19772 = pi14 ? n19264 : n19166;
  assign n19773 = pi20 ? n14286 : n32;
  assign n19774 = pi19 ? n19773 : n32;
  assign n19775 = pi18 ? n19774 : n32;
  assign n19776 = pi17 ? n19775 : n1943;
  assign n19777 = pi16 ? n1135 : ~n19776;
  assign n19778 = pi16 ? n1233 : ~n1944;
  assign n19779 = pi18 ? n19750 : n32;
  assign n19780 = pi17 ? n19779 : n2325;
  assign n19781 = pi16 ? n19652 : ~n19780;
  assign n19782 = pi15 ? n19778 : n19781;
  assign n19783 = pi14 ? n19777 : n19782;
  assign n19784 = pi13 ? n19772 : n19783;
  assign n19785 = pi18 ? n880 : ~n237;
  assign n19786 = pi17 ? n32 : n19785;
  assign n19787 = pi16 ? n32 : n19786;
  assign n19788 = pi15 ? n19787 : n18142;
  assign n19789 = pi14 ? n19788 : n18008;
  assign n19790 = pi14 ? n19668 : n17885;
  assign n19791 = pi13 ? n19789 : n19790;
  assign n19792 = pi12 ? n19784 : n19791;
  assign n19793 = pi11 ? n19771 : n19792;
  assign n19794 = pi10 ? n19762 : n19793;
  assign n19795 = pi09 ? n32 : n19794;
  assign n19796 = pi14 ? n32 : n19744;
  assign n19797 = pi13 ? n32 : n19796;
  assign n19798 = pi12 ? n32 : n19797;
  assign n19799 = pi15 ? n19753 : n116;
  assign n19800 = pi14 ? n19799 : n19755;
  assign n19801 = pi13 ? n19800 : n32;
  assign n19802 = pi15 ? n156 : n19503;
  assign n19803 = pi18 ? n32 : n248;
  assign n19804 = pi17 ? n32 : n19803;
  assign n19805 = pi16 ? n32 : n19804;
  assign n19806 = pi15 ? n19384 : n19805;
  assign n19807 = pi14 ? n19802 : n19806;
  assign n19808 = pi13 ? n32 : n19807;
  assign n19809 = pi12 ? n19801 : n19808;
  assign n19810 = pi11 ? n19798 : n19809;
  assign n19811 = pi19 ? n9724 : n32;
  assign n19812 = pi18 ? n32 : n19811;
  assign n19813 = pi17 ? n32 : n19812;
  assign n19814 = pi16 ? n32 : n19813;
  assign n19815 = pi15 ? n32 : n19814;
  assign n19816 = pi14 ? n91 : n19815;
  assign n19817 = pi13 ? n19816 : n19814;
  assign n19818 = pi15 ? n19691 : n19694;
  assign n19819 = pi18 ? n209 : ~n3336;
  assign n19820 = pi17 ? n32 : n19819;
  assign n19821 = pi16 ? n32 : n19820;
  assign n19822 = pi15 ? n19691 : n19821;
  assign n19823 = pi14 ? n19818 : n19822;
  assign n19824 = pi18 ? n684 : ~n350;
  assign n19825 = pi17 ? n32 : n19824;
  assign n19826 = pi16 ? n32 : n19825;
  assign n19827 = pi15 ? n19826 : n19628;
  assign n19828 = pi14 ? n19827 : n19398;
  assign n19829 = pi13 ? n19823 : n19828;
  assign n19830 = pi12 ? n19817 : n19829;
  assign n19831 = pi16 ? n1135 : ~n1944;
  assign n19832 = pi16 ? n1214 : ~n19780;
  assign n19833 = pi15 ? n19831 : n19832;
  assign n19834 = pi14 ? n19777 : n19833;
  assign n19835 = pi13 ? n19772 : n19834;
  assign n19836 = pi15 ? n19787 : n18294;
  assign n19837 = pi14 ? n19836 : n18297;
  assign n19838 = pi15 ? n18008 : n19184;
  assign n19839 = pi14 ? n19838 : n17876;
  assign n19840 = pi13 ? n19837 : n19839;
  assign n19841 = pi12 ? n19835 : n19840;
  assign n19842 = pi11 ? n19830 : n19841;
  assign n19843 = pi10 ? n19810 : n19842;
  assign n19844 = pi09 ? n32 : n19843;
  assign n19845 = pi08 ? n19795 : n19844;
  assign n19846 = pi07 ? n19727 : n19845;
  assign n19847 = pi20 ? n17654 : n32;
  assign n19848 = pi19 ? n19847 : n32;
  assign n19849 = pi18 ? n32 : n19848;
  assign n19850 = pi17 ? n32 : n19849;
  assign n19851 = pi16 ? n32 : n19850;
  assign n19852 = pi20 ? n18158 : n32;
  assign n19853 = pi19 ? n19852 : n32;
  assign n19854 = pi18 ? n32 : n19853;
  assign n19855 = pi17 ? n32 : n19854;
  assign n19856 = pi16 ? n32 : n19855;
  assign n19857 = pi15 ? n19851 : n19856;
  assign n19858 = pi14 ? n32 : n19857;
  assign n19859 = pi13 ? n32 : n19858;
  assign n19860 = pi12 ? n32 : n19859;
  assign n19861 = pi15 ? n19856 : n180;
  assign n19862 = pi15 ? n180 : n32;
  assign n19863 = pi14 ? n19861 : n19862;
  assign n19864 = pi13 ? n19863 : n32;
  assign n19865 = pi19 ? n7881 : n32;
  assign n19866 = pi18 ? n32 : n19865;
  assign n19867 = pi17 ? n32 : n19866;
  assign n19868 = pi16 ? n32 : n19867;
  assign n19869 = pi15 ? n32 : n19868;
  assign n19870 = pi14 ? n19869 : n117;
  assign n19871 = pi19 ? n16651 : n32;
  assign n19872 = pi18 ? n32 : n19871;
  assign n19873 = pi17 ? n32 : n19872;
  assign n19874 = pi16 ? n32 : n19873;
  assign n19875 = pi15 ? n19874 : n19805;
  assign n19876 = pi14 ? n19875 : n19758;
  assign n19877 = pi13 ? n19870 : n19876;
  assign n19878 = pi12 ? n19864 : n19877;
  assign n19879 = pi11 ? n19860 : n19878;
  assign n19880 = pi15 ? n19235 : n19814;
  assign n19881 = pi14 ? n19447 : n19880;
  assign n19882 = pi13 ? n19881 : n19814;
  assign n19883 = pi18 ? n4380 : n19688;
  assign n19884 = pi17 ? n32 : n19883;
  assign n19885 = pi16 ? n32 : n19884;
  assign n19886 = pi18 ? n32 : n6145;
  assign n19887 = pi18 ? n496 : ~n350;
  assign n19888 = pi17 ? n19886 : n19887;
  assign n19889 = pi16 ? n32 : n19888;
  assign n19890 = pi15 ? n19885 : n19889;
  assign n19891 = pi14 ? n19691 : n19890;
  assign n19892 = pi20 ? n14159 : n32;
  assign n19893 = pi19 ? n19892 : n32;
  assign n19894 = pi18 ? n32 : n19893;
  assign n19895 = pi17 ? n32 : n19894;
  assign n19896 = pi16 ? n32 : n19895;
  assign n19897 = pi15 ? n19628 : n19896;
  assign n19898 = pi14 ? n19628 : n19897;
  assign n19899 = pi13 ? n19891 : n19898;
  assign n19900 = pi12 ? n19882 : n19899;
  assign n19901 = pi15 ? n19398 : n19706;
  assign n19902 = pi15 ? n19264 : n18535;
  assign n19903 = pi14 ? n19901 : n19902;
  assign n19904 = pi18 ? n13945 : n32;
  assign n19905 = pi17 ? n19904 : n2136;
  assign n19906 = pi16 ? n1135 : ~n19905;
  assign n19907 = pi18 ? n5009 : n32;
  assign n19908 = pi17 ? n19907 : n1943;
  assign n19909 = pi16 ? n1471 : ~n19908;
  assign n19910 = pi15 ? n19778 : n19909;
  assign n19911 = pi14 ? n19906 : n19910;
  assign n19912 = pi13 ? n19903 : n19911;
  assign n19913 = pi15 ? n18142 : n18297;
  assign n19914 = pi14 ? n18694 : n19913;
  assign n19915 = pi15 ? n18008 : n17894;
  assign n19916 = pi14 ? n19915 : n17894;
  assign n19917 = pi13 ? n19914 : n19916;
  assign n19918 = pi12 ? n19912 : n19917;
  assign n19919 = pi11 ? n19900 : n19918;
  assign n19920 = pi10 ? n19879 : n19919;
  assign n19921 = pi09 ? n32 : n19920;
  assign n19922 = pi15 ? n19856 : n72;
  assign n19923 = pi14 ? n19922 : n19862;
  assign n19924 = pi13 ? n19923 : n32;
  assign n19925 = pi15 ? n32 : n19805;
  assign n19926 = pi14 ? n19925 : n32;
  assign n19927 = pi15 ? n116 : n19805;
  assign n19928 = pi14 ? n19927 : n156;
  assign n19929 = pi13 ? n19926 : n19928;
  assign n19930 = pi12 ? n19924 : n19929;
  assign n19931 = pi11 ? n19860 : n19930;
  assign n19932 = pi15 ? n156 : n32;
  assign n19933 = pi19 ? n7468 : n32;
  assign n19934 = pi18 ? n32 : n19933;
  assign n19935 = pi17 ? n32 : n19934;
  assign n19936 = pi16 ? n32 : n19935;
  assign n19937 = pi15 ? n19384 : n19936;
  assign n19938 = pi14 ? n19932 : n19937;
  assign n19939 = pi13 ? n19938 : n19936;
  assign n19940 = pi18 ? n4380 : n19811;
  assign n19941 = pi17 ? n32 : n19940;
  assign n19942 = pi16 ? n32 : n19941;
  assign n19943 = pi18 ? n496 : ~n3336;
  assign n19944 = pi17 ? n19886 : n19943;
  assign n19945 = pi16 ? n32 : n19944;
  assign n19946 = pi15 ? n19942 : n19945;
  assign n19947 = pi14 ? n19814 : n19946;
  assign n19948 = pi15 ? n19694 : n19628;
  assign n19949 = pi14 ? n19948 : n19897;
  assign n19950 = pi13 ? n19947 : n19949;
  assign n19951 = pi12 ? n19939 : n19950;
  assign n19952 = pi15 ? n19831 : n19909;
  assign n19953 = pi14 ? n19906 : n19952;
  assign n19954 = pi13 ? n19903 : n19953;
  assign n19955 = pi15 ? n18428 : n18294;
  assign n19956 = pi15 ? n18294 : n18297;
  assign n19957 = pi14 ? n19955 : n19956;
  assign n19958 = pi15 ? n18297 : n18008;
  assign n19959 = pi14 ? n19958 : n18008;
  assign n19960 = pi13 ? n19957 : n19959;
  assign n19961 = pi12 ? n19954 : n19960;
  assign n19962 = pi11 ? n19951 : n19961;
  assign n19963 = pi10 ? n19931 : n19962;
  assign n19964 = pi09 ? n32 : n19963;
  assign n19965 = pi08 ? n19921 : n19964;
  assign n19966 = pi19 ? n16969 : n32;
  assign n19967 = pi18 ? n32 : n19966;
  assign n19968 = pi17 ? n32 : n19967;
  assign n19969 = pi16 ? n32 : n19968;
  assign n19970 = pi15 ? n32 : n19969;
  assign n19971 = pi17 ? n32 : n18395;
  assign n19972 = pi16 ? n32 : n19971;
  assign n19973 = pi14 ? n19970 : n19972;
  assign n19974 = pi13 ? n32 : n19973;
  assign n19975 = pi12 ? n32 : n19974;
  assign n19976 = pi15 ? n19972 : n19969;
  assign n19977 = pi15 ? n19969 : n32;
  assign n19978 = pi14 ? n19976 : n19977;
  assign n19979 = pi13 ? n19978 : n32;
  assign n19980 = pi15 ? n180 : n19805;
  assign n19981 = pi14 ? n19980 : n180;
  assign n19982 = pi15 ? n180 : n19868;
  assign n19983 = pi15 ? n19868 : n19805;
  assign n19984 = pi14 ? n19982 : n19983;
  assign n19985 = pi13 ? n19981 : n19984;
  assign n19986 = pi12 ? n19979 : n19985;
  assign n19987 = pi11 ? n19975 : n19986;
  assign n19988 = pi18 ? n463 : n19933;
  assign n19989 = pi17 ? n32 : n19988;
  assign n19990 = pi16 ? n32 : n19989;
  assign n19991 = pi15 ? n19990 : n19936;
  assign n19992 = pi14 ? n19932 : n19991;
  assign n19993 = pi19 ? n7853 : n32;
  assign n19994 = pi18 ? n32 : n19993;
  assign n19995 = pi17 ? n32 : n19994;
  assign n19996 = pi16 ? n32 : n19995;
  assign n19997 = pi18 ? n32 : ~n2318;
  assign n19998 = pi17 ? n32 : n19997;
  assign n19999 = pi16 ? n32 : n19998;
  assign n20000 = pi15 ? n19996 : n19999;
  assign n20001 = pi14 ? n19936 : n20000;
  assign n20002 = pi13 ? n19992 : n20001;
  assign n20003 = pi18 ? n17118 : n19811;
  assign n20004 = pi17 ? n32 : n20003;
  assign n20005 = pi16 ? n32 : n20004;
  assign n20006 = pi20 ? n32 : ~n206;
  assign n20007 = pi19 ? n32 : n20006;
  assign n20008 = pi18 ? n20007 : n19811;
  assign n20009 = pi17 ? n32 : n20008;
  assign n20010 = pi16 ? n32 : n20009;
  assign n20011 = pi18 ? n32 : n5667;
  assign n20012 = pi17 ? n20011 : n19943;
  assign n20013 = pi16 ? n32 : n20012;
  assign n20014 = pi15 ? n20010 : n20013;
  assign n20015 = pi14 ? n20005 : n20014;
  assign n20016 = pi15 ? n19628 : n19531;
  assign n20017 = pi14 ? n19694 : n20016;
  assign n20018 = pi13 ? n20015 : n20017;
  assign n20019 = pi12 ? n20002 : n20018;
  assign n20020 = pi19 ? n1464 : n32;
  assign n20021 = pi18 ? n32 : n20020;
  assign n20022 = pi20 ? n11048 : ~n32;
  assign n20023 = pi19 ? n20022 : ~n32;
  assign n20024 = pi18 ? n32 : ~n20023;
  assign n20025 = pi17 ? n20021 : n20024;
  assign n20026 = pi16 ? n32 : n20025;
  assign n20027 = pi17 ? n20021 : n18529;
  assign n20028 = pi16 ? n32 : n20027;
  assign n20029 = pi15 ? n20026 : n20028;
  assign n20030 = pi14 ? n19628 : n20029;
  assign n20031 = pi18 ? n9865 : n32;
  assign n20032 = pi17 ? n20031 : n1814;
  assign n20033 = pi16 ? n1214 : ~n20032;
  assign n20034 = pi16 ? n1135 : ~n2137;
  assign n20035 = pi17 ? n19907 : n2136;
  assign n20036 = pi16 ? n1471 : ~n20035;
  assign n20037 = pi15 ? n20034 : n20036;
  assign n20038 = pi14 ? n20033 : n20037;
  assign n20039 = pi13 ? n20030 : n20038;
  assign n20040 = pi14 ? n57 : n42;
  assign n20041 = pi15 ? n41 : n18142;
  assign n20042 = pi14 ? n20041 : n18142;
  assign n20043 = pi13 ? n20040 : n20042;
  assign n20044 = pi12 ? n20039 : n20043;
  assign n20045 = pi11 ? n20019 : n20044;
  assign n20046 = pi10 ? n19987 : n20045;
  assign n20047 = pi09 ? n32 : n20046;
  assign n20048 = pi16 ? n32 : n18083;
  assign n20049 = pi15 ? n32 : n20048;
  assign n20050 = pi14 ? n20049 : n20048;
  assign n20051 = pi13 ? n32 : n20050;
  assign n20052 = pi12 ? n32 : n20051;
  assign n20053 = pi15 ? n20048 : n19969;
  assign n20054 = pi14 ? n20053 : n19977;
  assign n20055 = pi13 ? n20054 : n32;
  assign n20056 = pi14 ? n19980 : n19862;
  assign n20057 = pi15 ? n72 : n19868;
  assign n20058 = pi14 ? n20057 : n19868;
  assign n20059 = pi13 ? n20056 : n20058;
  assign n20060 = pi12 ? n20055 : n20059;
  assign n20061 = pi11 ? n20052 : n20060;
  assign n20062 = pi18 ? n463 : n4689;
  assign n20063 = pi17 ? n32 : n20062;
  assign n20064 = pi16 ? n32 : n20063;
  assign n20065 = pi18 ? n32 : n4689;
  assign n20066 = pi17 ? n32 : n20065;
  assign n20067 = pi16 ? n32 : n20066;
  assign n20068 = pi15 ? n20064 : n20067;
  assign n20069 = pi14 ? n19755 : n20068;
  assign n20070 = pi18 ? n32 : ~n344;
  assign n20071 = pi17 ? n32 : n20070;
  assign n20072 = pi16 ? n32 : n20071;
  assign n20073 = pi15 ? n19805 : n20072;
  assign n20074 = pi14 ? n20067 : n20073;
  assign n20075 = pi13 ? n20069 : n20074;
  assign n20076 = pi18 ? n17118 : n19933;
  assign n20077 = pi17 ? n32 : n20076;
  assign n20078 = pi16 ? n32 : n20077;
  assign n20079 = pi18 ? n20007 : n19933;
  assign n20080 = pi17 ? n32 : n20079;
  assign n20081 = pi16 ? n32 : n20080;
  assign n20082 = pi18 ? n496 : ~n1548;
  assign n20083 = pi17 ? n20011 : n20082;
  assign n20084 = pi16 ? n32 : n20083;
  assign n20085 = pi15 ? n20081 : n20084;
  assign n20086 = pi14 ? n20078 : n20085;
  assign n20087 = pi18 ? n32 : ~n1548;
  assign n20088 = pi17 ? n32 : n20087;
  assign n20089 = pi16 ? n32 : n20088;
  assign n20090 = pi15 ? n20089 : n19694;
  assign n20091 = pi15 ? n19694 : n19691;
  assign n20092 = pi14 ? n20090 : n20091;
  assign n20093 = pi13 ? n20086 : n20092;
  assign n20094 = pi12 ? n20075 : n20093;
  assign n20095 = pi18 ? n32 : ~n1353;
  assign n20096 = pi17 ? n20021 : n20095;
  assign n20097 = pi16 ? n32 : n20096;
  assign n20098 = pi17 ? n20021 : n19529;
  assign n20099 = pi16 ? n32 : n20098;
  assign n20100 = pi15 ? n20097 : n20099;
  assign n20101 = pi14 ? n19694 : n20100;
  assign n20102 = pi17 ? n20031 : n1807;
  assign n20103 = pi16 ? n1214 : ~n20102;
  assign n20104 = pi16 ? n1135 : ~n1815;
  assign n20105 = pi17 ? n19907 : n1814;
  assign n20106 = pi16 ? n1471 : ~n20105;
  assign n20107 = pi15 ? n20104 : n20106;
  assign n20108 = pi14 ? n20103 : n20107;
  assign n20109 = pi13 ? n20101 : n20108;
  assign n20110 = pi15 ? n18535 : n57;
  assign n20111 = pi15 ? n57 : n18294;
  assign n20112 = pi14 ? n20110 : n20111;
  assign n20113 = pi14 ? n18435 : n18142;
  assign n20114 = pi13 ? n20112 : n20113;
  assign n20115 = pi12 ? n20109 : n20114;
  assign n20116 = pi11 ? n20094 : n20115;
  assign n20117 = pi10 ? n20061 : n20116;
  assign n20118 = pi09 ? n32 : n20117;
  assign n20119 = pi08 ? n20047 : n20118;
  assign n20120 = pi07 ? n19965 : n20119;
  assign n20121 = pi06 ? n19846 : n20120;
  assign n20122 = pi05 ? n19576 : n20121;
  assign n20123 = pi14 ? n20049 : n13684;
  assign n20124 = pi13 ? n32 : n20123;
  assign n20125 = pi12 ? n32 : n20124;
  assign n20126 = pi15 ? n13684 : n20048;
  assign n20127 = pi15 ? n20048 : n32;
  assign n20128 = pi14 ? n20126 : n20127;
  assign n20129 = pi13 ? n20128 : n32;
  assign n20130 = pi22 ? n34 : ~n34;
  assign n20131 = pi21 ? n32 : n20130;
  assign n20132 = pi20 ? n20131 : n32;
  assign n20133 = pi19 ? n20132 : n32;
  assign n20134 = pi18 ? n32 : n20133;
  assign n20135 = pi17 ? n32 : n20134;
  assign n20136 = pi16 ? n32 : n20135;
  assign n20137 = pi15 ? n32 : n20136;
  assign n20138 = pi14 ? n32 : n20137;
  assign n20139 = pi15 ? n13392 : n180;
  assign n20140 = pi15 ? n180 : n116;
  assign n20141 = pi14 ? n20139 : n20140;
  assign n20142 = pi13 ? n20138 : n20141;
  assign n20143 = pi12 ? n20129 : n20142;
  assign n20144 = pi11 ? n20125 : n20143;
  assign n20145 = pi18 ? n17819 : n248;
  assign n20146 = pi17 ? n32 : n20145;
  assign n20147 = pi16 ? n32 : n20146;
  assign n20148 = pi15 ? n116 : n20147;
  assign n20149 = pi18 ? n684 : ~n344;
  assign n20150 = pi17 ? n32 : n20149;
  assign n20151 = pi16 ? n32 : n20150;
  assign n20152 = pi15 ? n20151 : n20067;
  assign n20153 = pi14 ? n20148 : n20152;
  assign n20154 = pi13 ? n20153 : n20067;
  assign n20155 = pi18 ? n4380 : n19933;
  assign n20156 = pi17 ? n32 : n20155;
  assign n20157 = pi16 ? n32 : n20156;
  assign n20158 = pi17 ? n16103 : n20155;
  assign n20159 = pi16 ? n32 : n20158;
  assign n20160 = pi15 ? n20157 : n20159;
  assign n20161 = pi18 ? n4380 : n19318;
  assign n20162 = pi17 ? n32 : n20161;
  assign n20163 = pi16 ? n32 : n20162;
  assign n20164 = pi19 ? n32 : ~n349;
  assign n20165 = pi18 ? n32 : n20164;
  assign n20166 = pi19 ? n32 : n5741;
  assign n20167 = pi18 ? n20166 : ~n289;
  assign n20168 = pi17 ? n20165 : n20167;
  assign n20169 = pi16 ? n32 : n20168;
  assign n20170 = pi15 ? n20163 : n20169;
  assign n20171 = pi14 ? n20160 : n20170;
  assign n20172 = pi19 ? n32 : ~n236;
  assign n20173 = pi18 ? n32 : n20172;
  assign n20174 = pi17 ? n20173 : n20087;
  assign n20175 = pi16 ? n32 : n20174;
  assign n20176 = pi15 ? n19235 : n20175;
  assign n20177 = pi14 ? n19235 : n20176;
  assign n20178 = pi13 ? n20171 : n20177;
  assign n20179 = pi12 ? n20154 : n20178;
  assign n20180 = pi17 ? n20173 : n19812;
  assign n20181 = pi16 ? n32 : n20180;
  assign n20182 = pi19 ? n507 : ~n6988;
  assign n20183 = pi18 ? n32 : n20182;
  assign n20184 = pi18 ? n19350 : ~n1548;
  assign n20185 = pi17 ? n20183 : n20184;
  assign n20186 = pi16 ? n32 : n20185;
  assign n20187 = pi15 ? n20181 : n20186;
  assign n20188 = pi18 ? n18532 : n323;
  assign n20189 = pi19 ? n6307 : ~n11879;
  assign n20190 = pi18 ? n20189 : ~n3336;
  assign n20191 = pi17 ? n20188 : n20190;
  assign n20192 = pi16 ? n32 : n20191;
  assign n20193 = pi19 ? n32 : ~n4342;
  assign n20194 = pi19 ? n9368 : ~n32;
  assign n20195 = pi18 ? n20193 : n20194;
  assign n20196 = pi17 ? n10245 : n20195;
  assign n20197 = pi16 ? n32 : ~n20196;
  assign n20198 = pi15 ? n20192 : n20197;
  assign n20199 = pi14 ? n20187 : n20198;
  assign n20200 = pi18 ? n6145 : n32;
  assign n20201 = pi17 ? n20200 : n3337;
  assign n20202 = pi16 ? n1214 : ~n20201;
  assign n20203 = pi18 ? n32 : ~n19688;
  assign n20204 = pi17 ? n20200 : n20203;
  assign n20205 = pi16 ? n1214 : ~n20204;
  assign n20206 = pi15 ? n20202 : n20205;
  assign n20207 = pi18 ? n18710 : ~n32;
  assign n20208 = pi17 ? n32 : n20207;
  assign n20209 = pi18 ? n6145 : n863;
  assign n20210 = pi18 ? n863 : n350;
  assign n20211 = pi17 ? n20209 : n20210;
  assign n20212 = pi16 ? n20208 : ~n20211;
  assign n20213 = pi15 ? n20212 : n18531;
  assign n20214 = pi14 ? n20206 : n20213;
  assign n20215 = pi13 ? n20199 : n20214;
  assign n20216 = pi15 ? n18531 : n18535;
  assign n20217 = pi14 ? n20216 : n20110;
  assign n20218 = pi14 ? n18694 : n18294;
  assign n20219 = pi13 ? n20217 : n20218;
  assign n20220 = pi12 ? n20215 : n20219;
  assign n20221 = pi11 ? n20179 : n20220;
  assign n20222 = pi10 ? n20144 : n20221;
  assign n20223 = pi09 ? n32 : n20222;
  assign n20224 = pi15 ? n32 : n13684;
  assign n20225 = pi14 ? n20224 : n13684;
  assign n20226 = pi13 ? n32 : n20225;
  assign n20227 = pi12 ? n32 : n20226;
  assign n20228 = pi14 ? n20126 : n107;
  assign n20229 = pi13 ? n20228 : n32;
  assign n20230 = pi15 ? n32 : n13392;
  assign n20231 = pi14 ? n32 : n20230;
  assign n20232 = pi15 ? n13392 : n72;
  assign n20233 = pi19 ? n16998 : n32;
  assign n20234 = pi18 ? n32 : n20233;
  assign n20235 = pi17 ? n32 : n20234;
  assign n20236 = pi16 ? n32 : n20235;
  assign n20237 = pi15 ? n20236 : n72;
  assign n20238 = pi14 ? n20232 : n20237;
  assign n20239 = pi13 ? n20231 : n20238;
  assign n20240 = pi12 ? n20229 : n20239;
  assign n20241 = pi11 ? n20227 : n20240;
  assign n20242 = pi18 ? n17819 : n19865;
  assign n20243 = pi17 ? n32 : n20242;
  assign n20244 = pi16 ? n32 : n20243;
  assign n20245 = pi15 ? n32 : n20244;
  assign n20246 = pi18 ? n684 : ~n2304;
  assign n20247 = pi17 ? n32 : n20246;
  assign n20248 = pi16 ? n32 : n20247;
  assign n20249 = pi19 ? n7443 : n32;
  assign n20250 = pi18 ? n32 : n20249;
  assign n20251 = pi17 ? n32 : n20250;
  assign n20252 = pi16 ? n32 : n20251;
  assign n20253 = pi15 ? n20248 : n20252;
  assign n20254 = pi14 ? n20245 : n20253;
  assign n20255 = pi13 ? n20254 : n20252;
  assign n20256 = pi18 ? n4380 : n4689;
  assign n20257 = pi17 ? n32 : n20256;
  assign n20258 = pi16 ? n32 : n20257;
  assign n20259 = pi17 ? n16103 : n20256;
  assign n20260 = pi16 ? n32 : n20259;
  assign n20261 = pi15 ? n20258 : n20260;
  assign n20262 = pi18 ? n4380 : n248;
  assign n20263 = pi17 ? n32 : n20262;
  assign n20264 = pi16 ? n32 : n20263;
  assign n20265 = pi21 ? n206 : n242;
  assign n20266 = pi20 ? n20265 : ~n32;
  assign n20267 = pi19 ? n20266 : ~n32;
  assign n20268 = pi18 ? n20166 : ~n20267;
  assign n20269 = pi17 ? n20165 : n20268;
  assign n20270 = pi16 ? n32 : n20269;
  assign n20271 = pi15 ? n20264 : n20270;
  assign n20272 = pi14 ? n20261 : n20271;
  assign n20273 = pi14 ? n19621 : n20176;
  assign n20274 = pi13 ? n20272 : n20273;
  assign n20275 = pi12 ? n20255 : n20274;
  assign n20276 = pi16 ? n19652 : ~n20201;
  assign n20277 = pi16 ? n19652 : ~n20204;
  assign n20278 = pi15 ? n20276 : n20277;
  assign n20279 = pi19 ? n15696 : n32;
  assign n20280 = pi18 ? n32 : n20279;
  assign n20281 = pi17 ? n32 : n20280;
  assign n20282 = pi16 ? n32 : n20281;
  assign n20283 = pi15 ? n20212 : n20282;
  assign n20284 = pi14 ? n20278 : n20283;
  assign n20285 = pi13 ? n20199 : n20284;
  assign n20286 = pi15 ? n18657 : n18805;
  assign n20287 = pi14 ? n20286 : n18535;
  assign n20288 = pi15 ? n19267 : n18294;
  assign n20289 = pi15 ? n18294 : n41;
  assign n20290 = pi14 ? n20288 : n20289;
  assign n20291 = pi13 ? n20287 : n20290;
  assign n20292 = pi12 ? n20285 : n20291;
  assign n20293 = pi11 ? n20275 : n20292;
  assign n20294 = pi10 ? n20241 : n20293;
  assign n20295 = pi09 ? n32 : n20294;
  assign n20296 = pi08 ? n20223 : n20295;
  assign n20297 = pi15 ? n32 : n146;
  assign n20298 = pi19 ? n17062 : n32;
  assign n20299 = pi18 ? n32 : n20298;
  assign n20300 = pi17 ? n32 : n20299;
  assign n20301 = pi16 ? n32 : n20300;
  assign n20302 = pi15 ? n20301 : n13952;
  assign n20303 = pi14 ? n20297 : n20302;
  assign n20304 = pi13 ? n32 : n20303;
  assign n20305 = pi12 ? n32 : n20304;
  assign n20306 = pi15 ? n13952 : n146;
  assign n20307 = pi14 ? n20306 : n147;
  assign n20308 = pi13 ? n20307 : n32;
  assign n20309 = pi14 ? n32 : n20049;
  assign n20310 = pi13 ? n20309 : n20054;
  assign n20311 = pi12 ? n20308 : n20310;
  assign n20312 = pi11 ? n20305 : n20311;
  assign n20313 = pi18 ? n32 : n19774;
  assign n20314 = pi17 ? n32 : n20313;
  assign n20315 = pi16 ? n32 : n20314;
  assign n20316 = pi15 ? n32 : n20315;
  assign n20317 = pi18 ? n880 : ~n430;
  assign n20318 = pi17 ? n32 : n20317;
  assign n20319 = pi16 ? n32 : n20318;
  assign n20320 = pi19 ? n10645 : n32;
  assign n20321 = pi18 ? n32 : n20320;
  assign n20322 = pi17 ? n32 : n20321;
  assign n20323 = pi16 ? n32 : n20322;
  assign n20324 = pi15 ? n20319 : n20323;
  assign n20325 = pi14 ? n20316 : n20324;
  assign n20326 = pi20 ? n18624 : n32;
  assign n20327 = pi19 ? n20326 : n32;
  assign n20328 = pi18 ? n32 : n20327;
  assign n20329 = pi17 ? n32 : n20328;
  assign n20330 = pi16 ? n32 : n20329;
  assign n20331 = pi15 ? n20323 : n20330;
  assign n20332 = pi18 ? n17848 : n20327;
  assign n20333 = pi17 ? n32 : n20332;
  assign n20334 = pi16 ? n32 : n20333;
  assign n20335 = pi15 ? n20323 : n20334;
  assign n20336 = pi14 ? n20331 : n20335;
  assign n20337 = pi13 ? n20325 : n20336;
  assign n20338 = pi19 ? n16597 : n32;
  assign n20339 = pi18 ? n4380 : n20338;
  assign n20340 = pi17 ? n32 : n20339;
  assign n20341 = pi16 ? n32 : n20340;
  assign n20342 = pi15 ? n20341 : n19503;
  assign n20343 = pi14 ? n20341 : n20342;
  assign n20344 = pi15 ? n19805 : n91;
  assign n20345 = pi19 ? n14552 : ~n32;
  assign n20346 = pi18 ? n4380 : ~n20345;
  assign n20347 = pi17 ? n16099 : n20346;
  assign n20348 = pi16 ? n32 : n20347;
  assign n20349 = pi15 ? n91 : n20348;
  assign n20350 = pi14 ? n20344 : n20349;
  assign n20351 = pi13 ? n20343 : n20350;
  assign n20352 = pi12 ? n20337 : n20351;
  assign n20353 = pi21 ? n259 : ~n242;
  assign n20354 = pi20 ? n20353 : n32;
  assign n20355 = pi19 ? n20354 : n32;
  assign n20356 = pi18 ? n32 : n20355;
  assign n20357 = pi17 ? n16103 : n20356;
  assign n20358 = pi16 ? n32 : n20357;
  assign n20359 = pi19 ? n32 : ~n5694;
  assign n20360 = pi18 ? n32 : n20359;
  assign n20361 = pi19 ? n349 : ~n1464;
  assign n20362 = pi18 ? n20361 : n2318;
  assign n20363 = pi17 ? n20360 : ~n20362;
  assign n20364 = pi16 ? n32 : n20363;
  assign n20365 = pi15 ? n20358 : n20364;
  assign n20366 = pi19 ? n16294 : n32;
  assign n20367 = pi18 ? n20366 : n323;
  assign n20368 = pi20 ? n266 : n915;
  assign n20369 = pi19 ? n32 : n20368;
  assign n20370 = pi18 ? n20369 : n1548;
  assign n20371 = pi17 ? n20367 : ~n20370;
  assign n20372 = pi16 ? n32 : n20371;
  assign n20373 = pi18 ? n4689 : n323;
  assign n20374 = pi19 ? n10890 : ~n32;
  assign n20375 = pi18 ? n20193 : n20374;
  assign n20376 = pi17 ? n20373 : ~n20375;
  assign n20377 = pi16 ? n32 : n20376;
  assign n20378 = pi15 ? n20372 : n20377;
  assign n20379 = pi14 ? n20365 : n20378;
  assign n20380 = pi19 ? n32 : n440;
  assign n20381 = pi18 ? n20380 : n32;
  assign n20382 = pi17 ? n20381 : n2537;
  assign n20383 = pi16 ? n1214 : ~n20382;
  assign n20384 = pi19 ? n507 : ~n813;
  assign n20385 = pi18 ? n20384 : n32;
  assign n20386 = pi19 ? n16304 : n32;
  assign n20387 = pi18 ? n32 : ~n20386;
  assign n20388 = pi17 ? n20385 : n20387;
  assign n20389 = pi16 ? n1214 : ~n20388;
  assign n20390 = pi15 ? n20383 : n20389;
  assign n20391 = pi20 ? n17665 : n1817;
  assign n20392 = pi19 ? n20391 : n1817;
  assign n20393 = pi18 ? n463 : n20392;
  assign n20394 = pi17 ? n32 : n20393;
  assign n20395 = pi19 ? n19547 : n19129;
  assign n20396 = pi21 ? n313 : ~n405;
  assign n20397 = pi20 ? n1817 : ~n20396;
  assign n20398 = pi19 ? n19551 : n20397;
  assign n20399 = pi18 ? n20395 : n20398;
  assign n20400 = pi20 ? n18129 : n309;
  assign n20401 = pi20 ? n18415 : ~n333;
  assign n20402 = pi19 ? n20400 : ~n20401;
  assign n20403 = pi18 ? n20402 : n18894;
  assign n20404 = pi17 ? n20399 : n20403;
  assign n20405 = pi16 ? n20394 : n20404;
  assign n20406 = pi15 ? n20405 : n18657;
  assign n20407 = pi14 ? n20390 : n20406;
  assign n20408 = pi13 ? n20379 : n20407;
  assign n20409 = pi14 ? n18662 : n19333;
  assign n20410 = pi14 ? n20110 : n57;
  assign n20411 = pi13 ? n20409 : n20410;
  assign n20412 = pi12 ? n20408 : n20411;
  assign n20413 = pi11 ? n20352 : n20412;
  assign n20414 = pi10 ? n20312 : n20413;
  assign n20415 = pi09 ? n32 : n20414;
  assign n20416 = pi15 ? n32 : n13952;
  assign n20417 = pi14 ? n20416 : n13952;
  assign n20418 = pi13 ? n32 : n20417;
  assign n20419 = pi12 ? n32 : n20418;
  assign n20420 = pi13 ? n20309 : n20127;
  assign n20421 = pi12 ? n20308 : n20420;
  assign n20422 = pi11 ? n20419 : n20421;
  assign n20423 = pi15 ? n19969 : n19856;
  assign n20424 = pi18 ? n880 : ~n2298;
  assign n20425 = pi17 ? n32 : n20424;
  assign n20426 = pi16 ? n32 : n20425;
  assign n20427 = pi15 ? n20426 : n13089;
  assign n20428 = pi14 ? n20423 : n20427;
  assign n20429 = pi21 ? n206 : n14158;
  assign n20430 = pi20 ? n20429 : n32;
  assign n20431 = pi19 ? n20430 : n32;
  assign n20432 = pi18 ? n32 : n20431;
  assign n20433 = pi17 ? n32 : n20432;
  assign n20434 = pi16 ? n32 : n20433;
  assign n20435 = pi15 ? n13089 : n20434;
  assign n20436 = pi18 ? n17848 : n20431;
  assign n20437 = pi17 ? n32 : n20436;
  assign n20438 = pi16 ? n32 : n20437;
  assign n20439 = pi15 ? n13089 : n20438;
  assign n20440 = pi14 ? n20435 : n20439;
  assign n20441 = pi13 ? n20428 : n20440;
  assign n20442 = pi18 ? n4380 : n19774;
  assign n20443 = pi17 ? n32 : n20442;
  assign n20444 = pi16 ? n32 : n20443;
  assign n20445 = pi15 ? n20444 : n19503;
  assign n20446 = pi14 ? n20444 : n20445;
  assign n20447 = pi15 ? n19805 : n19503;
  assign n20448 = pi18 ? n4380 : ~n350;
  assign n20449 = pi17 ? n16099 : n20448;
  assign n20450 = pi16 ? n32 : n20449;
  assign n20451 = pi15 ? n19503 : n20450;
  assign n20452 = pi14 ? n20447 : n20451;
  assign n20453 = pi13 ? n20446 : n20452;
  assign n20454 = pi12 ? n20441 : n20453;
  assign n20455 = pi20 ? n1817 : ~n831;
  assign n20456 = pi19 ? n358 : n20455;
  assign n20457 = pi18 ? n20395 : n20456;
  assign n20458 = pi20 ? n18129 : n3523;
  assign n20459 = pi19 ? n20458 : n334;
  assign n20460 = pi18 ? n20459 : n18894;
  assign n20461 = pi17 ? n20457 : n20460;
  assign n20462 = pi16 ? n32 : n20461;
  assign n20463 = pi15 ? n20462 : n19030;
  assign n20464 = pi14 ? n20390 : n20463;
  assign n20465 = pi13 ? n20379 : n20464;
  assign n20466 = pi14 ? n18662 : n18947;
  assign n20467 = pi13 ? n20466 : n20410;
  assign n20468 = pi12 ? n20465 : n20467;
  assign n20469 = pi11 ? n20454 : n20468;
  assign n20470 = pi10 ? n20422 : n20469;
  assign n20471 = pi09 ? n32 : n20470;
  assign n20472 = pi08 ? n20415 : n20471;
  assign n20473 = pi07 ? n20296 : n20472;
  assign n20474 = pi19 ? n8035 : n32;
  assign n20475 = pi18 ? n32 : n20474;
  assign n20476 = pi17 ? n32 : n20475;
  assign n20477 = pi16 ? n32 : n20476;
  assign n20478 = pi15 ? n32 : n20477;
  assign n20479 = pi14 ? n20478 : n20477;
  assign n20480 = pi13 ? n32 : n20479;
  assign n20481 = pi12 ? n32 : n20480;
  assign n20482 = pi20 ? n32 : n15660;
  assign n20483 = pi19 ? n20482 : n32;
  assign n20484 = pi18 ? n32 : n20483;
  assign n20485 = pi17 ? n32 : n20484;
  assign n20486 = pi16 ? n32 : n20485;
  assign n20487 = pi15 ? n20486 : n671;
  assign n20488 = pi14 ? n20487 : n32;
  assign n20489 = pi13 ? n20488 : n32;
  assign n20490 = pi19 ? n16949 : n32;
  assign n20491 = pi18 ? n32 : n20490;
  assign n20492 = pi17 ? n32 : n20491;
  assign n20493 = pi16 ? n32 : n20492;
  assign n20494 = pi15 ? n32 : n20493;
  assign n20495 = pi14 ? n20049 : n20494;
  assign n20496 = pi15 ? n20493 : n20048;
  assign n20497 = pi14 ? n20496 : n107;
  assign n20498 = pi13 ? n20495 : n20497;
  assign n20499 = pi12 ? n20489 : n20498;
  assign n20500 = pi11 ? n20481 : n20499;
  assign n20501 = pi21 ? n174 : ~n7107;
  assign n20502 = pi20 ? n20501 : ~n32;
  assign n20503 = pi19 ? n20502 : ~n32;
  assign n20504 = pi18 ? n268 : ~n20503;
  assign n20505 = pi17 ? n32 : n20504;
  assign n20506 = pi16 ? n32 : n20505;
  assign n20507 = pi21 ? n206 : n7107;
  assign n20508 = pi20 ? n20507 : n32;
  assign n20509 = pi19 ? n20508 : n32;
  assign n20510 = pi18 ? n32 : n20509;
  assign n20511 = pi17 ? n32 : n20510;
  assign n20512 = pi16 ? n32 : n20511;
  assign n20513 = pi15 ? n20506 : n20512;
  assign n20514 = pi15 ? n20434 : n19856;
  assign n20515 = pi14 ? n20513 : n20514;
  assign n20516 = pi21 ? n32 : ~n14158;
  assign n20517 = pi20 ? n20516 : ~n32;
  assign n20518 = pi19 ? n20517 : ~n32;
  assign n20519 = pi18 ? n751 : ~n20518;
  assign n20520 = pi17 ? n32 : n20519;
  assign n20521 = pi16 ? n32 : n20520;
  assign n20522 = pi15 ? n19856 : n20521;
  assign n20523 = pi14 ? n19856 : n20522;
  assign n20524 = pi13 ? n20515 : n20523;
  assign n20525 = pi19 ? n11108 : ~n32;
  assign n20526 = pi18 ? n32 : ~n20525;
  assign n20527 = pi17 ? n32 : n20526;
  assign n20528 = pi16 ? n32 : n20527;
  assign n20529 = pi18 ? n32 : n19750;
  assign n20530 = pi17 ? n32 : n20529;
  assign n20531 = pi16 ? n32 : n20530;
  assign n20532 = pi15 ? n20528 : n20531;
  assign n20533 = pi18 ? n940 : n19750;
  assign n20534 = pi17 ? n32 : n20533;
  assign n20535 = pi16 ? n32 : n20534;
  assign n20536 = pi18 ? n32 : n20338;
  assign n20537 = pi17 ? n32 : n20536;
  assign n20538 = pi16 ? n32 : n20537;
  assign n20539 = pi15 ? n20535 : n20538;
  assign n20540 = pi14 ? n20532 : n20539;
  assign n20541 = pi18 ? n4380 : ~n344;
  assign n20542 = pi17 ? n32 : n20541;
  assign n20543 = pi16 ? n32 : n20542;
  assign n20544 = pi15 ? n20258 : n20543;
  assign n20545 = pi17 ? n15850 : n20541;
  assign n20546 = pi16 ? n32 : n20545;
  assign n20547 = pi19 ? n4342 : n208;
  assign n20548 = pi18 ? n20547 : ~n344;
  assign n20549 = pi17 ? n3067 : n20548;
  assign n20550 = pi16 ? n32 : n20549;
  assign n20551 = pi15 ? n20546 : n20550;
  assign n20552 = pi14 ? n20544 : n20551;
  assign n20553 = pi13 ? n20540 : n20552;
  assign n20554 = pi12 ? n20524 : n20553;
  assign n20555 = pi20 ? n321 : ~n246;
  assign n20556 = pi19 ? n343 : n20555;
  assign n20557 = pi18 ? n20556 : n344;
  assign n20558 = pi17 ? n3067 : ~n20557;
  assign n20559 = pi16 ? n32 : n20558;
  assign n20560 = pi18 ? n13668 : n496;
  assign n20561 = pi18 ? n16847 : n344;
  assign n20562 = pi17 ? n20560 : ~n20561;
  assign n20563 = pi16 ? n32 : n20562;
  assign n20564 = pi15 ? n20559 : n20563;
  assign n20565 = pi19 ? n32 : n19749;
  assign n20566 = pi18 ? n20565 : n32;
  assign n20567 = pi18 ? n16847 : n2318;
  assign n20568 = pi17 ? n20566 : n20567;
  assign n20569 = pi16 ? n1471 : ~n20568;
  assign n20570 = pi18 ? n16449 : n32;
  assign n20571 = pi17 ? n20570 : n2319;
  assign n20572 = pi16 ? n1471 : ~n20571;
  assign n20573 = pi15 ? n20569 : n20572;
  assign n20574 = pi14 ? n20564 : n20573;
  assign n20575 = pi18 ? n268 : n19933;
  assign n20576 = pi17 ? n32 : n20575;
  assign n20577 = pi16 ? n32 : n20576;
  assign n20578 = pi15 ? n20572 : n20577;
  assign n20579 = pi15 ? n18904 : n19030;
  assign n20580 = pi14 ? n20578 : n20579;
  assign n20581 = pi13 ? n20574 : n20580;
  assign n20582 = pi15 ? n19030 : n32;
  assign n20583 = pi15 ? n32 : n18661;
  assign n20584 = pi14 ? n20582 : n20583;
  assign n20585 = pi14 ? n20216 : n18948;
  assign n20586 = pi13 ? n20584 : n20585;
  assign n20587 = pi12 ? n20581 : n20586;
  assign n20588 = pi11 ? n20554 : n20587;
  assign n20589 = pi10 ? n20500 : n20588;
  assign n20590 = pi09 ? n32 : n20589;
  assign n20591 = pi15 ? n20477 : n32;
  assign n20592 = pi14 ? n20591 : n32;
  assign n20593 = pi13 ? n20592 : n32;
  assign n20594 = pi15 ? n32 : n20301;
  assign n20595 = pi14 ? n20049 : n20594;
  assign n20596 = pi15 ? n20301 : n13684;
  assign n20597 = pi14 ? n20596 : n147;
  assign n20598 = pi13 ? n20595 : n20597;
  assign n20599 = pi12 ? n20593 : n20598;
  assign n20600 = pi11 ? n20481 : n20599;
  assign n20601 = pi19 ? n6619 : ~n32;
  assign n20602 = pi18 ? n268 : ~n20601;
  assign n20603 = pi17 ? n32 : n20602;
  assign n20604 = pi16 ? n32 : n20603;
  assign n20605 = pi19 ? n7642 : n32;
  assign n20606 = pi18 ? n32 : n20605;
  assign n20607 = pi17 ? n32 : n20606;
  assign n20608 = pi16 ? n32 : n20607;
  assign n20609 = pi15 ? n20604 : n20608;
  assign n20610 = pi20 ? n287 : n32;
  assign n20611 = pi19 ? n20610 : n32;
  assign n20612 = pi18 ? n32 : n20611;
  assign n20613 = pi17 ? n32 : n20612;
  assign n20614 = pi16 ? n32 : n20613;
  assign n20615 = pi19 ? n16542 : n32;
  assign n20616 = pi18 ? n32 : n20615;
  assign n20617 = pi17 ? n32 : n20616;
  assign n20618 = pi16 ? n32 : n20617;
  assign n20619 = pi15 ? n20614 : n20618;
  assign n20620 = pi14 ? n20609 : n20619;
  assign n20621 = pi19 ? n11531 : ~n32;
  assign n20622 = pi18 ? n751 : ~n20621;
  assign n20623 = pi17 ? n32 : n20622;
  assign n20624 = pi16 ? n32 : n20623;
  assign n20625 = pi15 ? n20618 : n20624;
  assign n20626 = pi14 ? n20618 : n20625;
  assign n20627 = pi13 ? n20620 : n20626;
  assign n20628 = pi19 ? n11561 : ~n32;
  assign n20629 = pi18 ? n32 : ~n20628;
  assign n20630 = pi17 ? n32 : n20629;
  assign n20631 = pi16 ? n32 : n20630;
  assign n20632 = pi15 ? n20631 : n19851;
  assign n20633 = pi14 ? n20632 : n20539;
  assign n20634 = pi18 ? n4380 : n20249;
  assign n20635 = pi17 ? n32 : n20634;
  assign n20636 = pi16 ? n32 : n20635;
  assign n20637 = pi18 ? n4380 : ~n2304;
  assign n20638 = pi17 ? n32 : n20637;
  assign n20639 = pi16 ? n32 : n20638;
  assign n20640 = pi15 ? n20636 : n20639;
  assign n20641 = pi14 ? n20640 : n20551;
  assign n20642 = pi13 ? n20633 : n20641;
  assign n20643 = pi12 ? n20627 : n20642;
  assign n20644 = pi18 ? n32 : n20386;
  assign n20645 = pi17 ? n32 : n20644;
  assign n20646 = pi16 ? n32 : n20645;
  assign n20647 = pi15 ? n20646 : n19235;
  assign n20648 = pi14 ? n20578 : n20647;
  assign n20649 = pi13 ? n20574 : n20648;
  assign n20650 = pi14 ? n18905 : n18657;
  assign n20651 = pi14 ? n20216 : n18535;
  assign n20652 = pi13 ? n20650 : n20651;
  assign n20653 = pi12 ? n20649 : n20652;
  assign n20654 = pi11 ? n20643 : n20653;
  assign n20655 = pi10 ? n20600 : n20654;
  assign n20656 = pi09 ? n32 : n20655;
  assign n20657 = pi08 ? n20590 : n20656;
  assign n20658 = pi18 ? n32 : n7221;
  assign n20659 = pi17 ? n32 : n20658;
  assign n20660 = pi16 ? n32 : n20659;
  assign n20661 = pi15 ? n32 : n20660;
  assign n20662 = pi14 ? n20661 : n20660;
  assign n20663 = pi13 ? n32 : n20662;
  assign n20664 = pi12 ? n32 : n20663;
  assign n20665 = pi15 ? n20660 : n32;
  assign n20666 = pi14 ? n20665 : n32;
  assign n20667 = pi13 ? n20666 : n32;
  assign n20668 = pi15 ? n486 : n20477;
  assign n20669 = pi14 ? n487 : n20668;
  assign n20670 = pi15 ? n20477 : n146;
  assign n20671 = pi19 ? n16828 : n32;
  assign n20672 = pi18 ? n863 : n20671;
  assign n20673 = pi17 ? n32 : n20672;
  assign n20674 = pi16 ? n32 : n20673;
  assign n20675 = pi15 ? n146 : n20674;
  assign n20676 = pi14 ? n20670 : n20675;
  assign n20677 = pi13 ? n20669 : n20676;
  assign n20678 = pi12 ? n20667 : n20677;
  assign n20679 = pi11 ? n20664 : n20678;
  assign n20680 = pi19 ? n9903 : ~n32;
  assign n20681 = pi18 ? n4127 : ~n20680;
  assign n20682 = pi17 ? n32 : n20681;
  assign n20683 = pi16 ? n32 : n20682;
  assign n20684 = pi18 ? n863 : n20605;
  assign n20685 = pi17 ? n32 : n20684;
  assign n20686 = pi16 ? n32 : n20685;
  assign n20687 = pi15 ? n20683 : n20686;
  assign n20688 = pi15 ? n20608 : n19972;
  assign n20689 = pi14 ? n20687 : n20688;
  assign n20690 = pi18 ? n32 : n4343;
  assign n20691 = pi17 ? n32 : n20690;
  assign n20692 = pi16 ? n32 : n20691;
  assign n20693 = pi18 ? n940 : ~n532;
  assign n20694 = pi17 ? n32 : n20693;
  assign n20695 = pi16 ? n32 : n20694;
  assign n20696 = pi15 ? n20692 : n20695;
  assign n20697 = pi14 ? n19972 : n20696;
  assign n20698 = pi13 ? n20689 : n20697;
  assign n20699 = pi18 ? n4380 : ~n20628;
  assign n20700 = pi17 ? n32 : n20699;
  assign n20701 = pi16 ? n32 : n20700;
  assign n20702 = pi18 ? n940 : n20431;
  assign n20703 = pi17 ? n32 : n20702;
  assign n20704 = pi16 ? n32 : n20703;
  assign n20705 = pi15 ? n20701 : n20704;
  assign n20706 = pi18 ? n17848 : n20338;
  assign n20707 = pi17 ? n32 : n20706;
  assign n20708 = pi16 ? n32 : n20707;
  assign n20709 = pi15 ? n13392 : n20708;
  assign n20710 = pi14 ? n20705 : n20709;
  assign n20711 = pi18 ? n4380 : n19865;
  assign n20712 = pi17 ? n32 : n20711;
  assign n20713 = pi16 ? n32 : n20712;
  assign n20714 = pi15 ? n20713 : n20639;
  assign n20715 = pi17 ? n16848 : n20637;
  assign n20716 = pi16 ? n32 : n20715;
  assign n20717 = pi19 ? n5004 : n208;
  assign n20718 = pi18 ? n20717 : ~n2304;
  assign n20719 = pi17 ? n2726 : n20718;
  assign n20720 = pi16 ? n32 : n20719;
  assign n20721 = pi15 ? n20716 : n20720;
  assign n20722 = pi14 ? n20714 : n20721;
  assign n20723 = pi13 ? n20710 : n20722;
  assign n20724 = pi12 ? n20698 : n20723;
  assign n20725 = pi19 ? n208 : n4964;
  assign n20726 = pi18 ? n20725 : n2304;
  assign n20727 = pi17 ? n2733 : ~n20726;
  assign n20728 = pi16 ? n32 : n20727;
  assign n20729 = pi19 ? n916 : n32;
  assign n20730 = pi18 ? n20729 : n496;
  assign n20731 = pi18 ? n16847 : n2304;
  assign n20732 = pi17 ? n20730 : ~n20731;
  assign n20733 = pi16 ? n32 : n20732;
  assign n20734 = pi15 ? n20728 : n20733;
  assign n20735 = pi18 ? n16234 : n32;
  assign n20736 = pi17 ? n20735 : n20561;
  assign n20737 = pi16 ? n1471 : ~n20736;
  assign n20738 = pi18 ? n17063 : n32;
  assign n20739 = pi17 ? n20738 : n1933;
  assign n20740 = pi16 ? n1471 : ~n20739;
  assign n20741 = pi15 ? n20737 : n20740;
  assign n20742 = pi14 ? n20734 : n20741;
  assign n20743 = pi15 ? n20740 : n19384;
  assign n20744 = pi14 ? n20743 : n19235;
  assign n20745 = pi13 ? n20742 : n20744;
  assign n20746 = pi15 ? n165 : n32;
  assign n20747 = pi14 ? n20746 : n19626;
  assign n20748 = pi13 ? n20747 : n20466;
  assign n20749 = pi12 ? n20745 : n20748;
  assign n20750 = pi11 ? n20724 : n20749;
  assign n20751 = pi10 ? n20679 : n20750;
  assign n20752 = pi09 ? n32 : n20751;
  assign n20753 = pi19 ? n17294 : n32;
  assign n20754 = pi18 ? n32 : n20753;
  assign n20755 = pi17 ? n32 : n20754;
  assign n20756 = pi16 ? n32 : n20755;
  assign n20757 = pi15 ? n32 : n20756;
  assign n20758 = pi15 ? n20756 : n20660;
  assign n20759 = pi14 ? n20757 : n20758;
  assign n20760 = pi13 ? n32 : n20759;
  assign n20761 = pi12 ? n32 : n20760;
  assign n20762 = pi14 ? n32 : n20668;
  assign n20763 = pi15 ? n32 : n20674;
  assign n20764 = pi14 ? n20487 : n20763;
  assign n20765 = pi13 ? n20762 : n20764;
  assign n20766 = pi12 ? n20667 : n20765;
  assign n20767 = pi11 ? n20761 : n20766;
  assign n20768 = pi20 ? n206 : ~n141;
  assign n20769 = pi19 ? n20768 : n32;
  assign n20770 = pi18 ? n863 : n20769;
  assign n20771 = pi17 ? n32 : n20770;
  assign n20772 = pi16 ? n32 : n20771;
  assign n20773 = pi15 ? n20683 : n20772;
  assign n20774 = pi18 ? n32 : n20769;
  assign n20775 = pi17 ? n32 : n20774;
  assign n20776 = pi16 ? n32 : n20775;
  assign n20777 = pi18 ? n32 : n20671;
  assign n20778 = pi17 ? n32 : n20777;
  assign n20779 = pi16 ? n32 : n20778;
  assign n20780 = pi15 ? n20776 : n20779;
  assign n20781 = pi14 ? n20773 : n20780;
  assign n20782 = pi18 ? n940 : ~n3786;
  assign n20783 = pi17 ? n32 : n20782;
  assign n20784 = pi16 ? n32 : n20783;
  assign n20785 = pi15 ? n13380 : n20784;
  assign n20786 = pi14 ? n20779 : n20785;
  assign n20787 = pi13 ? n20781 : n20786;
  assign n20788 = pi19 ? n8818 : ~n32;
  assign n20789 = pi18 ? n4380 : ~n20788;
  assign n20790 = pi17 ? n32 : n20789;
  assign n20791 = pi16 ? n32 : n20790;
  assign n20792 = pi18 ? n940 : n20611;
  assign n20793 = pi17 ? n32 : n20792;
  assign n20794 = pi16 ? n32 : n20793;
  assign n20795 = pi15 ? n20791 : n20794;
  assign n20796 = pi18 ? n17848 : n19774;
  assign n20797 = pi17 ? n32 : n20796;
  assign n20798 = pi16 ? n32 : n20797;
  assign n20799 = pi15 ? n13392 : n20798;
  assign n20800 = pi14 ? n20795 : n20799;
  assign n20801 = pi18 ? n4380 : n19750;
  assign n20802 = pi17 ? n32 : n20801;
  assign n20803 = pi16 ? n32 : n20802;
  assign n20804 = pi18 ? n4380 : ~n430;
  assign n20805 = pi17 ? n32 : n20804;
  assign n20806 = pi16 ? n32 : n20805;
  assign n20807 = pi15 ? n20803 : n20806;
  assign n20808 = pi17 ? n16848 : n20541;
  assign n20809 = pi16 ? n32 : n20808;
  assign n20810 = pi18 ? n20717 : ~n344;
  assign n20811 = pi17 ? n2726 : n20810;
  assign n20812 = pi16 ? n32 : n20811;
  assign n20813 = pi15 ? n20809 : n20812;
  assign n20814 = pi14 ? n20807 : n20813;
  assign n20815 = pi13 ? n20800 : n20814;
  assign n20816 = pi12 ? n20787 : n20815;
  assign n20817 = pi15 ? n20740 : n19805;
  assign n20818 = pi14 ? n20817 : n19621;
  assign n20819 = pi13 ? n20742 : n20818;
  assign n20820 = pi13 ? n19627 : n20466;
  assign n20821 = pi12 ? n20819 : n20820;
  assign n20822 = pi11 ? n20816 : n20821;
  assign n20823 = pi10 ? n20767 : n20822;
  assign n20824 = pi09 ? n32 : n20823;
  assign n20825 = pi08 ? n20752 : n20824;
  assign n20826 = pi07 ? n20657 : n20825;
  assign n20827 = pi06 ? n20473 : n20826;
  assign n20828 = pi19 ? n17332 : n32;
  assign n20829 = pi18 ? n32 : n20828;
  assign n20830 = pi17 ? n32 : n20829;
  assign n20831 = pi16 ? n32 : n20830;
  assign n20832 = pi15 ? n32 : n20831;
  assign n20833 = pi14 ? n32 : n20832;
  assign n20834 = pi18 ? n32 : n5158;
  assign n20835 = pi17 ? n32 : n20834;
  assign n20836 = pi16 ? n32 : n20835;
  assign n20837 = pi15 ? n20831 : n20836;
  assign n20838 = pi15 ? n20831 : n32;
  assign n20839 = pi14 ? n20837 : n20838;
  assign n20840 = pi13 ? n20833 : n20839;
  assign n20841 = pi12 ? n32 : n20840;
  assign n20842 = pi14 ? n20838 : n32;
  assign n20843 = pi13 ? n20842 : n32;
  assign n20844 = pi15 ? n32 : n13948;
  assign n20845 = pi15 ? n13948 : n20660;
  assign n20846 = pi14 ? n20844 : n20845;
  assign n20847 = pi15 ? n486 : n13952;
  assign n20848 = pi19 ? n7405 : n32;
  assign n20849 = pi18 ? n863 : n20848;
  assign n20850 = pi17 ? n32 : n20849;
  assign n20851 = pi16 ? n32 : n20850;
  assign n20852 = pi18 ? n863 : n13668;
  assign n20853 = pi17 ? n32 : n20852;
  assign n20854 = pi16 ? n32 : n20853;
  assign n20855 = pi15 ? n20851 : n20854;
  assign n20856 = pi14 ? n20847 : n20855;
  assign n20857 = pi13 ? n20846 : n20856;
  assign n20858 = pi12 ? n20843 : n20857;
  assign n20859 = pi11 ? n20841 : n20858;
  assign n20860 = pi18 ? n4722 : n20605;
  assign n20861 = pi17 ? n32 : n20860;
  assign n20862 = pi16 ? n32 : n20861;
  assign n20863 = pi18 ? n940 : n4671;
  assign n20864 = pi17 ? n32 : n20863;
  assign n20865 = pi16 ? n32 : n20864;
  assign n20866 = pi15 ? n20862 : n20865;
  assign n20867 = pi14 ? n20866 : n19972;
  assign n20868 = pi18 ? n17848 : n4671;
  assign n20869 = pi17 ? n32 : n20868;
  assign n20870 = pi16 ? n32 : n20869;
  assign n20871 = pi18 ? n4380 : n4343;
  assign n20872 = pi17 ? n32 : n20871;
  assign n20873 = pi16 ? n32 : n20872;
  assign n20874 = pi15 ? n20870 : n20873;
  assign n20875 = pi18 ? n4380 : n13377;
  assign n20876 = pi17 ? n32 : n20875;
  assign n20877 = pi16 ? n32 : n20876;
  assign n20878 = pi15 ? n20877 : n20784;
  assign n20879 = pi14 ? n20874 : n20878;
  assign n20880 = pi13 ? n20867 : n20879;
  assign n20881 = pi18 ? n880 : ~n532;
  assign n20882 = pi17 ? n32 : n20881;
  assign n20883 = pi16 ? n32 : n20882;
  assign n20884 = pi20 ? n4279 : n32;
  assign n20885 = pi19 ? n20884 : n32;
  assign n20886 = pi18 ? n32 : n20885;
  assign n20887 = pi17 ? n32 : n20886;
  assign n20888 = pi16 ? n32 : n20887;
  assign n20889 = pi15 ? n20883 : n20888;
  assign n20890 = pi18 ? n17848 : n177;
  assign n20891 = pi17 ? n32 : n20890;
  assign n20892 = pi16 ? n32 : n20891;
  assign n20893 = pi15 ? n20870 : n20892;
  assign n20894 = pi14 ? n20889 : n20893;
  assign n20895 = pi18 ? n940 : ~n430;
  assign n20896 = pi17 ? n32 : n20895;
  assign n20897 = pi16 ? n32 : n20896;
  assign n20898 = pi15 ? n20806 : n20897;
  assign n20899 = pi18 ? n209 : ~n430;
  assign n20900 = pi17 ? n17463 : n20899;
  assign n20901 = pi16 ? n32 : n20900;
  assign n20902 = pi18 ? n14413 : n430;
  assign n20903 = pi17 ? n2959 : ~n20902;
  assign n20904 = pi16 ? n32 : n20903;
  assign n20905 = pi15 ? n20901 : n20904;
  assign n20906 = pi14 ? n20898 : n20905;
  assign n20907 = pi13 ? n20894 : n20906;
  assign n20908 = pi12 ? n20880 : n20907;
  assign n20909 = pi18 ? n6581 : n430;
  assign n20910 = pi17 ? n2959 : ~n20909;
  assign n20911 = pi16 ? n32 : n20910;
  assign n20912 = pi19 ? n4518 : n32;
  assign n20913 = pi18 ? n20912 : n880;
  assign n20914 = pi18 ? n32 : n20525;
  assign n20915 = pi17 ? n20913 : ~n20914;
  assign n20916 = pi16 ? n32 : n20915;
  assign n20917 = pi15 ? n20911 : n20916;
  assign n20918 = pi17 ? n17734 : n2305;
  assign n20919 = pi16 ? n1683 : ~n20918;
  assign n20920 = pi19 ? n207 : n342;
  assign n20921 = pi18 ? n32 : n20920;
  assign n20922 = pi17 ? n32 : n20921;
  assign n20923 = pi20 ? n342 : n220;
  assign n20924 = pi19 ? n20923 : ~n267;
  assign n20925 = pi20 ? n220 : n342;
  assign n20926 = pi19 ? n20925 : n32;
  assign n20927 = pi18 ? n20924 : ~n20926;
  assign n20928 = pi18 ? n940 : ~n19865;
  assign n20929 = pi17 ? n20927 : ~n20928;
  assign n20930 = pi16 ? n20922 : n20929;
  assign n20931 = pi15 ? n20919 : n20930;
  assign n20932 = pi14 ? n20917 : n20931;
  assign n20933 = pi20 ? n1331 : n18129;
  assign n20934 = pi19 ? n20933 : n175;
  assign n20935 = pi18 ? n32 : n20934;
  assign n20936 = pi17 ? n32 : n20935;
  assign n20937 = pi20 ? n175 : n1331;
  assign n20938 = pi20 ? n18073 : n9641;
  assign n20939 = pi19 ? n20937 : n20938;
  assign n20940 = pi20 ? n428 : n274;
  assign n20941 = pi20 ? n18415 : ~n309;
  assign n20942 = pi19 ? n20940 : ~n20941;
  assign n20943 = pi18 ? n20939 : n20942;
  assign n20944 = pi21 ? n259 : n313;
  assign n20945 = pi20 ? n309 : ~n20944;
  assign n20946 = pi19 ? n20945 : n18789;
  assign n20947 = pi18 ? n20946 : n19865;
  assign n20948 = pi17 ? n20943 : n20947;
  assign n20949 = pi16 ? n20936 : n20948;
  assign n20950 = pi15 ? n20949 : n19805;
  assign n20951 = pi20 ? n17724 : n32;
  assign n20952 = pi19 ? n20951 : n32;
  assign n20953 = pi18 ? n32 : n20952;
  assign n20954 = pi17 ? n32 : n20953;
  assign n20955 = pi16 ? n32 : n20954;
  assign n20956 = pi15 ? n20955 : n19384;
  assign n20957 = pi14 ? n20950 : n20956;
  assign n20958 = pi13 ? n20932 : n20957;
  assign n20959 = pi14 ? n19326 : n166;
  assign n20960 = pi15 ? n18657 : n19531;
  assign n20961 = pi14 ? n18905 : n20960;
  assign n20962 = pi13 ? n20959 : n20961;
  assign n20963 = pi12 ? n20958 : n20962;
  assign n20964 = pi11 ? n20908 : n20963;
  assign n20965 = pi10 ? n20859 : n20964;
  assign n20966 = pi09 ? n32 : n20965;
  assign n20967 = pi15 ? n32 : n20836;
  assign n20968 = pi14 ? n32 : n20967;
  assign n20969 = pi15 ? n20836 : n32;
  assign n20970 = pi14 ? n20836 : n20969;
  assign n20971 = pi13 ? n20968 : n20970;
  assign n20972 = pi12 ? n32 : n20971;
  assign n20973 = pi14 ? n20832 : n20838;
  assign n20974 = pi13 ? n20973 : n32;
  assign n20975 = pi15 ? n20660 : n13952;
  assign n20976 = pi14 ? n20975 : n20855;
  assign n20977 = pi13 ? n20846 : n20976;
  assign n20978 = pi12 ? n20974 : n20977;
  assign n20979 = pi11 ? n20972 : n20978;
  assign n20980 = pi18 ? n4722 : n20848;
  assign n20981 = pi17 ? n32 : n20980;
  assign n20982 = pi16 ? n32 : n20981;
  assign n20983 = pi18 ? n940 : n13668;
  assign n20984 = pi17 ? n32 : n20983;
  assign n20985 = pi16 ? n32 : n20984;
  assign n20986 = pi15 ? n20982 : n20985;
  assign n20987 = pi14 ? n20986 : n13671;
  assign n20988 = pi18 ? n17848 : n13668;
  assign n20989 = pi17 ? n32 : n20988;
  assign n20990 = pi16 ? n32 : n20989;
  assign n20991 = pi18 ? n4380 : n13372;
  assign n20992 = pi17 ? n32 : n20991;
  assign n20993 = pi16 ? n32 : n20992;
  assign n20994 = pi15 ? n20990 : n20993;
  assign n20995 = pi18 ? n940 : ~n418;
  assign n20996 = pi17 ? n32 : n20995;
  assign n20997 = pi16 ? n32 : n20996;
  assign n20998 = pi15 ? n20993 : n20997;
  assign n20999 = pi14 ? n20994 : n20998;
  assign n21000 = pi13 ? n20987 : n20999;
  assign n21001 = pi18 ? n880 : ~n3786;
  assign n21002 = pi17 ? n32 : n21001;
  assign n21003 = pi16 ? n32 : n21002;
  assign n21004 = pi15 ? n21003 : n19972;
  assign n21005 = pi18 ? n17848 : n13389;
  assign n21006 = pi17 ? n32 : n21005;
  assign n21007 = pi16 ? n32 : n21006;
  assign n21008 = pi14 ? n21004 : n21007;
  assign n21009 = pi13 ? n21008 : n20906;
  assign n21010 = pi12 ? n21000 : n21009;
  assign n21011 = pi20 ? n18415 : ~n357;
  assign n21012 = pi19 ? n32 : ~n21011;
  assign n21013 = pi18 ? n177 : n21012;
  assign n21014 = pi19 ? n9169 : n1844;
  assign n21015 = pi18 ? n21014 : n19865;
  assign n21016 = pi17 ? n21013 : n21015;
  assign n21017 = pi16 ? n20936 : n21016;
  assign n21018 = pi15 ? n21017 : n19805;
  assign n21019 = pi14 ? n21018 : n19384;
  assign n21020 = pi13 ? n20932 : n21019;
  assign n21021 = pi15 ? n18657 : n18531;
  assign n21022 = pi14 ? n18905 : n21021;
  assign n21023 = pi13 ? n20959 : n21022;
  assign n21024 = pi12 ? n21020 : n21023;
  assign n21025 = pi11 ? n21010 : n21024;
  assign n21026 = pi10 ? n20979 : n21025;
  assign n21027 = pi09 ? n32 : n21026;
  assign n21028 = pi08 ? n20966 : n21027;
  assign n21029 = pi20 ? n32 : n7487;
  assign n21030 = pi19 ? n21029 : n32;
  assign n21031 = pi18 ? n32 : n21030;
  assign n21032 = pi17 ? n32 : n21031;
  assign n21033 = pi16 ? n32 : n21032;
  assign n21034 = pi15 ? n20836 : n21033;
  assign n21035 = pi15 ? n21033 : n20836;
  assign n21036 = pi14 ? n21034 : n21035;
  assign n21037 = pi13 ? n32 : n21036;
  assign n21038 = pi12 ? n32 : n21037;
  assign n21039 = pi15 ? n20831 : n20756;
  assign n21040 = pi14 ? n20832 : n21039;
  assign n21041 = pi15 ? n20660 : n486;
  assign n21042 = pi20 ? n206 : ~n243;
  assign n21043 = pi19 ? n21042 : n32;
  assign n21044 = pi18 ? n863 : n21043;
  assign n21045 = pi17 ? n32 : n21044;
  assign n21046 = pi16 ? n32 : n21045;
  assign n21047 = pi20 ? n428 : ~n243;
  assign n21048 = pi19 ? n21047 : n32;
  assign n21049 = pi18 ? n863 : n21048;
  assign n21050 = pi17 ? n32 : n21049;
  assign n21051 = pi16 ? n32 : n21050;
  assign n21052 = pi15 ? n21046 : n21051;
  assign n21053 = pi14 ? n21041 : n21052;
  assign n21054 = pi13 ? n21040 : n21053;
  assign n21055 = pi12 ? n32 : n21054;
  assign n21056 = pi11 ? n21038 : n21055;
  assign n21057 = pi15 ? n12098 : n20985;
  assign n21058 = pi14 ? n21057 : n13671;
  assign n21059 = pi18 ? n4380 : n13668;
  assign n21060 = pi17 ? n32 : n21059;
  assign n21061 = pi16 ? n32 : n21060;
  assign n21062 = pi15 ? n21061 : n20993;
  assign n21063 = pi14 ? n21062 : n20998;
  assign n21064 = pi13 ? n21058 : n21063;
  assign n21065 = pi20 ? n32 : ~n9641;
  assign n21066 = pi19 ? n32 : n21065;
  assign n21067 = pi20 ? n1385 : n141;
  assign n21068 = pi19 ? n21067 : ~n32;
  assign n21069 = pi18 ? n21066 : ~n21068;
  assign n21070 = pi17 ? n32 : n21069;
  assign n21071 = pi16 ? n32 : n21070;
  assign n21072 = pi15 ? n21071 : n20779;
  assign n21073 = pi14 ? n21072 : n20053;
  assign n21074 = pi18 ? n4380 : ~n2298;
  assign n21075 = pi17 ? n32 : n21074;
  assign n21076 = pi16 ? n32 : n21075;
  assign n21077 = pi18 ? n940 : ~n2298;
  assign n21078 = pi17 ? n32 : n21077;
  assign n21079 = pi16 ? n32 : n21078;
  assign n21080 = pi15 ? n21076 : n21079;
  assign n21081 = pi19 ? n507 : n208;
  assign n21082 = pi18 ? n21081 : ~n2298;
  assign n21083 = pi17 ? n4261 : n21082;
  assign n21084 = pi16 ? n32 : n21083;
  assign n21085 = pi18 ? n14982 : n2298;
  assign n21086 = pi17 ? n2954 : ~n21085;
  assign n21087 = pi16 ? n32 : n21086;
  assign n21088 = pi15 ? n21084 : n21087;
  assign n21089 = pi14 ? n21080 : n21088;
  assign n21090 = pi13 ? n21073 : n21089;
  assign n21091 = pi12 ? n21064 : n21090;
  assign n21092 = pi18 ? n15241 : n2298;
  assign n21093 = pi17 ? n3164 : ~n21092;
  assign n21094 = pi16 ? n32 : n21093;
  assign n21095 = pi18 ? n18474 : n880;
  assign n21096 = pi18 ? n32 : n20628;
  assign n21097 = pi17 ? n21095 : ~n21096;
  assign n21098 = pi16 ? n32 : n21097;
  assign n21099 = pi15 ? n21094 : n21098;
  assign n21100 = pi17 ? n210 : n2410;
  assign n21101 = pi16 ? n1683 : ~n21100;
  assign n21102 = pi19 ? n342 : n357;
  assign n21103 = pi18 ? n32 : n21102;
  assign n21104 = pi17 ? n32 : n21103;
  assign n21105 = pi20 ? n357 : n6085;
  assign n21106 = pi19 ? n21105 : n18574;
  assign n21107 = pi20 ? n274 : n333;
  assign n21108 = pi20 ? n2385 : n12884;
  assign n21109 = pi19 ? n21107 : n21108;
  assign n21110 = pi18 ? n21106 : n21109;
  assign n21111 = pi21 ? n174 : ~n405;
  assign n21112 = pi20 ? n259 : n21111;
  assign n21113 = pi20 ? n4279 : n309;
  assign n21114 = pi19 ? n21112 : ~n21113;
  assign n21115 = pi18 ? n21114 : ~n19750;
  assign n21116 = pi17 ? n21110 : ~n21115;
  assign n21117 = pi16 ? n21104 : n21116;
  assign n21118 = pi15 ? n21101 : n21117;
  assign n21119 = pi14 ? n21099 : n21118;
  assign n21120 = pi14 ? n20538 : n19758;
  assign n21121 = pi13 ? n21119 : n21120;
  assign n21122 = pi14 ? n32 : n19236;
  assign n21123 = pi15 ? n19235 : n18904;
  assign n21124 = pi15 ? n19691 : n18657;
  assign n21125 = pi14 ? n21123 : n21124;
  assign n21126 = pi13 ? n21122 : n21125;
  assign n21127 = pi12 ? n21121 : n21126;
  assign n21128 = pi11 ? n21091 : n21127;
  assign n21129 = pi10 ? n21056 : n21128;
  assign n21130 = pi09 ? n32 : n21129;
  assign n21131 = pi15 ? n32 : n14613;
  assign n21132 = pi14 ? n32 : n21131;
  assign n21133 = pi15 ? n14613 : n21033;
  assign n21134 = pi14 ? n21133 : n21035;
  assign n21135 = pi13 ? n21132 : n21134;
  assign n21136 = pi12 ? n32 : n21135;
  assign n21137 = pi20 ? n32 : n1629;
  assign n21138 = pi19 ? n21137 : n32;
  assign n21139 = pi18 ? n32 : n21138;
  assign n21140 = pi17 ? n32 : n21139;
  assign n21141 = pi16 ? n32 : n21140;
  assign n21142 = pi15 ? n21141 : n32;
  assign n21143 = pi14 ? n20967 : n21142;
  assign n21144 = pi13 ? n21143 : n32;
  assign n21145 = pi14 ? n32 : n21039;
  assign n21146 = pi15 ? n20756 : n32;
  assign n21147 = pi14 ? n21146 : n21052;
  assign n21148 = pi13 ? n21145 : n21147;
  assign n21149 = pi12 ? n21144 : n21148;
  assign n21150 = pi11 ? n21136 : n21149;
  assign n21151 = pi18 ? n880 : ~n2424;
  assign n21152 = pi17 ? n32 : n21151;
  assign n21153 = pi16 ? n32 : n21152;
  assign n21154 = pi20 ? n342 : ~n243;
  assign n21155 = pi19 ? n21154 : n32;
  assign n21156 = pi18 ? n940 : n21155;
  assign n21157 = pi17 ? n32 : n21156;
  assign n21158 = pi16 ? n32 : n21157;
  assign n21159 = pi15 ? n21153 : n21158;
  assign n21160 = pi18 ? n32 : n21155;
  assign n21161 = pi17 ? n32 : n21160;
  assign n21162 = pi16 ? n32 : n21161;
  assign n21163 = pi14 ? n21159 : n21162;
  assign n21164 = pi18 ? n4380 : n21155;
  assign n21165 = pi17 ? n32 : n21164;
  assign n21166 = pi16 ? n32 : n21165;
  assign n21167 = pi20 ? n321 : ~n243;
  assign n21168 = pi19 ? n21167 : n32;
  assign n21169 = pi18 ? n4380 : n21168;
  assign n21170 = pi17 ? n32 : n21169;
  assign n21171 = pi16 ? n32 : n21170;
  assign n21172 = pi15 ? n21166 : n21171;
  assign n21173 = pi18 ? n940 : ~n2424;
  assign n21174 = pi17 ? n32 : n21173;
  assign n21175 = pi16 ? n32 : n21174;
  assign n21176 = pi15 ? n21171 : n21175;
  assign n21177 = pi14 ? n21172 : n21176;
  assign n21178 = pi13 ? n21163 : n21177;
  assign n21179 = pi20 ? n1385 : n339;
  assign n21180 = pi19 ? n21179 : ~n32;
  assign n21181 = pi18 ? n21066 : ~n21180;
  assign n21182 = pi17 ? n32 : n21181;
  assign n21183 = pi16 ? n32 : n21182;
  assign n21184 = pi15 ? n21183 : n20779;
  assign n21185 = pi14 ? n21184 : n20048;
  assign n21186 = pi15 ? n20806 : n21079;
  assign n21187 = pi18 ? n21081 : ~n430;
  assign n21188 = pi17 ? n32 : n21187;
  assign n21189 = pi16 ? n32 : n21188;
  assign n21190 = pi15 ? n21189 : n21087;
  assign n21191 = pi14 ? n21186 : n21190;
  assign n21192 = pi13 ? n21185 : n21191;
  assign n21193 = pi12 ? n21178 : n21192;
  assign n21194 = pi19 ? n357 : n32;
  assign n21195 = pi19 ? n32 : n21108;
  assign n21196 = pi18 ? n21194 : n21195;
  assign n21197 = pi20 ? n342 : n3523;
  assign n21198 = pi19 ? n9007 : n21197;
  assign n21199 = pi18 ? n21198 : n19750;
  assign n21200 = pi17 ? n21196 : n21199;
  assign n21201 = pi16 ? n21104 : n21200;
  assign n21202 = pi15 ? n21101 : n21201;
  assign n21203 = pi14 ? n21099 : n21202;
  assign n21204 = pi15 ? n20315 : n20538;
  assign n21205 = pi14 ? n21204 : n19758;
  assign n21206 = pi13 ? n21203 : n21205;
  assign n21207 = pi15 ? n32 : n19240;
  assign n21208 = pi14 ? n19447 : n21207;
  assign n21209 = pi13 ? n21208 : n21125;
  assign n21210 = pi12 ? n21206 : n21209;
  assign n21211 = pi11 ? n21193 : n21210;
  assign n21212 = pi10 ? n21150 : n21211;
  assign n21213 = pi09 ? n32 : n21212;
  assign n21214 = pi08 ? n21130 : n21213;
  assign n21215 = pi07 ? n21028 : n21214;
  assign n21216 = pi15 ? n14613 : n14397;
  assign n21217 = pi15 ? n14397 : n32;
  assign n21218 = pi14 ? n21216 : n21217;
  assign n21219 = pi13 ? n21132 : n21218;
  assign n21220 = pi12 ? n32 : n21219;
  assign n21221 = pi21 ? n13784 : n32;
  assign n21222 = pi20 ? n32 : n21221;
  assign n21223 = pi19 ? n21222 : n32;
  assign n21224 = pi18 ? n32 : n21223;
  assign n21225 = pi17 ? n32 : n21224;
  assign n21226 = pi16 ? n32 : n21225;
  assign n21227 = pi15 ? n20836 : n21226;
  assign n21228 = pi14 ? n20836 : n21227;
  assign n21229 = pi19 ? n17257 : n32;
  assign n21230 = pi18 ? n32 : n21229;
  assign n21231 = pi17 ? n32 : n21230;
  assign n21232 = pi16 ? n32 : n21231;
  assign n21233 = pi20 ? n266 : n36;
  assign n21234 = pi19 ? n21233 : n32;
  assign n21235 = pi18 ? n863 : n21234;
  assign n21236 = pi17 ? n32 : n21235;
  assign n21237 = pi16 ? n32 : n21236;
  assign n21238 = pi15 ? n21232 : n21237;
  assign n21239 = pi18 ? n863 : n19194;
  assign n21240 = pi17 ? n32 : n21239;
  assign n21241 = pi16 ? n32 : n21240;
  assign n21242 = pi18 ? n863 : n20474;
  assign n21243 = pi17 ? n32 : n21242;
  assign n21244 = pi16 ? n32 : n21243;
  assign n21245 = pi15 ? n21241 : n21244;
  assign n21246 = pi14 ? n21238 : n21245;
  assign n21247 = pi13 ? n21228 : n21246;
  assign n21248 = pi12 ? n32 : n21247;
  assign n21249 = pi11 ? n21220 : n21248;
  assign n21250 = pi15 ? n486 : n21162;
  assign n21251 = pi14 ? n20668 : n21250;
  assign n21252 = pi18 ? n32 : n21168;
  assign n21253 = pi17 ? n32 : n21252;
  assign n21254 = pi16 ? n32 : n21253;
  assign n21255 = pi19 ? n507 : n1464;
  assign n21256 = pi20 ? n266 : n243;
  assign n21257 = pi19 ? n21256 : ~n32;
  assign n21258 = pi18 ? n21255 : ~n21257;
  assign n21259 = pi17 ? n32 : n21258;
  assign n21260 = pi16 ? n32 : n21259;
  assign n21261 = pi15 ? n21254 : n21260;
  assign n21262 = pi14 ? n21254 : n21261;
  assign n21263 = pi13 ? n21251 : n21262;
  assign n21264 = pi15 ? n20779 : n19972;
  assign n21265 = pi14 ? n20301 : n21264;
  assign n21266 = pi18 ? n20172 : n4343;
  assign n21267 = pi17 ? n32 : n21266;
  assign n21268 = pi16 ? n32 : n21267;
  assign n21269 = pi15 ? n13083 : n21268;
  assign n21270 = pi19 ? n531 : ~n4964;
  assign n21271 = pi18 ? n21270 : ~n532;
  assign n21272 = pi17 ? n32 : n21271;
  assign n21273 = pi16 ? n32 : n21272;
  assign n21274 = pi19 ? n531 : ~n4342;
  assign n21275 = pi18 ? n21274 : ~n532;
  assign n21276 = pi17 ? n32 : n21275;
  assign n21277 = pi16 ? n32 : n21276;
  assign n21278 = pi15 ? n21273 : n21277;
  assign n21279 = pi14 ? n21269 : n21278;
  assign n21280 = pi13 ? n21265 : n21279;
  assign n21281 = pi12 ? n21263 : n21280;
  assign n21282 = pi20 ? n206 : ~n321;
  assign n21283 = pi19 ? n7642 : n21282;
  assign n21284 = pi18 ? n21283 : n532;
  assign n21285 = pi17 ? n32 : ~n21284;
  assign n21286 = pi16 ? n32 : n21285;
  assign n21287 = pi19 ? n32 : n9724;
  assign n21288 = pi18 ? n21287 : n32;
  assign n21289 = pi17 ? n21288 : ~n2531;
  assign n21290 = pi16 ? n32 : n21289;
  assign n21291 = pi15 ? n21286 : n21290;
  assign n21292 = pi19 ? n5694 : ~n5694;
  assign n21293 = pi18 ? n463 : n21292;
  assign n21294 = pi17 ? n32 : n21293;
  assign n21295 = pi19 ? n321 : n6308;
  assign n21296 = pi20 ? n749 : n342;
  assign n21297 = pi19 ? n21296 : ~n247;
  assign n21298 = pi18 ? n21295 : n21297;
  assign n21299 = pi19 ? n1464 : n4126;
  assign n21300 = pi18 ? n21299 : n20628;
  assign n21301 = pi17 ? n21298 : ~n21300;
  assign n21302 = pi16 ? n21294 : n21301;
  assign n21303 = pi15 ? n21302 : n20315;
  assign n21304 = pi14 ? n21291 : n21303;
  assign n21305 = pi15 ? n20538 : n156;
  assign n21306 = pi14 ? n20315 : n21305;
  assign n21307 = pi13 ? n21304 : n21306;
  assign n21308 = pi15 ? n19996 : n19814;
  assign n21309 = pi15 ? n20646 : n18904;
  assign n21310 = pi14 ? n21308 : n21309;
  assign n21311 = pi13 ? n93 : n21310;
  assign n21312 = pi12 ? n21307 : n21311;
  assign n21313 = pi11 ? n21281 : n21312;
  assign n21314 = pi10 ? n21249 : n21313;
  assign n21315 = pi09 ? n32 : n21314;
  assign n21316 = pi19 ? n6057 : n32;
  assign n21317 = pi18 ? n32 : n21316;
  assign n21318 = pi17 ? n32 : n21317;
  assign n21319 = pi16 ? n32 : n21318;
  assign n21320 = pi15 ? n32 : n21319;
  assign n21321 = pi14 ? n32 : n21320;
  assign n21322 = pi15 ? n21319 : n14397;
  assign n21323 = pi14 ? n21322 : n21217;
  assign n21324 = pi13 ? n21321 : n21323;
  assign n21325 = pi12 ? n32 : n21324;
  assign n21326 = pi15 ? n14613 : n32;
  assign n21327 = pi14 ? n21131 : n21326;
  assign n21328 = pi13 ? n21327 : n32;
  assign n21329 = pi20 ? n266 : n357;
  assign n21330 = pi19 ? n21329 : n32;
  assign n21331 = pi18 ? n863 : n21330;
  assign n21332 = pi17 ? n32 : n21331;
  assign n21333 = pi16 ? n32 : n21332;
  assign n21334 = pi15 ? n13943 : n21333;
  assign n21335 = pi18 ? n863 : n13945;
  assign n21336 = pi17 ? n32 : n21335;
  assign n21337 = pi16 ? n32 : n21336;
  assign n21338 = pi15 ? n21241 : n21337;
  assign n21339 = pi14 ? n21334 : n21338;
  assign n21340 = pi13 ? n20836 : n21339;
  assign n21341 = pi12 ? n21328 : n21340;
  assign n21342 = pi11 ? n21325 : n21341;
  assign n21343 = pi15 ? n20660 : n13948;
  assign n21344 = pi18 ? n32 : n5749;
  assign n21345 = pi17 ? n32 : n21344;
  assign n21346 = pi16 ? n32 : n21345;
  assign n21347 = pi15 ? n20660 : n21346;
  assign n21348 = pi14 ? n21343 : n21347;
  assign n21349 = pi20 ? n266 : n207;
  assign n21350 = pi19 ? n21349 : ~n32;
  assign n21351 = pi18 ? n21255 : ~n21350;
  assign n21352 = pi17 ? n32 : n21351;
  assign n21353 = pi16 ? n32 : n21352;
  assign n21354 = pi15 ? n13369 : n21353;
  assign n21355 = pi14 ? n13369 : n21354;
  assign n21356 = pi13 ? n21348 : n21355;
  assign n21357 = pi15 ? n20477 : n13952;
  assign n21358 = pi14 ? n21357 : n20779;
  assign n21359 = pi13 ? n21358 : n21279;
  assign n21360 = pi12 ? n21356 : n21359;
  assign n21361 = pi20 ? n12884 : ~n32;
  assign n21362 = pi19 ? n21361 : ~n21282;
  assign n21363 = pi18 ? n21362 : ~n532;
  assign n21364 = pi17 ? n32 : n21363;
  assign n21365 = pi16 ? n32 : n21364;
  assign n21366 = pi15 ? n21365 : n21290;
  assign n21367 = pi15 ? n21302 : n13392;
  assign n21368 = pi14 ? n21366 : n21367;
  assign n21369 = pi20 ? n13785 : n32;
  assign n21370 = pi19 ? n21369 : n32;
  assign n21371 = pi18 ? n32 : n21370;
  assign n21372 = pi17 ? n32 : n21371;
  assign n21373 = pi16 ? n32 : n21372;
  assign n21374 = pi15 ? n13392 : n21373;
  assign n21375 = pi15 ? n19874 : n156;
  assign n21376 = pi14 ? n21374 : n21375;
  assign n21377 = pi13 ? n21368 : n21376;
  assign n21378 = pi15 ? n32 : n20955;
  assign n21379 = pi14 ? n19932 : n21378;
  assign n21380 = pi13 ? n21379 : n21310;
  assign n21381 = pi12 ? n21377 : n21380;
  assign n21382 = pi11 ? n21360 : n21381;
  assign n21383 = pi10 ? n21342 : n21382;
  assign n21384 = pi09 ? n32 : n21383;
  assign n21385 = pi08 ? n21315 : n21384;
  assign n21386 = pi19 ? n18218 : n32;
  assign n21387 = pi18 ? n32 : n21386;
  assign n21388 = pi17 ? n32 : n21387;
  assign n21389 = pi16 ? n32 : n21388;
  assign n21390 = pi15 ? n21319 : n21389;
  assign n21391 = pi15 ? n21389 : n32;
  assign n21392 = pi14 ? n21390 : n21391;
  assign n21393 = pi13 ? n21321 : n21392;
  assign n21394 = pi12 ? n32 : n21393;
  assign n21395 = pi14 ? n14613 : n21133;
  assign n21396 = pi20 ? n266 : ~n1940;
  assign n21397 = pi19 ? n21396 : n32;
  assign n21398 = pi18 ? n863 : n21397;
  assign n21399 = pi17 ? n32 : n21398;
  assign n21400 = pi16 ? n32 : n21399;
  assign n21401 = pi15 ? n13943 : n21400;
  assign n21402 = pi15 ? n21400 : n32;
  assign n21403 = pi14 ? n21401 : n21402;
  assign n21404 = pi13 ? n21395 : n21403;
  assign n21405 = pi12 ? n32 : n21404;
  assign n21406 = pi11 ? n21394 : n21405;
  assign n21407 = pi15 ? n13948 : n21346;
  assign n21408 = pi14 ? n13948 : n21407;
  assign n21409 = pi18 ? n16316 : n5005;
  assign n21410 = pi17 ? n32 : n21409;
  assign n21411 = pi16 ? n32 : n21410;
  assign n21412 = pi20 ? n32 : n174;
  assign n21413 = pi20 ? n357 : n428;
  assign n21414 = pi19 ? n21412 : n21413;
  assign n21415 = pi20 ? n2385 : ~n207;
  assign n21416 = pi19 ? n21415 : n32;
  assign n21417 = pi18 ? n21414 : n21416;
  assign n21418 = pi17 ? n32 : n21417;
  assign n21419 = pi16 ? n32 : n21418;
  assign n21420 = pi15 ? n21411 : n21419;
  assign n21421 = pi14 ? n13369 : n21420;
  assign n21422 = pi13 ? n21408 : n21421;
  assign n21423 = pi15 ? n20477 : n21162;
  assign n21424 = pi14 ? n21423 : n20779;
  assign n21425 = pi19 ? n507 : n358;
  assign n21426 = pi18 ? n21425 : n13075;
  assign n21427 = pi17 ? n32 : n21426;
  assign n21428 = pi16 ? n32 : n21427;
  assign n21429 = pi18 ? n20172 : n13377;
  assign n21430 = pi17 ? n32 : n21429;
  assign n21431 = pi16 ? n32 : n21430;
  assign n21432 = pi15 ? n21428 : n21431;
  assign n21433 = pi18 ? n21270 : ~n3786;
  assign n21434 = pi17 ? n32 : n21433;
  assign n21435 = pi16 ? n32 : n21434;
  assign n21436 = pi18 ? n21274 : ~n3786;
  assign n21437 = pi17 ? n32 : n21436;
  assign n21438 = pi16 ? n32 : n21437;
  assign n21439 = pi15 ? n21435 : n21438;
  assign n21440 = pi14 ? n21432 : n21439;
  assign n21441 = pi13 ? n21424 : n21440;
  assign n21442 = pi12 ? n21422 : n21441;
  assign n21443 = pi19 ? n6298 : ~n6988;
  assign n21444 = pi18 ? n21443 : ~n3786;
  assign n21445 = pi17 ? n32 : n21444;
  assign n21446 = pi16 ? n32 : n21445;
  assign n21447 = pi18 ? n532 : ~n3786;
  assign n21448 = pi17 ? n32 : n21447;
  assign n21449 = pi16 ? n32 : n21448;
  assign n21450 = pi15 ? n21446 : n21449;
  assign n21451 = pi15 ? n19969 : n13392;
  assign n21452 = pi14 ? n21450 : n21451;
  assign n21453 = pi14 ? n20139 : n19862;
  assign n21454 = pi13 ? n21452 : n21453;
  assign n21455 = pi14 ? n32 : n19925;
  assign n21456 = pi15 ? n19805 : n19384;
  assign n21457 = pi15 ? n19996 : n18904;
  assign n21458 = pi14 ? n21456 : n21457;
  assign n21459 = pi13 ? n21455 : n21458;
  assign n21460 = pi12 ? n21454 : n21459;
  assign n21461 = pi11 ? n21442 : n21460;
  assign n21462 = pi10 ? n21406 : n21461;
  assign n21463 = pi09 ? n32 : n21462;
  assign n21464 = pi16 ? n32 : n2280;
  assign n21465 = pi15 ? n32 : n21464;
  assign n21466 = pi14 ? n32 : n21465;
  assign n21467 = pi15 ? n21464 : n32;
  assign n21468 = pi14 ? n21464 : n21467;
  assign n21469 = pi13 ? n21466 : n21468;
  assign n21470 = pi12 ? n32 : n21469;
  assign n21471 = pi14 ? n21320 : n32;
  assign n21472 = pi13 ? n21471 : n32;
  assign n21473 = pi15 ? n14613 : n14405;
  assign n21474 = pi14 ? n21131 : n21473;
  assign n21475 = pi20 ? n32 : ~n16176;
  assign n21476 = pi19 ? n21475 : n32;
  assign n21477 = pi18 ? n32 : n21476;
  assign n21478 = pi17 ? n32 : n21477;
  assign n21479 = pi16 ? n32 : n21478;
  assign n21480 = pi15 ? n21479 : n21400;
  assign n21481 = pi15 ? n21400 : n20831;
  assign n21482 = pi14 ? n21480 : n21481;
  assign n21483 = pi13 ? n21474 : n21482;
  assign n21484 = pi12 ? n21472 : n21483;
  assign n21485 = pi11 ? n21470 : n21484;
  assign n21486 = pi20 ? n342 : ~n1940;
  assign n21487 = pi19 ? n21486 : n32;
  assign n21488 = pi18 ? n32 : n21487;
  assign n21489 = pi17 ? n32 : n21488;
  assign n21490 = pi16 ? n32 : n21489;
  assign n21491 = pi15 ? n21232 : n21490;
  assign n21492 = pi14 ? n21232 : n21491;
  assign n21493 = pi20 ? n321 : ~n1940;
  assign n21494 = pi19 ? n21493 : n32;
  assign n21495 = pi18 ? n32 : n21494;
  assign n21496 = pi17 ? n32 : n21495;
  assign n21497 = pi16 ? n32 : n21496;
  assign n21498 = pi18 ? n16316 : n21494;
  assign n21499 = pi17 ? n32 : n21498;
  assign n21500 = pi16 ? n32 : n21499;
  assign n21501 = pi20 ? n2385 : n17449;
  assign n21502 = pi19 ? n21501 : n32;
  assign n21503 = pi18 ? n8106 : n21502;
  assign n21504 = pi17 ? n32 : n21503;
  assign n21505 = pi16 ? n32 : n21504;
  assign n21506 = pi15 ? n21500 : n21505;
  assign n21507 = pi14 ? n21497 : n21506;
  assign n21508 = pi13 ? n21492 : n21507;
  assign n21509 = pi15 ? n20486 : n21162;
  assign n21510 = pi14 ? n21509 : n13671;
  assign n21511 = pi18 ? n21425 : n13080;
  assign n21512 = pi17 ? n32 : n21511;
  assign n21513 = pi16 ? n32 : n21512;
  assign n21514 = pi15 ? n21513 : n21268;
  assign n21515 = pi14 ? n21514 : n21278;
  assign n21516 = pi13 ? n21510 : n21515;
  assign n21517 = pi12 ? n21508 : n21516;
  assign n21518 = pi19 ? n6324 : n32;
  assign n21519 = pi18 ? n32 : n21518;
  assign n21520 = pi17 ? n32 : n21519;
  assign n21521 = pi16 ? n32 : n21520;
  assign n21522 = pi15 ? n20048 : n21521;
  assign n21523 = pi14 ? n21450 : n21522;
  assign n21524 = pi15 ? n19972 : n180;
  assign n21525 = pi14 ? n21524 : n20140;
  assign n21526 = pi13 ? n21523 : n21525;
  assign n21527 = pi14 ? n19755 : n19925;
  assign n21528 = pi15 ? n19996 : n20646;
  assign n21529 = pi14 ? n21456 : n21528;
  assign n21530 = pi13 ? n21527 : n21529;
  assign n21531 = pi12 ? n21526 : n21530;
  assign n21532 = pi11 ? n21517 : n21531;
  assign n21533 = pi10 ? n21485 : n21532;
  assign n21534 = pi09 ? n32 : n21533;
  assign n21535 = pi08 ? n21463 : n21534;
  assign n21536 = pi07 ? n21385 : n21535;
  assign n21537 = pi06 ? n21215 : n21536;
  assign n21538 = pi05 ? n20827 : n21537;
  assign n21539 = pi04 ? n20122 : n21538;
  assign n21540 = pi03 ? n18881 : n21539;
  assign n21541 = pi18 ? n32 : n9578;
  assign n21542 = pi17 ? n32 : n21541;
  assign n21543 = pi16 ? n32 : n21542;
  assign n21544 = pi14 ? n21543 : n21467;
  assign n21545 = pi13 ? n21466 : n21544;
  assign n21546 = pi12 ? n32 : n21545;
  assign n21547 = pi14 ? n14397 : n21322;
  assign n21548 = pi19 ? n17212 : n32;
  assign n21549 = pi18 ? n32 : n21548;
  assign n21550 = pi17 ? n32 : n21549;
  assign n21551 = pi16 ? n32 : n21550;
  assign n21552 = pi15 ? n21551 : n13943;
  assign n21553 = pi15 ? n13943 : n32;
  assign n21554 = pi14 ? n21552 : n21553;
  assign n21555 = pi13 ? n21547 : n21554;
  assign n21556 = pi12 ? n32 : n21555;
  assign n21557 = pi11 ? n21546 : n21556;
  assign n21558 = pi15 ? n13948 : n32;
  assign n21559 = pi14 ? n21558 : n21346;
  assign n21560 = pi15 ? n21490 : n21497;
  assign n21561 = pi20 ? n428 : ~n1940;
  assign n21562 = pi19 ? n21561 : n32;
  assign n21563 = pi18 ? n32 : n21562;
  assign n21564 = pi17 ? n32 : n21563;
  assign n21565 = pi16 ? n32 : n21564;
  assign n21566 = pi14 ? n21560 : n21565;
  assign n21567 = pi13 ? n21559 : n21566;
  assign n21568 = pi19 ? n7349 : n32;
  assign n21569 = pi18 ? n32 : n21568;
  assign n21570 = pi17 ? n32 : n21569;
  assign n21571 = pi16 ? n32 : n21570;
  assign n21572 = pi15 ? n21571 : n13948;
  assign n21573 = pi18 ? n16449 : n13668;
  assign n21574 = pi17 ? n32 : n21573;
  assign n21575 = pi16 ? n32 : n21574;
  assign n21576 = pi19 ? n32 : ~n4406;
  assign n21577 = pi18 ? n21576 : n13668;
  assign n21578 = pi17 ? n32 : n21577;
  assign n21579 = pi16 ? n32 : n21578;
  assign n21580 = pi15 ? n21575 : n21579;
  assign n21581 = pi14 ? n21572 : n21580;
  assign n21582 = pi18 ? n17058 : n32;
  assign n21583 = pi18 ? n350 : ~n418;
  assign n21584 = pi17 ? n21582 : n21583;
  assign n21585 = pi16 ? n32 : n21584;
  assign n21586 = pi20 ? n32 : ~n354;
  assign n21587 = pi19 ? n32 : n21586;
  assign n21588 = pi20 ? n9641 : n32;
  assign n21589 = pi19 ? n17665 : n21588;
  assign n21590 = pi18 ? n21587 : n21589;
  assign n21591 = pi18 ? n6063 : ~n418;
  assign n21592 = pi17 ? n21590 : n21591;
  assign n21593 = pi16 ? n32 : n21592;
  assign n21594 = pi15 ? n21585 : n21593;
  assign n21595 = pi19 ? n322 : ~n4670;
  assign n21596 = pi20 ? n207 : ~n339;
  assign n21597 = pi19 ? n21596 : n32;
  assign n21598 = pi18 ? n21595 : n21597;
  assign n21599 = pi17 ? n32 : n21598;
  assign n21600 = pi16 ? n32 : n21599;
  assign n21601 = pi18 ? n323 : ~n418;
  assign n21602 = pi17 ? n32 : n21601;
  assign n21603 = pi16 ? n32 : n21602;
  assign n21604 = pi15 ? n21600 : n21603;
  assign n21605 = pi14 ? n21594 : n21604;
  assign n21606 = pi13 ? n21581 : n21605;
  assign n21607 = pi12 ? n21567 : n21606;
  assign n21608 = pi15 ? n13375 : n20301;
  assign n21609 = pi14 ? n21608 : n19972;
  assign n21610 = pi14 ? n21524 : n19862;
  assign n21611 = pi13 ? n21609 : n21610;
  assign n21612 = pi15 ? n116 : n19868;
  assign n21613 = pi14 ? n32 : n21612;
  assign n21614 = pi14 ? n19983 : n19621;
  assign n21615 = pi13 ? n21613 : n21614;
  assign n21616 = pi12 ? n21611 : n21615;
  assign n21617 = pi11 ? n21607 : n21616;
  assign n21618 = pi10 ? n21557 : n21617;
  assign n21619 = pi09 ? n32 : n21618;
  assign n21620 = pi15 ? n32 : n387;
  assign n21621 = pi14 ? n32 : n21620;
  assign n21622 = pi14 ? n21543 : n388;
  assign n21623 = pi13 ? n21621 : n21622;
  assign n21624 = pi12 ? n32 : n21623;
  assign n21625 = pi14 ? n21465 : n32;
  assign n21626 = pi13 ? n21625 : n32;
  assign n21627 = pi15 ? n658 : n21319;
  assign n21628 = pi14 ? n14397 : n21627;
  assign n21629 = pi15 ? n14156 : n13943;
  assign n21630 = pi15 ? n13943 : n20836;
  assign n21631 = pi14 ? n21629 : n21630;
  assign n21632 = pi13 ? n21628 : n21631;
  assign n21633 = pi12 ? n21626 : n21632;
  assign n21634 = pi11 ? n21624 : n21633;
  assign n21635 = pi14 ? n21630 : n13660;
  assign n21636 = pi15 ? n13660 : n13360;
  assign n21637 = pi20 ? n428 : ~n749;
  assign n21638 = pi19 ? n21637 : n32;
  assign n21639 = pi18 ? n32 : n21638;
  assign n21640 = pi17 ? n32 : n21639;
  assign n21641 = pi16 ? n32 : n21640;
  assign n21642 = pi14 ? n21636 : n21641;
  assign n21643 = pi13 ? n21635 : n21642;
  assign n21644 = pi18 ? n16449 : n21155;
  assign n21645 = pi17 ? n32 : n21644;
  assign n21646 = pi16 ? n32 : n21645;
  assign n21647 = pi18 ? n21576 : n21155;
  assign n21648 = pi17 ? n32 : n21647;
  assign n21649 = pi16 ? n32 : n21648;
  assign n21650 = pi15 ? n21646 : n21649;
  assign n21651 = pi14 ? n21572 : n21650;
  assign n21652 = pi19 ? n32 : ~n19246;
  assign n21653 = pi18 ? n858 : n21652;
  assign n21654 = pi17 ? n32 : n21653;
  assign n21655 = pi20 ? n1331 : ~n6050;
  assign n21656 = pi19 ? n1331 : n21655;
  assign n21657 = pi20 ? n9641 : n3523;
  assign n21658 = pi19 ? n17665 : n21657;
  assign n21659 = pi18 ? n21656 : n21658;
  assign n21660 = pi20 ? n13171 : ~n207;
  assign n21661 = pi19 ? n21660 : n32;
  assign n21662 = pi18 ? n21661 : n418;
  assign n21663 = pi17 ? n21659 : ~n21662;
  assign n21664 = pi16 ? n21654 : n21663;
  assign n21665 = pi15 ? n21585 : n21664;
  assign n21666 = pi14 ? n21665 : n21604;
  assign n21667 = pi13 ? n21651 : n21666;
  assign n21668 = pi12 ? n21643 : n21667;
  assign n21669 = pi14 ? n21608 : n20779;
  assign n21670 = pi15 ? n20779 : n13392;
  assign n21671 = pi14 ? n21670 : n20139;
  assign n21672 = pi13 ? n21669 : n21671;
  assign n21673 = pi14 ? n32 : n19869;
  assign n21674 = pi14 ? n19983 : n21456;
  assign n21675 = pi13 ? n21673 : n21674;
  assign n21676 = pi12 ? n21672 : n21675;
  assign n21677 = pi11 ? n21668 : n21676;
  assign n21678 = pi10 ? n21634 : n21677;
  assign n21679 = pi09 ? n32 : n21678;
  assign n21680 = pi08 ? n21619 : n21679;
  assign n21681 = pi15 ? n32 : n21543;
  assign n21682 = pi14 ? n32 : n21681;
  assign n21683 = pi19 ? n17713 : n32;
  assign n21684 = pi18 ? n32 : n21683;
  assign n21685 = pi17 ? n32 : n21684;
  assign n21686 = pi16 ? n32 : n21685;
  assign n21687 = pi15 ? n21686 : n21543;
  assign n21688 = pi14 ? n21687 : n388;
  assign n21689 = pi13 ? n21682 : n21688;
  assign n21690 = pi12 ? n32 : n21689;
  assign n21691 = pi13 ? n32 : n21466;
  assign n21692 = pi19 ? n17982 : n32;
  assign n21693 = pi18 ? n32 : n21692;
  assign n21694 = pi17 ? n32 : n21693;
  assign n21695 = pi16 ? n32 : n21694;
  assign n21696 = pi15 ? n21695 : n21464;
  assign n21697 = pi15 ? n21695 : n14397;
  assign n21698 = pi14 ? n21696 : n21697;
  assign n21699 = pi20 ? n32 : ~n11048;
  assign n21700 = pi19 ? n21699 : n32;
  assign n21701 = pi18 ? n32 : n21700;
  assign n21702 = pi17 ? n32 : n21701;
  assign n21703 = pi16 ? n32 : n21702;
  assign n21704 = pi15 ? n14156 : n21703;
  assign n21705 = pi14 ? n21704 : n21326;
  assign n21706 = pi13 ? n21698 : n21705;
  assign n21707 = pi12 ? n21691 : n21706;
  assign n21708 = pi11 ? n21690 : n21707;
  assign n21709 = pi18 ? n17767 : n13657;
  assign n21710 = pi17 ? n32 : n21709;
  assign n21711 = pi16 ? n32 : n21710;
  assign n21712 = pi18 ? n16389 : n13940;
  assign n21713 = pi17 ? n32 : n21712;
  assign n21714 = pi16 ? n32 : n21713;
  assign n21715 = pi15 ? n21711 : n21714;
  assign n21716 = pi14 ? n21630 : n21715;
  assign n21717 = pi18 ? n16603 : n5164;
  assign n21718 = pi17 ? n32 : n21717;
  assign n21719 = pi16 ? n32 : n21718;
  assign n21720 = pi15 ? n21641 : n21719;
  assign n21721 = pi14 ? n21720 : n13943;
  assign n21722 = pi13 ? n21716 : n21721;
  assign n21723 = pi20 ? n342 : n481;
  assign n21724 = pi19 ? n21723 : n32;
  assign n21725 = pi18 ? n16449 : n21724;
  assign n21726 = pi17 ? n32 : n21725;
  assign n21727 = pi16 ? n32 : n21726;
  assign n21728 = pi18 ? n15227 : n21155;
  assign n21729 = pi17 ? n32 : n21728;
  assign n21730 = pi16 ? n32 : n21729;
  assign n21731 = pi15 ? n21727 : n21730;
  assign n21732 = pi14 ? n13948 : n21731;
  assign n21733 = pi18 ? n350 : ~n2424;
  assign n21734 = pi17 ? n17734 : n21733;
  assign n21735 = pi16 ? n32 : n21734;
  assign n21736 = pi20 ? n357 : n12884;
  assign n21737 = pi19 ? n32 : n21736;
  assign n21738 = pi18 ? n936 : n21737;
  assign n21739 = pi17 ? n32 : n21738;
  assign n21740 = pi20 ? n246 : n220;
  assign n21741 = pi19 ? n246 : n21740;
  assign n21742 = pi20 ? n246 : ~n2385;
  assign n21743 = pi19 ? n21742 : ~n7089;
  assign n21744 = pi18 ? n21741 : ~n21743;
  assign n21745 = pi18 ? n6059 : n2424;
  assign n21746 = pi17 ? n21744 : ~n21745;
  assign n21747 = pi16 ? n21739 : n21746;
  assign n21748 = pi15 ? n21735 : n21747;
  assign n21749 = pi19 ? n11991 : ~n32;
  assign n21750 = pi18 ? n323 : ~n21749;
  assign n21751 = pi17 ? n32 : n21750;
  assign n21752 = pi16 ? n32 : n21751;
  assign n21753 = pi18 ? n323 : ~n2424;
  assign n21754 = pi17 ? n32 : n21753;
  assign n21755 = pi16 ? n32 : n21754;
  assign n21756 = pi15 ? n21752 : n21755;
  assign n21757 = pi14 ? n21748 : n21756;
  assign n21758 = pi13 ? n21732 : n21757;
  assign n21759 = pi12 ? n21722 : n21758;
  assign n21760 = pi18 ? n16389 : n21168;
  assign n21761 = pi17 ? n32 : n21760;
  assign n21762 = pi16 ? n32 : n21761;
  assign n21763 = pi15 ? n21762 : n13671;
  assign n21764 = pi14 ? n21763 : n13684;
  assign n21765 = pi15 ? n13684 : n19969;
  assign n21766 = pi14 ? n21765 : n19977;
  assign n21767 = pi13 ? n21764 : n21766;
  assign n21768 = pi15 ? n180 : n20531;
  assign n21769 = pi14 ? n181 : n21768;
  assign n21770 = pi15 ? n20531 : n19805;
  assign n21771 = pi19 ? n16511 : n32;
  assign n21772 = pi18 ? n32 : n21771;
  assign n21773 = pi17 ? n32 : n21772;
  assign n21774 = pi16 ? n32 : n21773;
  assign n21775 = pi19 ? n1740 : ~n6308;
  assign n21776 = pi18 ? n21775 : ~n2318;
  assign n21777 = pi17 ? n464 : n21776;
  assign n21778 = pi16 ? n32 : n21777;
  assign n21779 = pi15 ? n21774 : n21778;
  assign n21780 = pi14 ? n21770 : n21779;
  assign n21781 = pi13 ? n21769 : n21780;
  assign n21782 = pi12 ? n21767 : n21781;
  assign n21783 = pi11 ? n21759 : n21782;
  assign n21784 = pi10 ? n21708 : n21783;
  assign n21785 = pi09 ? n32 : n21784;
  assign n21786 = pi16 ? n32 : n2095;
  assign n21787 = pi15 ? n32 : n21786;
  assign n21788 = pi14 ? n32 : n21787;
  assign n21789 = pi15 ? n21686 : n21786;
  assign n21790 = pi15 ? n21786 : n32;
  assign n21791 = pi14 ? n21789 : n21790;
  assign n21792 = pi13 ? n21788 : n21791;
  assign n21793 = pi12 ? n32 : n21792;
  assign n21794 = pi14 ? n21543 : n32;
  assign n21795 = pi13 ? n21794 : n32;
  assign n21796 = pi15 ? n14397 : n21464;
  assign n21797 = pi14 ? n21796 : n21695;
  assign n21798 = pi19 ? n7795 : n32;
  assign n21799 = pi18 ? n32 : n21798;
  assign n21800 = pi17 ? n32 : n21799;
  assign n21801 = pi16 ? n32 : n21800;
  assign n21802 = pi15 ? n21801 : n21703;
  assign n21803 = pi14 ? n21802 : n14613;
  assign n21804 = pi13 ? n21797 : n21803;
  assign n21805 = pi12 ? n21795 : n21804;
  assign n21806 = pi11 ? n21793 : n21805;
  assign n21807 = pi15 ? n21551 : n21033;
  assign n21808 = pi19 ? n16820 : n32;
  assign n21809 = pi18 ? n17767 : n21808;
  assign n21810 = pi17 ? n32 : n21809;
  assign n21811 = pi16 ? n32 : n21810;
  assign n21812 = pi18 ? n16389 : n21548;
  assign n21813 = pi17 ? n32 : n21812;
  assign n21814 = pi16 ? n32 : n21813;
  assign n21815 = pi15 ? n21811 : n21814;
  assign n21816 = pi14 ? n21807 : n21815;
  assign n21817 = pi20 ? n321 : ~n1475;
  assign n21818 = pi19 ? n21817 : n32;
  assign n21819 = pi18 ? n16603 : n21818;
  assign n21820 = pi17 ? n32 : n21819;
  assign n21821 = pi16 ? n32 : n21820;
  assign n21822 = pi15 ? n13930 : n21821;
  assign n21823 = pi14 ? n21822 : n21551;
  assign n21824 = pi13 ? n21816 : n21823;
  assign n21825 = pi18 ? n16449 : n17650;
  assign n21826 = pi17 ? n32 : n21825;
  assign n21827 = pi16 ? n32 : n21826;
  assign n21828 = pi18 ? n15227 : n13668;
  assign n21829 = pi17 ? n32 : n21828;
  assign n21830 = pi16 ? n32 : n21829;
  assign n21831 = pi15 ? n21827 : n21830;
  assign n21832 = pi14 ? n21232 : n21831;
  assign n21833 = pi13 ? n21832 : n21757;
  assign n21834 = pi12 ? n21824 : n21833;
  assign n21835 = pi15 ? n21762 : n21162;
  assign n21836 = pi14 ? n21835 : n20301;
  assign n21837 = pi14 ? n20126 : n19977;
  assign n21838 = pi13 ? n21836 : n21837;
  assign n21839 = pi15 ? n20531 : n19868;
  assign n21840 = pi18 ? n21775 : ~n344;
  assign n21841 = pi17 ? n464 : n21840;
  assign n21842 = pi16 ? n32 : n21841;
  assign n21843 = pi15 ? n19868 : n21842;
  assign n21844 = pi14 ? n21839 : n21843;
  assign n21845 = pi13 ? n21769 : n21844;
  assign n21846 = pi12 ? n21838 : n21845;
  assign n21847 = pi11 ? n21834 : n21846;
  assign n21848 = pi10 ? n21806 : n21847;
  assign n21849 = pi09 ? n32 : n21848;
  assign n21850 = pi08 ? n21785 : n21849;
  assign n21851 = pi07 ? n21680 : n21850;
  assign n21852 = pi17 ? n32 : n20021;
  assign n21853 = pi16 ? n32 : n21852;
  assign n21854 = pi15 ? n21853 : n21786;
  assign n21855 = pi14 ? n21854 : n32;
  assign n21856 = pi13 ? n21788 : n21855;
  assign n21857 = pi12 ? n32 : n21856;
  assign n21858 = pi15 ? n387 : n21543;
  assign n21859 = pi20 ? n32 : ~n1377;
  assign n21860 = pi19 ? n21859 : n32;
  assign n21861 = pi18 ? n32 : n21860;
  assign n21862 = pi17 ? n32 : n21861;
  assign n21863 = pi16 ? n32 : n21862;
  assign n21864 = pi15 ? n14394 : n21863;
  assign n21865 = pi14 ? n21858 : n21864;
  assign n21866 = pi15 ? n21319 : n14613;
  assign n21867 = pi14 ? n21697 : n21866;
  assign n21868 = pi13 ? n21865 : n21867;
  assign n21869 = pi12 ? n32 : n21868;
  assign n21870 = pi11 ? n21857 : n21869;
  assign n21871 = pi14 ? n14613 : n21035;
  assign n21872 = pi18 ? n15844 : n21548;
  assign n21873 = pi17 ? n32 : n21872;
  assign n21874 = pi16 ? n32 : n21873;
  assign n21875 = pi18 ? n16316 : n14161;
  assign n21876 = pi17 ? n32 : n21875;
  assign n21877 = pi16 ? n32 : n21876;
  assign n21878 = pi15 ? n21874 : n21877;
  assign n21879 = pi14 ? n21878 : n21551;
  assign n21880 = pi13 ? n21871 : n21879;
  assign n21881 = pi18 ? n15844 : n20753;
  assign n21882 = pi17 ? n32 : n21881;
  assign n21883 = pi16 ? n32 : n21882;
  assign n21884 = pi15 ? n20756 : n21883;
  assign n21885 = pi18 ? n16234 : n5749;
  assign n21886 = pi17 ? n32 : n21885;
  assign n21887 = pi16 ? n32 : n21886;
  assign n21888 = pi19 ? n32 : ~n208;
  assign n21889 = pi18 ? n21888 : n13945;
  assign n21890 = pi17 ? n32 : n21889;
  assign n21891 = pi16 ? n32 : n21890;
  assign n21892 = pi15 ? n21887 : n21891;
  assign n21893 = pi14 ? n21884 : n21892;
  assign n21894 = pi18 ? n532 : ~n605;
  assign n21895 = pi17 ? n18316 : n21894;
  assign n21896 = pi16 ? n32 : n21895;
  assign n21897 = pi18 ? n605 : ~n605;
  assign n21898 = pi17 ? n18316 : n21897;
  assign n21899 = pi16 ? n32 : n21898;
  assign n21900 = pi15 ? n21896 : n21899;
  assign n21901 = pi18 ? n21595 : ~n605;
  assign n21902 = pi17 ? n32 : n21901;
  assign n21903 = pi16 ? n32 : n21902;
  assign n21904 = pi15 ? n11426 : n21903;
  assign n21905 = pi14 ? n21900 : n21904;
  assign n21906 = pi13 ? n21893 : n21905;
  assign n21907 = pi12 ? n21880 : n21906;
  assign n21908 = pi14 ? n20477 : n20301;
  assign n21909 = pi14 ? n20126 : n32;
  assign n21910 = pi13 ? n21908 : n21909;
  assign n21911 = pi14 ? n19970 : n21451;
  assign n21912 = pi15 ? n19856 : n20538;
  assign n21913 = pi18 ? n16432 : n19865;
  assign n21914 = pi17 ? n32 : n21913;
  assign n21915 = pi16 ? n32 : n21914;
  assign n21916 = pi18 ? n15844 : n248;
  assign n21917 = pi17 ? n32 : n21916;
  assign n21918 = pi16 ? n32 : n21917;
  assign n21919 = pi15 ? n21915 : n21918;
  assign n21920 = pi14 ? n21912 : n21919;
  assign n21921 = pi13 ? n21911 : n21920;
  assign n21922 = pi12 ? n21910 : n21921;
  assign n21923 = pi11 ? n21907 : n21922;
  assign n21924 = pi10 ? n21870 : n21923;
  assign n21925 = pi09 ? n32 : n21924;
  assign n21926 = pi18 ? n32 : n6399;
  assign n21927 = pi17 ? n32 : n21926;
  assign n21928 = pi16 ? n32 : n21927;
  assign n21929 = pi15 ? n32 : n21928;
  assign n21930 = pi14 ? n32 : n21929;
  assign n21931 = pi15 ? n21853 : n476;
  assign n21932 = pi14 ? n21931 : n32;
  assign n21933 = pi13 ? n21930 : n21932;
  assign n21934 = pi12 ? n32 : n21933;
  assign n21935 = pi14 ? n21786 : n32;
  assign n21936 = pi13 ? n21935 : n32;
  assign n21937 = pi20 ? n32 : ~n6886;
  assign n21938 = pi19 ? n21937 : n32;
  assign n21939 = pi18 ? n32 : n21938;
  assign n21940 = pi17 ? n32 : n21939;
  assign n21941 = pi16 ? n32 : n21940;
  assign n21942 = pi15 ? n14394 : n21941;
  assign n21943 = pi14 ? n21543 : n21942;
  assign n21944 = pi14 ? n21697 : n21319;
  assign n21945 = pi13 ? n21943 : n21944;
  assign n21946 = pi12 ? n21936 : n21945;
  assign n21947 = pi11 ? n21934 : n21946;
  assign n21948 = pi14 ? n21319 : n14397;
  assign n21949 = pi18 ? n15844 : n14153;
  assign n21950 = pi17 ? n32 : n21949;
  assign n21951 = pi16 ? n32 : n21950;
  assign n21952 = pi18 ? n32 : n20729;
  assign n21953 = pi17 ? n32 : n21952;
  assign n21954 = pi16 ? n32 : n21953;
  assign n21955 = pi15 ? n21951 : n21954;
  assign n21956 = pi15 ? n14156 : n21551;
  assign n21957 = pi14 ? n21955 : n21956;
  assign n21958 = pi13 ? n21948 : n21957;
  assign n21959 = pi18 ? n15844 : n20828;
  assign n21960 = pi17 ? n32 : n21959;
  assign n21961 = pi16 ? n32 : n21960;
  assign n21962 = pi15 ? n20836 : n21961;
  assign n21963 = pi14 ? n21962 : n21892;
  assign n21964 = pi13 ? n21963 : n21905;
  assign n21965 = pi12 ? n21958 : n21964;
  assign n21966 = pi18 ? n32 : n21048;
  assign n21967 = pi17 ? n32 : n21966;
  assign n21968 = pi16 ? n32 : n21967;
  assign n21969 = pi20 ? n101 : ~n243;
  assign n21970 = pi19 ? n21969 : n32;
  assign n21971 = pi18 ? n32 : n21970;
  assign n21972 = pi17 ? n32 : n21971;
  assign n21973 = pi16 ? n32 : n21972;
  assign n21974 = pi15 ? n21968 : n21973;
  assign n21975 = pi14 ? n21343 : n21974;
  assign n21976 = pi19 ? n17166 : n32;
  assign n21977 = pi18 ? n32 : n21976;
  assign n21978 = pi17 ? n32 : n21977;
  assign n21979 = pi16 ? n32 : n21978;
  assign n21980 = pi19 ? n17086 : n32;
  assign n21981 = pi18 ? n32 : n21980;
  assign n21982 = pi17 ? n32 : n21981;
  assign n21983 = pi16 ? n32 : n21982;
  assign n21984 = pi15 ? n21979 : n21983;
  assign n21985 = pi14 ? n21984 : n107;
  assign n21986 = pi13 ? n21975 : n21985;
  assign n21987 = pi18 ? n16432 : n19750;
  assign n21988 = pi17 ? n32 : n21987;
  assign n21989 = pi16 ? n32 : n21988;
  assign n21990 = pi18 ? n15844 : n19865;
  assign n21991 = pi17 ? n32 : n21990;
  assign n21992 = pi16 ? n32 : n21991;
  assign n21993 = pi15 ? n21989 : n21992;
  assign n21994 = pi14 ? n21374 : n21993;
  assign n21995 = pi13 ? n20231 : n21994;
  assign n21996 = pi12 ? n21986 : n21995;
  assign n21997 = pi11 ? n21965 : n21996;
  assign n21998 = pi10 ? n21947 : n21997;
  assign n21999 = pi09 ? n32 : n21998;
  assign n22000 = pi08 ? n21925 : n21999;
  assign n22001 = pi13 ? n32 : n478;
  assign n22002 = pi12 ? n32 : n22001;
  assign n22003 = pi19 ? n17718 : n32;
  assign n22004 = pi18 ? n32 : n22003;
  assign n22005 = pi17 ? n32 : n22004;
  assign n22006 = pi16 ? n32 : n22005;
  assign n22007 = pi15 ? n22006 : n14394;
  assign n22008 = pi14 ? n21786 : n22007;
  assign n22009 = pi15 ? n21543 : n21464;
  assign n22010 = pi14 ? n22009 : n32;
  assign n22011 = pi13 ? n22008 : n22010;
  assign n22012 = pi12 ? n32 : n22011;
  assign n22013 = pi11 ? n22002 : n22012;
  assign n22014 = pi15 ? n21951 : n14397;
  assign n22015 = pi15 ? n14156 : n21033;
  assign n22016 = pi14 ? n22014 : n22015;
  assign n22017 = pi13 ? n14397 : n22016;
  assign n22018 = pi15 ? n13943 : n21961;
  assign n22019 = pi20 ? n342 : n52;
  assign n22020 = pi19 ? n22019 : n32;
  assign n22021 = pi18 ? n16234 : n22020;
  assign n22022 = pi17 ? n32 : n22021;
  assign n22023 = pi16 ? n32 : n22022;
  assign n22024 = pi20 ? n207 : n1940;
  assign n22025 = pi19 ? n22024 : ~n32;
  assign n22026 = pi18 ? n21888 : ~n22025;
  assign n22027 = pi17 ? n32 : n22026;
  assign n22028 = pi16 ? n32 : n22027;
  assign n22029 = pi15 ? n22023 : n22028;
  assign n22030 = pi14 ? n22018 : n22029;
  assign n22031 = pi18 ? n532 : ~n2413;
  assign n22032 = pi17 ? n19262 : n22031;
  assign n22033 = pi16 ? n32 : n22032;
  assign n22034 = pi18 ? n702 : ~n2413;
  assign n22035 = pi17 ? n32 : n22034;
  assign n22036 = pi16 ? n32 : n22035;
  assign n22037 = pi15 ? n22033 : n22036;
  assign n22038 = pi20 ? n1324 : n428;
  assign n22039 = pi19 ? n32 : n22038;
  assign n22040 = pi18 ? n22039 : n20753;
  assign n22041 = pi17 ? n32 : n22040;
  assign n22042 = pi16 ? n32 : n22041;
  assign n22043 = pi15 ? n22036 : n22042;
  assign n22044 = pi14 ? n22037 : n22043;
  assign n22045 = pi13 ? n22030 : n22044;
  assign n22046 = pi12 ? n22017 : n22045;
  assign n22047 = pi14 ? n21343 : n21357;
  assign n22048 = pi14 ? n147 : n32;
  assign n22049 = pi13 ? n22047 : n22048;
  assign n22050 = pi15 ? n19972 : n13392;
  assign n22051 = pi14 ? n19972 : n22050;
  assign n22052 = pi15 ? n13392 : n20315;
  assign n22053 = pi15 ? n21992 : n21918;
  assign n22054 = pi14 ? n22052 : n22053;
  assign n22055 = pi13 ? n22051 : n22054;
  assign n22056 = pi12 ? n22049 : n22055;
  assign n22057 = pi11 ? n22046 : n22056;
  assign n22058 = pi10 ? n22013 : n22057;
  assign n22059 = pi09 ? n32 : n22058;
  assign n22060 = pi14 ? n648 : n649;
  assign n22061 = pi13 ? n32 : n22060;
  assign n22062 = pi12 ? n32 : n22061;
  assign n22063 = pi14 ? n476 : n32;
  assign n22064 = pi13 ? n22063 : n32;
  assign n22065 = pi14 ? n22009 : n21464;
  assign n22066 = pi13 ? n22008 : n22065;
  assign n22067 = pi12 ? n22064 : n22066;
  assign n22068 = pi11 ? n22062 : n22067;
  assign n22069 = pi18 ? n15844 : n21798;
  assign n22070 = pi17 ? n32 : n22069;
  assign n22071 = pi16 ? n32 : n22070;
  assign n22072 = pi20 ? n32 : n16210;
  assign n22073 = pi19 ? n22072 : n32;
  assign n22074 = pi18 ? n32 : n22073;
  assign n22075 = pi17 ? n32 : n22074;
  assign n22076 = pi16 ? n32 : n22075;
  assign n22077 = pi15 ? n22071 : n22076;
  assign n22078 = pi21 ? n51 : n140;
  assign n22079 = pi20 ? n32 : ~n22078;
  assign n22080 = pi19 ? n22079 : n32;
  assign n22081 = pi18 ? n32 : n22080;
  assign n22082 = pi17 ? n32 : n22081;
  assign n22083 = pi16 ? n32 : n22082;
  assign n22084 = pi19 ? n17859 : n32;
  assign n22085 = pi18 ? n32 : n22084;
  assign n22086 = pi17 ? n32 : n22085;
  assign n22087 = pi16 ? n32 : n22086;
  assign n22088 = pi15 ? n22083 : n22087;
  assign n22089 = pi14 ? n22077 : n22088;
  assign n22090 = pi13 ? n21695 : n22089;
  assign n22091 = pi18 ? n15844 : n5158;
  assign n22092 = pi17 ? n32 : n22091;
  assign n22093 = pi16 ? n32 : n22092;
  assign n22094 = pi15 ? n21551 : n22093;
  assign n22095 = pi18 ? n16234 : n4671;
  assign n22096 = pi17 ? n32 : n22095;
  assign n22097 = pi16 ? n32 : n22096;
  assign n22098 = pi18 ? n21888 : ~n18891;
  assign n22099 = pi17 ? n32 : n22098;
  assign n22100 = pi16 ? n32 : n22099;
  assign n22101 = pi15 ? n22097 : n22100;
  assign n22102 = pi14 ? n22094 : n22101;
  assign n22103 = pi17 ? n19262 : n21894;
  assign n22104 = pi16 ? n32 : n22103;
  assign n22105 = pi15 ? n22104 : n11426;
  assign n22106 = pi20 ? n246 : n428;
  assign n22107 = pi19 ? n32 : n22106;
  assign n22108 = pi18 ? n22107 : n32;
  assign n22109 = pi17 ? n32 : n22108;
  assign n22110 = pi16 ? n32 : n22109;
  assign n22111 = pi15 ? n11426 : n22110;
  assign n22112 = pi14 ? n22105 : n22111;
  assign n22113 = pi13 ? n22102 : n22112;
  assign n22114 = pi12 ? n22090 : n22113;
  assign n22115 = pi15 ? n13948 : n20477;
  assign n22116 = pi14 ? n20756 : n22115;
  assign n22117 = pi14 ? n20306 : n32;
  assign n22118 = pi13 ? n22116 : n22117;
  assign n22119 = pi15 ? n19972 : n20315;
  assign n22120 = pi18 ? n15844 : n19750;
  assign n22121 = pi17 ? n32 : n22120;
  assign n22122 = pi16 ? n32 : n22121;
  assign n22123 = pi15 ? n22122 : n21992;
  assign n22124 = pi14 ? n22119 : n22123;
  assign n22125 = pi13 ? n19972 : n22124;
  assign n22126 = pi12 ? n22118 : n22125;
  assign n22127 = pi11 ? n22114 : n22126;
  assign n22128 = pi10 ? n22068 : n22127;
  assign n22129 = pi09 ? n32 : n22128;
  assign n22130 = pi08 ? n22059 : n22129;
  assign n22131 = pi07 ? n22000 : n22130;
  assign n22132 = pi06 ? n21851 : n22131;
  assign n22133 = pi15 ? n21928 : n32;
  assign n22134 = pi14 ? n22133 : n32;
  assign n22135 = pi13 ? n22134 : n32;
  assign n22136 = pi15 ? n21853 : n21686;
  assign n22137 = pi14 ? n21928 : n22136;
  assign n22138 = pi14 ? n21687 : n32;
  assign n22139 = pi13 ? n22137 : n22138;
  assign n22140 = pi12 ? n22135 : n22139;
  assign n22141 = pi11 ? n22062 : n22140;
  assign n22142 = pi15 ? n32 : n21801;
  assign n22143 = pi18 ? n222 : n21798;
  assign n22144 = pi17 ? n32 : n22143;
  assign n22145 = pi16 ? n32 : n22144;
  assign n22146 = pi18 ? n4127 : n21692;
  assign n22147 = pi17 ? n32 : n22146;
  assign n22148 = pi16 ? n32 : n22147;
  assign n22149 = pi15 ? n22145 : n22148;
  assign n22150 = pi14 ? n22142 : n22149;
  assign n22151 = pi14 ? n21695 : n21697;
  assign n22152 = pi13 ? n22150 : n22151;
  assign n22153 = pi15 ? n14405 : n21141;
  assign n22154 = pi20 ? n206 : n274;
  assign n22155 = pi19 ? n22154 : n32;
  assign n22156 = pi18 ? n15844 : n22155;
  assign n22157 = pi17 ? n32 : n22156;
  assign n22158 = pi16 ? n32 : n22157;
  assign n22159 = pi19 ? n1053 : ~n32;
  assign n22160 = pi18 ? n496 : ~n22159;
  assign n22161 = pi17 ? n32 : n22160;
  assign n22162 = pi16 ? n32 : n22161;
  assign n22163 = pi15 ? n22158 : n22162;
  assign n22164 = pi14 ? n22153 : n22163;
  assign n22165 = pi18 ? n702 : ~n797;
  assign n22166 = pi17 ? n32 : n22165;
  assign n22167 = pi16 ? n32 : n22166;
  assign n22168 = pi18 ? n697 : ~n797;
  assign n22169 = pi17 ? n32 : n22168;
  assign n22170 = pi16 ? n32 : n22169;
  assign n22171 = pi15 ? n22167 : n22170;
  assign n22172 = pi18 ? n15406 : n13058;
  assign n22173 = pi17 ? n32 : n22172;
  assign n22174 = pi16 ? n32 : n22173;
  assign n22175 = pi15 ? n22174 : n32;
  assign n22176 = pi14 ? n22171 : n22175;
  assign n22177 = pi13 ? n22164 : n22176;
  assign n22178 = pi12 ? n22152 : n22177;
  assign n22179 = pi14 ? n21232 : n22115;
  assign n22180 = pi14 ? n672 : n20297;
  assign n22181 = pi13 ? n22179 : n22180;
  assign n22182 = pi14 ? n146 : n19972;
  assign n22183 = pi19 ? n18211 : n20925;
  assign n22184 = pi18 ? n6059 : n22183;
  assign n22185 = pi20 ? n207 : ~n246;
  assign n22186 = pi19 ? n3692 : n22185;
  assign n22187 = pi18 ? n22186 : ~n19750;
  assign n22188 = pi17 ? n22184 : ~n22187;
  assign n22189 = pi16 ? n32 : n22188;
  assign n22190 = pi15 ? n19972 : n22189;
  assign n22191 = pi18 ? n16801 : ~n20525;
  assign n22192 = pi17 ? n32 : n22191;
  assign n22193 = pi16 ? n32 : n22192;
  assign n22194 = pi19 ? n8286 : ~n32;
  assign n22195 = pi18 ? n16801 : ~n22194;
  assign n22196 = pi17 ? n32 : n22195;
  assign n22197 = pi16 ? n32 : n22196;
  assign n22198 = pi15 ? n22193 : n22197;
  assign n22199 = pi14 ? n22190 : n22198;
  assign n22200 = pi13 ? n22182 : n22199;
  assign n22201 = pi12 ? n22181 : n22200;
  assign n22202 = pi11 ? n22178 : n22201;
  assign n22203 = pi10 ? n22141 : n22202;
  assign n22204 = pi09 ? n32 : n22203;
  assign n22205 = pi15 ? n32 : n15263;
  assign n22206 = pi14 ? n32 : n22205;
  assign n22207 = pi14 ? n15263 : n15267;
  assign n22208 = pi13 ? n22206 : n22207;
  assign n22209 = pi12 ? n32 : n22208;
  assign n22210 = pi14 ? n648 : n32;
  assign n22211 = pi14 ? n32 : n737;
  assign n22212 = pi13 ? n22210 : n22211;
  assign n22213 = pi15 ? n21928 : n476;
  assign n22214 = pi14 ? n22213 : n22136;
  assign n22215 = pi14 ? n21687 : n21543;
  assign n22216 = pi13 ? n22214 : n22215;
  assign n22217 = pi12 ? n22212 : n22216;
  assign n22218 = pi11 ? n22209 : n22217;
  assign n22219 = pi15 ? n21543 : n14152;
  assign n22220 = pi18 ? n222 : n5731;
  assign n22221 = pi17 ? n32 : n22220;
  assign n22222 = pi16 ? n32 : n22221;
  assign n22223 = pi18 ? n4127 : n5351;
  assign n22224 = pi17 ? n32 : n22223;
  assign n22225 = pi16 ? n32 : n22224;
  assign n22226 = pi15 ? n22222 : n22225;
  assign n22227 = pi14 ? n22219 : n22226;
  assign n22228 = pi15 ? n14394 : n21695;
  assign n22229 = pi14 ? n14394 : n22228;
  assign n22230 = pi13 ? n22227 : n22229;
  assign n22231 = pi14 ? n21866 : n22163;
  assign n22232 = pi15 ? n22174 : n20836;
  assign n22233 = pi14 ? n22171 : n22232;
  assign n22234 = pi13 ? n22231 : n22233;
  assign n22235 = pi12 ? n22230 : n22234;
  assign n22236 = pi15 ? n13943 : n21232;
  assign n22237 = pi14 ? n22236 : n13948;
  assign n22238 = pi14 ? n21357 : n32;
  assign n22239 = pi13 ? n22237 : n22238;
  assign n22240 = pi14 ? n32 : n20779;
  assign n22241 = pi18 ? n22186 : ~n19848;
  assign n22242 = pi17 ? n22184 : ~n22241;
  assign n22243 = pi16 ? n32 : n22242;
  assign n22244 = pi15 ? n20779 : n22243;
  assign n22245 = pi14 ? n22244 : n22198;
  assign n22246 = pi13 ? n22240 : n22245;
  assign n22247 = pi12 ? n22239 : n22246;
  assign n22248 = pi11 ? n22235 : n22247;
  assign n22249 = pi10 ? n22218 : n22248;
  assign n22250 = pi09 ? n32 : n22249;
  assign n22251 = pi08 ? n22204 : n22250;
  assign n22252 = pi15 ? n32 : n15123;
  assign n22253 = pi14 ? n32 : n22252;
  assign n22254 = pi14 ? n15123 : n15127;
  assign n22255 = pi13 ? n22253 : n22254;
  assign n22256 = pi12 ? n32 : n22255;
  assign n22257 = pi15 ? n32 : n648;
  assign n22258 = pi14 ? n32 : n22257;
  assign n22259 = pi13 ? n650 : n22258;
  assign n22260 = pi15 ? n648 : n14790;
  assign n22261 = pi15 ? n14790 : n21853;
  assign n22262 = pi14 ? n22260 : n22261;
  assign n22263 = pi13 ? n22262 : n21855;
  assign n22264 = pi12 ? n22259 : n22263;
  assign n22265 = pi11 ? n22256 : n22264;
  assign n22266 = pi18 ? n222 : n9578;
  assign n22267 = pi17 ? n32 : n22266;
  assign n22268 = pi16 ? n32 : n22267;
  assign n22269 = pi20 ? n339 : n518;
  assign n22270 = pi19 ? n22269 : ~n32;
  assign n22271 = pi18 ? n4127 : ~n22270;
  assign n22272 = pi17 ? n32 : n22271;
  assign n22273 = pi16 ? n32 : n22272;
  assign n22274 = pi15 ? n22268 : n22273;
  assign n22275 = pi18 ? n209 : ~n22270;
  assign n22276 = pi17 ? n32 : n22275;
  assign n22277 = pi16 ? n32 : n22276;
  assign n22278 = pi20 ? n9641 : n9863;
  assign n22279 = pi19 ? n22278 : n32;
  assign n22280 = pi18 ? n32 : n22279;
  assign n22281 = pi17 ? n32 : n22280;
  assign n22282 = pi16 ? n32 : n22281;
  assign n22283 = pi15 ? n22277 : n22282;
  assign n22284 = pi14 ? n22274 : n22283;
  assign n22285 = pi15 ? n14394 : n21389;
  assign n22286 = pi14 ? n14394 : n22285;
  assign n22287 = pi13 ? n22284 : n22286;
  assign n22288 = pi20 ? n266 : n6229;
  assign n22289 = pi19 ? n22288 : n32;
  assign n22290 = pi18 ? n4380 : n22289;
  assign n22291 = pi17 ? n32 : n22290;
  assign n22292 = pi16 ? n32 : n22291;
  assign n22293 = pi15 ? n21319 : n22292;
  assign n22294 = pi20 ? n206 : n6229;
  assign n22295 = pi19 ? n22294 : n32;
  assign n22296 = pi18 ? n15844 : n22295;
  assign n22297 = pi17 ? n32 : n22296;
  assign n22298 = pi16 ? n32 : n22297;
  assign n22299 = pi19 ? n15460 : ~n32;
  assign n22300 = pi18 ? n496 : ~n22299;
  assign n22301 = pi17 ? n32 : n22300;
  assign n22302 = pi16 ? n32 : n22301;
  assign n22303 = pi15 ? n22298 : n22302;
  assign n22304 = pi14 ? n22293 : n22303;
  assign n22305 = pi19 ? n5694 : ~n18502;
  assign n22306 = pi18 ? n5158 : n22305;
  assign n22307 = pi19 ? n342 : ~n32;
  assign n22308 = pi18 ? n22307 : ~n2291;
  assign n22309 = pi17 ? n22306 : n22308;
  assign n22310 = pi16 ? n32 : n22309;
  assign n22311 = pi18 ? n684 : ~n2291;
  assign n22312 = pi17 ? n32 : n22311;
  assign n22313 = pi16 ? n32 : n22312;
  assign n22314 = pi15 ? n22310 : n22313;
  assign n22315 = pi14 ? n22314 : n20836;
  assign n22316 = pi13 ? n22304 : n22315;
  assign n22317 = pi12 ? n22287 : n22316;
  assign n22318 = pi15 ? n21226 : n20756;
  assign n22319 = pi14 ? n22318 : n20660;
  assign n22320 = pi15 ? n486 : n32;
  assign n22321 = pi14 ? n22320 : n13952;
  assign n22322 = pi13 ? n22319 : n22321;
  assign n22323 = pi14 ? n13952 : n20779;
  assign n22324 = pi18 ? n1464 : n19848;
  assign n22325 = pi17 ? n18560 : n22324;
  assign n22326 = pi16 ? n32 : n22325;
  assign n22327 = pi15 ? n20779 : n22326;
  assign n22328 = pi18 ? n16801 : n20320;
  assign n22329 = pi17 ? n32 : n22328;
  assign n22330 = pi16 ? n32 : n22329;
  assign n22331 = pi21 ? n174 : ~n1939;
  assign n22332 = pi20 ? n22331 : n32;
  assign n22333 = pi19 ? n22332 : n32;
  assign n22334 = pi18 ? n16389 : n22333;
  assign n22335 = pi17 ? n32 : n22334;
  assign n22336 = pi16 ? n32 : n22335;
  assign n22337 = pi15 ? n22330 : n22336;
  assign n22338 = pi14 ? n22327 : n22337;
  assign n22339 = pi13 ? n22323 : n22338;
  assign n22340 = pi12 ? n22322 : n22339;
  assign n22341 = pi11 ? n22317 : n22340;
  assign n22342 = pi10 ? n22265 : n22341;
  assign n22343 = pi09 ? n32 : n22342;
  assign n22344 = pi19 ? n17685 : n32;
  assign n22345 = pi18 ? n32 : n22344;
  assign n22346 = pi17 ? n32 : n22345;
  assign n22347 = pi16 ? n32 : n22346;
  assign n22348 = pi15 ? n32 : n22347;
  assign n22349 = pi14 ? n32 : n22348;
  assign n22350 = pi15 ? n22347 : n32;
  assign n22351 = pi14 ? n22347 : n22350;
  assign n22352 = pi13 ? n22349 : n22351;
  assign n22353 = pi12 ? n32 : n22352;
  assign n22354 = pi14 ? n15123 : n32;
  assign n22355 = pi13 ? n22354 : n22258;
  assign n22356 = pi14 ? n21854 : n21786;
  assign n22357 = pi13 ? n22262 : n22356;
  assign n22358 = pi12 ? n22355 : n22357;
  assign n22359 = pi11 ? n22353 : n22358;
  assign n22360 = pi18 ? n222 : n21683;
  assign n22361 = pi17 ? n32 : n22360;
  assign n22362 = pi16 ? n32 : n22361;
  assign n22363 = pi20 ? n339 : n1319;
  assign n22364 = pi19 ? n22363 : ~n32;
  assign n22365 = pi18 ? n4127 : ~n22364;
  assign n22366 = pi17 ? n32 : n22365;
  assign n22367 = pi16 ? n32 : n22366;
  assign n22368 = pi15 ? n22362 : n22367;
  assign n22369 = pi18 ? n209 : ~n22364;
  assign n22370 = pi17 ? n32 : n22369;
  assign n22371 = pi16 ? n32 : n22370;
  assign n22372 = pi20 ? n32 : n7852;
  assign n22373 = pi19 ? n22372 : n32;
  assign n22374 = pi18 ? n32 : n22373;
  assign n22375 = pi17 ? n32 : n22374;
  assign n22376 = pi16 ? n32 : n22375;
  assign n22377 = pi15 ? n22371 : n22376;
  assign n22378 = pi14 ? n22368 : n22377;
  assign n22379 = pi18 ? n32 : n9865;
  assign n22380 = pi17 ? n32 : n22379;
  assign n22381 = pi16 ? n32 : n22380;
  assign n22382 = pi15 ? n14394 : n22381;
  assign n22383 = pi14 ? n22007 : n22382;
  assign n22384 = pi13 ? n22378 : n22383;
  assign n22385 = pi19 ? n17769 : n32;
  assign n22386 = pi18 ? n4380 : n22385;
  assign n22387 = pi17 ? n32 : n22386;
  assign n22388 = pi16 ? n32 : n22387;
  assign n22389 = pi15 ? n21389 : n22388;
  assign n22390 = pi18 ? n15844 : n20605;
  assign n22391 = pi17 ? n32 : n22390;
  assign n22392 = pi16 ? n32 : n22391;
  assign n22393 = pi15 ? n22392 : n22302;
  assign n22394 = pi14 ? n22389 : n22393;
  assign n22395 = pi14 ? n22314 : n21133;
  assign n22396 = pi13 ? n22394 : n22395;
  assign n22397 = pi12 ? n22384 : n22396;
  assign n22398 = pi15 ? n21033 : n14168;
  assign n22399 = pi14 ? n22398 : n20758;
  assign n22400 = pi14 ? n21041 : n13952;
  assign n22401 = pi13 ? n22399 : n22400;
  assign n22402 = pi14 ? n13952 : n13671;
  assign n22403 = pi18 ? n1464 : n4343;
  assign n22404 = pi17 ? n18560 : n22403;
  assign n22405 = pi16 ? n32 : n22404;
  assign n22406 = pi15 ? n20779 : n22405;
  assign n22407 = pi18 ? n16801 : n13086;
  assign n22408 = pi17 ? n32 : n22407;
  assign n22409 = pi16 ? n32 : n22408;
  assign n22410 = pi20 ? n21111 : n32;
  assign n22411 = pi19 ? n22410 : n32;
  assign n22412 = pi18 ? n16389 : n22411;
  assign n22413 = pi17 ? n32 : n22412;
  assign n22414 = pi16 ? n32 : n22413;
  assign n22415 = pi15 ? n22409 : n22414;
  assign n22416 = pi14 ? n22406 : n22415;
  assign n22417 = pi13 ? n22402 : n22416;
  assign n22418 = pi12 ? n22401 : n22417;
  assign n22419 = pi11 ? n22397 : n22418;
  assign n22420 = pi10 ? n22359 : n22419;
  assign n22421 = pi09 ? n32 : n22420;
  assign n22422 = pi08 ? n22343 : n22421;
  assign n22423 = pi07 ? n22251 : n22422;
  assign n22424 = pi15 ? n32 : n15389;
  assign n22425 = pi14 ? n32 : n22424;
  assign n22426 = pi14 ? n15389 : n15390;
  assign n22427 = pi13 ? n22425 : n22426;
  assign n22428 = pi12 ? n32 : n22427;
  assign n22429 = pi13 ? n15268 : n22253;
  assign n22430 = pi20 ? n32 : ~n11107;
  assign n22431 = pi19 ? n22430 : n32;
  assign n22432 = pi18 ? n32 : n22431;
  assign n22433 = pi17 ? n32 : n22432;
  assign n22434 = pi16 ? n32 : n22433;
  assign n22435 = pi18 ? n32 : n20912;
  assign n22436 = pi17 ? n32 : n22435;
  assign n22437 = pi16 ? n32 : n22436;
  assign n22438 = pi15 ? n22434 : n22437;
  assign n22439 = pi15 ? n22437 : n14973;
  assign n22440 = pi14 ? n22438 : n22439;
  assign n22441 = pi15 ? n14973 : n476;
  assign n22442 = pi14 ? n22441 : n21787;
  assign n22443 = pi13 ? n22440 : n22442;
  assign n22444 = pi12 ? n22429 : n22443;
  assign n22445 = pi11 ? n22428 : n22444;
  assign n22446 = pi18 ? n751 : n9012;
  assign n22447 = pi17 ? n32 : n22446;
  assign n22448 = pi16 ? n32 : n22447;
  assign n22449 = pi20 ? n32 : ~n17509;
  assign n22450 = pi19 ? n22449 : ~n32;
  assign n22451 = pi18 ? n940 : ~n22450;
  assign n22452 = pi17 ? n32 : n22451;
  assign n22453 = pi16 ? n32 : n22452;
  assign n22454 = pi15 ? n22448 : n22453;
  assign n22455 = pi18 ? n4380 : ~n2747;
  assign n22456 = pi17 ? n32 : n22455;
  assign n22457 = pi16 ? n32 : n22456;
  assign n22458 = pi21 ? n309 : ~n242;
  assign n22459 = pi20 ? n266 : n22458;
  assign n22460 = pi19 ? n22459 : n32;
  assign n22461 = pi18 ? n32 : n22460;
  assign n22462 = pi17 ? n32 : n22461;
  assign n22463 = pi16 ? n32 : n22462;
  assign n22464 = pi15 ? n22457 : n22463;
  assign n22465 = pi14 ? n22454 : n22464;
  assign n22466 = pi19 ? n17941 : n32;
  assign n22467 = pi18 ? n32 : n22466;
  assign n22468 = pi17 ? n32 : n22467;
  assign n22469 = pi16 ? n32 : n22468;
  assign n22470 = pi15 ? n22469 : n14394;
  assign n22471 = pi18 ? n268 : n9865;
  assign n22472 = pi17 ? n32 : n22471;
  assign n22473 = pi16 ? n32 : n22472;
  assign n22474 = pi15 ? n14394 : n22473;
  assign n22475 = pi14 ? n22470 : n22474;
  assign n22476 = pi13 ? n22465 : n22475;
  assign n22477 = pi18 ? n4380 : n21938;
  assign n22478 = pi17 ? n32 : n22477;
  assign n22479 = pi16 ? n32 : n22478;
  assign n22480 = pi20 ? n207 : ~n1331;
  assign n22481 = pi19 ? n22480 : ~n32;
  assign n22482 = pi18 ? n880 : ~n22481;
  assign n22483 = pi17 ? n32 : n22482;
  assign n22484 = pi16 ? n32 : n22483;
  assign n22485 = pi15 ? n22479 : n22484;
  assign n22486 = pi19 ? n7168 : ~n32;
  assign n22487 = pi18 ? n684 : ~n22486;
  assign n22488 = pi17 ? n32 : n22487;
  assign n22489 = pi16 ? n32 : n22488;
  assign n22490 = pi20 ? n266 : ~n1331;
  assign n22491 = pi19 ? n22490 : ~n32;
  assign n22492 = pi18 ? n496 : ~n22491;
  assign n22493 = pi17 ? n32 : n22492;
  assign n22494 = pi16 ? n32 : n22493;
  assign n22495 = pi15 ? n22489 : n22494;
  assign n22496 = pi14 ? n22485 : n22495;
  assign n22497 = pi19 ? n5435 : n342;
  assign n22498 = pi20 ? n6621 : n321;
  assign n22499 = pi19 ? n18396 : n22498;
  assign n22500 = pi18 ? n22497 : n22499;
  assign n22501 = pi20 ? n207 : n206;
  assign n22502 = pi19 ? n22501 : n32;
  assign n22503 = pi18 ? n22502 : n323;
  assign n22504 = pi17 ? n22500 : ~n22503;
  assign n22505 = pi16 ? n16104 : n22504;
  assign n22506 = pi20 ? n246 : ~n501;
  assign n22507 = pi19 ? n22506 : n32;
  assign n22508 = pi18 ? n1379 : n22507;
  assign n22509 = pi17 ? n32 : n22508;
  assign n22510 = pi16 ? n32 : n22509;
  assign n22511 = pi15 ? n22505 : n22510;
  assign n22512 = pi14 ? n22511 : n21133;
  assign n22513 = pi13 ? n22496 : n22512;
  assign n22514 = pi12 ? n22476 : n22513;
  assign n22515 = pi14 ? n21041 : n486;
  assign n22516 = pi13 ? n22399 : n22515;
  assign n22517 = pi18 ? n4380 : n20298;
  assign n22518 = pi17 ? n32 : n22517;
  assign n22519 = pi16 ? n32 : n22518;
  assign n22520 = pi15 ? n13952 : n22519;
  assign n22521 = pi14 ? n21357 : n22520;
  assign n22522 = pi18 ? n880 : n13377;
  assign n22523 = pi17 ? n32 : n22522;
  assign n22524 = pi16 ? n32 : n22523;
  assign n22525 = pi20 ? n342 : ~n246;
  assign n22526 = pi19 ? n32 : n22525;
  assign n22527 = pi18 ? n22526 : n4343;
  assign n22528 = pi17 ? n32 : n22527;
  assign n22529 = pi16 ? n32 : n22528;
  assign n22530 = pi15 ? n22524 : n22529;
  assign n22531 = pi15 ? n19851 : n20531;
  assign n22532 = pi14 ? n22530 : n22531;
  assign n22533 = pi13 ? n22521 : n22532;
  assign n22534 = pi12 ? n22516 : n22533;
  assign n22535 = pi11 ? n22514 : n22534;
  assign n22536 = pi10 ? n22445 : n22535;
  assign n22537 = pi09 ? n32 : n22536;
  assign n22538 = pi18 ? n32 : n6118;
  assign n22539 = pi17 ? n32 : n22538;
  assign n22540 = pi16 ? n32 : n22539;
  assign n22541 = pi15 ? n32 : n22540;
  assign n22542 = pi14 ? n32 : n22541;
  assign n22543 = pi15 ? n22540 : n32;
  assign n22544 = pi14 ? n22540 : n22543;
  assign n22545 = pi13 ? n22542 : n22544;
  assign n22546 = pi12 ? n32 : n22545;
  assign n22547 = pi14 ? n15389 : n32;
  assign n22548 = pi13 ? n22547 : n22253;
  assign n22549 = pi15 ? n14973 : n21928;
  assign n22550 = pi14 ? n22549 : n21928;
  assign n22551 = pi13 ? n22440 : n22550;
  assign n22552 = pi12 ? n22548 : n22551;
  assign n22553 = pi11 ? n22546 : n22552;
  assign n22554 = pi19 ? n311 : n32;
  assign n22555 = pi18 ? n751 : n22554;
  assign n22556 = pi17 ? n32 : n22555;
  assign n22557 = pi16 ? n32 : n22556;
  assign n22558 = pi20 ? n32 : ~n310;
  assign n22559 = pi19 ? n22558 : ~n32;
  assign n22560 = pi18 ? n940 : ~n22559;
  assign n22561 = pi17 ? n32 : n22560;
  assign n22562 = pi16 ? n32 : n22561;
  assign n22563 = pi15 ? n22557 : n22562;
  assign n22564 = pi18 ? n4380 : ~n508;
  assign n22565 = pi17 ? n32 : n22564;
  assign n22566 = pi16 ? n32 : n22565;
  assign n22567 = pi20 ? n266 : n12884;
  assign n22568 = pi19 ? n22567 : n32;
  assign n22569 = pi18 ? n32 : n22568;
  assign n22570 = pi17 ? n32 : n22569;
  assign n22571 = pi16 ? n32 : n22570;
  assign n22572 = pi15 ? n22566 : n22571;
  assign n22573 = pi14 ? n22563 : n22572;
  assign n22574 = pi15 ? n14147 : n22006;
  assign n22575 = pi18 ? n268 : n21683;
  assign n22576 = pi17 ? n32 : n22575;
  assign n22577 = pi16 ? n32 : n22576;
  assign n22578 = pi15 ? n22006 : n22577;
  assign n22579 = pi14 ? n22574 : n22578;
  assign n22580 = pi13 ? n22573 : n22579;
  assign n22581 = pi18 ? n4380 : n21860;
  assign n22582 = pi17 ? n32 : n22581;
  assign n22583 = pi16 ? n32 : n22582;
  assign n22584 = pi20 ? n207 : ~n160;
  assign n22585 = pi19 ? n22584 : ~n32;
  assign n22586 = pi18 ? n880 : ~n22585;
  assign n22587 = pi17 ? n32 : n22586;
  assign n22588 = pi16 ? n32 : n22587;
  assign n22589 = pi15 ? n22583 : n22588;
  assign n22590 = pi14 ? n22589 : n22495;
  assign n22591 = pi20 ? n3523 : ~n501;
  assign n22592 = pi19 ? n22591 : n32;
  assign n22593 = pi18 ? n863 : n22592;
  assign n22594 = pi17 ? n32 : n22593;
  assign n22595 = pi16 ? n32 : n22594;
  assign n22596 = pi15 ? n22505 : n22595;
  assign n22597 = pi14 ? n22596 : n21322;
  assign n22598 = pi13 ? n22590 : n22597;
  assign n22599 = pi12 ? n22580 : n22598;
  assign n22600 = pi15 ? n21033 : n14164;
  assign n22601 = pi15 ? n14168 : n20756;
  assign n22602 = pi14 ? n22600 : n22601;
  assign n22603 = pi20 ? n32 : n18423;
  assign n22604 = pi19 ? n22603 : n32;
  assign n22605 = pi18 ? n32 : n22604;
  assign n22606 = pi17 ? n32 : n22605;
  assign n22607 = pi16 ? n32 : n22606;
  assign n22608 = pi15 ? n22607 : n32;
  assign n22609 = pi14 ? n22608 : n487;
  assign n22610 = pi13 ? n22602 : n22609;
  assign n22611 = pi15 ? n20477 : n22519;
  assign n22612 = pi14 ? n20477 : n22611;
  assign n22613 = pi18 ? n880 : n13372;
  assign n22614 = pi17 ? n32 : n22613;
  assign n22615 = pi16 ? n32 : n22614;
  assign n22616 = pi18 ? n22526 : n13377;
  assign n22617 = pi17 ? n32 : n22616;
  assign n22618 = pi16 ? n32 : n22617;
  assign n22619 = pi15 ? n22615 : n22618;
  assign n22620 = pi15 ? n20692 : n19851;
  assign n22621 = pi14 ? n22619 : n22620;
  assign n22622 = pi13 ? n22612 : n22621;
  assign n22623 = pi12 ? n22610 : n22622;
  assign n22624 = pi11 ? n22599 : n22623;
  assign n22625 = pi10 ? n22553 : n22624;
  assign n22626 = pi09 ? n32 : n22625;
  assign n22627 = pi08 ? n22537 : n22626;
  assign n22628 = pi14 ? n22424 : n15389;
  assign n22629 = pi13 ? n15391 : n22628;
  assign n22630 = pi19 ? n18022 : n32;
  assign n22631 = pi18 ? n32 : n22630;
  assign n22632 = pi17 ? n32 : n22631;
  assign n22633 = pi16 ? n32 : n22632;
  assign n22634 = pi15 ? n22633 : n22437;
  assign n22635 = pi15 ? n15123 : n14967;
  assign n22636 = pi14 ? n22634 : n22635;
  assign n22637 = pi15 ? n15123 : n14973;
  assign n22638 = pi15 ? n21928 : n21853;
  assign n22639 = pi14 ? n22637 : n22638;
  assign n22640 = pi13 ? n22636 : n22639;
  assign n22641 = pi12 ? n22629 : n22640;
  assign n22642 = pi11 ? n22546 : n22641;
  assign n22643 = pi20 ? n310 : ~n206;
  assign n22644 = pi19 ? n22643 : n32;
  assign n22645 = pi18 ? n940 : n22644;
  assign n22646 = pi17 ? n32 : n22645;
  assign n22647 = pi16 ? n32 : n22646;
  assign n22648 = pi18 ? n940 : ~n508;
  assign n22649 = pi17 ? n32 : n22648;
  assign n22650 = pi16 ? n32 : n22649;
  assign n22651 = pi15 ? n22647 : n22650;
  assign n22652 = pi20 ? n266 : n220;
  assign n22653 = pi19 ? n22652 : n32;
  assign n22654 = pi18 ? n32 : n22653;
  assign n22655 = pi17 ? n32 : n22654;
  assign n22656 = pi16 ? n32 : n22655;
  assign n22657 = pi15 ? n13338 : n22656;
  assign n22658 = pi14 ? n22651 : n22657;
  assign n22659 = pi18 ? n268 : n9578;
  assign n22660 = pi17 ? n32 : n22659;
  assign n22661 = pi16 ? n32 : n22660;
  assign n22662 = pi15 ? n22006 : n22661;
  assign n22663 = pi14 ? n22574 : n22662;
  assign n22664 = pi13 ? n22658 : n22663;
  assign n22665 = pi18 ? n4380 : n5351;
  assign n22666 = pi17 ? n32 : n22665;
  assign n22667 = pi16 ? n32 : n22666;
  assign n22668 = pi17 ? n17119 : n22586;
  assign n22669 = pi16 ? n32 : n22668;
  assign n22670 = pi15 ? n22667 : n22669;
  assign n22671 = pi20 ? n321 : ~n7388;
  assign n22672 = pi19 ? n22671 : ~n32;
  assign n22673 = pi18 ? n209 : ~n22672;
  assign n22674 = pi17 ? n17433 : n22673;
  assign n22675 = pi16 ? n32 : n22674;
  assign n22676 = pi20 ? n32 : ~n7388;
  assign n22677 = pi19 ? n22676 : ~n32;
  assign n22678 = pi18 ? n209 : ~n22677;
  assign n22679 = pi17 ? n32 : n22678;
  assign n22680 = pi16 ? n32 : n22679;
  assign n22681 = pi15 ? n22675 : n22680;
  assign n22682 = pi14 ? n22670 : n22681;
  assign n22683 = pi20 ? n357 : ~n9367;
  assign n22684 = pi19 ? n22683 : n32;
  assign n22685 = pi18 ? n17848 : n22684;
  assign n22686 = pi17 ? n32 : n22685;
  assign n22687 = pi16 ? n32 : n22686;
  assign n22688 = pi15 ? n22687 : n21319;
  assign n22689 = pi14 ? n22688 : n21319;
  assign n22690 = pi13 ? n22682 : n22689;
  assign n22691 = pi12 ? n22664 : n22690;
  assign n22692 = pi15 ? n20836 : n20831;
  assign n22693 = pi14 ? n21033 : n22692;
  assign n22694 = pi14 ? n20758 : n20660;
  assign n22695 = pi13 ? n22693 : n22694;
  assign n22696 = pi19 ? n246 : ~n339;
  assign n22697 = pi20 ? n339 : n7939;
  assign n22698 = pi20 ? n6621 : n175;
  assign n22699 = pi19 ? n22697 : ~n22698;
  assign n22700 = pi18 ? n22696 : ~n22699;
  assign n22701 = pi20 ? n207 : n287;
  assign n22702 = pi20 ? n5854 : ~n7939;
  assign n22703 = pi19 ? n22701 : ~n22702;
  assign n22704 = pi20 ? n266 : n339;
  assign n22705 = pi19 ? n22704 : ~n32;
  assign n22706 = pi18 ? n22703 : n22705;
  assign n22707 = pi17 ? n22700 : ~n22706;
  assign n22708 = pi16 ? n32 : n22707;
  assign n22709 = pi15 ? n20477 : n22708;
  assign n22710 = pi14 ? n486 : n22709;
  assign n22711 = pi18 ? n880 : ~n22705;
  assign n22712 = pi17 ? n32 : n22711;
  assign n22713 = pi16 ? n32 : n22712;
  assign n22714 = pi18 ? n4722 : n13377;
  assign n22715 = pi17 ? n32 : n22714;
  assign n22716 = pi16 ? n32 : n22715;
  assign n22717 = pi15 ? n22713 : n22716;
  assign n22718 = pi15 ? n19972 : n19851;
  assign n22719 = pi14 ? n22717 : n22718;
  assign n22720 = pi13 ? n22710 : n22719;
  assign n22721 = pi12 ? n22695 : n22720;
  assign n22722 = pi11 ? n22691 : n22721;
  assign n22723 = pi10 ? n22642 : n22722;
  assign n22724 = pi09 ? n32 : n22723;
  assign n22725 = pi19 ? n594 : ~n1105;
  assign n22726 = pi18 ? n32 : n22725;
  assign n22727 = pi17 ? n32 : n22726;
  assign n22728 = pi16 ? n32 : n22727;
  assign n22729 = pi15 ? n22728 : n32;
  assign n22730 = pi14 ? n1109 : n22729;
  assign n22731 = pi13 ? n1111 : n22730;
  assign n22732 = pi12 ? n32 : n22731;
  assign n22733 = pi16 ? n32 : n2074;
  assign n22734 = pi15 ? n22540 : n22733;
  assign n22735 = pi14 ? n22734 : n32;
  assign n22736 = pi13 ? n22735 : n22628;
  assign n22737 = pi15 ? n14973 : n14790;
  assign n22738 = pi14 ? n22637 : n22737;
  assign n22739 = pi13 ? n22636 : n22738;
  assign n22740 = pi12 ? n22736 : n22739;
  assign n22741 = pi11 ? n22732 : n22740;
  assign n22742 = pi20 ? n310 : ~n8285;
  assign n22743 = pi19 ? n22742 : n32;
  assign n22744 = pi18 ? n940 : n22743;
  assign n22745 = pi17 ? n32 : n22744;
  assign n22746 = pi16 ? n32 : n22745;
  assign n22747 = pi18 ? n940 : ~n2627;
  assign n22748 = pi17 ? n32 : n22747;
  assign n22749 = pi16 ? n32 : n22748;
  assign n22750 = pi15 ? n22746 : n22749;
  assign n22751 = pi20 ? n207 : ~n2140;
  assign n22752 = pi19 ? n22751 : n32;
  assign n22753 = pi18 ? n32 : n22752;
  assign n22754 = pi17 ? n32 : n22753;
  assign n22755 = pi16 ? n32 : n22754;
  assign n22756 = pi20 ? n266 : n7442;
  assign n22757 = pi19 ? n22756 : n32;
  assign n22758 = pi18 ? n32 : n22757;
  assign n22759 = pi17 ? n32 : n22758;
  assign n22760 = pi16 ? n32 : n22759;
  assign n22761 = pi15 ? n22755 : n22760;
  assign n22762 = pi14 ? n22750 : n22761;
  assign n22763 = pi15 ? n14147 : n14389;
  assign n22764 = pi15 ? n14389 : n22577;
  assign n22765 = pi14 ? n22763 : n22764;
  assign n22766 = pi13 ? n22762 : n22765;
  assign n22767 = pi18 ? n4380 : n22003;
  assign n22768 = pi17 ? n32 : n22767;
  assign n22769 = pi16 ? n32 : n22768;
  assign n22770 = pi17 ? n17119 : n19785;
  assign n22771 = pi16 ? n32 : n22770;
  assign n22772 = pi15 ? n22769 : n22771;
  assign n22773 = pi18 ? n209 : ~n5372;
  assign n22774 = pi17 ? n17433 : n22773;
  assign n22775 = pi16 ? n32 : n22774;
  assign n22776 = pi15 ? n22775 : n22680;
  assign n22777 = pi14 ? n22772 : n22776;
  assign n22778 = pi20 ? n32 : ~n7013;
  assign n22779 = pi19 ? n22778 : n32;
  assign n22780 = pi18 ? n17848 : n22779;
  assign n22781 = pi17 ? n32 : n22780;
  assign n22782 = pi16 ? n32 : n22781;
  assign n22783 = pi15 ? n22782 : n21389;
  assign n22784 = pi15 ? n21389 : n21319;
  assign n22785 = pi14 ? n22783 : n22784;
  assign n22786 = pi13 ? n22777 : n22785;
  assign n22787 = pi12 ? n22766 : n22786;
  assign n22788 = pi14 ? n14397 : n21035;
  assign n22789 = pi13 ? n22788 : n22694;
  assign n22790 = pi18 ? n22703 : n21257;
  assign n22791 = pi17 ? n22700 : ~n22790;
  assign n22792 = pi16 ? n32 : n22791;
  assign n22793 = pi15 ? n13948 : n22792;
  assign n22794 = pi14 ? n20660 : n22793;
  assign n22795 = pi18 ? n880 : ~n21257;
  assign n22796 = pi17 ? n32 : n22795;
  assign n22797 = pi16 ? n32 : n22796;
  assign n22798 = pi18 ? n4722 : n13372;
  assign n22799 = pi17 ? n32 : n22798;
  assign n22800 = pi16 ? n32 : n22799;
  assign n22801 = pi15 ? n22797 : n22800;
  assign n22802 = pi14 ? n22801 : n22718;
  assign n22803 = pi13 ? n22794 : n22802;
  assign n22804 = pi12 ? n22789 : n22803;
  assign n22805 = pi11 ? n22787 : n22804;
  assign n22806 = pi10 ? n22741 : n22805;
  assign n22807 = pi09 ? n32 : n22806;
  assign n22808 = pi08 ? n22724 : n22807;
  assign n22809 = pi07 ? n22627 : n22808;
  assign n22810 = pi06 ? n22423 : n22809;
  assign n22811 = pi05 ? n22132 : n22810;
  assign n22812 = pi15 ? n1109 : n32;
  assign n22813 = pi14 ? n1109 : n22812;
  assign n22814 = pi13 ? n1111 : n22813;
  assign n22815 = pi12 ? n32 : n22814;
  assign n22816 = pi17 ? n32 : n19886;
  assign n22817 = pi16 ? n32 : n22816;
  assign n22818 = pi15 ? n32 : n22817;
  assign n22819 = pi19 ? n1490 : n32;
  assign n22820 = pi18 ? n32 : n22819;
  assign n22821 = pi17 ? n32 : n22820;
  assign n22822 = pi16 ? n32 : n22821;
  assign n22823 = pi18 ? n32 : n5715;
  assign n22824 = pi17 ? n32 : n22823;
  assign n22825 = pi16 ? n32 : n22824;
  assign n22826 = pi15 ? n22822 : n22825;
  assign n22827 = pi14 ? n22818 : n22826;
  assign n22828 = pi13 ? n32 : n22827;
  assign n22829 = pi15 ? n22817 : n22347;
  assign n22830 = pi14 ? n22829 : n22347;
  assign n22831 = pi15 ? n22347 : n22437;
  assign n22832 = pi14 ? n22831 : n21853;
  assign n22833 = pi13 ? n22830 : n22832;
  assign n22834 = pi12 ? n22828 : n22833;
  assign n22835 = pi11 ? n22815 : n22834;
  assign n22836 = pi18 ? n4380 : ~n2627;
  assign n22837 = pi17 ? n32 : n22836;
  assign n22838 = pi16 ? n32 : n22837;
  assign n22839 = pi20 ? n10644 : ~n22331;
  assign n22840 = pi19 ? n22839 : ~n32;
  assign n22841 = pi18 ? n936 : ~n22840;
  assign n22842 = pi17 ? n32 : n22841;
  assign n22843 = pi16 ? n32 : n22842;
  assign n22844 = pi15 ? n22838 : n22843;
  assign n22845 = pi20 ? n342 : n7442;
  assign n22846 = pi19 ? n22845 : n32;
  assign n22847 = pi18 ? n32 : n22846;
  assign n22848 = pi17 ? n32 : n22847;
  assign n22849 = pi16 ? n32 : n22848;
  assign n22850 = pi19 ? n17842 : n32;
  assign n22851 = pi18 ? n4380 : n22850;
  assign n22852 = pi17 ? n32 : n22851;
  assign n22853 = pi16 ? n32 : n22852;
  assign n22854 = pi15 ? n22849 : n22853;
  assign n22855 = pi14 ? n22844 : n22854;
  assign n22856 = pi15 ? n14389 : n21853;
  assign n22857 = pi19 ? n20555 : ~n32;
  assign n22858 = pi18 ? n32 : ~n22857;
  assign n22859 = pi17 ? n32 : n22858;
  assign n22860 = pi16 ? n32 : n22859;
  assign n22861 = pi15 ? n22860 : n12524;
  assign n22862 = pi14 ? n22856 : n22861;
  assign n22863 = pi13 ? n22855 : n22862;
  assign n22864 = pi20 ? n342 : ~n266;
  assign n22865 = pi19 ? n32 : n22864;
  assign n22866 = pi18 ? n22865 : ~n520;
  assign n22867 = pi17 ? n32 : n22866;
  assign n22868 = pi16 ? n32 : n22867;
  assign n22869 = pi15 ? n12524 : n22868;
  assign n22870 = pi17 ? n17346 : n12074;
  assign n22871 = pi16 ? n32 : n22870;
  assign n22872 = pi19 ? n17964 : ~n32;
  assign n22873 = pi18 ? n209 : ~n22872;
  assign n22874 = pi17 ? n17346 : n22873;
  assign n22875 = pi16 ? n32 : n22874;
  assign n22876 = pi15 ? n22871 : n22875;
  assign n22877 = pi14 ? n22869 : n22876;
  assign n22878 = pi15 ? n21464 : n14397;
  assign n22879 = pi14 ? n21464 : n22878;
  assign n22880 = pi13 ? n22877 : n22879;
  assign n22881 = pi12 ? n22863 : n22880;
  assign n22882 = pi15 ? n20831 : n13948;
  assign n22883 = pi14 ? n20831 : n22882;
  assign n22884 = pi13 ? n22788 : n22883;
  assign n22885 = pi19 ? n32 : n4982;
  assign n22886 = pi18 ? n22885 : n5005;
  assign n22887 = pi17 ? n32 : n22886;
  assign n22888 = pi16 ? n32 : n22887;
  assign n22889 = pi19 ? n507 : n247;
  assign n22890 = pi18 ? n8106 : n22889;
  assign n22891 = pi20 ? n339 : ~n6621;
  assign n22892 = pi20 ? n18129 : ~n32;
  assign n22893 = pi19 ? n22891 : ~n22892;
  assign n22894 = pi20 ? n1331 : n243;
  assign n22895 = pi19 ? n22894 : ~n32;
  assign n22896 = pi18 ? n22893 : n22895;
  assign n22897 = pi17 ? n22890 : ~n22896;
  assign n22898 = pi16 ? n32 : n22897;
  assign n22899 = pi15 ? n22888 : n22898;
  assign n22900 = pi14 ? n13948 : n22899;
  assign n22901 = pi20 ? n220 : n243;
  assign n22902 = pi19 ? n22901 : ~n32;
  assign n22903 = pi18 ? n4380 : ~n22902;
  assign n22904 = pi17 ? n32 : n22903;
  assign n22905 = pi16 ? n32 : n22904;
  assign n22906 = pi18 ? n17118 : n20298;
  assign n22907 = pi17 ? n32 : n22906;
  assign n22908 = pi16 ? n32 : n22907;
  assign n22909 = pi15 ? n22905 : n22908;
  assign n22910 = pi21 ? n32 : ~n2076;
  assign n22911 = pi20 ? n22910 : ~n32;
  assign n22912 = pi19 ? n22911 : ~n32;
  assign n22913 = pi18 ? n32 : ~n22912;
  assign n22914 = pi17 ? n32 : n22913;
  assign n22915 = pi16 ? n32 : n22914;
  assign n22916 = pi15 ? n20048 : n22915;
  assign n22917 = pi14 ? n22909 : n22916;
  assign n22918 = pi13 ? n22900 : n22917;
  assign n22919 = pi12 ? n22884 : n22918;
  assign n22920 = pi11 ? n22881 : n22919;
  assign n22921 = pi10 ? n22835 : n22920;
  assign n22922 = pi09 ? n32 : n22921;
  assign n22923 = pi16 ? n32 : n1543;
  assign n22924 = pi14 ? n32 : n22923;
  assign n22925 = pi15 ? n22923 : n32;
  assign n22926 = pi14 ? n22925 : n32;
  assign n22927 = pi13 ? n22924 : n22926;
  assign n22928 = pi12 ? n32 : n22927;
  assign n22929 = pi14 ? n1109 : n32;
  assign n22930 = pi13 ? n22929 : n22827;
  assign n22931 = pi15 ? n22817 : n15123;
  assign n22932 = pi14 ? n22931 : n22347;
  assign n22933 = pi14 ? n22831 : n22437;
  assign n22934 = pi13 ? n22932 : n22933;
  assign n22935 = pi12 ? n22930 : n22934;
  assign n22936 = pi11 ? n22928 : n22935;
  assign n22937 = pi18 ? n4380 : ~n595;
  assign n22938 = pi17 ? n32 : n22937;
  assign n22939 = pi16 ? n32 : n22938;
  assign n22940 = pi20 ? n10644 : ~n1385;
  assign n22941 = pi19 ? n22940 : ~n32;
  assign n22942 = pi18 ? n32 : ~n22941;
  assign n22943 = pi17 ? n32 : n22942;
  assign n22944 = pi16 ? n32 : n22943;
  assign n22945 = pi15 ? n22939 : n22944;
  assign n22946 = pi20 ? n342 : n10644;
  assign n22947 = pi19 ? n22946 : n32;
  assign n22948 = pi18 ? n32 : n22947;
  assign n22949 = pi17 ? n32 : n22948;
  assign n22950 = pi16 ? n32 : n22949;
  assign n22951 = pi18 ? n4380 : n14590;
  assign n22952 = pi17 ? n32 : n22951;
  assign n22953 = pi16 ? n32 : n22952;
  assign n22954 = pi15 ? n22950 : n22953;
  assign n22955 = pi14 ? n22945 : n22954;
  assign n22956 = pi18 ? n32 : n22850;
  assign n22957 = pi17 ? n32 : n22956;
  assign n22958 = pi16 ? n32 : n22957;
  assign n22959 = pi15 ? n22958 : n14790;
  assign n22960 = pi20 ? n321 : ~n7880;
  assign n22961 = pi19 ? n22960 : ~n32;
  assign n22962 = pi18 ? n32 : ~n22961;
  assign n22963 = pi17 ? n32 : n22962;
  assign n22964 = pi16 ? n32 : n22963;
  assign n22965 = pi15 ? n22964 : n22650;
  assign n22966 = pi14 ? n22959 : n22965;
  assign n22967 = pi13 ? n22955 : n22966;
  assign n22968 = pi15 ? n22650 : n22868;
  assign n22969 = pi14 ? n22968 : n22876;
  assign n22970 = pi15 ? n21543 : n21695;
  assign n22971 = pi14 ? n21543 : n22970;
  assign n22972 = pi13 ? n22969 : n22971;
  assign n22973 = pi12 ? n22967 : n22972;
  assign n22974 = pi15 ? n14397 : n21033;
  assign n22975 = pi14 ? n21695 : n22974;
  assign n22976 = pi15 ? n20831 : n21232;
  assign n22977 = pi14 ? n20969 : n22976;
  assign n22978 = pi13 ? n22975 : n22977;
  assign n22979 = pi20 ? n1331 : n207;
  assign n22980 = pi19 ? n22979 : ~n32;
  assign n22981 = pi18 ? n22893 : n22980;
  assign n22982 = pi17 ? n22890 : ~n22981;
  assign n22983 = pi16 ? n32 : n22982;
  assign n22984 = pi15 ? n22888 : n22983;
  assign n22985 = pi14 ? n21232 : n22984;
  assign n22986 = pi18 ? n4380 : ~n6019;
  assign n22987 = pi17 ? n32 : n22986;
  assign n22988 = pi16 ? n32 : n22987;
  assign n22989 = pi20 ? n2140 : ~n243;
  assign n22990 = pi19 ? n22989 : n32;
  assign n22991 = pi18 ? n17118 : n22990;
  assign n22992 = pi17 ? n32 : n22991;
  assign n22993 = pi16 ? n32 : n22992;
  assign n22994 = pi15 ? n22988 : n22993;
  assign n22995 = pi20 ? n7880 : ~n32;
  assign n22996 = pi19 ? n22995 : ~n32;
  assign n22997 = pi18 ? n32 : ~n22996;
  assign n22998 = pi17 ? n32 : n22997;
  assign n22999 = pi16 ? n32 : n22998;
  assign n23000 = pi15 ? n20493 : n22999;
  assign n23001 = pi14 ? n22994 : n23000;
  assign n23002 = pi13 ? n22985 : n23001;
  assign n23003 = pi12 ? n22978 : n23002;
  assign n23004 = pi11 ? n22973 : n23003;
  assign n23005 = pi10 ? n22936 : n23004;
  assign n23006 = pi09 ? n32 : n23005;
  assign n23007 = pi08 ? n22922 : n23006;
  assign n23008 = pi19 ? n507 : ~n1105;
  assign n23009 = pi18 ? n32 : n23008;
  assign n23010 = pi17 ? n32 : n23009;
  assign n23011 = pi16 ? n32 : n23010;
  assign n23012 = pi15 ? n32 : n23011;
  assign n23013 = pi19 ? n1490 : ~n1105;
  assign n23014 = pi18 ? n32 : n23013;
  assign n23015 = pi17 ? n32 : n23014;
  assign n23016 = pi16 ? n32 : n23015;
  assign n23017 = pi19 ? n1325 : ~n1105;
  assign n23018 = pi18 ? n32 : n23017;
  assign n23019 = pi17 ? n32 : n23018;
  assign n23020 = pi16 ? n32 : n23019;
  assign n23021 = pi15 ? n23016 : n23020;
  assign n23022 = pi14 ? n23012 : n23021;
  assign n23023 = pi13 ? n32 : n23022;
  assign n23024 = pi14 ? n22540 : n22817;
  assign n23025 = pi15 ? n22817 : n22437;
  assign n23026 = pi20 ? n246 : n1385;
  assign n23027 = pi19 ? n23026 : n32;
  assign n23028 = pi18 ? n32 : n23027;
  assign n23029 = pi17 ? n32 : n23028;
  assign n23030 = pi16 ? n32 : n23029;
  assign n23031 = pi14 ? n23025 : n23030;
  assign n23032 = pi13 ? n23024 : n23031;
  assign n23033 = pi12 ? n23023 : n23032;
  assign n23034 = pi11 ? n22928 : n23033;
  assign n23035 = pi18 ? n32 : ~n595;
  assign n23036 = pi17 ? n32 : n23035;
  assign n23037 = pi16 ? n32 : n23036;
  assign n23038 = pi15 ? n23037 : n22437;
  assign n23039 = pi20 ? n246 : n7880;
  assign n23040 = pi19 ? n23039 : n32;
  assign n23041 = pi18 ? n32 : n23040;
  assign n23042 = pi17 ? n32 : n23041;
  assign n23043 = pi16 ? n32 : n23042;
  assign n23044 = pi15 ? n22950 : n23043;
  assign n23045 = pi14 ? n23038 : n23044;
  assign n23046 = pi18 ? n4380 : ~n22961;
  assign n23047 = pi17 ? n32 : n23046;
  assign n23048 = pi16 ? n32 : n23047;
  assign n23049 = pi15 ? n23048 : n22650;
  assign n23050 = pi14 ? n22959 : n23049;
  assign n23051 = pi13 ? n23045 : n23050;
  assign n23052 = pi18 ? n32 : n4380;
  assign n23053 = pi17 ? n23052 : n12522;
  assign n23054 = pi16 ? n32 : n23053;
  assign n23055 = pi17 ? n17346 : n12522;
  assign n23056 = pi16 ? n32 : n23055;
  assign n23057 = pi15 ? n23056 : n21543;
  assign n23058 = pi14 ? n23054 : n23057;
  assign n23059 = pi15 ? n387 : n21464;
  assign n23060 = pi14 ? n387 : n23059;
  assign n23061 = pi13 ? n23058 : n23060;
  assign n23062 = pi12 ? n23051 : n23061;
  assign n23063 = pi15 ? n14613 : n20836;
  assign n23064 = pi14 ? n21389 : n23063;
  assign n23065 = pi14 ? n21141 : n20831;
  assign n23066 = pi13 ? n23064 : n23065;
  assign n23067 = pi15 ? n12095 : n12538;
  assign n23068 = pi14 ? n20838 : n23067;
  assign n23069 = pi18 ? n4380 : n5749;
  assign n23070 = pi17 ? n32 : n23069;
  assign n23071 = pi16 ? n32 : n23070;
  assign n23072 = pi15 ? n23071 : n21162;
  assign n23073 = pi19 ? n6298 : ~n32;
  assign n23074 = pi18 ? n4380 : ~n23073;
  assign n23075 = pi17 ? n32 : n23074;
  assign n23076 = pi16 ? n32 : n23075;
  assign n23077 = pi15 ? n20776 : n23076;
  assign n23078 = pi14 ? n23072 : n23077;
  assign n23079 = pi13 ? n23068 : n23078;
  assign n23080 = pi12 ? n23066 : n23079;
  assign n23081 = pi11 ? n23062 : n23080;
  assign n23082 = pi10 ? n23034 : n23081;
  assign n23083 = pi09 ? n32 : n23082;
  assign n23084 = pi14 ? n32 : n15518;
  assign n23085 = pi15 ? n15518 : n32;
  assign n23086 = pi14 ? n23085 : n32;
  assign n23087 = pi13 ? n23084 : n23086;
  assign n23088 = pi12 ? n32 : n23087;
  assign n23089 = pi14 ? n22923 : n32;
  assign n23090 = pi13 ? n23089 : n23022;
  assign n23091 = pi19 ? n17655 : n32;
  assign n23092 = pi18 ? n32 : n23091;
  assign n23093 = pi17 ? n32 : n23092;
  assign n23094 = pi16 ? n32 : n23093;
  assign n23095 = pi15 ? n22817 : n23094;
  assign n23096 = pi20 ? n246 : n17654;
  assign n23097 = pi19 ? n23096 : n32;
  assign n23098 = pi18 ? n32 : n23097;
  assign n23099 = pi17 ? n32 : n23098;
  assign n23100 = pi16 ? n32 : n23099;
  assign n23101 = pi14 ? n23095 : n23100;
  assign n23102 = pi13 ? n23024 : n23101;
  assign n23103 = pi12 ? n23090 : n23102;
  assign n23104 = pi11 ? n23088 : n23103;
  assign n23105 = pi15 ? n13035 : n23094;
  assign n23106 = pi20 ? n342 : n13084;
  assign n23107 = pi19 ? n23106 : n32;
  assign n23108 = pi18 ? n32 : n23107;
  assign n23109 = pi17 ? n32 : n23108;
  assign n23110 = pi16 ? n32 : n23109;
  assign n23111 = pi15 ? n23110 : n23030;
  assign n23112 = pi14 ? n23105 : n23111;
  assign n23113 = pi15 ? n14593 : n22437;
  assign n23114 = pi20 ? n321 : ~n1385;
  assign n23115 = pi19 ? n23114 : ~n32;
  assign n23116 = pi18 ? n4380 : ~n23115;
  assign n23117 = pi17 ? n32 : n23116;
  assign n23118 = pi16 ? n32 : n23117;
  assign n23119 = pi15 ? n23118 : n22749;
  assign n23120 = pi14 ? n23113 : n23119;
  assign n23121 = pi13 ? n23112 : n23120;
  assign n23122 = pi21 ? n32 : n7410;
  assign n23123 = pi20 ? n32 : n23122;
  assign n23124 = pi19 ? n23123 : ~n32;
  assign n23125 = pi18 ? n940 : ~n23124;
  assign n23126 = pi17 ? n23052 : n23125;
  assign n23127 = pi16 ? n32 : n23126;
  assign n23128 = pi18 ? n940 : ~n520;
  assign n23129 = pi17 ? n23052 : n23128;
  assign n23130 = pi16 ? n32 : n23129;
  assign n23131 = pi15 ? n23127 : n23130;
  assign n23132 = pi17 ? n17346 : n23128;
  assign n23133 = pi16 ? n32 : n23132;
  assign n23134 = pi15 ? n23133 : n21686;
  assign n23135 = pi14 ? n23131 : n23134;
  assign n23136 = pi14 ? n21786 : n21681;
  assign n23137 = pi13 ? n23135 : n23136;
  assign n23138 = pi12 ? n23121 : n23137;
  assign n23139 = pi15 ? n21319 : n21033;
  assign n23140 = pi14 ? n22381 : n23139;
  assign n23141 = pi14 ? n20967 : n20836;
  assign n23142 = pi13 ? n23140 : n23141;
  assign n23143 = pi15 ? n12091 : n12535;
  assign n23144 = pi14 ? n32 : n23143;
  assign n23145 = pi18 ? n4380 : n21487;
  assign n23146 = pi17 ? n32 : n23145;
  assign n23147 = pi16 ? n32 : n23146;
  assign n23148 = pi15 ? n23147 : n21162;
  assign n23149 = pi14 ? n23148 : n23077;
  assign n23150 = pi13 ? n23144 : n23149;
  assign n23151 = pi12 ? n23142 : n23150;
  assign n23152 = pi11 ? n23138 : n23151;
  assign n23153 = pi10 ? n23104 : n23152;
  assign n23154 = pi09 ? n32 : n23153;
  assign n23155 = pi08 ? n23083 : n23154;
  assign n23156 = pi07 ? n23007 : n23155;
  assign n23157 = pi19 ? n32 : n5626;
  assign n23158 = pi18 ? n32 : n23157;
  assign n23159 = pi17 ? n32 : n23158;
  assign n23160 = pi16 ? n32 : n23159;
  assign n23161 = pi14 ? n32 : n23160;
  assign n23162 = pi15 ? n23160 : n32;
  assign n23163 = pi14 ? n23162 : n32;
  assign n23164 = pi13 ? n23161 : n23163;
  assign n23165 = pi12 ? n32 : n23164;
  assign n23166 = pi19 ? n1464 : ~n617;
  assign n23167 = pi18 ? n32 : n23166;
  assign n23168 = pi17 ? n32 : n23167;
  assign n23169 = pi16 ? n32 : n23168;
  assign n23170 = pi15 ? n32 : n23169;
  assign n23171 = pi14 ? n23170 : n22923;
  assign n23172 = pi13 ? n32 : n23171;
  assign n23173 = pi14 ? n1109 : n23011;
  assign n23174 = pi15 ? n22728 : n22347;
  assign n23175 = pi14 ? n23174 : n15389;
  assign n23176 = pi13 ? n23173 : n23175;
  assign n23177 = pi12 ? n23172 : n23176;
  assign n23178 = pi11 ? n23165 : n23177;
  assign n23179 = pi15 ? n15389 : n22347;
  assign n23180 = pi20 ? n266 : n175;
  assign n23181 = pi19 ? n23180 : n32;
  assign n23182 = pi18 ? n936 : n23181;
  assign n23183 = pi17 ? n32 : n23182;
  assign n23184 = pi16 ? n32 : n23183;
  assign n23185 = pi15 ? n15389 : n23184;
  assign n23186 = pi14 ? n23179 : n23185;
  assign n23187 = pi18 ? n32 : ~n2627;
  assign n23188 = pi17 ? n32 : n23187;
  assign n23189 = pi16 ? n32 : n23188;
  assign n23190 = pi15 ? n23037 : n23189;
  assign n23191 = pi14 ? n22437 : n23190;
  assign n23192 = pi13 ? n23186 : n23191;
  assign n23193 = pi20 ? n32 : n12884;
  assign n23194 = pi19 ? n32 : n23193;
  assign n23195 = pi18 ? n23194 : ~n508;
  assign n23196 = pi17 ? n32 : n23195;
  assign n23197 = pi16 ? n32 : n23196;
  assign n23198 = pi15 ? n13040 : n23197;
  assign n23199 = pi20 ? n207 : ~n3523;
  assign n23200 = pi19 ? n23199 : ~n32;
  assign n23201 = pi18 ? n463 : ~n23200;
  assign n23202 = pi17 ? n32 : n23201;
  assign n23203 = pi16 ? n32 : n23202;
  assign n23204 = pi15 ? n23203 : n21786;
  assign n23205 = pi14 ? n23198 : n23204;
  assign n23206 = pi13 ? n23205 : n23136;
  assign n23207 = pi12 ? n23192 : n23206;
  assign n23208 = pi20 ? n32 : n16369;
  assign n23209 = pi19 ? n23208 : n32;
  assign n23210 = pi18 ? n32 : n23209;
  assign n23211 = pi17 ? n32 : n23210;
  assign n23212 = pi16 ? n32 : n23211;
  assign n23213 = pi14 ? n23212 : n21866;
  assign n23214 = pi14 ? n23063 : n20836;
  assign n23215 = pi13 ? n23213 : n23214;
  assign n23216 = pi15 ? n20836 : n12538;
  assign n23217 = pi19 ? n7823 : ~n32;
  assign n23218 = pi18 ? n863 : ~n23217;
  assign n23219 = pi17 ? n32 : n23218;
  assign n23220 = pi16 ? n32 : n23219;
  assign n23221 = pi15 ? n12535 : n23220;
  assign n23222 = pi14 ? n23216 : n23221;
  assign n23223 = pi19 ? n9874 : ~n32;
  assign n23224 = pi18 ? n32 : ~n23223;
  assign n23225 = pi17 ? n32 : n23224;
  assign n23226 = pi16 ? n32 : n23225;
  assign n23227 = pi20 ? n1324 : ~n243;
  assign n23228 = pi19 ? n23227 : n32;
  assign n23229 = pi18 ? n863 : n23228;
  assign n23230 = pi17 ? n32 : n23229;
  assign n23231 = pi16 ? n32 : n23230;
  assign n23232 = pi15 ? n23226 : n23231;
  assign n23233 = pi20 ? n220 : ~n141;
  assign n23234 = pi19 ? n23233 : n32;
  assign n23235 = pi18 ? n863 : n23234;
  assign n23236 = pi17 ? n32 : n23235;
  assign n23237 = pi16 ? n32 : n23236;
  assign n23238 = pi18 ? n863 : ~n344;
  assign n23239 = pi17 ? n32 : n23238;
  assign n23240 = pi16 ? n32 : n23239;
  assign n23241 = pi15 ? n23237 : n23240;
  assign n23242 = pi14 ? n23232 : n23241;
  assign n23243 = pi13 ? n23222 : n23242;
  assign n23244 = pi12 ? n23215 : n23243;
  assign n23245 = pi11 ? n23207 : n23244;
  assign n23246 = pi10 ? n23178 : n23245;
  assign n23247 = pi09 ? n32 : n23246;
  assign n23248 = pi18 ? n32 : n6114;
  assign n23249 = pi17 ? n32 : n23248;
  assign n23250 = pi16 ? n32 : n23249;
  assign n23251 = pi14 ? n32 : n23250;
  assign n23252 = pi15 ? n23250 : n32;
  assign n23253 = pi14 ? n23252 : n32;
  assign n23254 = pi13 ? n23251 : n23253;
  assign n23255 = pi12 ? n32 : n23254;
  assign n23256 = pi14 ? n23160 : n32;
  assign n23257 = pi13 ? n23256 : n23171;
  assign n23258 = pi14 ? n32 : n23011;
  assign n23259 = pi15 ? n22728 : n22817;
  assign n23260 = pi14 ? n23259 : n22540;
  assign n23261 = pi13 ? n23258 : n23260;
  assign n23262 = pi12 ? n23257 : n23261;
  assign n23263 = pi11 ? n23255 : n23262;
  assign n23264 = pi15 ? n22540 : n22817;
  assign n23265 = pi20 ? n266 : n13387;
  assign n23266 = pi19 ? n23265 : n32;
  assign n23267 = pi18 ? n936 : n23266;
  assign n23268 = pi17 ? n32 : n23267;
  assign n23269 = pi16 ? n32 : n23268;
  assign n23270 = pi15 ? n22540 : n23269;
  assign n23271 = pi14 ? n23264 : n23270;
  assign n23272 = pi15 ? n13035 : n23037;
  assign n23273 = pi14 ? n23094 : n23272;
  assign n23274 = pi13 ? n23271 : n23273;
  assign n23275 = pi15 ? n23189 : n23197;
  assign n23276 = pi20 ? n207 : ~n151;
  assign n23277 = pi19 ? n23276 : ~n32;
  assign n23278 = pi18 ? n32 : ~n23277;
  assign n23279 = pi17 ? n32 : n23278;
  assign n23280 = pi16 ? n32 : n23279;
  assign n23281 = pi15 ? n23280 : n476;
  assign n23282 = pi14 ? n23275 : n23281;
  assign n23283 = pi14 ? n477 : n21787;
  assign n23284 = pi13 ? n23282 : n23283;
  assign n23285 = pi12 ? n23274 : n23284;
  assign n23286 = pi15 ? n21389 : n658;
  assign n23287 = pi14 ? n22376 : n23286;
  assign n23288 = pi14 ? n20967 : n21033;
  assign n23289 = pi13 ? n23287 : n23288;
  assign n23290 = pi15 ? n21033 : n12531;
  assign n23291 = pi19 ? n7813 : ~n32;
  assign n23292 = pi18 ? n863 : ~n23291;
  assign n23293 = pi17 ? n32 : n23292;
  assign n23294 = pi16 ? n32 : n23293;
  assign n23295 = pi15 ? n12531 : n23294;
  assign n23296 = pi14 ? n23290 : n23295;
  assign n23297 = pi19 ? n13512 : ~n32;
  assign n23298 = pi18 ? n32 : ~n23297;
  assign n23299 = pi17 ? n32 : n23298;
  assign n23300 = pi16 ? n32 : n23299;
  assign n23301 = pi20 ? n1324 : ~n207;
  assign n23302 = pi19 ? n23301 : n32;
  assign n23303 = pi18 ? n863 : n23302;
  assign n23304 = pi17 ? n32 : n23303;
  assign n23305 = pi16 ? n32 : n23304;
  assign n23306 = pi15 ? n23300 : n23305;
  assign n23307 = pi20 ? n220 : ~n339;
  assign n23308 = pi19 ? n23307 : n32;
  assign n23309 = pi18 ? n863 : n23308;
  assign n23310 = pi17 ? n32 : n23309;
  assign n23311 = pi16 ? n32 : n23310;
  assign n23312 = pi19 ? n10072 : ~n32;
  assign n23313 = pi18 ? n863 : ~n23312;
  assign n23314 = pi17 ? n32 : n23313;
  assign n23315 = pi16 ? n32 : n23314;
  assign n23316 = pi15 ? n23311 : n23315;
  assign n23317 = pi14 ? n23306 : n23316;
  assign n23318 = pi13 ? n23296 : n23317;
  assign n23319 = pi12 ? n23289 : n23318;
  assign n23320 = pi11 ? n23285 : n23319;
  assign n23321 = pi10 ? n23263 : n23320;
  assign n23322 = pi09 ? n32 : n23321;
  assign n23323 = pi08 ? n23247 : n23322;
  assign n23324 = pi15 ? n32 : n15836;
  assign n23325 = pi14 ? n23324 : n15836;
  assign n23326 = pi15 ? n15836 : n32;
  assign n23327 = pi14 ? n23326 : n32;
  assign n23328 = pi13 ? n23325 : n23327;
  assign n23329 = pi12 ? n32 : n23328;
  assign n23330 = pi19 ? n1464 : ~n2614;
  assign n23331 = pi18 ? n32 : n23330;
  assign n23332 = pi17 ? n32 : n23331;
  assign n23333 = pi16 ? n32 : n23332;
  assign n23334 = pi15 ? n23160 : n23333;
  assign n23335 = pi14 ? n23334 : n15518;
  assign n23336 = pi13 ? n32 : n23335;
  assign n23337 = pi14 ? n22923 : n15119;
  assign n23338 = pi18 ? n32 : n6380;
  assign n23339 = pi17 ? n32 : n23338;
  assign n23340 = pi16 ? n32 : n23339;
  assign n23341 = pi15 ? n23340 : n22817;
  assign n23342 = pi14 ? n23341 : n22540;
  assign n23343 = pi13 ? n23337 : n23342;
  assign n23344 = pi12 ? n23336 : n23343;
  assign n23345 = pi11 ? n23329 : n23344;
  assign n23346 = pi20 ? n206 : n175;
  assign n23347 = pi19 ? n23346 : n32;
  assign n23348 = pi18 ? n32 : n23347;
  assign n23349 = pi17 ? n32 : n23348;
  assign n23350 = pi16 ? n32 : n23349;
  assign n23351 = pi15 ? n22817 : n23350;
  assign n23352 = pi14 ? n23264 : n23351;
  assign n23353 = pi15 ? n23094 : n22347;
  assign n23354 = pi18 ? n19082 : ~n4098;
  assign n23355 = pi17 ? n32 : n23354;
  assign n23356 = pi16 ? n32 : n23355;
  assign n23357 = pi18 ? n19082 : ~n595;
  assign n23358 = pi17 ? n32 : n23357;
  assign n23359 = pi16 ? n32 : n23358;
  assign n23360 = pi15 ? n23356 : n23359;
  assign n23361 = pi14 ? n23353 : n23360;
  assign n23362 = pi13 ? n23352 : n23361;
  assign n23363 = pi19 ? n247 : n6057;
  assign n23364 = pi18 ? n23363 : ~n2627;
  assign n23365 = pi17 ? n4282 : n23364;
  assign n23366 = pi16 ? n32 : n23365;
  assign n23367 = pi18 ? n9170 : ~n2627;
  assign n23368 = pi17 ? n3282 : n23367;
  assign n23369 = pi16 ? n32 : n23368;
  assign n23370 = pi15 ? n23366 : n23369;
  assign n23371 = pi14 ? n23370 : n21928;
  assign n23372 = pi14 ? n22213 : n21681;
  assign n23373 = pi13 ? n23371 : n23372;
  assign n23374 = pi12 ? n23362 : n23373;
  assign n23375 = pi21 ? n100 : ~n242;
  assign n23376 = pi20 ? n32 : n23375;
  assign n23377 = pi19 ? n23376 : n32;
  assign n23378 = pi18 ? n32 : n23377;
  assign n23379 = pi17 ? n32 : n23378;
  assign n23380 = pi16 ? n32 : n23379;
  assign n23381 = pi15 ? n21686 : n23380;
  assign n23382 = pi15 ? n23212 : n658;
  assign n23383 = pi14 ? n23381 : n23382;
  assign n23384 = pi13 ? n23383 : n32;
  assign n23385 = pi18 ? n940 : ~n2291;
  assign n23386 = pi17 ? n17119 : n23385;
  assign n23387 = pi16 ? n32 : n23386;
  assign n23388 = pi15 ? n20836 : n23387;
  assign n23389 = pi17 ? n32 : n23385;
  assign n23390 = pi16 ? n32 : n23389;
  assign n23391 = pi18 ? n936 : ~n2291;
  assign n23392 = pi17 ? n32 : n23391;
  assign n23393 = pi16 ? n32 : n23392;
  assign n23394 = pi15 ? n23390 : n23393;
  assign n23395 = pi14 ? n23388 : n23394;
  assign n23396 = pi20 ? n342 : n1475;
  assign n23397 = pi19 ? n23396 : ~n32;
  assign n23398 = pi18 ? n936 : ~n23397;
  assign n23399 = pi17 ? n32 : n23398;
  assign n23400 = pi16 ? n32 : n23399;
  assign n23401 = pi19 ? n17766 : n32;
  assign n23402 = pi18 ? n863 : n23401;
  assign n23403 = pi17 ? n32 : n23402;
  assign n23404 = pi16 ? n32 : n23403;
  assign n23405 = pi15 ? n23400 : n23404;
  assign n23406 = pi20 ? n220 : ~n243;
  assign n23407 = pi19 ? n23406 : n32;
  assign n23408 = pi18 ? n863 : n23407;
  assign n23409 = pi17 ? n32 : n23408;
  assign n23410 = pi16 ? n32 : n23409;
  assign n23411 = pi18 ? n863 : ~n3786;
  assign n23412 = pi17 ? n32 : n23411;
  assign n23413 = pi16 ? n32 : n23412;
  assign n23414 = pi15 ? n23410 : n23413;
  assign n23415 = pi14 ? n23405 : n23414;
  assign n23416 = pi13 ? n23395 : n23415;
  assign n23417 = pi12 ? n23384 : n23416;
  assign n23418 = pi11 ? n23374 : n23417;
  assign n23419 = pi10 ? n23345 : n23418;
  assign n23420 = pi09 ? n32 : n23419;
  assign n23421 = pi15 ? n32 : n16108;
  assign n23422 = pi14 ? n23421 : n16108;
  assign n23423 = pi14 ? n16110 : n32;
  assign n23424 = pi13 ? n23422 : n23423;
  assign n23425 = pi12 ? n32 : n23424;
  assign n23426 = pi14 ? n23250 : n32;
  assign n23427 = pi13 ? n23426 : n23335;
  assign n23428 = pi15 ? n23340 : n23011;
  assign n23429 = pi14 ? n23428 : n22728;
  assign n23430 = pi13 ? n23337 : n23429;
  assign n23431 = pi12 ? n23427 : n23430;
  assign n23432 = pi11 ? n23425 : n23431;
  assign n23433 = pi15 ? n22728 : n23011;
  assign n23434 = pi19 ? n19151 : n32;
  assign n23435 = pi18 ? n32 : n23434;
  assign n23436 = pi17 ? n32 : n23435;
  assign n23437 = pi16 ? n32 : n23436;
  assign n23438 = pi15 ? n22817 : n23437;
  assign n23439 = pi14 ? n23433 : n23438;
  assign n23440 = pi19 ? n322 : n32;
  assign n23441 = pi18 ? n32 : n23440;
  assign n23442 = pi17 ? n32 : n23441;
  assign n23443 = pi16 ? n32 : n23442;
  assign n23444 = pi19 ? n2141 : n32;
  assign n23445 = pi18 ? n32 : n23444;
  assign n23446 = pi17 ? n32 : n23445;
  assign n23447 = pi16 ? n32 : n23446;
  assign n23448 = pi15 ? n23443 : n23447;
  assign n23449 = pi18 ? n19082 : ~n702;
  assign n23450 = pi17 ? n32 : n23449;
  assign n23451 = pi16 ? n32 : n23450;
  assign n23452 = pi15 ? n23451 : n23356;
  assign n23453 = pi14 ? n23448 : n23452;
  assign n23454 = pi13 ? n23439 : n23453;
  assign n23455 = pi18 ? n23363 : ~n508;
  assign n23456 = pi17 ? n4282 : n23455;
  assign n23457 = pi16 ? n32 : n23456;
  assign n23458 = pi18 ? n9170 : ~n508;
  assign n23459 = pi17 ? n3282 : n23458;
  assign n23460 = pi16 ? n32 : n23459;
  assign n23461 = pi15 ? n23457 : n23460;
  assign n23462 = pi14 ? n23461 : n648;
  assign n23463 = pi14 ? n648 : n22638;
  assign n23464 = pi13 ? n23462 : n23463;
  assign n23465 = pi12 ? n23454 : n23464;
  assign n23466 = pi15 ? n21543 : n32;
  assign n23467 = pi14 ? n21853 : n23466;
  assign n23468 = pi14 ? n21319 : n21627;
  assign n23469 = pi13 ? n23467 : n23468;
  assign n23470 = pi18 ? n863 : ~n418;
  assign n23471 = pi17 ? n32 : n23470;
  assign n23472 = pi16 ? n32 : n23471;
  assign n23473 = pi15 ? n23311 : n23472;
  assign n23474 = pi14 ? n23405 : n23473;
  assign n23475 = pi13 ? n23395 : n23474;
  assign n23476 = pi12 ? n23469 : n23475;
  assign n23477 = pi11 ? n23465 : n23476;
  assign n23478 = pi10 ? n23432 : n23477;
  assign n23479 = pi09 ? n32 : n23478;
  assign n23480 = pi08 ? n23420 : n23479;
  assign n23481 = pi07 ? n23323 : n23480;
  assign n23482 = pi06 ? n23156 : n23481;
  assign n23483 = pi17 ? n32 : n20173;
  assign n23484 = pi16 ? n32 : n23483;
  assign n23485 = pi15 ? n23250 : n23484;
  assign n23486 = pi14 ? n23485 : n23484;
  assign n23487 = pi13 ? n32 : n23486;
  assign n23488 = pi14 ? n23160 : n15518;
  assign n23489 = pi20 ? n32 : ~n10644;
  assign n23490 = pi19 ? n23489 : ~n2614;
  assign n23491 = pi18 ? n32 : n23490;
  assign n23492 = pi17 ? n32 : n23491;
  assign n23493 = pi16 ? n32 : n23492;
  assign n23494 = pi19 ? n23489 : n32;
  assign n23495 = pi18 ? n32 : n23494;
  assign n23496 = pi17 ? n32 : n23495;
  assign n23497 = pi16 ? n32 : n23496;
  assign n23498 = pi15 ? n23493 : n23497;
  assign n23499 = pi14 ? n23498 : n1109;
  assign n23500 = pi13 ? n23488 : n23499;
  assign n23501 = pi12 ? n23487 : n23500;
  assign n23502 = pi11 ? n23425 : n23501;
  assign n23503 = pi15 ? n1109 : n23011;
  assign n23504 = pi19 ? n20555 : n32;
  assign n23505 = pi18 ? n32 : n23504;
  assign n23506 = pi17 ? n32 : n23505;
  assign n23507 = pi16 ? n32 : n23506;
  assign n23508 = pi19 ? n4391 : n32;
  assign n23509 = pi18 ? n32 : n23508;
  assign n23510 = pi17 ? n32 : n23509;
  assign n23511 = pi16 ? n32 : n23510;
  assign n23512 = pi15 ? n23507 : n23511;
  assign n23513 = pi14 ? n23503 : n23512;
  assign n23514 = pi19 ? n236 : n32;
  assign n23515 = pi18 ? n32 : n23514;
  assign n23516 = pi17 ? n32 : n23515;
  assign n23517 = pi16 ? n32 : n23516;
  assign n23518 = pi18 ? n863 : n23514;
  assign n23519 = pi17 ? n32 : n23518;
  assign n23520 = pi16 ? n32 : n23519;
  assign n23521 = pi15 ? n23517 : n23520;
  assign n23522 = pi14 ? n23264 : n23521;
  assign n23523 = pi13 ? n23513 : n23522;
  assign n23524 = pi20 ? n220 : ~n11107;
  assign n23525 = pi19 ? n23524 : n32;
  assign n23526 = pi18 ? n4380 : n23525;
  assign n23527 = pi17 ? n32 : n23526;
  assign n23528 = pi16 ? n32 : n23527;
  assign n23529 = pi15 ? n23528 : n32;
  assign n23530 = pi14 ? n23529 : n32;
  assign n23531 = pi14 ? n32 : n14973;
  assign n23532 = pi13 ? n23530 : n23531;
  assign n23533 = pi12 ? n23523 : n23532;
  assign n23534 = pi15 ? n21686 : n21464;
  assign n23535 = pi14 ? n14790 : n23534;
  assign n23536 = pi13 ? n23535 : n32;
  assign n23537 = pi19 ? n6398 : n349;
  assign n23538 = pi18 ? n32 : n23537;
  assign n23539 = pi19 ? n5694 : n247;
  assign n23540 = pi18 ? n23539 : n323;
  assign n23541 = pi17 ? n23538 : ~n23540;
  assign n23542 = pi16 ? n32 : n23541;
  assign n23543 = pi19 ? n9037 : ~n32;
  assign n23544 = pi18 ? n940 : ~n23543;
  assign n23545 = pi17 ? n32 : n23544;
  assign n23546 = pi16 ? n32 : n23545;
  assign n23547 = pi15 ? n23542 : n23546;
  assign n23548 = pi19 ? n15405 : n32;
  assign n23549 = pi18 ? n32 : n23548;
  assign n23550 = pi17 ? n32 : n23549;
  assign n23551 = pi16 ? n32 : n23550;
  assign n23552 = pi14 ? n23547 : n23551;
  assign n23553 = pi20 ? n207 : ~n1475;
  assign n23554 = pi19 ? n23553 : n32;
  assign n23555 = pi18 ? n32 : n23554;
  assign n23556 = pi17 ? n32 : n23555;
  assign n23557 = pi16 ? n32 : n23556;
  assign n23558 = pi15 ? n23557 : n13948;
  assign n23559 = pi18 ? n32 : ~n418;
  assign n23560 = pi17 ? n32 : n23559;
  assign n23561 = pi16 ? n32 : n23560;
  assign n23562 = pi15 ? n13375 : n23561;
  assign n23563 = pi14 ? n23558 : n23562;
  assign n23564 = pi13 ? n23552 : n23563;
  assign n23565 = pi12 ? n23536 : n23564;
  assign n23566 = pi11 ? n23533 : n23565;
  assign n23567 = pi10 ? n23502 : n23566;
  assign n23568 = pi09 ? n32 : n23567;
  assign n23569 = pi16 ? n32 : n1633;
  assign n23570 = pi15 ? n32 : n23569;
  assign n23571 = pi19 ? n32 : n5614;
  assign n23572 = pi18 ? n32 : n23571;
  assign n23573 = pi17 ? n32 : n23572;
  assign n23574 = pi16 ? n32 : n23573;
  assign n23575 = pi14 ? n23570 : n23574;
  assign n23576 = pi15 ? n23574 : n32;
  assign n23577 = pi14 ? n23576 : n32;
  assign n23578 = pi13 ? n23575 : n23577;
  assign n23579 = pi12 ? n32 : n23578;
  assign n23580 = pi14 ? n16108 : n32;
  assign n23581 = pi13 ? n23580 : n23486;
  assign n23582 = pi15 ? n32 : n23160;
  assign n23583 = pi14 ? n23582 : n15518;
  assign n23584 = pi19 ? n23489 : ~n617;
  assign n23585 = pi18 ? n32 : n23584;
  assign n23586 = pi17 ? n32 : n23585;
  assign n23587 = pi16 ? n32 : n23586;
  assign n23588 = pi15 ? n23493 : n23587;
  assign n23589 = pi14 ? n23588 : n22923;
  assign n23590 = pi13 ? n23583 : n23589;
  assign n23591 = pi12 ? n23581 : n23590;
  assign n23592 = pi11 ? n23579 : n23591;
  assign n23593 = pi15 ? n22923 : n15119;
  assign n23594 = pi19 ? n20555 : ~n617;
  assign n23595 = pi18 ? n32 : n23594;
  assign n23596 = pi17 ? n32 : n23595;
  assign n23597 = pi16 ? n32 : n23596;
  assign n23598 = pi15 ? n23597 : n23511;
  assign n23599 = pi14 ? n23593 : n23598;
  assign n23600 = pi15 ? n13321 : n23520;
  assign n23601 = pi14 ? n23433 : n23600;
  assign n23602 = pi13 ? n23599 : n23601;
  assign n23603 = pi15 ? n23528 : n15263;
  assign n23604 = pi15 ? n15123 : n15263;
  assign n23605 = pi14 ? n23603 : n23604;
  assign n23606 = pi14 ? n15127 : n14973;
  assign n23607 = pi13 ? n23605 : n23606;
  assign n23608 = pi12 ? n23602 : n23607;
  assign n23609 = pi15 ? n21686 : n32;
  assign n23610 = pi14 ? n14790 : n23609;
  assign n23611 = pi13 ? n23610 : n21464;
  assign n23612 = pi18 ? n32 : ~n2424;
  assign n23613 = pi17 ? n32 : n23612;
  assign n23614 = pi16 ? n32 : n23613;
  assign n23615 = pi15 ? n21254 : n23614;
  assign n23616 = pi14 ? n23558 : n23615;
  assign n23617 = pi13 ? n23552 : n23616;
  assign n23618 = pi12 ? n23611 : n23617;
  assign n23619 = pi11 ? n23608 : n23618;
  assign n23620 = pi10 ? n23592 : n23619;
  assign n23621 = pi09 ? n32 : n23620;
  assign n23622 = pi08 ? n23568 : n23621;
  assign n23623 = pi15 ? n32 : n23574;
  assign n23624 = pi14 ? n23623 : n23574;
  assign n23625 = pi13 ? n23624 : n23577;
  assign n23626 = pi12 ? n32 : n23625;
  assign n23627 = pi14 ? n32 : n23421;
  assign n23628 = pi19 ? n32 : n7502;
  assign n23629 = pi18 ? n32 : n23628;
  assign n23630 = pi17 ? n32 : n23629;
  assign n23631 = pi16 ? n32 : n23630;
  assign n23632 = pi15 ? n23631 : n23250;
  assign n23633 = pi14 ? n23631 : n23632;
  assign n23634 = pi13 ? n23627 : n23633;
  assign n23635 = pi19 ? n23489 : ~n236;
  assign n23636 = pi18 ? n32 : n23635;
  assign n23637 = pi17 ? n32 : n23636;
  assign n23638 = pi16 ? n32 : n23637;
  assign n23639 = pi15 ? n23638 : n23340;
  assign n23640 = pi14 ? n23639 : n22923;
  assign n23641 = pi13 ? n23486 : n23640;
  assign n23642 = pi12 ? n23634 : n23641;
  assign n23643 = pi11 ? n23626 : n23642;
  assign n23644 = pi20 ? n266 : n246;
  assign n23645 = pi19 ? n23644 : n617;
  assign n23646 = pi18 ? n863 : ~n23645;
  assign n23647 = pi17 ? n32 : n23646;
  assign n23648 = pi16 ? n32 : n23647;
  assign n23649 = pi19 ? n4391 : ~n617;
  assign n23650 = pi18 ? n32 : n23649;
  assign n23651 = pi17 ? n32 : n23650;
  assign n23652 = pi16 ? n32 : n23651;
  assign n23653 = pi15 ? n23648 : n23652;
  assign n23654 = pi14 ? n23593 : n23653;
  assign n23655 = pi19 ? n22106 : ~n617;
  assign n23656 = pi18 ? n32 : n23655;
  assign n23657 = pi17 ? n32 : n23656;
  assign n23658 = pi16 ? n32 : n23657;
  assign n23659 = pi15 ? n23658 : n13025;
  assign n23660 = pi19 ? n321 : ~n18489;
  assign n23661 = pi19 ? n617 : ~n1105;
  assign n23662 = pi18 ? n23660 : ~n23661;
  assign n23663 = pi17 ? n32 : ~n23662;
  assign n23664 = pi16 ? n32 : n23663;
  assign n23665 = pi15 ? n13025 : n23664;
  assign n23666 = pi14 ? n23659 : n23665;
  assign n23667 = pi13 ? n23654 : n23666;
  assign n23668 = pi21 ? n174 : n100;
  assign n23669 = pi20 ? n749 : ~n23668;
  assign n23670 = pi19 ? n23669 : n32;
  assign n23671 = pi18 ? n32 : n23670;
  assign n23672 = pi17 ? n32 : n23671;
  assign n23673 = pi16 ? n32 : n23672;
  assign n23674 = pi15 ? n23673 : n32;
  assign n23675 = pi14 ? n23674 : n32;
  assign n23676 = pi14 ? n22252 : n22635;
  assign n23677 = pi13 ? n23675 : n23676;
  assign n23678 = pi12 ? n23667 : n23677;
  assign n23679 = pi15 ? n22437 : n14790;
  assign n23680 = pi20 ? n321 : n7467;
  assign n23681 = pi19 ? n23680 : n32;
  assign n23682 = pi18 ? n32 : n23681;
  assign n23683 = pi17 ? n32 : n23682;
  assign n23684 = pi16 ? n32 : n23683;
  assign n23685 = pi15 ? n23684 : n32;
  assign n23686 = pi14 ? n23679 : n23685;
  assign n23687 = pi13 ? n23686 : n21466;
  assign n23688 = pi20 ? n321 : n428;
  assign n23689 = pi19 ? n23688 : ~n4342;
  assign n23690 = pi18 ? n23689 : ~n2754;
  assign n23691 = pi17 ? n2733 : n23690;
  assign n23692 = pi16 ? n32 : n23691;
  assign n23693 = pi20 ? n246 : n1839;
  assign n23694 = pi19 ? n23693 : ~n32;
  assign n23695 = pi18 ? n940 : ~n23694;
  assign n23696 = pi17 ? n32 : n23695;
  assign n23697 = pi16 ? n32 : n23696;
  assign n23698 = pi15 ? n23692 : n23697;
  assign n23699 = pi20 ? n207 : ~n1839;
  assign n23700 = pi19 ? n23699 : n32;
  assign n23701 = pi18 ? n32 : n23700;
  assign n23702 = pi17 ? n32 : n23701;
  assign n23703 = pi16 ? n32 : n23702;
  assign n23704 = pi15 ? n23703 : n23551;
  assign n23705 = pi14 ? n23698 : n23704;
  assign n23706 = pi18 ? n32 : n21724;
  assign n23707 = pi17 ? n32 : n23706;
  assign n23708 = pi16 ? n32 : n23707;
  assign n23709 = pi20 ? n274 : n220;
  assign n23710 = pi19 ? n23709 : n32;
  assign n23711 = pi18 ? n32 : n23710;
  assign n23712 = pi18 ? n32 : ~n21749;
  assign n23713 = pi17 ? n23711 : n23712;
  assign n23714 = pi16 ? n32 : n23713;
  assign n23715 = pi15 ? n23708 : n23714;
  assign n23716 = pi14 ? n23558 : n23715;
  assign n23717 = pi13 ? n23705 : n23716;
  assign n23718 = pi12 ? n23687 : n23717;
  assign n23719 = pi11 ? n23678 : n23718;
  assign n23720 = pi10 ? n23643 : n23719;
  assign n23721 = pi09 ? n32 : n23720;
  assign n23722 = pi19 ? n32 : n6230;
  assign n23723 = pi18 ? n32 : n23722;
  assign n23724 = pi17 ? n32 : n23723;
  assign n23725 = pi16 ? n32 : n23724;
  assign n23726 = pi15 ? n32 : n23725;
  assign n23727 = pi19 ? n32 : n7488;
  assign n23728 = pi18 ? n32 : n23727;
  assign n23729 = pi17 ? n32 : n23728;
  assign n23730 = pi16 ? n32 : n23729;
  assign n23731 = pi14 ? n23726 : n23730;
  assign n23732 = pi15 ? n23730 : n32;
  assign n23733 = pi14 ? n23732 : n32;
  assign n23734 = pi13 ? n23731 : n23733;
  assign n23735 = pi12 ? n32 : n23734;
  assign n23736 = pi15 ? n23574 : n23569;
  assign n23737 = pi14 ? n23736 : n23421;
  assign n23738 = pi19 ? n32 : n18424;
  assign n23739 = pi18 ? n32 : n23738;
  assign n23740 = pi17 ? n32 : n23739;
  assign n23741 = pi16 ? n32 : n23740;
  assign n23742 = pi15 ? n16108 : n23741;
  assign n23743 = pi15 ? n16108 : n15836;
  assign n23744 = pi14 ? n23742 : n23743;
  assign n23745 = pi13 ? n23737 : n23744;
  assign n23746 = pi19 ? n32 : ~n1941;
  assign n23747 = pi18 ? n32 : n23746;
  assign n23748 = pi17 ? n32 : n23747;
  assign n23749 = pi16 ? n32 : n23748;
  assign n23750 = pi15 ? n32 : n23749;
  assign n23751 = pi14 ? n23750 : n23749;
  assign n23752 = pi19 ? n23489 : ~n1941;
  assign n23753 = pi18 ? n32 : n23752;
  assign n23754 = pi17 ? n32 : n23753;
  assign n23755 = pi16 ? n32 : n23754;
  assign n23756 = pi15 ? n23755 : n15386;
  assign n23757 = pi14 ? n23756 : n15518;
  assign n23758 = pi13 ? n23751 : n23757;
  assign n23759 = pi12 ? n23745 : n23758;
  assign n23760 = pi11 ? n23735 : n23759;
  assign n23761 = pi15 ? n15518 : n15255;
  assign n23762 = pi14 ? n23761 : n23653;
  assign n23763 = pi13 ? n23762 : n23666;
  assign n23764 = pi20 ? n8943 : ~n206;
  assign n23765 = pi19 ? n23764 : n32;
  assign n23766 = pi18 ? n32 : n23765;
  assign n23767 = pi17 ? n32 : n23766;
  assign n23768 = pi16 ? n32 : n23767;
  assign n23769 = pi15 ? n23768 : n15389;
  assign n23770 = pi14 ? n23769 : n15389;
  assign n23771 = pi15 ? n15389 : n15123;
  assign n23772 = pi14 ? n23771 : n22635;
  assign n23773 = pi13 ? n23770 : n23772;
  assign n23774 = pi12 ? n23763 : n23773;
  assign n23775 = pi15 ? n23684 : n387;
  assign n23776 = pi14 ? n14974 : n23775;
  assign n23777 = pi14 ? n387 : n22009;
  assign n23778 = pi13 ? n23776 : n23777;
  assign n23779 = pi17 ? n32 : n17651;
  assign n23780 = pi16 ? n32 : n23779;
  assign n23781 = pi18 ? n32 : ~n805;
  assign n23782 = pi17 ? n23711 : n23781;
  assign n23783 = pi16 ? n32 : n23782;
  assign n23784 = pi15 ? n23780 : n23783;
  assign n23785 = pi14 ? n23558 : n23784;
  assign n23786 = pi13 ? n23705 : n23785;
  assign n23787 = pi12 ? n23778 : n23786;
  assign n23788 = pi11 ? n23774 : n23787;
  assign n23789 = pi10 ? n23760 : n23788;
  assign n23790 = pi09 ? n32 : n23789;
  assign n23791 = pi08 ? n23721 : n23790;
  assign n23792 = pi07 ? n23622 : n23791;
  assign n23793 = pi14 ? n23726 : n23725;
  assign n23794 = pi15 ? n23725 : n32;
  assign n23795 = pi14 ? n23794 : n32;
  assign n23796 = pi13 ? n23793 : n23795;
  assign n23797 = pi12 ? n32 : n23796;
  assign n23798 = pi14 ? n23794 : n23623;
  assign n23799 = pi19 ? n267 : n5614;
  assign n23800 = pi18 ? n32 : n23799;
  assign n23801 = pi17 ? n32 : n23800;
  assign n23802 = pi16 ? n32 : n23801;
  assign n23803 = pi15 ? n23574 : n23802;
  assign n23804 = pi14 ? n23574 : n23803;
  assign n23805 = pi13 ? n23798 : n23804;
  assign n23806 = pi20 ? n428 : ~n1385;
  assign n23807 = pi19 ? n23806 : ~n1941;
  assign n23808 = pi18 ? n32 : n23807;
  assign n23809 = pi17 ? n32 : n23808;
  assign n23810 = pi16 ? n32 : n23809;
  assign n23811 = pi15 ? n23749 : n23810;
  assign n23812 = pi14 ? n23749 : n23811;
  assign n23813 = pi20 ? n342 : ~n1385;
  assign n23814 = pi19 ? n23813 : ~n1941;
  assign n23815 = pi18 ? n32 : n23814;
  assign n23816 = pi17 ? n32 : n23815;
  assign n23817 = pi16 ? n32 : n23816;
  assign n23818 = pi20 ? n3523 : n11107;
  assign n23819 = pi19 ? n23818 : n5626;
  assign n23820 = pi18 ? n32 : n23819;
  assign n23821 = pi17 ? n32 : n23820;
  assign n23822 = pi16 ? n32 : n23821;
  assign n23823 = pi15 ? n23817 : n23822;
  assign n23824 = pi14 ? n23823 : n23160;
  assign n23825 = pi13 ? n23812 : n23824;
  assign n23826 = pi12 ? n23805 : n23825;
  assign n23827 = pi11 ? n23797 : n23826;
  assign n23828 = pi15 ? n23160 : n15518;
  assign n23829 = pi19 ? n3524 : ~n2614;
  assign n23830 = pi18 ? n32 : n23829;
  assign n23831 = pi17 ? n32 : n23830;
  assign n23832 = pi16 ? n32 : n23831;
  assign n23833 = pi19 ? n343 : ~n2614;
  assign n23834 = pi18 ? n32 : n23833;
  assign n23835 = pi17 ? n32 : n23834;
  assign n23836 = pi16 ? n32 : n23835;
  assign n23837 = pi15 ? n23832 : n23836;
  assign n23838 = pi14 ? n23828 : n23837;
  assign n23839 = pi19 ? n1757 : n2614;
  assign n23840 = pi18 ? n32 : ~n23839;
  assign n23841 = pi17 ? n32 : n23840;
  assign n23842 = pi16 ? n32 : n23841;
  assign n23843 = pi15 ? n23836 : n23842;
  assign n23844 = pi19 ? n1757 : n617;
  assign n23845 = pi18 ? n32 : ~n23844;
  assign n23846 = pi17 ? n32 : n23845;
  assign n23847 = pi16 ? n32 : n23846;
  assign n23848 = pi19 ? n247 : n1105;
  assign n23849 = pi18 ? n32 : ~n23848;
  assign n23850 = pi17 ? n32 : n23849;
  assign n23851 = pi16 ? n32 : n23850;
  assign n23852 = pi15 ? n23847 : n23851;
  assign n23853 = pi14 ? n23843 : n23852;
  assign n23854 = pi13 ? n23838 : n23853;
  assign n23855 = pi20 ? n32 : ~n20516;
  assign n23856 = pi19 ? n23855 : n32;
  assign n23857 = pi18 ? n32 : n23856;
  assign n23858 = pi17 ? n32 : n23857;
  assign n23859 = pi16 ? n32 : n23858;
  assign n23860 = pi15 ? n22347 : n23859;
  assign n23861 = pi14 ? n23179 : n23860;
  assign n23862 = pi13 ? n32 : n23861;
  assign n23863 = pi12 ? n23854 : n23862;
  assign n23864 = pi20 ? n32 : ~n19604;
  assign n23865 = pi19 ? n23864 : n32;
  assign n23866 = pi18 ? n32 : n23865;
  assign n23867 = pi17 ? n32 : n23866;
  assign n23868 = pi16 ? n32 : n23867;
  assign n23869 = pi15 ? n22437 : n23868;
  assign n23870 = pi14 ? n23869 : n21790;
  assign n23871 = pi19 ? n18041 : n32;
  assign n23872 = pi18 ? n32 : n23871;
  assign n23873 = pi17 ? n32 : n23872;
  assign n23874 = pi16 ? n32 : n23873;
  assign n23875 = pi19 ? n349 : ~n18478;
  assign n23876 = pi18 ? n23875 : n520;
  assign n23877 = pi17 ? n17463 : ~n23876;
  assign n23878 = pi16 ? n32 : n23877;
  assign n23879 = pi15 ? n23874 : n23878;
  assign n23880 = pi14 ? n32 : n23879;
  assign n23881 = pi13 ? n23870 : n23880;
  assign n23882 = pi19 ? n236 : ~n5688;
  assign n23883 = pi18 ? n23882 : n520;
  assign n23884 = pi17 ? n32 : ~n23883;
  assign n23885 = pi16 ? n32 : n23884;
  assign n23886 = pi15 ? n23885 : n13046;
  assign n23887 = pi18 ? n32 : ~n2754;
  assign n23888 = pi17 ? n32 : n23887;
  assign n23889 = pi16 ? n32 : n23888;
  assign n23890 = pi18 ? n32 : ~n323;
  assign n23891 = pi17 ? n32 : n23890;
  assign n23892 = pi16 ? n32 : n23891;
  assign n23893 = pi15 ? n23889 : n23892;
  assign n23894 = pi14 ? n23886 : n23893;
  assign n23895 = pi20 ? n266 : ~n321;
  assign n23896 = pi19 ? n5694 : ~n23895;
  assign n23897 = pi18 ? n20164 : n23896;
  assign n23898 = pi20 ? n206 : ~n1324;
  assign n23899 = pi19 ? n16431 : n23898;
  assign n23900 = pi18 ? n23899 : ~n2291;
  assign n23901 = pi17 ? n23897 : n23900;
  assign n23902 = pi16 ? n32 : n23901;
  assign n23903 = pi15 ? n23902 : n13369;
  assign n23904 = pi19 ? n267 : ~n15405;
  assign n23905 = pi18 ? n32 : n23904;
  assign n23906 = pi19 ? n9037 : n1757;
  assign n23907 = pi18 ? n23906 : n5005;
  assign n23908 = pi17 ? n23905 : n23907;
  assign n23909 = pi16 ? n32 : n23908;
  assign n23910 = pi20 ? n274 : ~n321;
  assign n23911 = pi19 ? n23910 : ~n1464;
  assign n23912 = pi18 ? n268 : n23911;
  assign n23913 = pi19 ? n16282 : n32;
  assign n23914 = pi18 ? n16432 : ~n23913;
  assign n23915 = pi17 ? n23912 : ~n23914;
  assign n23916 = pi16 ? n32 : n23915;
  assign n23917 = pi15 ? n23909 : n23916;
  assign n23918 = pi14 ? n23903 : n23917;
  assign n23919 = pi13 ? n23894 : n23918;
  assign n23920 = pi12 ? n23881 : n23919;
  assign n23921 = pi11 ? n23863 : n23920;
  assign n23922 = pi10 ? n23827 : n23921;
  assign n23923 = pi09 ? n32 : n23922;
  assign n23924 = pi15 ? n32 : n16319;
  assign n23925 = pi14 ? n23924 : n16319;
  assign n23926 = pi13 ? n23925 : n16322;
  assign n23927 = pi12 ? n32 : n23926;
  assign n23928 = pi14 ? n23725 : n23623;
  assign n23929 = pi13 ? n23928 : n23804;
  assign n23930 = pi19 ? n32 : ~n813;
  assign n23931 = pi18 ? n32 : n23930;
  assign n23932 = pi17 ? n32 : n23931;
  assign n23933 = pi16 ? n32 : n23932;
  assign n23934 = pi19 ? n23806 : ~n813;
  assign n23935 = pi18 ? n32 : n23934;
  assign n23936 = pi17 ? n32 : n23935;
  assign n23937 = pi16 ? n32 : n23936;
  assign n23938 = pi15 ? n23933 : n23937;
  assign n23939 = pi14 ? n23933 : n23938;
  assign n23940 = pi19 ? n23813 : ~n813;
  assign n23941 = pi18 ? n32 : n23940;
  assign n23942 = pi17 ? n32 : n23941;
  assign n23943 = pi16 ? n32 : n23942;
  assign n23944 = pi20 ? n32 : n11107;
  assign n23945 = pi19 ? n23944 : n358;
  assign n23946 = pi18 ? n32 : n23945;
  assign n23947 = pi17 ? n32 : n23946;
  assign n23948 = pi16 ? n32 : n23947;
  assign n23949 = pi15 ? n23943 : n23948;
  assign n23950 = pi14 ? n23949 : n23250;
  assign n23951 = pi13 ? n23939 : n23950;
  assign n23952 = pi12 ? n23929 : n23951;
  assign n23953 = pi11 ? n23927 : n23952;
  assign n23954 = pi14 ? n23485 : n23837;
  assign n23955 = pi13 ? n23954 : n23853;
  assign n23956 = pi13 ? n22540 : n23861;
  assign n23957 = pi12 ? n23955 : n23956;
  assign n23958 = pi14 ? n23869 : n21786;
  assign n23959 = pi14 ? n21786 : n23879;
  assign n23960 = pi13 ? n23958 : n23959;
  assign n23961 = pi15 ? n23902 : n21497;
  assign n23962 = pi18 ? n23906 : n21494;
  assign n23963 = pi17 ? n23905 : n23962;
  assign n23964 = pi16 ? n32 : n23963;
  assign n23965 = pi20 ? n749 : ~n1940;
  assign n23966 = pi19 ? n23965 : n32;
  assign n23967 = pi18 ? n16432 : ~n23966;
  assign n23968 = pi17 ? n23912 : ~n23967;
  assign n23969 = pi16 ? n32 : n23968;
  assign n23970 = pi15 ? n23964 : n23969;
  assign n23971 = pi14 ? n23961 : n23970;
  assign n23972 = pi13 ? n23894 : n23971;
  assign n23973 = pi12 ? n23960 : n23972;
  assign n23974 = pi11 ? n23957 : n23973;
  assign n23975 = pi10 ? n23953 : n23974;
  assign n23976 = pi09 ? n32 : n23975;
  assign n23977 = pi08 ? n23923 : n23976;
  assign n23978 = pi19 ? n32 : n5446;
  assign n23979 = pi18 ? n32 : n23978;
  assign n23980 = pi17 ? n32 : n23979;
  assign n23981 = pi16 ? n32 : n23980;
  assign n23982 = pi15 ? n32 : n23981;
  assign n23983 = pi14 ? n23982 : n16319;
  assign n23984 = pi13 ? n23983 : n32;
  assign n23985 = pi12 ? n32 : n23984;
  assign n23986 = pi14 ? n16105 : n23726;
  assign n23987 = pi15 ? n23725 : n14389;
  assign n23988 = pi14 ? n23725 : n23987;
  assign n23989 = pi13 ? n23986 : n23988;
  assign n23990 = pi19 ? n5694 : ~n813;
  assign n23991 = pi18 ? n32 : n23990;
  assign n23992 = pi17 ? n32 : n23991;
  assign n23993 = pi16 ? n32 : n23992;
  assign n23994 = pi15 ? n23933 : n23993;
  assign n23995 = pi14 ? n23933 : n23994;
  assign n23996 = pi19 ? n5694 : ~n1941;
  assign n23997 = pi18 ? n32 : n23996;
  assign n23998 = pi17 ? n32 : n23997;
  assign n23999 = pi16 ? n32 : n23998;
  assign n24000 = pi15 ? n23999 : n23484;
  assign n24001 = pi14 ? n24000 : n23485;
  assign n24002 = pi13 ? n23995 : n24001;
  assign n24003 = pi12 ? n23989 : n24002;
  assign n24004 = pi11 ? n23985 : n24003;
  assign n24005 = pi19 ? n462 : ~n236;
  assign n24006 = pi18 ? n32 : n24005;
  assign n24007 = pi17 ? n32 : n24006;
  assign n24008 = pi16 ? n32 : n24007;
  assign n24009 = pi15 ? n23250 : n24008;
  assign n24010 = pi20 ? n17665 : ~n32;
  assign n24011 = pi19 ? n24010 : ~n236;
  assign n24012 = pi18 ? n32 : n24011;
  assign n24013 = pi17 ? n32 : n24012;
  assign n24014 = pi16 ? n32 : n24013;
  assign n24015 = pi19 ? n343 : ~n236;
  assign n24016 = pi18 ? n32 : n24015;
  assign n24017 = pi17 ? n32 : n24016;
  assign n24018 = pi16 ? n32 : n24017;
  assign n24019 = pi15 ? n24014 : n24018;
  assign n24020 = pi14 ? n24009 : n24019;
  assign n24021 = pi15 ? n24018 : n23842;
  assign n24022 = pi15 ? n23847 : n22923;
  assign n24023 = pi14 ? n24021 : n24022;
  assign n24024 = pi13 ? n24020 : n24023;
  assign n24025 = pi19 ? n1508 : n32;
  assign n24026 = pi18 ? n32 : n24025;
  assign n24027 = pi17 ? n32 : n24026;
  assign n24028 = pi16 ? n32 : n24027;
  assign n24029 = pi15 ? n22817 : n24028;
  assign n24030 = pi14 ? n22817 : n24029;
  assign n24031 = pi13 ? n32 : n24030;
  assign n24032 = pi12 ? n24024 : n24031;
  assign n24033 = pi15 ? n23094 : n22434;
  assign n24034 = pi14 ? n24033 : n32;
  assign n24035 = pi20 ? n32 : n14490;
  assign n24036 = pi19 ? n24035 : ~n32;
  assign n24037 = pi18 ? n32 : ~n24036;
  assign n24038 = pi17 ? n32 : n24037;
  assign n24039 = pi16 ? n32 : n24038;
  assign n24040 = pi15 ? n24039 : n12767;
  assign n24041 = pi14 ? n32 : n24040;
  assign n24042 = pi13 ? n24034 : n24041;
  assign n24043 = pi20 ? n266 : n1319;
  assign n24044 = pi19 ? n24043 : ~n32;
  assign n24045 = pi18 ? n16603 : ~n24044;
  assign n24046 = pi17 ? n32 : n24045;
  assign n24047 = pi16 ? n32 : n24046;
  assign n24048 = pi15 ? n24047 : n13043;
  assign n24049 = pi18 ? n15844 : ~n520;
  assign n24050 = pi17 ? n32 : n24049;
  assign n24051 = pi16 ? n32 : n24050;
  assign n24052 = pi15 ? n24051 : n23889;
  assign n24053 = pi14 ? n24048 : n24052;
  assign n24054 = pi19 ? n32 : ~n6298;
  assign n24055 = pi20 ? n207 : n246;
  assign n24056 = pi19 ? n24055 : n266;
  assign n24057 = pi18 ? n24054 : ~n24056;
  assign n24058 = pi19 ? n16002 : n22185;
  assign n24059 = pi18 ? n24058 : ~n323;
  assign n24060 = pi17 ? n24057 : n24059;
  assign n24061 = pi16 ? n32 : n24060;
  assign n24062 = pi15 ? n24061 : n21497;
  assign n24063 = pi19 ? n32 : n18678;
  assign n24064 = pi19 ? n3692 : n1757;
  assign n24065 = pi18 ? n24063 : ~n24064;
  assign n24066 = pi19 ? n4670 : n221;
  assign n24067 = pi18 ? n24066 : n2413;
  assign n24068 = pi17 ? n24065 : ~n24067;
  assign n24069 = pi16 ? n32 : n24068;
  assign n24070 = pi19 ? n5730 : ~n5688;
  assign n24071 = pi18 ? n32 : n24070;
  assign n24072 = pi19 ? n342 : n16431;
  assign n24073 = pi18 ? n24072 : ~n13063;
  assign n24074 = pi17 ? n24071 : ~n24073;
  assign n24075 = pi16 ? n32 : n24074;
  assign n24076 = pi15 ? n24069 : n24075;
  assign n24077 = pi14 ? n24062 : n24076;
  assign n24078 = pi13 ? n24053 : n24077;
  assign n24079 = pi12 ? n24042 : n24078;
  assign n24080 = pi11 ? n24032 : n24079;
  assign n24081 = pi10 ? n24004 : n24080;
  assign n24082 = pi09 ? n32 : n24081;
  assign n24083 = pi14 ? n32 : n16314;
  assign n24084 = pi14 ? n16378 : n32;
  assign n24085 = pi13 ? n24083 : n24084;
  assign n24086 = pi12 ? n32 : n24085;
  assign n24087 = pi19 ? n221 : n6230;
  assign n24088 = pi18 ? n32 : n24087;
  assign n24089 = pi17 ? n32 : n24088;
  assign n24090 = pi16 ? n32 : n24089;
  assign n24091 = pi15 ? n23725 : n24090;
  assign n24092 = pi14 ? n23725 : n24091;
  assign n24093 = pi13 ? n23986 : n24092;
  assign n24094 = pi19 ? n32 : ~n1812;
  assign n24095 = pi18 ? n32 : n24094;
  assign n24096 = pi17 ? n32 : n24095;
  assign n24097 = pi16 ? n32 : n24096;
  assign n24098 = pi15 ? n24097 : n23993;
  assign n24099 = pi14 ? n24097 : n24098;
  assign n24100 = pi15 ? n23993 : n23749;
  assign n24101 = pi15 ? n23631 : n23749;
  assign n24102 = pi14 ? n24100 : n24101;
  assign n24103 = pi13 ? n24099 : n24102;
  assign n24104 = pi12 ? n24093 : n24103;
  assign n24105 = pi11 ? n24086 : n24104;
  assign n24106 = pi15 ? n23631 : n24008;
  assign n24107 = pi14 ? n24106 : n24019;
  assign n24108 = pi15 ? n23847 : n32;
  assign n24109 = pi14 ? n24021 : n24108;
  assign n24110 = pi13 ? n24107 : n24109;
  assign n24111 = pi20 ? n32 : ~n11782;
  assign n24112 = pi19 ? n24111 : n32;
  assign n24113 = pi18 ? n32 : n24112;
  assign n24114 = pi17 ? n32 : n24113;
  assign n24115 = pi16 ? n32 : n24114;
  assign n24116 = pi15 ? n22817 : n24115;
  assign n24117 = pi14 ? n22817 : n24116;
  assign n24118 = pi13 ? n22813 : n24117;
  assign n24119 = pi12 ? n24110 : n24118;
  assign n24120 = pi20 ? n32 : ~n8285;
  assign n24121 = pi19 ? n24120 : n32;
  assign n24122 = pi18 ? n32 : n24121;
  assign n24123 = pi17 ? n32 : n24122;
  assign n24124 = pi16 ? n32 : n24123;
  assign n24125 = pi15 ? n22437 : n24124;
  assign n24126 = pi14 ? n24125 : n21928;
  assign n24127 = pi14 ? n22133 : n24040;
  assign n24128 = pi13 ? n24126 : n24127;
  assign n24129 = pi15 ? n24047 : n13046;
  assign n24130 = pi18 ? n15844 : ~n2754;
  assign n24131 = pi17 ? n32 : n24130;
  assign n24132 = pi16 ? n32 : n24131;
  assign n24133 = pi15 ? n24132 : n23892;
  assign n24134 = pi14 ? n24129 : n24133;
  assign n24135 = pi18 ? n24058 : ~n2291;
  assign n24136 = pi17 ? n24057 : n24135;
  assign n24137 = pi16 ? n32 : n24136;
  assign n24138 = pi15 ? n24137 : n13360;
  assign n24139 = pi18 ? n24066 : n605;
  assign n24140 = pi17 ? n24065 : ~n24139;
  assign n24141 = pi16 ? n32 : n24140;
  assign n24142 = pi18 ? n24072 : ~n13070;
  assign n24143 = pi17 ? n24071 : ~n24142;
  assign n24144 = pi16 ? n32 : n24143;
  assign n24145 = pi15 ? n24141 : n24144;
  assign n24146 = pi14 ? n24138 : n24145;
  assign n24147 = pi13 ? n24134 : n24146;
  assign n24148 = pi12 ? n24128 : n24147;
  assign n24149 = pi11 ? n24119 : n24148;
  assign n24150 = pi10 ? n24105 : n24149;
  assign n24151 = pi09 ? n32 : n24150;
  assign n24152 = pi08 ? n24082 : n24151;
  assign n24153 = pi07 ? n23977 : n24152;
  assign n24154 = pi06 ? n23792 : n24153;
  assign n24155 = pi05 ? n23482 : n24154;
  assign n24156 = pi04 ? n22811 : n24155;
  assign n24157 = pi14 ? n32 : n16377;
  assign n24158 = pi13 ? n24157 : n24084;
  assign n24159 = pi12 ? n32 : n24158;
  assign n24160 = pi14 ? n16377 : n16105;
  assign n24161 = pi15 ? n16105 : n32;
  assign n24162 = pi14 ? n16105 : n24161;
  assign n24163 = pi13 ? n24160 : n24162;
  assign n24164 = pi19 ? n221 : ~n813;
  assign n24165 = pi18 ? n32 : n24164;
  assign n24166 = pi17 ? n32 : n24165;
  assign n24167 = pi16 ? n32 : n24166;
  assign n24168 = pi15 ? n24097 : n24167;
  assign n24169 = pi14 ? n24097 : n24168;
  assign n24170 = pi15 ? n23933 : n23749;
  assign n24171 = pi15 ? n23631 : n16108;
  assign n24172 = pi14 ? n24170 : n24171;
  assign n24173 = pi13 ? n24169 : n24172;
  assign n24174 = pi12 ? n24163 : n24173;
  assign n24175 = pi11 ? n24159 : n24174;
  assign n24176 = pi19 ? n531 : ~n1941;
  assign n24177 = pi18 ? n32 : n24176;
  assign n24178 = pi17 ? n32 : n24177;
  assign n24179 = pi16 ? n32 : n24178;
  assign n24180 = pi14 ? n24101 : n24179;
  assign n24181 = pi15 ? n24179 : n24018;
  assign n24182 = pi19 ? n4126 : ~n2614;
  assign n24183 = pi18 ? n32 : n24182;
  assign n24184 = pi17 ? n32 : n24183;
  assign n24185 = pi16 ? n32 : n24184;
  assign n24186 = pi15 ? n24185 : n32;
  assign n24187 = pi14 ? n24181 : n24186;
  assign n24188 = pi13 ? n24180 : n24187;
  assign n24189 = pi15 ? n23011 : n22817;
  assign n24190 = pi14 ? n23503 : n24189;
  assign n24191 = pi13 ? n32 : n24190;
  assign n24192 = pi12 ? n24188 : n24191;
  assign n24193 = pi15 ? n22347 : n15123;
  assign n24194 = pi14 ? n24193 : n32;
  assign n24195 = pi19 ? n20923 : n32;
  assign n24196 = pi18 ? n32 : n24195;
  assign n24197 = pi17 ? n32 : n24196;
  assign n24198 = pi16 ? n32 : n24197;
  assign n24199 = pi15 ? n32 : n24198;
  assign n24200 = pi15 ? n13040 : n13338;
  assign n24201 = pi14 ? n24199 : n24200;
  assign n24202 = pi13 ? n24194 : n24201;
  assign n24203 = pi15 ? n13338 : n13344;
  assign n24204 = pi20 ? n32 : n10889;
  assign n24205 = pi19 ? n24204 : ~n32;
  assign n24206 = pi18 ? n32 : ~n24205;
  assign n24207 = pi17 ? n32 : n24206;
  assign n24208 = pi16 ? n32 : n24207;
  assign n24209 = pi20 ? n342 : ~n1839;
  assign n24210 = pi19 ? n24209 : n32;
  assign n24211 = pi18 ? n32 : n24210;
  assign n24212 = pi17 ? n32 : n24211;
  assign n24213 = pi16 ? n32 : n24212;
  assign n24214 = pi15 ? n24208 : n24213;
  assign n24215 = pi14 ? n24203 : n24214;
  assign n24216 = pi17 ? n1470 : ~n2519;
  assign n24217 = pi16 ? n32 : n24216;
  assign n24218 = pi20 ? n266 : n749;
  assign n24219 = pi19 ? n24218 : ~n32;
  assign n24220 = pi18 ? n32 : ~n24219;
  assign n24221 = pi17 ? n32 : n24220;
  assign n24222 = pi16 ? n32 : n24221;
  assign n24223 = pi15 ? n24217 : n24222;
  assign n24224 = pi19 ? n321 : ~n9007;
  assign n24225 = pi18 ? n268 : n24224;
  assign n24226 = pi18 ? n247 : ~n13058;
  assign n24227 = pi17 ? n24225 : ~n24226;
  assign n24228 = pi16 ? n32 : n24227;
  assign n24229 = pi15 ? n24228 : n13360;
  assign n24230 = pi14 ? n24223 : n24229;
  assign n24231 = pi13 ? n24215 : n24230;
  assign n24232 = pi12 ? n24202 : n24231;
  assign n24233 = pi11 ? n24192 : n24232;
  assign n24234 = pi10 ? n24175 : n24233;
  assign n24235 = pi09 ? n32 : n24234;
  assign n24236 = pi17 ? n32 : n3497;
  assign n24237 = pi16 ? n32 : n24236;
  assign n24238 = pi14 ? n32 : n24237;
  assign n24239 = pi15 ? n24237 : n32;
  assign n24240 = pi14 ? n24239 : n32;
  assign n24241 = pi13 ? n24238 : n24240;
  assign n24242 = pi12 ? n32 : n24241;
  assign n24243 = pi15 ? n16105 : n16319;
  assign n24244 = pi14 ? n16105 : n24243;
  assign n24245 = pi13 ? n24160 : n24244;
  assign n24246 = pi17 ? n32 : n20165;
  assign n24247 = pi16 ? n32 : n24246;
  assign n24248 = pi19 ? n221 : ~n1812;
  assign n24249 = pi18 ? n32 : n24248;
  assign n24250 = pi17 ? n32 : n24249;
  assign n24251 = pi16 ? n32 : n24250;
  assign n24252 = pi15 ? n24247 : n24251;
  assign n24253 = pi14 ? n24247 : n24252;
  assign n24254 = pi18 ? n32 : n20380;
  assign n24255 = pi17 ? n32 : n24254;
  assign n24256 = pi16 ? n32 : n24255;
  assign n24257 = pi15 ? n24256 : n23574;
  assign n24258 = pi14 ? n23933 : n24257;
  assign n24259 = pi13 ? n24253 : n24258;
  assign n24260 = pi12 ? n24245 : n24259;
  assign n24261 = pi11 ? n24242 : n24260;
  assign n24262 = pi15 ? n24256 : n23484;
  assign n24263 = pi14 ? n24262 : n24179;
  assign n24264 = pi19 ? n23944 : ~n2614;
  assign n24265 = pi18 ? n32 : n24264;
  assign n24266 = pi17 ? n32 : n24265;
  assign n24267 = pi16 ? n32 : n24266;
  assign n24268 = pi15 ? n24267 : n32;
  assign n24269 = pi14 ? n24181 : n24268;
  assign n24270 = pi13 ? n24263 : n24269;
  assign n24271 = pi19 ? n32 : n5635;
  assign n24272 = pi18 ? n32 : n24271;
  assign n24273 = pi17 ? n32 : n24272;
  assign n24274 = pi16 ? n32 : n24273;
  assign n24275 = pi15 ? n22923 : n24274;
  assign n24276 = pi14 ? n24275 : n22925;
  assign n24277 = pi13 ? n24276 : n24190;
  assign n24278 = pi12 ? n24270 : n24277;
  assign n24279 = pi14 ? n24193 : n648;
  assign n24280 = pi13 ? n24279 : n24201;
  assign n24281 = pi12 ? n24280 : n24231;
  assign n24282 = pi11 ? n24278 : n24281;
  assign n24283 = pi10 ? n24261 : n24282;
  assign n24284 = pi09 ? n32 : n24283;
  assign n24285 = pi08 ? n24235 : n24284;
  assign n24286 = pi19 ? n32 : n7693;
  assign n24287 = pi18 ? n32 : n24286;
  assign n24288 = pi17 ? n32 : n24287;
  assign n24289 = pi16 ? n32 : n24288;
  assign n24290 = pi15 ? n24289 : n16377;
  assign n24291 = pi14 ? n24237 : n24290;
  assign n24292 = pi15 ? n16377 : n16105;
  assign n24293 = pi14 ? n16377 : n24292;
  assign n24294 = pi13 ? n24291 : n24293;
  assign n24295 = pi15 ? n24247 : n24097;
  assign n24296 = pi14 ? n24247 : n24295;
  assign n24297 = pi14 ? n23933 : n23574;
  assign n24298 = pi13 ? n24296 : n24297;
  assign n24299 = pi12 ? n24294 : n24298;
  assign n24300 = pi11 ? n24242 : n24299;
  assign n24301 = pi19 ? n1464 : ~n813;
  assign n24302 = pi18 ? n32 : n24301;
  assign n24303 = pi17 ? n32 : n24302;
  assign n24304 = pi16 ? n32 : n24303;
  assign n24305 = pi15 ? n23574 : n24304;
  assign n24306 = pi19 ? n1464 : n1757;
  assign n24307 = pi18 ? n24306 : n14567;
  assign n24308 = pi17 ? n32 : n24307;
  assign n24309 = pi16 ? n32 : n24308;
  assign n24310 = pi19 ? n349 : ~n813;
  assign n24311 = pi18 ? n32 : n24310;
  assign n24312 = pi17 ? n32 : n24311;
  assign n24313 = pi16 ? n32 : n24312;
  assign n24314 = pi15 ? n24309 : n24313;
  assign n24315 = pi14 ? n24305 : n24314;
  assign n24316 = pi19 ? n343 : ~n813;
  assign n24317 = pi18 ? n32 : n24316;
  assign n24318 = pi17 ? n32 : n24317;
  assign n24319 = pi16 ? n32 : n24318;
  assign n24320 = pi19 ? n3507 : ~n1941;
  assign n24321 = pi18 ? n32 : n24320;
  assign n24322 = pi17 ? n32 : n24321;
  assign n24323 = pi16 ? n32 : n24322;
  assign n24324 = pi15 ? n24319 : n24323;
  assign n24325 = pi14 ? n24324 : n23252;
  assign n24326 = pi13 ? n24315 : n24325;
  assign n24327 = pi15 ? n32 : n22923;
  assign n24328 = pi14 ? n32 : n24327;
  assign n24329 = pi15 ? n15119 : n23011;
  assign n24330 = pi14 ? n23593 : n24329;
  assign n24331 = pi13 ? n24328 : n24330;
  assign n24332 = pi12 ? n24326 : n24331;
  assign n24333 = pi14 ? n22829 : n32;
  assign n24334 = pi15 ? n32 : n13910;
  assign n24335 = pi15 ? n23189 : n22755;
  assign n24336 = pi14 ? n24334 : n24335;
  assign n24337 = pi13 ? n24333 : n24336;
  assign n24338 = pi15 ? n13338 : n13913;
  assign n24339 = pi15 ? n13043 : n13920;
  assign n24340 = pi14 ? n24338 : n24339;
  assign n24341 = pi17 ? n1470 : ~n2755;
  assign n24342 = pi16 ? n32 : n24341;
  assign n24343 = pi20 ? n220 : ~n266;
  assign n24344 = pi19 ? n24343 : ~n32;
  assign n24345 = pi18 ? n32 : n24344;
  assign n24346 = pi17 ? n24345 : ~n2408;
  assign n24347 = pi16 ? n32 : n24346;
  assign n24348 = pi15 ? n24342 : n24347;
  assign n24349 = pi20 ? n206 : n207;
  assign n24350 = pi19 ? n18678 : n24349;
  assign n24351 = pi18 ? n32 : n24350;
  assign n24352 = pi19 ? n3692 : ~n8818;
  assign n24353 = pi20 ? n357 : n749;
  assign n24354 = pi19 ? n24353 : ~n32;
  assign n24355 = pi18 ? n24352 : n24354;
  assign n24356 = pi17 ? n24351 : ~n24355;
  assign n24357 = pi16 ? n32 : n24356;
  assign n24358 = pi15 ? n24357 : n13360;
  assign n24359 = pi14 ? n24348 : n24358;
  assign n24360 = pi13 ? n24340 : n24359;
  assign n24361 = pi12 ? n24337 : n24360;
  assign n24362 = pi11 ? n24332 : n24361;
  assign n24363 = pi10 ? n24300 : n24362;
  assign n24364 = pi09 ? n32 : n24363;
  assign n24365 = pi18 ? n32 : n5267;
  assign n24366 = pi17 ? n32 : n24365;
  assign n24367 = pi16 ? n32 : n24366;
  assign n24368 = pi15 ? n32 : n24367;
  assign n24369 = pi14 ? n24368 : n24367;
  assign n24370 = pi15 ? n24367 : n32;
  assign n24371 = pi14 ? n24370 : n32;
  assign n24372 = pi13 ? n24369 : n24371;
  assign n24373 = pi12 ? n32 : n24372;
  assign n24374 = pi15 ? n16105 : n16377;
  assign n24375 = pi14 ? n24239 : n24374;
  assign n24376 = pi15 ? n16377 : n24289;
  assign n24377 = pi14 ? n16377 : n24376;
  assign n24378 = pi13 ? n24375 : n24377;
  assign n24379 = pi19 ? n32 : ~n2848;
  assign n24380 = pi18 ? n32 : n24379;
  assign n24381 = pi17 ? n32 : n24380;
  assign n24382 = pi16 ? n32 : n24381;
  assign n24383 = pi15 ? n24382 : n24247;
  assign n24384 = pi14 ? n24382 : n24383;
  assign n24385 = pi19 ? n32 : ~n20022;
  assign n24386 = pi18 ? n32 : n24385;
  assign n24387 = pi17 ? n32 : n24386;
  assign n24388 = pi16 ? n32 : n24387;
  assign n24389 = pi15 ? n24097 : n24388;
  assign n24390 = pi15 ? n23730 : n23725;
  assign n24391 = pi14 ? n24389 : n24390;
  assign n24392 = pi13 ? n24384 : n24391;
  assign n24393 = pi12 ? n24378 : n24392;
  assign n24394 = pi11 ? n24373 : n24393;
  assign n24395 = pi15 ? n23730 : n24304;
  assign n24396 = pi14 ? n24395 : n24314;
  assign n24397 = pi15 ? n23250 : n23160;
  assign n24398 = pi14 ? n24324 : n24397;
  assign n24399 = pi13 ? n24396 : n24398;
  assign n24400 = pi14 ? n23160 : n24327;
  assign n24401 = pi13 ? n24400 : n24330;
  assign n24402 = pi12 ? n24399 : n24401;
  assign n24403 = pi19 ? n19370 : n32;
  assign n24404 = pi18 ? n32 : n24403;
  assign n24405 = pi17 ? n32 : n24404;
  assign n24406 = pi16 ? n32 : n24405;
  assign n24407 = pi15 ? n22817 : n24406;
  assign n24408 = pi14 ? n24407 : n32;
  assign n24409 = pi13 ? n24408 : n24336;
  assign n24410 = pi17 ? n24345 : ~n2292;
  assign n24411 = pi16 ? n32 : n24410;
  assign n24412 = pi15 ? n24342 : n24411;
  assign n24413 = pi20 ? n357 : n1475;
  assign n24414 = pi19 ? n24413 : ~n32;
  assign n24415 = pi18 ? n24352 : n24414;
  assign n24416 = pi17 ? n24351 : ~n24415;
  assign n24417 = pi16 ? n32 : n24416;
  assign n24418 = pi18 ? n32 : n21818;
  assign n24419 = pi17 ? n32 : n24418;
  assign n24420 = pi16 ? n32 : n24419;
  assign n24421 = pi15 ? n24417 : n24420;
  assign n24422 = pi14 ? n24412 : n24421;
  assign n24423 = pi13 ? n24340 : n24422;
  assign n24424 = pi12 ? n24409 : n24423;
  assign n24425 = pi11 ? n24402 : n24424;
  assign n24426 = pi10 ? n24394 : n24425;
  assign n24427 = pi09 ? n32 : n24426;
  assign n24428 = pi08 ? n24364 : n24427;
  assign n24429 = pi07 ? n24285 : n24428;
  assign n24430 = pi15 ? n24367 : n24237;
  assign n24431 = pi14 ? n24430 : n24237;
  assign n24432 = pi15 ? n24237 : n24289;
  assign n24433 = pi14 ? n24237 : n24432;
  assign n24434 = pi13 ? n24431 : n24433;
  assign n24435 = pi15 ? n24382 : n16105;
  assign n24436 = pi14 ? n24382 : n24435;
  assign n24437 = pi13 ? n24436 : n23793;
  assign n24438 = pi12 ? n24434 : n24437;
  assign n24439 = pi11 ? n24373 : n24438;
  assign n24440 = pi19 ? n208 : ~n1812;
  assign n24441 = pi18 ? n32 : n24440;
  assign n24442 = pi17 ? n32 : n24441;
  assign n24443 = pi16 ? n32 : n24442;
  assign n24444 = pi15 ? n23725 : n24443;
  assign n24445 = pi19 ? n422 : ~n1812;
  assign n24446 = pi18 ? n16449 : n24445;
  assign n24447 = pi17 ? n32 : n24446;
  assign n24448 = pi16 ? n32 : n24447;
  assign n24449 = pi18 ? n32 : n24445;
  assign n24450 = pi17 ? n32 : n24449;
  assign n24451 = pi16 ? n32 : n24450;
  assign n24452 = pi15 ? n24448 : n24451;
  assign n24453 = pi14 ? n24444 : n24452;
  assign n24454 = pi19 ? n1818 : n15923;
  assign n24455 = pi18 ? n24454 : n24440;
  assign n24456 = pi17 ? n32 : n24455;
  assign n24457 = pi16 ? n32 : n24456;
  assign n24458 = pi15 ? n24457 : n23631;
  assign n24459 = pi14 ? n24458 : n23252;
  assign n24460 = pi13 ? n24453 : n24459;
  assign n24461 = pi14 ? n32 : n23828;
  assign n24462 = pi15 ? n15119 : n22728;
  assign n24463 = pi14 ? n23761 : n24462;
  assign n24464 = pi13 ? n24461 : n24463;
  assign n24465 = pi12 ? n24460 : n24464;
  assign n24466 = pi15 ? n14389 : n24124;
  assign n24467 = pi15 ? n13910 : n14143;
  assign n24468 = pi14 ? n24466 : n24467;
  assign n24469 = pi13 ? n24333 : n24468;
  assign n24470 = pi15 ? n13626 : n14147;
  assign n24471 = pi20 ? n321 : n1319;
  assign n24472 = pi19 ? n24471 : ~n32;
  assign n24473 = pi18 ? n32 : ~n24472;
  assign n24474 = pi17 ? n32 : n24473;
  assign n24475 = pi16 ? n32 : n24474;
  assign n24476 = pi19 ? n8196 : ~n32;
  assign n24477 = pi18 ? n32 : ~n24476;
  assign n24478 = pi17 ? n32 : n24477;
  assign n24479 = pi16 ? n32 : n24478;
  assign n24480 = pi15 ? n24475 : n24479;
  assign n24481 = pi14 ? n24470 : n24480;
  assign n24482 = pi17 ? n1470 : ~n2408;
  assign n24483 = pi16 ? n32 : n24482;
  assign n24484 = pi15 ? n24217 : n24483;
  assign n24485 = pi15 ? n14164 : n21551;
  assign n24486 = pi14 ? n24484 : n24485;
  assign n24487 = pi13 ? n24481 : n24486;
  assign n24488 = pi12 ? n24469 : n24487;
  assign n24489 = pi11 ? n24465 : n24488;
  assign n24490 = pi10 ? n24439 : n24489;
  assign n24491 = pi09 ? n32 : n24490;
  assign n24492 = pi19 ? n32 : n152;
  assign n24493 = pi18 ? n32 : n24492;
  assign n24494 = pi17 ? n32 : n24493;
  assign n24495 = pi16 ? n32 : n24494;
  assign n24496 = pi15 ? n32 : n24495;
  assign n24497 = pi14 ? n24496 : n16606;
  assign n24498 = pi15 ? n16606 : n32;
  assign n24499 = pi14 ? n24498 : n32;
  assign n24500 = pi13 ? n24497 : n24499;
  assign n24501 = pi12 ? n32 : n24500;
  assign n24502 = pi18 ? n32 : n21287;
  assign n24503 = pi17 ? n32 : n24502;
  assign n24504 = pi16 ? n32 : n24503;
  assign n24505 = pi15 ? n24237 : n24504;
  assign n24506 = pi14 ? n24237 : n24505;
  assign n24507 = pi13 ? n24431 : n24506;
  assign n24508 = pi19 ? n32 : ~n589;
  assign n24509 = pi18 ? n32 : n24508;
  assign n24510 = pi17 ? n32 : n24509;
  assign n24511 = pi16 ? n32 : n24510;
  assign n24512 = pi15 ? n24511 : n24289;
  assign n24513 = pi14 ? n24511 : n24512;
  assign n24514 = pi15 ? n16319 : n23981;
  assign n24515 = pi14 ? n24514 : n16319;
  assign n24516 = pi13 ? n24513 : n24515;
  assign n24517 = pi12 ? n24507 : n24516;
  assign n24518 = pi11 ? n24501 : n24517;
  assign n24519 = pi15 ? n32 : n24443;
  assign n24520 = pi14 ? n24519 : n24452;
  assign n24521 = pi15 ? n24457 : n24256;
  assign n24522 = pi15 ? n23741 : n15836;
  assign n24523 = pi14 ? n24521 : n24522;
  assign n24524 = pi13 ? n24520 : n24523;
  assign n24525 = pi19 ? n1574 : ~n617;
  assign n24526 = pi18 ? n32 : n24525;
  assign n24527 = pi17 ? n32 : n24526;
  assign n24528 = pi16 ? n32 : n24527;
  assign n24529 = pi15 ? n15119 : n24528;
  assign n24530 = pi14 ? n23761 : n24529;
  assign n24531 = pi13 ? n23161 : n24530;
  assign n24532 = pi12 ? n24524 : n24531;
  assign n24533 = pi15 ? n22728 : n22540;
  assign n24534 = pi14 ? n24533 : n32;
  assign n24535 = pi15 ? n14593 : n22434;
  assign n24536 = pi19 ? n12578 : n32;
  assign n24537 = pi18 ? n32 : n24536;
  assign n24538 = pi17 ? n32 : n24537;
  assign n24539 = pi16 ? n32 : n24538;
  assign n24540 = pi19 ? n17918 : n32;
  assign n24541 = pi18 ? n32 : n24540;
  assign n24542 = pi17 ? n32 : n24541;
  assign n24543 = pi16 ? n32 : n24542;
  assign n24544 = pi15 ? n24539 : n24543;
  assign n24545 = pi14 ? n24535 : n24544;
  assign n24546 = pi13 ? n24534 : n24545;
  assign n24547 = pi15 ? n13626 : n14143;
  assign n24548 = pi19 ? n9822 : ~n32;
  assign n24549 = pi18 ? n32 : ~n24548;
  assign n24550 = pi17 ? n32 : n24549;
  assign n24551 = pi16 ? n32 : n24550;
  assign n24552 = pi15 ? n24551 : n24479;
  assign n24553 = pi14 ? n24547 : n24552;
  assign n24554 = pi15 ? n24342 : n24217;
  assign n24555 = pi15 ? n14397 : n14156;
  assign n24556 = pi14 ? n24554 : n24555;
  assign n24557 = pi13 ? n24553 : n24556;
  assign n24558 = pi12 ? n24546 : n24557;
  assign n24559 = pi11 ? n24532 : n24558;
  assign n24560 = pi10 ? n24518 : n24559;
  assign n24561 = pi09 ? n32 : n24560;
  assign n24562 = pi08 ? n24491 : n24561;
  assign n24563 = pi15 ? n32 : n16606;
  assign n24564 = pi14 ? n24563 : n16606;
  assign n24565 = pi13 ? n24564 : n24499;
  assign n24566 = pi12 ? n32 : n24565;
  assign n24567 = pi15 ? n16452 : n24367;
  assign n24568 = pi14 ? n24567 : n24367;
  assign n24569 = pi19 ? n32 : n19317;
  assign n24570 = pi18 ? n32 : n24569;
  assign n24571 = pi17 ? n32 : n24570;
  assign n24572 = pi16 ? n32 : n24571;
  assign n24573 = pi15 ? n24572 : n24237;
  assign n24574 = pi14 ? n24367 : n24573;
  assign n24575 = pi13 ? n24568 : n24574;
  assign n24576 = pi15 ? n24511 : n16377;
  assign n24577 = pi14 ? n24511 : n24576;
  assign n24578 = pi15 ? n16319 : n16105;
  assign n24579 = pi19 ? n507 : n1757;
  assign n24580 = pi18 ? n32 : n24579;
  assign n24581 = pi17 ? n32 : n24580;
  assign n24582 = pi16 ? n32 : n24581;
  assign n24583 = pi15 ? n16105 : n24582;
  assign n24584 = pi14 ? n24578 : n24583;
  assign n24585 = pi13 ? n24577 : n24584;
  assign n24586 = pi12 ? n24575 : n24585;
  assign n24587 = pi11 ? n24566 : n24586;
  assign n24588 = pi19 ? n804 : ~n349;
  assign n24589 = pi18 ? n16389 : n24588;
  assign n24590 = pi17 ? n32 : n24589;
  assign n24591 = pi16 ? n32 : n24590;
  assign n24592 = pi15 ? n16105 : n24591;
  assign n24593 = pi18 ? n15844 : n24588;
  assign n24594 = pi17 ? n32 : n24593;
  assign n24595 = pi16 ? n32 : n24594;
  assign n24596 = pi15 ? n24595 : n12556;
  assign n24597 = pi14 ? n24592 : n24596;
  assign n24598 = pi20 ? n17669 : n266;
  assign n24599 = pi19 ? n857 : n24598;
  assign n24600 = pi20 ? n428 : n206;
  assign n24601 = pi19 ? n24600 : n7488;
  assign n24602 = pi18 ? n24599 : n24601;
  assign n24603 = pi17 ? n32 : n24602;
  assign n24604 = pi16 ? n32 : n24603;
  assign n24605 = pi15 ? n24604 : n24256;
  assign n24606 = pi14 ? n24605 : n23632;
  assign n24607 = pi13 ? n24597 : n24606;
  assign n24608 = pi14 ? n32 : n23582;
  assign n24609 = pi19 ? n322 : ~n2614;
  assign n24610 = pi18 ? n32 : n24609;
  assign n24611 = pi17 ? n32 : n24610;
  assign n24612 = pi16 ? n32 : n24611;
  assign n24613 = pi15 ? n15518 : n24612;
  assign n24614 = pi15 ? n15255 : n23340;
  assign n24615 = pi14 ? n24613 : n24614;
  assign n24616 = pi13 ? n24608 : n24615;
  assign n24617 = pi12 ? n24607 : n24616;
  assign n24618 = pi14 ? n23113 : n24543;
  assign n24619 = pi13 ? n24534 : n24618;
  assign n24620 = pi14 ? n14143 : n24552;
  assign n24621 = pi14 ? n24554 : n14397;
  assign n24622 = pi13 ? n24620 : n24621;
  assign n24623 = pi12 ? n24619 : n24622;
  assign n24624 = pi11 ? n24617 : n24623;
  assign n24625 = pi10 ? n24587 : n24624;
  assign n24626 = pi09 ? n32 : n24625;
  assign n24627 = pi15 ? n32 : n16786;
  assign n24628 = pi14 ? n24627 : n16601;
  assign n24629 = pi15 ? n16601 : n32;
  assign n24630 = pi14 ? n24629 : n32;
  assign n24631 = pi13 ? n24628 : n24630;
  assign n24632 = pi12 ? n32 : n24631;
  assign n24633 = pi15 ? n16452 : n32;
  assign n24634 = pi14 ? n24633 : n24368;
  assign n24635 = pi14 ? n24367 : n24572;
  assign n24636 = pi13 ? n24634 : n24635;
  assign n24637 = pi19 ? n32 : ~n2317;
  assign n24638 = pi18 ? n32 : n24637;
  assign n24639 = pi17 ? n32 : n24638;
  assign n24640 = pi16 ? n32 : n24639;
  assign n24641 = pi15 ? n24640 : n24237;
  assign n24642 = pi14 ? n24640 : n24641;
  assign n24643 = pi14 ? n24376 : n24583;
  assign n24644 = pi13 ? n24642 : n24643;
  assign n24645 = pi12 ? n24636 : n24644;
  assign n24646 = pi11 ? n24632 : n24645;
  assign n24647 = pi19 ? n32 : n18728;
  assign n24648 = pi20 ? n14400 : n32;
  assign n24649 = pi19 ? n24600 : n24648;
  assign n24650 = pi18 ? n24647 : n24649;
  assign n24651 = pi17 ? n32 : n24650;
  assign n24652 = pi16 ? n32 : n24651;
  assign n24653 = pi15 ? n24652 : n23730;
  assign n24654 = pi15 ? n23574 : n16108;
  assign n24655 = pi14 ? n24653 : n24654;
  assign n24656 = pi13 ? n24597 : n24655;
  assign n24657 = pi18 ? n32 : n6645;
  assign n24658 = pi17 ? n32 : n24657;
  assign n24659 = pi16 ? n32 : n24658;
  assign n24660 = pi15 ? n23484 : n24659;
  assign n24661 = pi15 ? n15255 : n15386;
  assign n24662 = pi14 ? n24660 : n24661;
  assign n24663 = pi13 ? n23251 : n24662;
  assign n24664 = pi12 ? n24656 : n24663;
  assign n24665 = pi15 ? n23340 : n22540;
  assign n24666 = pi14 ? n24665 : n22424;
  assign n24667 = pi19 ? n18031 : n32;
  assign n24668 = pi18 ? n32 : n24667;
  assign n24669 = pi17 ? n32 : n24668;
  assign n24670 = pi16 ? n32 : n24669;
  assign n24671 = pi15 ? n24670 : n23094;
  assign n24672 = pi15 ? n22633 : n24543;
  assign n24673 = pi14 ? n24671 : n24672;
  assign n24674 = pi13 ? n24666 : n24673;
  assign n24675 = pi15 ? n24543 : n14143;
  assign n24676 = pi15 ? n24551 : n24475;
  assign n24677 = pi14 ? n24675 : n24676;
  assign n24678 = pi17 ? n1470 : ~n2517;
  assign n24679 = pi16 ? n32 : n24678;
  assign n24680 = pi15 ? n24679 : n24342;
  assign n24681 = pi14 ? n24680 : n21697;
  assign n24682 = pi13 ? n24677 : n24681;
  assign n24683 = pi12 ? n24674 : n24682;
  assign n24684 = pi11 ? n24664 : n24683;
  assign n24685 = pi10 ? n24646 : n24684;
  assign n24686 = pi09 ? n32 : n24685;
  assign n24687 = pi08 ? n24626 : n24686;
  assign n24688 = pi07 ? n24562 : n24687;
  assign n24689 = pi06 ? n24429 : n24688;
  assign n24690 = pi14 ? n24627 : n16786;
  assign n24691 = pi15 ? n32 : n16452;
  assign n24692 = pi14 ? n16840 : n24691;
  assign n24693 = pi13 ? n24690 : n24692;
  assign n24694 = pi12 ? n32 : n24693;
  assign n24695 = pi15 ? n16520 : n16606;
  assign n24696 = pi14 ? n24695 : n16606;
  assign n24697 = pi19 ? n32 : ~n343;
  assign n24698 = pi18 ? n32 : n24697;
  assign n24699 = pi17 ? n32 : n24698;
  assign n24700 = pi16 ? n32 : n24699;
  assign n24701 = pi15 ? n16606 : n24700;
  assign n24702 = pi19 ? n507 : ~n2317;
  assign n24703 = pi18 ? n32 : n24702;
  assign n24704 = pi17 ? n32 : n24703;
  assign n24705 = pi16 ? n32 : n24704;
  assign n24706 = pi15 ? n24640 : n24705;
  assign n24707 = pi14 ? n24701 : n24706;
  assign n24708 = pi13 ? n24696 : n24707;
  assign n24709 = pi19 ? n32 : n7468;
  assign n24710 = pi18 ? n32 : n24709;
  assign n24711 = pi17 ? n32 : n24710;
  assign n24712 = pi16 ? n32 : n24711;
  assign n24713 = pi15 ? n24640 : n24712;
  assign n24714 = pi14 ? n24713 : n24573;
  assign n24715 = pi19 ? n32 : ~n7014;
  assign n24716 = pi18 ? n32 : n24715;
  assign n24717 = pi17 ? n32 : n24716;
  assign n24718 = pi16 ? n32 : n24717;
  assign n24719 = pi15 ? n24247 : n16105;
  assign n24720 = pi14 ? n24718 : n24719;
  assign n24721 = pi13 ? n24714 : n24720;
  assign n24722 = pi12 ? n24708 : n24721;
  assign n24723 = pi11 ? n24694 : n24722;
  assign n24724 = pi18 ? n22865 : n6669;
  assign n24725 = pi17 ? n32 : n24724;
  assign n24726 = pi16 ? n32 : n24725;
  assign n24727 = pi15 ? n24247 : n24726;
  assign n24728 = pi18 ? n16389 : n6669;
  assign n24729 = pi17 ? n32 : n24728;
  assign n24730 = pi16 ? n32 : n24729;
  assign n24731 = pi19 ? n1248 : ~n349;
  assign n24732 = pi18 ? n32 : n24731;
  assign n24733 = pi17 ? n32 : n24732;
  assign n24734 = pi16 ? n32 : n24733;
  assign n24735 = pi15 ? n24730 : n24734;
  assign n24736 = pi14 ? n24727 : n24735;
  assign n24737 = pi15 ? n16105 : n23730;
  assign n24738 = pi14 ? n24737 : n24654;
  assign n24739 = pi13 ? n24736 : n24738;
  assign n24740 = pi14 ? n32 : n23484;
  assign n24741 = pi17 ? n32 : n20011;
  assign n24742 = pi16 ? n32 : n24741;
  assign n24743 = pi15 ? n24742 : n23484;
  assign n24744 = pi14 ? n24743 : n15518;
  assign n24745 = pi13 ? n24740 : n24744;
  assign n24746 = pi12 ? n24739 : n24745;
  assign n24747 = pi15 ? n15119 : n22817;
  assign n24748 = pi15 ? n32 : n23094;
  assign n24749 = pi14 ? n24747 : n24748;
  assign n24750 = pi20 ? n342 : ~n101;
  assign n24751 = pi19 ? n24750 : n32;
  assign n24752 = pi18 ? n16603 : n24751;
  assign n24753 = pi17 ? n32 : n24752;
  assign n24754 = pi16 ? n32 : n24753;
  assign n24755 = pi20 ? n246 : n310;
  assign n24756 = pi19 ? n32 : n24755;
  assign n24757 = pi18 ? n24756 : n24540;
  assign n24758 = pi17 ? n32 : n24757;
  assign n24759 = pi16 ? n32 : n24758;
  assign n24760 = pi15 ? n24754 : n24759;
  assign n24761 = pi14 ? n23094 : n24760;
  assign n24762 = pi13 ? n24749 : n24761;
  assign n24763 = pi20 ? n266 : ~n428;
  assign n24764 = pi19 ? n24763 : n32;
  assign n24765 = pi18 ? n16098 : n24764;
  assign n24766 = pi17 ? n32 : n24765;
  assign n24767 = pi16 ? n32 : n24766;
  assign n24768 = pi18 ? n14982 : n22846;
  assign n24769 = pi17 ? n32 : n24768;
  assign n24770 = pi16 ? n32 : n24769;
  assign n24771 = pi15 ? n24767 : n24770;
  assign n24772 = pi18 ? n14153 : n4983;
  assign n24773 = pi17 ? n32 : n24772;
  assign n24774 = pi16 ? n32 : n24773;
  assign n24775 = pi19 ? n507 : n23895;
  assign n24776 = pi18 ? n24775 : n2747;
  assign n24777 = pi17 ? n2726 : ~n24776;
  assign n24778 = pi16 ? n32 : n24777;
  assign n24779 = pi15 ? n24774 : n24778;
  assign n24780 = pi14 ? n24771 : n24779;
  assign n24781 = pi18 ? n32 : n24063;
  assign n24782 = pi19 ? n18497 : n5694;
  assign n24783 = pi18 ? n24782 : ~n8908;
  assign n24784 = pi17 ? n24781 : ~n24783;
  assign n24785 = pi16 ? n32 : n24784;
  assign n24786 = pi18 ? n32 : n23073;
  assign n24787 = pi18 ? n16847 : n2754;
  assign n24788 = pi17 ? n24786 : ~n24787;
  assign n24789 = pi16 ? n32 : n24788;
  assign n24790 = pi15 ? n24785 : n24789;
  assign n24791 = pi14 ? n24790 : n21695;
  assign n24792 = pi13 ? n24780 : n24791;
  assign n24793 = pi12 ? n24762 : n24792;
  assign n24794 = pi11 ? n24746 : n24793;
  assign n24795 = pi10 ? n24723 : n24794;
  assign n24796 = pi09 ? n32 : n24795;
  assign n24797 = pi15 ? n32 : n16837;
  assign n24798 = pi14 ? n24797 : n16837;
  assign n24799 = pi15 ? n16837 : n32;
  assign n24800 = pi14 ? n24799 : n24691;
  assign n24801 = pi13 ? n24798 : n24800;
  assign n24802 = pi12 ? n32 : n24801;
  assign n24803 = pi15 ? n16520 : n24495;
  assign n24804 = pi14 ? n24803 : n24495;
  assign n24805 = pi15 ? n24700 : n15230;
  assign n24806 = pi14 ? n24701 : n24805;
  assign n24807 = pi13 ? n24804 : n24806;
  assign n24808 = pi15 ? n24700 : n16101;
  assign n24809 = pi14 ? n24808 : n24572;
  assign n24810 = pi19 ? n32 : ~n288;
  assign n24811 = pi18 ? n32 : n24810;
  assign n24812 = pi17 ? n32 : n24811;
  assign n24813 = pi16 ? n32 : n24812;
  assign n24814 = pi15 ? n24382 : n24289;
  assign n24815 = pi14 ? n24813 : n24814;
  assign n24816 = pi13 ? n24809 : n24815;
  assign n24817 = pi12 ? n24807 : n24816;
  assign n24818 = pi11 ? n24802 : n24817;
  assign n24819 = pi18 ? n22865 : n14329;
  assign n24820 = pi17 ? n32 : n24819;
  assign n24821 = pi16 ? n32 : n24820;
  assign n24822 = pi15 ? n24382 : n24821;
  assign n24823 = pi18 ? n16389 : n14329;
  assign n24824 = pi17 ? n32 : n24823;
  assign n24825 = pi16 ? n32 : n24824;
  assign n24826 = pi19 ? n1248 : ~n2848;
  assign n24827 = pi18 ? n32 : n24826;
  assign n24828 = pi17 ? n32 : n24827;
  assign n24829 = pi16 ? n32 : n24828;
  assign n24830 = pi15 ? n24825 : n24829;
  assign n24831 = pi14 ? n24822 : n24830;
  assign n24832 = pi14 ? n16105 : n23732;
  assign n24833 = pi13 ? n24831 : n24832;
  assign n24834 = pi14 ? n23421 : n23749;
  assign n24835 = pi19 ? n507 : ~n1941;
  assign n24836 = pi18 ? n32 : n24835;
  assign n24837 = pi17 ? n32 : n24836;
  assign n24838 = pi16 ? n32 : n24837;
  assign n24839 = pi15 ? n24838 : n23484;
  assign n24840 = pi15 ? n23484 : n15518;
  assign n24841 = pi14 ? n24839 : n24840;
  assign n24842 = pi13 ? n24834 : n24841;
  assign n24843 = pi12 ? n24833 : n24842;
  assign n24844 = pi15 ? n22540 : n23443;
  assign n24845 = pi14 ? n24329 : n24844;
  assign n24846 = pi15 ? n23443 : n23094;
  assign n24847 = pi18 ? n24756 : n22630;
  assign n24848 = pi17 ? n32 : n24847;
  assign n24849 = pi16 ? n32 : n24848;
  assign n24850 = pi15 ? n24754 : n24849;
  assign n24851 = pi14 ? n24846 : n24850;
  assign n24852 = pi13 ? n24845 : n24851;
  assign n24853 = pi18 ? n24775 : n508;
  assign n24854 = pi17 ? n2726 : ~n24853;
  assign n24855 = pi16 ? n32 : n24854;
  assign n24856 = pi15 ? n24774 : n24855;
  assign n24857 = pi14 ? n24771 : n24856;
  assign n24858 = pi18 ? n24782 : ~n13341;
  assign n24859 = pi17 ? n24781 : ~n24858;
  assign n24860 = pi16 ? n32 : n24859;
  assign n24861 = pi18 ? n16847 : n520;
  assign n24862 = pi17 ? n24786 : ~n24861;
  assign n24863 = pi16 ? n32 : n24862;
  assign n24864 = pi15 ? n24860 : n24863;
  assign n24865 = pi14 ? n24864 : n21695;
  assign n24866 = pi13 ? n24857 : n24865;
  assign n24867 = pi12 ? n24852 : n24866;
  assign n24868 = pi11 ? n24843 : n24867;
  assign n24869 = pi10 ? n24818 : n24868;
  assign n24870 = pi09 ? n32 : n24869;
  assign n24871 = pi08 ? n24796 : n24870;
  assign n24872 = pi18 ? n32 : n20565;
  assign n24873 = pi17 ? n32 : n24872;
  assign n24874 = pi16 ? n32 : n24873;
  assign n24875 = pi15 ? n32 : n24874;
  assign n24876 = pi14 ? n32 : n24875;
  assign n24877 = pi13 ? n32 : n24876;
  assign n24878 = pi12 ? n32 : n24877;
  assign n24879 = pi15 ? n24874 : n16786;
  assign n24880 = pi15 ? n16786 : n16520;
  assign n24881 = pi14 ? n24879 : n24880;
  assign n24882 = pi15 ? n16452 : n24700;
  assign n24883 = pi19 ? n4126 : ~n343;
  assign n24884 = pi18 ? n32 : n24883;
  assign n24885 = pi17 ? n32 : n24884;
  assign n24886 = pi16 ? n32 : n24885;
  assign n24887 = pi15 ? n24700 : n24886;
  assign n24888 = pi14 ? n24882 : n24887;
  assign n24889 = pi13 ? n24881 : n24888;
  assign n24890 = pi15 ? n16452 : n24572;
  assign n24891 = pi14 ? n24808 : n24890;
  assign n24892 = pi14 ? n24813 : n24435;
  assign n24893 = pi13 ? n24891 : n24892;
  assign n24894 = pi12 ? n24889 : n24893;
  assign n24895 = pi11 ? n24878 : n24894;
  assign n24896 = pi18 ? n17118 : n14329;
  assign n24897 = pi17 ? n32 : n24896;
  assign n24898 = pi16 ? n32 : n24897;
  assign n24899 = pi15 ? n24382 : n24898;
  assign n24900 = pi15 ? n14332 : n24289;
  assign n24901 = pi14 ? n24899 : n24900;
  assign n24902 = pi19 ? n32 : n24648;
  assign n24903 = pi18 ? n32 : n24902;
  assign n24904 = pi17 ? n32 : n24903;
  assign n24905 = pi16 ? n32 : n24904;
  assign n24906 = pi15 ? n24905 : n32;
  assign n24907 = pi14 ? n16105 : n24906;
  assign n24908 = pi13 ? n24901 : n24907;
  assign n24909 = pi15 ? n23749 : n23484;
  assign n24910 = pi14 ? n24909 : n15655;
  assign n24911 = pi13 ? n24834 : n24910;
  assign n24912 = pi12 ? n24908 : n24911;
  assign n24913 = pi15 ? n22923 : n1109;
  assign n24914 = pi15 ? n22817 : n23443;
  assign n24915 = pi14 ? n24913 : n24914;
  assign n24916 = pi19 ? n2359 : n32;
  assign n24917 = pi18 ? n32 : n24916;
  assign n24918 = pi17 ? n32 : n24917;
  assign n24919 = pi16 ? n32 : n24918;
  assign n24920 = pi15 ? n23443 : n24919;
  assign n24921 = pi18 ? n16389 : n24751;
  assign n24922 = pi17 ? n32 : n24921;
  assign n24923 = pi16 ? n32 : n24922;
  assign n24924 = pi20 ? n246 : n101;
  assign n24925 = pi19 ? n24924 : ~n32;
  assign n24926 = pi18 ? n1758 : ~n24925;
  assign n24927 = pi17 ? n32 : n24926;
  assign n24928 = pi16 ? n32 : n24927;
  assign n24929 = pi15 ? n24923 : n24928;
  assign n24930 = pi14 ? n24920 : n24929;
  assign n24931 = pi13 ? n24915 : n24930;
  assign n24932 = pi19 ? n32 : ~n267;
  assign n24933 = pi20 ? n321 : n101;
  assign n24934 = pi19 ? n24933 : ~n32;
  assign n24935 = pi18 ? n24932 : ~n24934;
  assign n24936 = pi17 ? n32 : n24935;
  assign n24937 = pi16 ? n32 : n24936;
  assign n24938 = pi18 ? n14982 : n20912;
  assign n24939 = pi17 ? n32 : n24938;
  assign n24940 = pi16 ? n32 : n24939;
  assign n24941 = pi15 ? n24937 : n24940;
  assign n24942 = pi19 ? n32 : n11879;
  assign n24943 = pi18 ? n24942 : n508;
  assign n24944 = pi17 ? n2726 : ~n24943;
  assign n24945 = pi16 ? n32 : n24944;
  assign n24946 = pi15 ? n24774 : n24945;
  assign n24947 = pi14 ? n24941 : n24946;
  assign n24948 = pi18 ? n32 : n276;
  assign n24949 = pi19 ? n3523 : ~n22480;
  assign n24950 = pi18 ? n24949 : n22003;
  assign n24951 = pi17 ? n24948 : n24950;
  assign n24952 = pi16 ? n32 : n24951;
  assign n24953 = pi17 ? n2119 : ~n24861;
  assign n24954 = pi16 ? n32 : n24953;
  assign n24955 = pi15 ? n24952 : n24954;
  assign n24956 = pi14 ? n24955 : n22228;
  assign n24957 = pi13 ? n24947 : n24956;
  assign n24958 = pi12 ? n24931 : n24957;
  assign n24959 = pi11 ? n24912 : n24958;
  assign n24960 = pi10 ? n24895 : n24959;
  assign n24961 = pi09 ? n32 : n24960;
  assign n24962 = pi15 ? n32 : n16973;
  assign n24963 = pi14 ? n24962 : n16973;
  assign n24964 = pi13 ? n24963 : n24876;
  assign n24965 = pi12 ? n32 : n24964;
  assign n24966 = pi15 ? n24874 : n16655;
  assign n24967 = pi15 ? n16655 : n16520;
  assign n24968 = pi14 ? n24966 : n24967;
  assign n24969 = pi13 ? n24968 : n24888;
  assign n24970 = pi14 ? n24808 : n16452;
  assign n24971 = pi19 ? n32 : ~n20266;
  assign n24972 = pi18 ? n32 : n24971;
  assign n24973 = pi17 ? n32 : n24972;
  assign n24974 = pi16 ? n32 : n24973;
  assign n24975 = pi15 ? n24974 : n24813;
  assign n24976 = pi15 ? n24511 : n24504;
  assign n24977 = pi14 ? n24975 : n24976;
  assign n24978 = pi13 ? n24970 : n24977;
  assign n24979 = pi12 ? n24969 : n24978;
  assign n24980 = pi11 ? n24965 : n24979;
  assign n24981 = pi19 ? n531 : ~n589;
  assign n24982 = pi18 ? n17118 : n24981;
  assign n24983 = pi17 ? n32 : n24982;
  assign n24984 = pi16 ? n32 : n24983;
  assign n24985 = pi15 ? n24511 : n24984;
  assign n24986 = pi18 ? n32 : n24981;
  assign n24987 = pi17 ? n32 : n24986;
  assign n24988 = pi16 ? n32 : n24987;
  assign n24989 = pi15 ? n24988 : n24289;
  assign n24990 = pi14 ? n24985 : n24989;
  assign n24991 = pi15 ? n24289 : n16105;
  assign n24992 = pi14 ? n24991 : n23794;
  assign n24993 = pi13 ? n24990 : n24992;
  assign n24994 = pi14 ? n23574 : n24170;
  assign n24995 = pi14 ? n23749 : n24397;
  assign n24996 = pi13 ? n24994 : n24995;
  assign n24997 = pi12 ? n24993 : n24996;
  assign n24998 = pi19 ? n322 : ~n1105;
  assign n24999 = pi18 ? n32 : n24998;
  assign n25000 = pi17 ? n32 : n24999;
  assign n25001 = pi16 ? n32 : n25000;
  assign n25002 = pi15 ? n23011 : n25001;
  assign n25003 = pi14 ? n22923 : n25002;
  assign n25004 = pi18 ? n16389 : n13901;
  assign n25005 = pi17 ? n32 : n25004;
  assign n25006 = pi16 ? n32 : n25005;
  assign n25007 = pi15 ? n25006 : n24928;
  assign n25008 = pi14 ? n24920 : n25007;
  assign n25009 = pi13 ? n25003 : n25008;
  assign n25010 = pi19 ? n23688 : ~n32;
  assign n25011 = pi18 ? n24932 : ~n25010;
  assign n25012 = pi17 ? n32 : n25011;
  assign n25013 = pi16 ? n32 : n25012;
  assign n25014 = pi18 ? n14982 : n14787;
  assign n25015 = pi17 ? n32 : n25014;
  assign n25016 = pi16 ? n32 : n25015;
  assign n25017 = pi15 ? n25013 : n25016;
  assign n25018 = pi18 ? n14153 : n14140;
  assign n25019 = pi17 ? n32 : n25018;
  assign n25020 = pi16 ? n32 : n25019;
  assign n25021 = pi15 ? n25020 : n24945;
  assign n25022 = pi14 ? n25017 : n25021;
  assign n25023 = pi19 ? n3523 : ~n236;
  assign n25024 = pi18 ? n25023 : n22003;
  assign n25025 = pi17 ? n32 : n25024;
  assign n25026 = pi16 ? n32 : n25025;
  assign n25027 = pi15 ? n25026 : n24954;
  assign n25028 = pi14 ? n25027 : n14394;
  assign n25029 = pi13 ? n25022 : n25028;
  assign n25030 = pi12 ? n25009 : n25029;
  assign n25031 = pi11 ? n24997 : n25030;
  assign n25032 = pi10 ? n24980 : n25031;
  assign n25033 = pi09 ? n32 : n25032;
  assign n25034 = pi08 ? n24961 : n25033;
  assign n25035 = pi07 ? n24871 : n25034;
  assign n25036 = pi14 ? n32 : n16973;
  assign n25037 = pi15 ? n24874 : n16899;
  assign n25038 = pi14 ? n16974 : n25037;
  assign n25039 = pi13 ? n25036 : n25038;
  assign n25040 = pi12 ? n32 : n25039;
  assign n25041 = pi19 ? n32 : n7443;
  assign n25042 = pi18 ? n32 : n25041;
  assign n25043 = pi17 ? n32 : n25042;
  assign n25044 = pi16 ? n32 : n25043;
  assign n25045 = pi14 ? n16520 : n25044;
  assign n25046 = pi13 ? n16837 : n25045;
  assign n25047 = pi19 ? n32 : n10632;
  assign n25048 = pi18 ? n32 : n25047;
  assign n25049 = pi17 ? n32 : n25048;
  assign n25050 = pi16 ? n32 : n25049;
  assign n25051 = pi15 ? n16101 : n25050;
  assign n25052 = pi14 ? n16520 : n25051;
  assign n25053 = pi15 ? n24572 : n24504;
  assign n25054 = pi15 ? n24237 : n16105;
  assign n25055 = pi14 ? n25053 : n25054;
  assign n25056 = pi13 ? n25052 : n25055;
  assign n25057 = pi12 ? n25046 : n25056;
  assign n25058 = pi11 ? n25040 : n25057;
  assign n25059 = pi19 ? n208 : n9724;
  assign n25060 = pi18 ? n32 : n25059;
  assign n25061 = pi17 ? n32 : n25060;
  assign n25062 = pi16 ? n32 : n25061;
  assign n25063 = pi19 ? n2386 : n9724;
  assign n25064 = pi18 ? n32 : n25063;
  assign n25065 = pi17 ? n32 : n25064;
  assign n25066 = pi16 ? n32 : n25065;
  assign n25067 = pi19 ? n32 : n19019;
  assign n25068 = pi18 ? n32 : n25067;
  assign n25069 = pi17 ? n32 : n25068;
  assign n25070 = pi16 ? n32 : n25069;
  assign n25071 = pi15 ? n25066 : n25070;
  assign n25072 = pi14 ? n25062 : n25071;
  assign n25073 = pi15 ? n25070 : n16314;
  assign n25074 = pi14 ? n25073 : n23794;
  assign n25075 = pi13 ? n25072 : n25074;
  assign n25076 = pi15 ? n23574 : n23933;
  assign n25077 = pi14 ? n23623 : n25076;
  assign n25078 = pi15 ? n23749 : n23250;
  assign n25079 = pi14 ? n23749 : n25078;
  assign n25080 = pi13 ? n25077 : n25079;
  assign n25081 = pi12 ? n25075 : n25080;
  assign n25082 = pi19 ? n4126 : ~n1105;
  assign n25083 = pi18 ? n32 : n25082;
  assign n25084 = pi17 ? n32 : n25083;
  assign n25085 = pi16 ? n32 : n25084;
  assign n25086 = pi15 ? n23011 : n25085;
  assign n25087 = pi14 ? n22923 : n25086;
  assign n25088 = pi15 ? n25001 : n23443;
  assign n25089 = pi20 ? n207 : ~n101;
  assign n25090 = pi19 ? n25089 : n32;
  assign n25091 = pi18 ? n17118 : n25090;
  assign n25092 = pi17 ? n32 : n25091;
  assign n25093 = pi16 ? n32 : n25092;
  assign n25094 = pi15 ? n14138 : n25093;
  assign n25095 = pi14 ? n25088 : n25094;
  assign n25096 = pi13 ? n25087 : n25095;
  assign n25097 = pi18 ? n15844 : n4098;
  assign n25098 = pi17 ? n2726 : ~n25097;
  assign n25099 = pi16 ? n32 : n25098;
  assign n25100 = pi20 ? n321 : ~n10878;
  assign n25101 = pi19 ? n25100 : ~n32;
  assign n25102 = pi18 ? n21274 : ~n25101;
  assign n25103 = pi17 ? n32 : n25102;
  assign n25104 = pi16 ? n32 : n25103;
  assign n25105 = pi15 ? n25099 : n25104;
  assign n25106 = pi18 ? n323 : n14603;
  assign n25107 = pi17 ? n32 : n25106;
  assign n25108 = pi16 ? n32 : n25107;
  assign n25109 = pi19 ? n6018 : n236;
  assign n25110 = pi19 ? n1508 : ~n32;
  assign n25111 = pi18 ? n25109 : ~n25110;
  assign n25112 = pi17 ? n32 : n25111;
  assign n25113 = pi16 ? n32 : n25112;
  assign n25114 = pi15 ? n25108 : n25113;
  assign n25115 = pi14 ? n25105 : n25114;
  assign n25116 = pi19 ? n9220 : n32;
  assign n25117 = pi18 ? n1965 : n25116;
  assign n25118 = pi17 ? n32 : n25117;
  assign n25119 = pi16 ? n32 : n25118;
  assign n25120 = pi20 ? n220 : n321;
  assign n25121 = pi19 ? n25120 : n22525;
  assign n25122 = pi18 ? n25121 : ~n24472;
  assign n25123 = pi17 ? n32 : n25122;
  assign n25124 = pi16 ? n32 : n25123;
  assign n25125 = pi15 ? n25119 : n25124;
  assign n25126 = pi15 ? n21543 : n14394;
  assign n25127 = pi14 ? n25125 : n25126;
  assign n25128 = pi13 ? n25115 : n25127;
  assign n25129 = pi12 ? n25096 : n25128;
  assign n25130 = pi11 ? n25081 : n25129;
  assign n25131 = pi10 ? n25058 : n25130;
  assign n25132 = pi09 ? n32 : n25131;
  assign n25133 = pi15 ? n17039 : n32;
  assign n25134 = pi14 ? n17039 : n25133;
  assign n25135 = pi14 ? n32 : n25037;
  assign n25136 = pi13 ? n25134 : n25135;
  assign n25137 = pi12 ? n32 : n25136;
  assign n25138 = pi15 ? n16899 : n16837;
  assign n25139 = pi14 ? n25138 : n16837;
  assign n25140 = pi15 ? n16101 : n25044;
  assign n25141 = pi14 ? n16452 : n25140;
  assign n25142 = pi13 ? n25139 : n25141;
  assign n25143 = pi20 ? n14374 : n32;
  assign n25144 = pi19 ? n32 : n25143;
  assign n25145 = pi18 ? n32 : n25144;
  assign n25146 = pi17 ? n32 : n25145;
  assign n25147 = pi16 ? n32 : n25146;
  assign n25148 = pi15 ? n25044 : n25147;
  assign n25149 = pi14 ? n16520 : n25148;
  assign n25150 = pi15 ? n16452 : n24712;
  assign n25151 = pi20 ? n17509 : n32;
  assign n25152 = pi19 ? n32 : n25151;
  assign n25153 = pi18 ? n32 : n25152;
  assign n25154 = pi17 ? n32 : n25153;
  assign n25155 = pi16 ? n32 : n25154;
  assign n25156 = pi15 ? n24572 : n25155;
  assign n25157 = pi14 ? n25150 : n25156;
  assign n25158 = pi13 ? n25149 : n25157;
  assign n25159 = pi12 ? n25142 : n25158;
  assign n25160 = pi11 ? n25137 : n25159;
  assign n25161 = pi19 ? n208 : n7468;
  assign n25162 = pi18 ? n32 : n25161;
  assign n25163 = pi17 ? n32 : n25162;
  assign n25164 = pi16 ? n32 : n25163;
  assign n25165 = pi15 ? n25066 : n24237;
  assign n25166 = pi14 ? n25164 : n25165;
  assign n25167 = pi15 ? n24237 : n16314;
  assign n25168 = pi14 ? n25167 : n16321;
  assign n25169 = pi13 ? n25166 : n25168;
  assign n25170 = pi15 ? n23725 : n23730;
  assign n25171 = pi15 ? n23730 : n23933;
  assign n25172 = pi14 ? n25170 : n25171;
  assign n25173 = pi14 ? n23933 : n25078;
  assign n25174 = pi13 ? n25172 : n25173;
  assign n25175 = pi12 ? n25169 : n25174;
  assign n25176 = pi15 ? n15119 : n25085;
  assign n25177 = pi14 ? n15518 : n25176;
  assign n25178 = pi18 ? n17118 : n23514;
  assign n25179 = pi17 ? n32 : n25178;
  assign n25180 = pi16 ? n32 : n25179;
  assign n25181 = pi15 ? n14131 : n25180;
  assign n25182 = pi14 ? n25001 : n25181;
  assign n25183 = pi13 ? n25177 : n25182;
  assign n25184 = pi20 ? n32 : n10878;
  assign n25185 = pi19 ? n25184 : n32;
  assign n25186 = pi18 ? n323 : n25185;
  assign n25187 = pi17 ? n32 : n25186;
  assign n25188 = pi16 ? n32 : n25187;
  assign n25189 = pi20 ? n32 : ~n7442;
  assign n25190 = pi19 ? n25189 : ~n32;
  assign n25191 = pi18 ? n25109 : ~n25190;
  assign n25192 = pi17 ? n32 : n25191;
  assign n25193 = pi16 ? n32 : n25192;
  assign n25194 = pi15 ? n25188 : n25193;
  assign n25195 = pi14 ? n25105 : n25194;
  assign n25196 = pi15 ? n21686 : n22006;
  assign n25197 = pi14 ? n25125 : n25196;
  assign n25198 = pi13 ? n25195 : n25197;
  assign n25199 = pi12 ? n25183 : n25198;
  assign n25200 = pi11 ? n25175 : n25199;
  assign n25201 = pi10 ? n25160 : n25200;
  assign n25202 = pi09 ? n32 : n25201;
  assign n25203 = pi08 ? n25132 : n25202;
  assign n25204 = pi15 ? n24874 : n16392;
  assign n25205 = pi14 ? n32 : n25204;
  assign n25206 = pi13 ? n25134 : n25205;
  assign n25207 = pi12 ? n32 : n25206;
  assign n25208 = pi19 ? n32 : n10645;
  assign n25209 = pi18 ? n32 : n25208;
  assign n25210 = pi17 ? n32 : n25209;
  assign n25211 = pi16 ? n32 : n25210;
  assign n25212 = pi14 ? n24874 : n25211;
  assign n25213 = pi13 ? n16899 : n25212;
  assign n25214 = pi14 ? n24874 : n16520;
  assign n25215 = pi15 ? n16298 : n16105;
  assign n25216 = pi19 ? n6398 : ~n349;
  assign n25217 = pi18 ? n32 : n25216;
  assign n25218 = pi17 ? n32 : n25217;
  assign n25219 = pi16 ? n32 : n25218;
  assign n25220 = pi15 ? n32 : n25219;
  assign n25221 = pi14 ? n25215 : n25220;
  assign n25222 = pi13 ? n25214 : n25221;
  assign n25223 = pi12 ? n25213 : n25222;
  assign n25224 = pi11 ? n25207 : n25223;
  assign n25225 = pi19 ? n1464 : ~n2317;
  assign n25226 = pi18 ? n32 : n25225;
  assign n25227 = pi17 ? n32 : n25226;
  assign n25228 = pi16 ? n32 : n25227;
  assign n25229 = pi14 ? n25228 : n24573;
  assign n25230 = pi15 ? n24237 : n16308;
  assign n25231 = pi14 ? n25230 : n16321;
  assign n25232 = pi13 ? n25229 : n25231;
  assign n25233 = pi14 ? n23726 : n25170;
  assign n25234 = pi15 ? n23574 : n24256;
  assign n25235 = pi14 ? n25234 : n23631;
  assign n25236 = pi13 ? n25233 : n25235;
  assign n25237 = pi12 ? n25232 : n25236;
  assign n25238 = pi19 ? n594 : n5626;
  assign n25239 = pi18 ? n32 : n25238;
  assign n25240 = pi17 ? n32 : n25239;
  assign n25241 = pi16 ? n32 : n25240;
  assign n25242 = pi15 ? n23160 : n25241;
  assign n25243 = pi14 ? n25242 : n23340;
  assign n25244 = pi19 ? n322 : ~n617;
  assign n25245 = pi18 ? n32 : n25244;
  assign n25246 = pi17 ? n32 : n25245;
  assign n25247 = pi16 ? n32 : n25246;
  assign n25248 = pi19 ? n208 : ~n1105;
  assign n25249 = pi18 ? n32 : n25248;
  assign n25250 = pi17 ? n32 : n25249;
  assign n25251 = pi16 ? n32 : n25250;
  assign n25252 = pi15 ? n25247 : n25251;
  assign n25253 = pi15 ? n14131 : n23517;
  assign n25254 = pi14 ? n25252 : n25253;
  assign n25255 = pi13 ? n25243 : n25254;
  assign n25256 = pi20 ? n321 : ~n17654;
  assign n25257 = pi19 ? n25256 : ~n32;
  assign n25258 = pi18 ? n21274 : ~n25257;
  assign n25259 = pi17 ? n32 : n25258;
  assign n25260 = pi16 ? n32 : n25259;
  assign n25261 = pi15 ? n25099 : n25260;
  assign n25262 = pi18 ? n323 : n24540;
  assign n25263 = pi17 ? n32 : n25262;
  assign n25264 = pi16 ? n32 : n25263;
  assign n25265 = pi20 ? n339 : n175;
  assign n25266 = pi19 ? n32 : ~n25265;
  assign n25267 = pi20 ? n357 : n7880;
  assign n25268 = pi19 ? n25267 : n32;
  assign n25269 = pi18 ? n25266 : n25268;
  assign n25270 = pi17 ? n32 : n25269;
  assign n25271 = pi16 ? n32 : n25270;
  assign n25272 = pi15 ? n25264 : n25271;
  assign n25273 = pi14 ? n25261 : n25272;
  assign n25274 = pi18 ? n880 : n14787;
  assign n25275 = pi17 ? n32 : n25274;
  assign n25276 = pi16 ? n32 : n25275;
  assign n25277 = pi19 ? n23644 : n4126;
  assign n25278 = pi18 ? n25277 : ~n24548;
  assign n25279 = pi17 ? n32 : n25278;
  assign n25280 = pi16 ? n32 : n25279;
  assign n25281 = pi15 ? n25276 : n25280;
  assign n25282 = pi14 ? n25281 : n25196;
  assign n25283 = pi13 ? n25273 : n25282;
  assign n25284 = pi12 ? n25255 : n25283;
  assign n25285 = pi11 ? n25237 : n25284;
  assign n25286 = pi10 ? n25224 : n25285;
  assign n25287 = pi09 ? n32 : n25286;
  assign n25288 = pi14 ? n32 : n17273;
  assign n25289 = pi13 ? n32 : n25288;
  assign n25290 = pi14 ? n17188 : n17189;
  assign n25291 = pi15 ? n15847 : n16392;
  assign n25292 = pi14 ? n32 : n25291;
  assign n25293 = pi13 ? n25290 : n25292;
  assign n25294 = pi12 ? n25289 : n25293;
  assign n25295 = pi15 ? n16392 : n16899;
  assign n25296 = pi14 ? n25295 : n16899;
  assign n25297 = pi13 ? n25296 : n25212;
  assign n25298 = pi19 ? n32 : n6314;
  assign n25299 = pi18 ? n32 : n25298;
  assign n25300 = pi17 ? n32 : n25299;
  assign n25301 = pi16 ? n32 : n25300;
  assign n25302 = pi15 ? n16298 : n25301;
  assign n25303 = pi19 ? n6398 : ~n1077;
  assign n25304 = pi18 ? n32 : n25303;
  assign n25305 = pi17 ? n32 : n25304;
  assign n25306 = pi16 ? n32 : n25305;
  assign n25307 = pi15 ? n16606 : n25306;
  assign n25308 = pi14 ? n25302 : n25307;
  assign n25309 = pi13 ? n24874 : n25308;
  assign n25310 = pi12 ? n25297 : n25309;
  assign n25311 = pi11 ? n25294 : n25310;
  assign n25312 = pi19 ? n1464 : ~n343;
  assign n25313 = pi18 ? n32 : n25312;
  assign n25314 = pi17 ? n32 : n25313;
  assign n25315 = pi16 ? n32 : n25314;
  assign n25316 = pi19 ? n32 : n20951;
  assign n25317 = pi18 ? n32 : n25316;
  assign n25318 = pi17 ? n32 : n25317;
  assign n25319 = pi16 ? n32 : n25318;
  assign n25320 = pi15 ? n24367 : n25319;
  assign n25321 = pi14 ? n25315 : n25320;
  assign n25322 = pi15 ? n25319 : n24237;
  assign n25323 = pi15 ? n16377 : n23981;
  assign n25324 = pi14 ? n25322 : n25323;
  assign n25325 = pi13 ? n25321 : n25324;
  assign n25326 = pi15 ? n32 : n24905;
  assign n25327 = pi14 ? n23981 : n25326;
  assign n25328 = pi19 ? n32 : n19892;
  assign n25329 = pi18 ? n32 : n25328;
  assign n25330 = pi17 ? n32 : n25329;
  assign n25331 = pi16 ? n32 : n25330;
  assign n25332 = pi15 ? n24905 : n25331;
  assign n25333 = pi15 ? n23574 : n23631;
  assign n25334 = pi14 ? n25332 : n25333;
  assign n25335 = pi13 ? n25327 : n25334;
  assign n25336 = pi12 ? n25325 : n25335;
  assign n25337 = pi19 ? n594 : n358;
  assign n25338 = pi18 ? n32 : n25337;
  assign n25339 = pi17 ? n32 : n25338;
  assign n25340 = pi16 ? n32 : n25339;
  assign n25341 = pi15 ? n23250 : n25340;
  assign n25342 = pi14 ? n25341 : n23340;
  assign n25343 = pi15 ? n25247 : n14580;
  assign n25344 = pi18 ? n32 : n6384;
  assign n25345 = pi17 ? n32 : n25344;
  assign n25346 = pi16 ? n32 : n25345;
  assign n25347 = pi15 ? n25346 : n13321;
  assign n25348 = pi14 ? n25343 : n25347;
  assign n25349 = pi13 ? n25342 : n25348;
  assign n25350 = pi18 ? n15844 : n702;
  assign n25351 = pi17 ? n2726 : ~n25350;
  assign n25352 = pi16 ? n32 : n25351;
  assign n25353 = pi15 ? n25352 : n25260;
  assign n25354 = pi18 ? n323 : n22630;
  assign n25355 = pi17 ? n32 : n25354;
  assign n25356 = pi16 ? n32 : n25355;
  assign n25357 = pi19 ? n32 : n12821;
  assign n25358 = pi18 ? n25357 : n20912;
  assign n25359 = pi17 ? n32 : n25358;
  assign n25360 = pi16 ? n32 : n25359;
  assign n25361 = pi15 ? n25356 : n25360;
  assign n25362 = pi14 ? n25353 : n25361;
  assign n25363 = pi15 ? n21853 : n22006;
  assign n25364 = pi14 ? n25281 : n25363;
  assign n25365 = pi13 ? n25362 : n25364;
  assign n25366 = pi12 ? n25349 : n25365;
  assign n25367 = pi11 ? n25336 : n25366;
  assign n25368 = pi10 ? n25311 : n25367;
  assign n25369 = pi09 ? n32 : n25368;
  assign n25370 = pi08 ? n25287 : n25369;
  assign n25371 = pi07 ? n25203 : n25370;
  assign n25372 = pi06 ? n25035 : n25371;
  assign n25373 = pi05 ? n24689 : n25372;
  assign n25374 = pi14 ? n32 : n16940;
  assign n25375 = pi13 ? n25290 : n25374;
  assign n25376 = pi12 ? n25289 : n25375;
  assign n25377 = pi15 ? n16392 : n17039;
  assign n25378 = pi15 ? n17039 : n16392;
  assign n25379 = pi14 ? n25377 : n25378;
  assign n25380 = pi13 ? n25379 : n16899;
  assign n25381 = pi19 ? n32 : n19847;
  assign n25382 = pi18 ? n32 : n25381;
  assign n25383 = pi17 ? n32 : n25382;
  assign n25384 = pi16 ? n32 : n25383;
  assign n25385 = pi15 ? n16899 : n25384;
  assign n25386 = pi14 ? n25385 : n24874;
  assign n25387 = pi15 ? n16452 : n16606;
  assign n25388 = pi14 ? n25387 : n16452;
  assign n25389 = pi13 ? n25386 : n25388;
  assign n25390 = pi12 ? n25380 : n25389;
  assign n25391 = pi11 ? n25376 : n25390;
  assign n25392 = pi15 ? n16298 : n16606;
  assign n25393 = pi14 ? n25392 : n24890;
  assign n25394 = pi14 ? n24573 : n16378;
  assign n25395 = pi13 ? n25393 : n25394;
  assign n25396 = pi14 ? n23730 : n16108;
  assign n25397 = pi13 ? n16105 : n25396;
  assign n25398 = pi12 ? n25395 : n25397;
  assign n25399 = pi14 ? n24659 : n23761;
  assign n25400 = pi15 ? n24612 : n25247;
  assign n25401 = pi15 ? n25346 : n14138;
  assign n25402 = pi14 ? n25400 : n25401;
  assign n25403 = pi13 ? n25399 : n25402;
  assign n25404 = pi18 ? n1249 : ~n702;
  assign n25405 = pi17 ? n32 : n25404;
  assign n25406 = pi16 ? n32 : n25405;
  assign n25407 = pi15 ? n25406 : n12059;
  assign n25408 = pi20 ? n266 : ~n101;
  assign n25409 = pi19 ? n25408 : n32;
  assign n25410 = pi18 ? n12368 : n25409;
  assign n25411 = pi17 ? n32 : n25410;
  assign n25412 = pi16 ? n32 : n25411;
  assign n25413 = pi18 ? n16389 : n22431;
  assign n25414 = pi17 ? n32 : n25413;
  assign n25415 = pi16 ? n32 : n25414;
  assign n25416 = pi15 ? n25412 : n25415;
  assign n25417 = pi14 ? n25407 : n25416;
  assign n25418 = pi20 ? n274 : n1385;
  assign n25419 = pi19 ? n25418 : n32;
  assign n25420 = pi18 ? n8192 : n25419;
  assign n25421 = pi17 ? n32 : n25420;
  assign n25422 = pi16 ? n32 : n25421;
  assign n25423 = pi18 ? n8192 : ~n508;
  assign n25424 = pi17 ? n32 : n25423;
  assign n25425 = pi16 ? n32 : n25424;
  assign n25426 = pi15 ? n25422 : n25425;
  assign n25427 = pi14 ? n25426 : n22136;
  assign n25428 = pi13 ? n25417 : n25427;
  assign n25429 = pi12 ? n25403 : n25428;
  assign n25430 = pi11 ? n25398 : n25429;
  assign n25431 = pi10 ? n25391 : n25430;
  assign n25432 = pi09 ? n32 : n25431;
  assign n25433 = pi14 ? n32 : n17112;
  assign n25434 = pi13 ? n32 : n25433;
  assign n25435 = pi14 ? n17111 : n17412;
  assign n25436 = pi13 ? n25435 : n25374;
  assign n25437 = pi12 ? n25434 : n25436;
  assign n25438 = pi15 ? n16832 : n17039;
  assign n25439 = pi14 ? n25438 : n25378;
  assign n25440 = pi13 ? n25439 : n16899;
  assign n25441 = pi15 ? n17002 : n25384;
  assign n25442 = pi14 ? n25441 : n25384;
  assign n25443 = pi15 ? n24874 : n16601;
  assign n25444 = pi14 ? n25443 : n16520;
  assign n25445 = pi13 ? n25442 : n25444;
  assign n25446 = pi12 ? n25440 : n25445;
  assign n25447 = pi11 ? n25437 : n25446;
  assign n25448 = pi20 ? n14601 : n32;
  assign n25449 = pi19 ? n32 : n25448;
  assign n25450 = pi18 ? n32 : n25449;
  assign n25451 = pi17 ? n32 : n25450;
  assign n25452 = pi16 ? n32 : n25451;
  assign n25453 = pi15 ? n25452 : n16606;
  assign n25454 = pi14 ? n25453 : n16606;
  assign n25455 = pi15 ? n16606 : n24237;
  assign n25456 = pi15 ? n24237 : n16377;
  assign n25457 = pi14 ? n25455 : n25456;
  assign n25458 = pi13 ? n25454 : n25457;
  assign n25459 = pi14 ? n24991 : n24578;
  assign n25460 = pi14 ? n15700 : n23574;
  assign n25461 = pi13 ? n25459 : n25460;
  assign n25462 = pi12 ? n25458 : n25461;
  assign n25463 = pi19 ? n322 : ~n1941;
  assign n25464 = pi18 ? n32 : n25463;
  assign n25465 = pi17 ? n32 : n25464;
  assign n25466 = pi16 ? n32 : n25465;
  assign n25467 = pi14 ? n25466 : n23761;
  assign n25468 = pi15 ? n25346 : n14131;
  assign n25469 = pi14 ? n24612 : n25468;
  assign n25470 = pi13 ? n25467 : n25469;
  assign n25471 = pi18 ? n1249 : ~n2622;
  assign n25472 = pi17 ? n32 : n25471;
  assign n25473 = pi16 ? n32 : n25472;
  assign n25474 = pi18 ? n684 : ~n702;
  assign n25475 = pi17 ? n32 : n25474;
  assign n25476 = pi16 ? n32 : n25475;
  assign n25477 = pi15 ? n25473 : n25476;
  assign n25478 = pi14 ? n25477 : n25416;
  assign n25479 = pi18 ? n8192 : ~n2627;
  assign n25480 = pi17 ? n32 : n25479;
  assign n25481 = pi16 ? n32 : n25480;
  assign n25482 = pi15 ? n25422 : n25481;
  assign n25483 = pi14 ? n25482 : n22136;
  assign n25484 = pi13 ? n25478 : n25483;
  assign n25485 = pi12 ? n25470 : n25484;
  assign n25486 = pi11 ? n25462 : n25485;
  assign n25487 = pi10 ? n25447 : n25486;
  assign n25488 = pi09 ? n32 : n25487;
  assign n25489 = pi08 ? n25432 : n25488;
  assign n25490 = pi13 ? n32 : n17313;
  assign n25491 = pi14 ? n16984 : n17412;
  assign n25492 = pi15 ? n32 : n17090;
  assign n25493 = pi15 ? n16832 : n17066;
  assign n25494 = pi14 ? n25492 : n25493;
  assign n25495 = pi13 ? n25491 : n25494;
  assign n25496 = pi12 ? n25490 : n25495;
  assign n25497 = pi15 ? n17066 : n17036;
  assign n25498 = pi15 ? n17188 : n16392;
  assign n25499 = pi14 ? n25497 : n25498;
  assign n25500 = pi14 ? n16392 : n25377;
  assign n25501 = pi13 ? n25499 : n25500;
  assign n25502 = pi15 ? n16392 : n15847;
  assign n25503 = pi14 ? n25502 : n25384;
  assign n25504 = pi15 ? n24874 : n32;
  assign n25505 = pi19 ? n507 : n7443;
  assign n25506 = pi18 ? n32 : n25505;
  assign n25507 = pi17 ? n32 : n25506;
  assign n25508 = pi16 ? n32 : n25507;
  assign n25509 = pi14 ? n25504 : n25508;
  assign n25510 = pi13 ? n25503 : n25509;
  assign n25511 = pi12 ? n25501 : n25510;
  assign n25512 = pi11 ? n25496 : n25511;
  assign n25513 = pi21 ? n206 : n7500;
  assign n25514 = pi20 ? n25513 : n32;
  assign n25515 = pi19 ? n594 : n25514;
  assign n25516 = pi18 ? n32 : n25515;
  assign n25517 = pi17 ? n32 : n25516;
  assign n25518 = pi16 ? n32 : n25517;
  assign n25519 = pi15 ? n25518 : n16601;
  assign n25520 = pi14 ? n25519 : n16607;
  assign n25521 = pi15 ? n16452 : n24237;
  assign n25522 = pi14 ? n25521 : n24239;
  assign n25523 = pi13 ? n25520 : n25522;
  assign n25524 = pi14 ? n24289 : n16314;
  assign n25525 = pi14 ? n16105 : n23574;
  assign n25526 = pi13 ? n25524 : n25525;
  assign n25527 = pi12 ? n25523 : n25526;
  assign n25528 = pi15 ? n25466 : n24838;
  assign n25529 = pi14 ? n25528 : n24742;
  assign n25530 = pi19 ? n1325 : ~n2614;
  assign n25531 = pi18 ? n32 : n25530;
  assign n25532 = pi17 ? n32 : n25531;
  assign n25533 = pi16 ? n32 : n25532;
  assign n25534 = pi15 ? n25533 : n24612;
  assign n25535 = pi14 ? n25534 : n25468;
  assign n25536 = pi13 ? n25529 : n25535;
  assign n25537 = pi18 ? n209 : ~n702;
  assign n25538 = pi17 ? n32 : n25537;
  assign n25539 = pi16 ? n32 : n25538;
  assign n25540 = pi15 ? n12753 : n25539;
  assign n25541 = pi15 ? n22825 : n23094;
  assign n25542 = pi14 ? n25540 : n25541;
  assign n25543 = pi18 ? n8192 : n22431;
  assign n25544 = pi17 ? n32 : n25543;
  assign n25545 = pi16 ? n32 : n25544;
  assign n25546 = pi15 ? n25545 : n25481;
  assign n25547 = pi14 ? n25546 : n22136;
  assign n25548 = pi13 ? n25542 : n25547;
  assign n25549 = pi12 ? n25536 : n25548;
  assign n25550 = pi11 ? n25527 : n25549;
  assign n25551 = pi10 ? n25512 : n25550;
  assign n25552 = pi09 ? n32 : n25551;
  assign n25553 = pi19 ? n32 : n482;
  assign n25554 = pi18 ? n32 : n25553;
  assign n25555 = pi17 ? n32 : n25554;
  assign n25556 = pi16 ? n32 : n25555;
  assign n25557 = pi15 ? n32 : n25556;
  assign n25558 = pi14 ? n32 : n25557;
  assign n25559 = pi13 ? n32 : n25558;
  assign n25560 = pi19 ? n32 : n8035;
  assign n25561 = pi18 ? n32 : n25560;
  assign n25562 = pi17 ? n32 : n25561;
  assign n25563 = pi16 ? n32 : n25562;
  assign n25564 = pi15 ? n25563 : n32;
  assign n25565 = pi14 ? n25556 : n25564;
  assign n25566 = pi15 ? n16392 : n17066;
  assign n25567 = pi14 ? n32 : n25566;
  assign n25568 = pi13 ? n25565 : n25567;
  assign n25569 = pi12 ? n25559 : n25568;
  assign n25570 = pi15 ? n16832 : n16485;
  assign n25571 = pi14 ? n25570 : n15847;
  assign n25572 = pi15 ? n24874 : n16837;
  assign n25573 = pi19 ? n507 : n10645;
  assign n25574 = pi18 ? n32 : n25573;
  assign n25575 = pi17 ? n32 : n25574;
  assign n25576 = pi16 ? n32 : n25575;
  assign n25577 = pi14 ? n25572 : n25576;
  assign n25578 = pi13 ? n25571 : n25577;
  assign n25579 = pi12 ? n25501 : n25578;
  assign n25580 = pi11 ? n25569 : n25579;
  assign n25581 = pi19 ? n594 : n1757;
  assign n25582 = pi18 ? n32 : n25581;
  assign n25583 = pi17 ? n32 : n25582;
  assign n25584 = pi16 ? n32 : n25583;
  assign n25585 = pi15 ? n25584 : n16601;
  assign n25586 = pi14 ? n25585 : n16601;
  assign n25587 = pi15 ? n16520 : n24572;
  assign n25588 = pi14 ? n25587 : n24573;
  assign n25589 = pi13 ? n25586 : n25588;
  assign n25590 = pi15 ? n24504 : n24289;
  assign n25591 = pi14 ? n25590 : n16314;
  assign n25592 = pi14 ? n24991 : n23730;
  assign n25593 = pi13 ? n25591 : n25592;
  assign n25594 = pi12 ? n25589 : n25593;
  assign n25595 = pi19 ? n322 : ~n813;
  assign n25596 = pi18 ? n32 : n25595;
  assign n25597 = pi17 ? n32 : n25596;
  assign n25598 = pi16 ? n32 : n25597;
  assign n25599 = pi15 ? n25598 : n24838;
  assign n25600 = pi14 ? n25599 : n24742;
  assign n25601 = pi19 ? n1325 : ~n236;
  assign n25602 = pi18 ? n32 : n25601;
  assign n25603 = pi17 ? n32 : n25602;
  assign n25604 = pi16 ? n32 : n25603;
  assign n25605 = pi15 ? n25604 : n24612;
  assign n25606 = pi14 ? n25605 : n25346;
  assign n25607 = pi13 ? n25600 : n25606;
  assign n25608 = pi20 ? n32 : ~n11560;
  assign n25609 = pi19 ? n25608 : n32;
  assign n25610 = pi18 ? n8192 : n25609;
  assign n25611 = pi17 ? n32 : n25610;
  assign n25612 = pi16 ? n32 : n25611;
  assign n25613 = pi18 ? n8192 : ~n595;
  assign n25614 = pi17 ? n32 : n25613;
  assign n25615 = pi16 ? n32 : n25614;
  assign n25616 = pi15 ? n25612 : n25615;
  assign n25617 = pi14 ? n25616 : n21853;
  assign n25618 = pi13 ? n25542 : n25617;
  assign n25619 = pi12 ? n25607 : n25618;
  assign n25620 = pi11 ? n25594 : n25619;
  assign n25621 = pi10 ? n25580 : n25620;
  assign n25622 = pi09 ? n32 : n25621;
  assign n25623 = pi08 ? n25552 : n25622;
  assign n25624 = pi07 ? n25489 : n25623;
  assign n25625 = pi15 ? n25556 : n32;
  assign n25626 = pi14 ? n25556 : n25625;
  assign n25627 = pi14 ? n32 : n25563;
  assign n25628 = pi13 ? n25626 : n25627;
  assign n25629 = pi12 ? n25559 : n25628;
  assign n25630 = pi15 ? n25563 : n16984;
  assign n25631 = pi15 ? n16984 : n17066;
  assign n25632 = pi14 ? n25630 : n25631;
  assign n25633 = pi15 ? n16832 : n16392;
  assign n25634 = pi15 ? n16832 : n17036;
  assign n25635 = pi14 ? n25633 : n25634;
  assign n25636 = pi13 ? n25632 : n25635;
  assign n25637 = pi15 ? n16629 : n16485;
  assign n25638 = pi15 ? n15403 : n16392;
  assign n25639 = pi14 ? n25637 : n25638;
  assign n25640 = pi15 ? n16837 : n24874;
  assign n25641 = pi14 ? n25640 : n16837;
  assign n25642 = pi13 ? n25639 : n25641;
  assign n25643 = pi12 ? n25636 : n25642;
  assign n25644 = pi11 ? n25629 : n25643;
  assign n25645 = pi15 ? n24874 : n16520;
  assign n25646 = pi14 ? n25640 : n25645;
  assign n25647 = pi15 ? n16520 : n24367;
  assign n25648 = pi14 ? n25647 : n24430;
  assign n25649 = pi13 ? n25646 : n25648;
  assign n25650 = pi15 ? n16308 : n24289;
  assign n25651 = pi14 ? n24237 : n25650;
  assign n25652 = pi14 ? n24991 : n25170;
  assign n25653 = pi13 ? n25651 : n25652;
  assign n25654 = pi12 ? n25649 : n25653;
  assign n25655 = pi18 ? n32 : n20384;
  assign n25656 = pi17 ? n32 : n25655;
  assign n25657 = pi16 ? n32 : n25656;
  assign n25658 = pi15 ? n24838 : n24742;
  assign n25659 = pi14 ? n25657 : n25658;
  assign n25660 = pi15 ? n24742 : n15255;
  assign n25661 = pi15 ? n14580 : n25247;
  assign n25662 = pi14 ? n25660 : n25661;
  assign n25663 = pi13 ? n25659 : n25662;
  assign n25664 = pi19 ? n5371 : ~n1105;
  assign n25665 = pi18 ? n32 : n25664;
  assign n25666 = pi17 ? n32 : n25665;
  assign n25667 = pi16 ? n32 : n25666;
  assign n25668 = pi15 ? n25667 : n25001;
  assign n25669 = pi19 ? n519 : ~n1105;
  assign n25670 = pi18 ? n32 : n25669;
  assign n25671 = pi17 ? n32 : n25670;
  assign n25672 = pi16 ? n32 : n25671;
  assign n25673 = pi19 ? n18159 : n32;
  assign n25674 = pi18 ? n32 : n25673;
  assign n25675 = pi17 ? n32 : n25674;
  assign n25676 = pi16 ? n32 : n25675;
  assign n25677 = pi15 ? n25672 : n25676;
  assign n25678 = pi14 ? n25668 : n25677;
  assign n25679 = pi20 ? n246 : ~n428;
  assign n25680 = pi19 ? n25679 : n32;
  assign n25681 = pi18 ? n32 : n25680;
  assign n25682 = pi17 ? n32 : n25681;
  assign n25683 = pi16 ? n32 : n25682;
  assign n25684 = pi15 ? n23859 : n25683;
  assign n25685 = pi14 ? n25684 : n22261;
  assign n25686 = pi13 ? n25678 : n25685;
  assign n25687 = pi12 ? n25663 : n25686;
  assign n25688 = pi11 ? n25654 : n25687;
  assign n25689 = pi10 ? n25644 : n25688;
  assign n25690 = pi09 ? n32 : n25689;
  assign n25691 = pi14 ? n32 : n17578;
  assign n25692 = pi13 ? n32 : n25691;
  assign n25693 = pi15 ? n17435 : n32;
  assign n25694 = pi14 ? n17435 : n25693;
  assign n25695 = pi14 ? n25557 : n25563;
  assign n25696 = pi13 ? n25694 : n25695;
  assign n25697 = pi12 ? n25692 : n25696;
  assign n25698 = pi14 ? n16832 : n25634;
  assign n25699 = pi13 ? n25632 : n25698;
  assign n25700 = pi20 ? n518 : ~n339;
  assign n25701 = pi19 ? n32 : n25700;
  assign n25702 = pi18 ? n32 : n25701;
  assign n25703 = pi17 ? n32 : n25702;
  assign n25704 = pi16 ? n32 : n25703;
  assign n25705 = pi19 ? n32 : n6420;
  assign n25706 = pi18 ? n32 : n25705;
  assign n25707 = pi17 ? n32 : n25706;
  assign n25708 = pi16 ? n32 : n25707;
  assign n25709 = pi15 ? n25704 : n25708;
  assign n25710 = pi19 ? n32 : n13074;
  assign n25711 = pi18 ? n32 : n25710;
  assign n25712 = pi17 ? n32 : n25711;
  assign n25713 = pi16 ? n32 : n25712;
  assign n25714 = pi15 ? n25713 : n16832;
  assign n25715 = pi14 ? n25709 : n25714;
  assign n25716 = pi14 ? n25385 : n16899;
  assign n25717 = pi13 ? n25715 : n25716;
  assign n25718 = pi12 ? n25699 : n25717;
  assign n25719 = pi11 ? n25697 : n25718;
  assign n25720 = pi14 ? n25640 : n24874;
  assign n25721 = pi15 ? n16606 : n24572;
  assign n25722 = pi14 ? n24695 : n25721;
  assign n25723 = pi13 ? n25720 : n25722;
  assign n25724 = pi15 ? n16308 : n24504;
  assign n25725 = pi14 ? n24237 : n25724;
  assign n25726 = pi15 ? n16319 : n23725;
  assign n25727 = pi14 ? n24991 : n25726;
  assign n25728 = pi13 ? n25725 : n25727;
  assign n25729 = pi12 ? n25723 : n25728;
  assign n25730 = pi14 ? n25657 : n24838;
  assign n25731 = pi15 ? n24838 : n15255;
  assign n25732 = pi19 ? n208 : ~n2614;
  assign n25733 = pi18 ? n32 : n25732;
  assign n25734 = pi17 ? n32 : n25733;
  assign n25735 = pi16 ? n32 : n25734;
  assign n25736 = pi15 ? n25735 : n25247;
  assign n25737 = pi14 ? n25731 : n25736;
  assign n25738 = pi13 ? n25730 : n25737;
  assign n25739 = pi14 ? n25684 : n14790;
  assign n25740 = pi13 ? n25678 : n25739;
  assign n25741 = pi12 ? n25738 : n25740;
  assign n25742 = pi11 ? n25729 : n25741;
  assign n25743 = pi10 ? n25719 : n25742;
  assign n25744 = pi09 ? n32 : n25743;
  assign n25745 = pi08 ? n25690 : n25744;
  assign n25746 = pi19 ? n32 : n662;
  assign n25747 = pi18 ? n32 : n25746;
  assign n25748 = pi17 ? n32 : n25747;
  assign n25749 = pi16 ? n32 : n25748;
  assign n25750 = pi15 ? n32 : n25749;
  assign n25751 = pi14 ? n32 : n25750;
  assign n25752 = pi13 ? n32 : n25751;
  assign n25753 = pi15 ? n17435 : n25749;
  assign n25754 = pi14 ? n25753 : n32;
  assign n25755 = pi14 ? n17271 : n17121;
  assign n25756 = pi13 ? n25754 : n25755;
  assign n25757 = pi12 ? n25752 : n25756;
  assign n25758 = pi15 ? n17121 : n25563;
  assign n25759 = pi14 ? n25758 : n25563;
  assign n25760 = pi19 ? n32 : n13667;
  assign n25761 = pi18 ? n32 : n25760;
  assign n25762 = pi17 ? n32 : n25761;
  assign n25763 = pi16 ? n32 : n25762;
  assign n25764 = pi14 ? n25763 : n16984;
  assign n25765 = pi13 ? n25759 : n25764;
  assign n25766 = pi14 ? n25763 : n16832;
  assign n25767 = pi15 ? n25384 : n16973;
  assign n25768 = pi14 ? n25385 : n25767;
  assign n25769 = pi13 ? n25766 : n25768;
  assign n25770 = pi12 ? n25765 : n25769;
  assign n25771 = pi11 ? n25757 : n25770;
  assign n25772 = pi15 ? n17002 : n16899;
  assign n25773 = pi14 ? n25772 : n16837;
  assign n25774 = pi15 ? n16786 : n16606;
  assign n25775 = pi15 ? n16606 : n24367;
  assign n25776 = pi14 ? n25774 : n25775;
  assign n25777 = pi13 ? n25773 : n25776;
  assign n25778 = pi14 ? n24572 : n24505;
  assign n25779 = pi15 ? n16105 : n24247;
  assign n25780 = pi14 ? n24991 : n25779;
  assign n25781 = pi13 ? n25778 : n25780;
  assign n25782 = pi12 ? n25777 : n25781;
  assign n25783 = pi15 ? n23749 : n24838;
  assign n25784 = pi14 ? n15248 : n25783;
  assign n25785 = pi14 ? n25658 : n24612;
  assign n25786 = pi13 ? n25784 : n25785;
  assign n25787 = pi19 ? n349 : ~n617;
  assign n25788 = pi18 ? n32 : n25787;
  assign n25789 = pi17 ? n32 : n25788;
  assign n25790 = pi16 ? n32 : n25789;
  assign n25791 = pi15 ? n25790 : n25247;
  assign n25792 = pi15 ? n25001 : n23094;
  assign n25793 = pi14 ? n25791 : n25792;
  assign n25794 = pi18 ? n32 : n25609;
  assign n25795 = pi17 ? n32 : n25794;
  assign n25796 = pi16 ? n32 : n25795;
  assign n25797 = pi15 ? n25796 : n22633;
  assign n25798 = pi15 ? n14606 : n14790;
  assign n25799 = pi14 ? n25797 : n25798;
  assign n25800 = pi13 ? n25793 : n25799;
  assign n25801 = pi12 ? n25786 : n25800;
  assign n25802 = pi11 ? n25782 : n25801;
  assign n25803 = pi10 ? n25771 : n25802;
  assign n25804 = pi09 ? n32 : n25803;
  assign n25805 = pi15 ? n17336 : n32;
  assign n25806 = pi14 ? n17336 : n25805;
  assign n25807 = pi13 ? n25806 : n25755;
  assign n25808 = pi12 ? n32 : n25807;
  assign n25809 = pi14 ? n25758 : n25630;
  assign n25810 = pi13 ? n25809 : n25764;
  assign n25811 = pi19 ? n32 : n21154;
  assign n25812 = pi18 ? n32 : n25811;
  assign n25813 = pi17 ? n32 : n25812;
  assign n25814 = pi16 ? n32 : n25813;
  assign n25815 = pi15 ? n25814 : n25763;
  assign n25816 = pi15 ? n25763 : n16832;
  assign n25817 = pi14 ? n25815 : n25816;
  assign n25818 = pi15 ? n15847 : n32;
  assign n25819 = pi14 ? n25502 : n25818;
  assign n25820 = pi13 ? n25817 : n25819;
  assign n25821 = pi12 ? n25810 : n25820;
  assign n25822 = pi11 ? n25808 : n25821;
  assign n25823 = pi15 ? n16973 : n16899;
  assign n25824 = pi14 ? n25823 : n25138;
  assign n25825 = pi15 ? n16786 : n16601;
  assign n25826 = pi14 ? n25825 : n24498;
  assign n25827 = pi13 ? n25824 : n25826;
  assign n25828 = pi15 ? n24237 : n24572;
  assign n25829 = pi15 ? n24572 : n24712;
  assign n25830 = pi14 ? n25828 : n25829;
  assign n25831 = pi15 ? n16105 : n24097;
  assign n25832 = pi14 ? n24289 : n25831;
  assign n25833 = pi13 ? n25830 : n25832;
  assign n25834 = pi12 ? n25827 : n25833;
  assign n25835 = pi14 ? n25658 : n24659;
  assign n25836 = pi13 ? n25784 : n25835;
  assign n25837 = pi19 ? n349 : ~n2614;
  assign n25838 = pi18 ? n32 : n25837;
  assign n25839 = pi17 ? n32 : n25838;
  assign n25840 = pi16 ? n32 : n25839;
  assign n25841 = pi15 ? n25840 : n25247;
  assign n25842 = pi14 ? n25841 : n25088;
  assign n25843 = pi19 ? n1248 : n32;
  assign n25844 = pi18 ? n32 : n25843;
  assign n25845 = pi17 ? n32 : n25844;
  assign n25846 = pi16 ? n32 : n25845;
  assign n25847 = pi15 ? n25846 : n22633;
  assign n25848 = pi18 ? n32 : n25185;
  assign n25849 = pi17 ? n32 : n25848;
  assign n25850 = pi16 ? n32 : n25849;
  assign n25851 = pi15 ? n25850 : n14790;
  assign n25852 = pi14 ? n25847 : n25851;
  assign n25853 = pi13 ? n25842 : n25852;
  assign n25854 = pi12 ? n25836 : n25853;
  assign n25855 = pi11 ? n25834 : n25854;
  assign n25856 = pi10 ? n25822 : n25855;
  assign n25857 = pi09 ? n32 : n25856;
  assign n25858 = pi08 ? n25804 : n25857;
  assign n25859 = pi07 ? n25745 : n25858;
  assign n25860 = pi06 ? n25624 : n25859;
  assign n25861 = pi15 ? n32 : n17336;
  assign n25862 = pi14 ? n25861 : n17261;
  assign n25863 = pi13 ? n25806 : n25862;
  assign n25864 = pi12 ? n32 : n25863;
  assign n25865 = pi15 ? n17261 : n17435;
  assign n25866 = pi14 ? n25865 : n25693;
  assign n25867 = pi15 ? n25556 : n25563;
  assign n25868 = pi14 ? n32 : n25867;
  assign n25869 = pi13 ? n25866 : n25868;
  assign n25870 = pi14 ? n16392 : n17039;
  assign n25871 = pi13 ? n25817 : n25870;
  assign n25872 = pi12 ? n25869 : n25871;
  assign n25873 = pi11 ? n25864 : n25872;
  assign n25874 = pi15 ? n17039 : n16899;
  assign n25875 = pi14 ? n25874 : n25138;
  assign n25876 = pi15 ? n16655 : n16452;
  assign n25877 = pi14 ? n24627 : n25876;
  assign n25878 = pi13 ? n25875 : n25877;
  assign n25879 = pi15 ? n24495 : n24367;
  assign n25880 = pi15 ? n24572 : n25319;
  assign n25881 = pi14 ? n25879 : n25880;
  assign n25882 = pi14 ? n25167 : n24383;
  assign n25883 = pi13 ? n25881 : n25882;
  assign n25884 = pi12 ? n25878 : n25883;
  assign n25885 = pi14 ? n24295 : n23749;
  assign n25886 = pi18 ? n32 : n18474;
  assign n25887 = pi17 ? n32 : n25886;
  assign n25888 = pi16 ? n32 : n25887;
  assign n25889 = pi15 ? n23749 : n25888;
  assign n25890 = pi14 ? n25889 : n25660;
  assign n25891 = pi13 ? n25885 : n25890;
  assign n25892 = pi14 ? n15119 : n25088;
  assign n25893 = pi14 ? n22347 : n23679;
  assign n25894 = pi13 ? n25892 : n25893;
  assign n25895 = pi12 ? n25891 : n25894;
  assign n25896 = pi11 ? n25884 : n25895;
  assign n25897 = pi10 ? n25873 : n25896;
  assign n25898 = pi09 ? n32 : n25897;
  assign n25899 = pi19 ? n32 : n21137;
  assign n25900 = pi18 ? n32 : n25899;
  assign n25901 = pi17 ? n32 : n25900;
  assign n25902 = pi16 ? n32 : n25901;
  assign n25903 = pi17 ? n32 : n24948;
  assign n25904 = pi16 ? n32 : n25903;
  assign n25905 = pi15 ? n25904 : n32;
  assign n25906 = pi14 ? n25902 : n25905;
  assign n25907 = pi15 ? n17121 : n17261;
  assign n25908 = pi14 ? n32 : n25907;
  assign n25909 = pi13 ? n25906 : n25908;
  assign n25910 = pi12 ? n32 : n25909;
  assign n25911 = pi15 ? n16804 : n25814;
  assign n25912 = pi14 ? n25911 : n25815;
  assign n25913 = pi14 ? n16832 : n32;
  assign n25914 = pi13 ? n25912 : n25913;
  assign n25915 = pi12 ? n25869 : n25914;
  assign n25916 = pi11 ? n25910 : n25915;
  assign n25917 = pi14 ? n16393 : n16392;
  assign n25918 = pi15 ? n16786 : n16452;
  assign n25919 = pi14 ? n16837 : n25918;
  assign n25920 = pi13 ? n25917 : n25919;
  assign n25921 = pi15 ? n24572 : n24367;
  assign n25922 = pi14 ? n16606 : n25921;
  assign n25923 = pi15 ? n24572 : n16308;
  assign n25924 = pi15 ? n24511 : n24382;
  assign n25925 = pi14 ? n25923 : n25924;
  assign n25926 = pi13 ? n25922 : n25925;
  assign n25927 = pi12 ? n25920 : n25926;
  assign n25928 = pi14 ? n24295 : n23933;
  assign n25929 = pi19 ? n594 : ~n1941;
  assign n25930 = pi18 ? n32 : n25929;
  assign n25931 = pi17 ? n32 : n25930;
  assign n25932 = pi16 ? n32 : n25931;
  assign n25933 = pi15 ? n23749 : n25932;
  assign n25934 = pi14 ? n25933 : n24742;
  assign n25935 = pi13 ? n25928 : n25934;
  assign n25936 = pi14 ? n15255 : n25247;
  assign n25937 = pi14 ? n22829 : n23679;
  assign n25938 = pi13 ? n25936 : n25937;
  assign n25939 = pi12 ? n25935 : n25938;
  assign n25940 = pi11 ? n25927 : n25939;
  assign n25941 = pi10 ? n25916 : n25940;
  assign n25942 = pi09 ? n32 : n25941;
  assign n25943 = pi08 ? n25898 : n25942;
  assign n25944 = pi14 ? n25904 : n25905;
  assign n25945 = pi15 ? n32 : n17431;
  assign n25946 = pi18 ? n32 : n19202;
  assign n25947 = pi17 ? n32 : n25946;
  assign n25948 = pi16 ? n32 : n25947;
  assign n25949 = pi14 ? n25945 : n25948;
  assign n25950 = pi13 ? n25944 : n25949;
  assign n25951 = pi12 ? n32 : n25950;
  assign n25952 = pi15 ? n25948 : n17336;
  assign n25953 = pi14 ? n25952 : n25805;
  assign n25954 = pi13 ? n25953 : n25755;
  assign n25955 = pi14 ? n16392 : n17188;
  assign n25956 = pi13 ? n25912 : n25955;
  assign n25957 = pi12 ? n25954 : n25956;
  assign n25958 = pi11 ? n25951 : n25957;
  assign n25959 = pi15 ? n17188 : n17039;
  assign n25960 = pi14 ? n25959 : n17039;
  assign n25961 = pi15 ? n16973 : n16837;
  assign n25962 = pi15 ? n16837 : n16601;
  assign n25963 = pi14 ? n25961 : n25962;
  assign n25964 = pi13 ? n25960 : n25963;
  assign n25965 = pi15 ? n16655 : n16606;
  assign n25966 = pi14 ? n25965 : n24367;
  assign n25967 = pi14 ? n24573 : n25924;
  assign n25968 = pi13 ? n25966 : n25967;
  assign n25969 = pi12 ? n25964 : n25968;
  assign n25970 = pi14 ? n24247 : n24257;
  assign n25971 = pi14 ? n23631 : n24909;
  assign n25972 = pi13 ? n25970 : n25971;
  assign n25973 = pi14 ? n24840 : n25247;
  assign n25974 = pi15 ? n23094 : n22437;
  assign n25975 = pi14 ? n24189 : n25974;
  assign n25976 = pi13 ? n25973 : n25975;
  assign n25977 = pi12 ? n25972 : n25976;
  assign n25978 = pi11 ? n25969 : n25977;
  assign n25979 = pi10 ? n25958 : n25978;
  assign n25980 = pi09 ? n32 : n25979;
  assign n25981 = pi19 ? n32 : n21029;
  assign n25982 = pi18 ? n32 : n25981;
  assign n25983 = pi17 ? n32 : n25982;
  assign n25984 = pi16 ? n32 : n25983;
  assign n25985 = pi19 ? n32 : n14609;
  assign n25986 = pi18 ? n32 : n25985;
  assign n25987 = pi17 ? n32 : n25986;
  assign n25988 = pi16 ? n32 : n25987;
  assign n25989 = pi15 ? n25984 : n25988;
  assign n25990 = pi15 ? n25984 : n32;
  assign n25991 = pi14 ? n25989 : n25990;
  assign n25992 = pi13 ? n25991 : n25949;
  assign n25993 = pi12 ? n32 : n25992;
  assign n25994 = pi19 ? n32 : n21486;
  assign n25995 = pi18 ? n32 : n25994;
  assign n25996 = pi17 ? n32 : n25995;
  assign n25997 = pi16 ? n32 : n25996;
  assign n25998 = pi15 ? n25997 : n16804;
  assign n25999 = pi14 ? n25998 : n16804;
  assign n26000 = pi14 ? n25763 : n17273;
  assign n26001 = pi13 ? n25999 : n26000;
  assign n26002 = pi12 ? n25954 : n26001;
  assign n26003 = pi11 ? n25993 : n26002;
  assign n26004 = pi15 ? n17188 : n17090;
  assign n26005 = pi14 ? n26004 : n17039;
  assign n26006 = pi19 ? n32 : n19773;
  assign n26007 = pi18 ? n32 : n26006;
  assign n26008 = pi17 ? n32 : n26007;
  assign n26009 = pi16 ? n32 : n26008;
  assign n26010 = pi15 ? n16899 : n26009;
  assign n26011 = pi14 ? n25874 : n26010;
  assign n26012 = pi13 ? n26005 : n26011;
  assign n26013 = pi14 ? n25774 : n16606;
  assign n26014 = pi14 ? n24573 : n24511;
  assign n26015 = pi13 ? n26013 : n26014;
  assign n26016 = pi12 ? n26012 : n26015;
  assign n26017 = pi15 ? n15834 : n16105;
  assign n26018 = pi14 ? n24382 : n26017;
  assign n26019 = pi15 ? n24256 : n23631;
  assign n26020 = pi14 ? n26019 : n24909;
  assign n26021 = pi13 ? n26018 : n26020;
  assign n26022 = pi14 ? n24840 : n25400;
  assign n26023 = pi14 ? n24747 : n25974;
  assign n26024 = pi13 ? n26022 : n26023;
  assign n26025 = pi12 ? n26021 : n26024;
  assign n26026 = pi11 ? n26016 : n26025;
  assign n26027 = pi10 ? n26003 : n26026;
  assign n26028 = pi09 ? n32 : n26027;
  assign n26029 = pi08 ? n25980 : n26028;
  assign n26030 = pi07 ? n25943 : n26029;
  assign n26031 = pi15 ? n32 : n25988;
  assign n26032 = pi14 ? n32 : n26031;
  assign n26033 = pi13 ? n32 : n26032;
  assign n26034 = pi15 ? n25988 : n32;
  assign n26035 = pi14 ? n25988 : n26034;
  assign n26036 = pi19 ? n32 : n14160;
  assign n26037 = pi18 ? n32 : n26036;
  assign n26038 = pi17 ? n32 : n26037;
  assign n26039 = pi16 ? n32 : n26038;
  assign n26040 = pi15 ? n32 : n26039;
  assign n26041 = pi15 ? n26039 : n25984;
  assign n26042 = pi14 ? n26040 : n26041;
  assign n26043 = pi13 ? n26035 : n26042;
  assign n26044 = pi12 ? n26033 : n26043;
  assign n26045 = pi15 ? n25984 : n25904;
  assign n26046 = pi14 ? n26045 : n25905;
  assign n26047 = pi15 ? n32 : n17261;
  assign n26048 = pi14 ? n26047 : n17261;
  assign n26049 = pi13 ? n26046 : n26048;
  assign n26050 = pi15 ? n17435 : n17061;
  assign n26051 = pi14 ? n25865 : n26050;
  assign n26052 = pi19 ? n32 : n22989;
  assign n26053 = pi18 ? n32 : n26052;
  assign n26054 = pi17 ? n32 : n26053;
  assign n26055 = pi16 ? n32 : n26054;
  assign n26056 = pi15 ? n26055 : n16984;
  assign n26057 = pi14 ? n26056 : n16984;
  assign n26058 = pi13 ? n26051 : n26057;
  assign n26059 = pi12 ? n26049 : n26058;
  assign n26060 = pi11 ? n26044 : n26059;
  assign n26061 = pi15 ? n16984 : n17036;
  assign n26062 = pi14 ? n26061 : n17039;
  assign n26063 = pi15 ? n32 : n16899;
  assign n26064 = pi14 ? n26063 : n25138;
  assign n26065 = pi13 ? n26062 : n26064;
  assign n26066 = pi15 ? n16601 : n24495;
  assign n26067 = pi15 ? n24495 : n16606;
  assign n26068 = pi14 ? n26066 : n26067;
  assign n26069 = pi21 ? n174 : ~n242;
  assign n26070 = pi20 ? n26069 : n32;
  assign n26071 = pi19 ? n32 : n26070;
  assign n26072 = pi18 ? n32 : n26071;
  assign n26073 = pi17 ? n32 : n26072;
  assign n26074 = pi16 ? n32 : n26073;
  assign n26075 = pi19 ? n32 : n8064;
  assign n26076 = pi18 ? n32 : n26075;
  assign n26077 = pi17 ? n32 : n26076;
  assign n26078 = pi16 ? n32 : n26077;
  assign n26079 = pi15 ? n26074 : n26078;
  assign n26080 = pi14 ? n24367 : n26079;
  assign n26081 = pi13 ? n26068 : n26080;
  assign n26082 = pi12 ? n26065 : n26081;
  assign n26083 = pi14 ? n25590 : n16105;
  assign n26084 = pi14 ? n23730 : n24170;
  assign n26085 = pi13 ? n26083 : n26084;
  assign n26086 = pi15 ? n25466 : n24612;
  assign n26087 = pi14 ? n26086 : n25247;
  assign n26088 = pi14 ? n25001 : n25974;
  assign n26089 = pi13 ? n26087 : n26088;
  assign n26090 = pi12 ? n26085 : n26089;
  assign n26091 = pi11 ? n26082 : n26090;
  assign n26092 = pi10 ? n26060 : n26091;
  assign n26093 = pi09 ? n32 : n26092;
  assign n26094 = pi18 ? n32 : n19082;
  assign n26095 = pi17 ? n32 : n26094;
  assign n26096 = pi16 ? n32 : n26095;
  assign n26097 = pi15 ? n32 : n26096;
  assign n26098 = pi14 ? n32 : n26097;
  assign n26099 = pi13 ? n32 : n26098;
  assign n26100 = pi15 ? n26096 : n32;
  assign n26101 = pi14 ? n26096 : n26100;
  assign n26102 = pi15 ? n17431 : n25984;
  assign n26103 = pi14 ? n25945 : n26102;
  assign n26104 = pi13 ? n26101 : n26103;
  assign n26105 = pi12 ? n26099 : n26104;
  assign n26106 = pi15 ? n25948 : n17298;
  assign n26107 = pi14 ? n26106 : n26050;
  assign n26108 = pi19 ? n32 : n21047;
  assign n26109 = pi18 ? n32 : n26108;
  assign n26110 = pi17 ? n32 : n26109;
  assign n26111 = pi16 ? n32 : n26110;
  assign n26112 = pi19 ? n32 : n20482;
  assign n26113 = pi18 ? n32 : n26112;
  assign n26114 = pi17 ? n32 : n26113;
  assign n26115 = pi16 ? n32 : n26114;
  assign n26116 = pi15 ? n26111 : n26115;
  assign n26117 = pi14 ? n26116 : n26115;
  assign n26118 = pi13 ? n26107 : n26117;
  assign n26119 = pi12 ? n26049 : n26118;
  assign n26120 = pi11 ? n26105 : n26119;
  assign n26121 = pi15 ? n17170 : n17090;
  assign n26122 = pi14 ? n26121 : n17090;
  assign n26123 = pi14 ? n24962 : n16974;
  assign n26124 = pi13 ? n26122 : n26123;
  assign n26125 = pi15 ? n24367 : n24572;
  assign n26126 = pi14 ? n26125 : n26079;
  assign n26127 = pi13 ? n26009 : n26126;
  assign n26128 = pi12 ? n26124 : n26127;
  assign n26129 = pi11 ? n26128 : n26090;
  assign n26130 = pi10 ? n26120 : n26129;
  assign n26131 = pi09 ? n32 : n26130;
  assign n26132 = pi08 ? n26093 : n26131;
  assign n26133 = pi15 ? n32 : n17348;
  assign n26134 = pi14 ? n32 : n26133;
  assign n26135 = pi13 ? n32 : n26134;
  assign n26136 = pi15 ? n26096 : n17348;
  assign n26137 = pi15 ? n17348 : n25904;
  assign n26138 = pi14 ? n26136 : n26137;
  assign n26139 = pi15 ? n25904 : n17428;
  assign n26140 = pi15 ? n17428 : n17348;
  assign n26141 = pi14 ? n26139 : n26140;
  assign n26142 = pi13 ? n26138 : n26141;
  assign n26143 = pi12 ? n26135 : n26142;
  assign n26144 = pi15 ? n17348 : n25988;
  assign n26145 = pi15 ? n25988 : n25984;
  assign n26146 = pi14 ? n26144 : n26145;
  assign n26147 = pi15 ? n32 : n25948;
  assign n26148 = pi14 ? n26147 : n25948;
  assign n26149 = pi13 ? n26146 : n26148;
  assign n26150 = pi20 ? n428 : n7501;
  assign n26151 = pi19 ? n32 : n26150;
  assign n26152 = pi18 ? n32 : n26151;
  assign n26153 = pi17 ? n32 : n26152;
  assign n26154 = pi16 ? n32 : n26153;
  assign n26155 = pi15 ? n25948 : n26154;
  assign n26156 = pi14 ? n26155 : n26050;
  assign n26157 = pi14 ? n25867 : n25563;
  assign n26158 = pi13 ? n26156 : n26157;
  assign n26159 = pi12 ? n26149 : n26158;
  assign n26160 = pi11 ? n26143 : n26159;
  assign n26161 = pi15 ? n17036 : n16832;
  assign n26162 = pi14 ? n25816 : n26161;
  assign n26163 = pi15 ? n32 : n17039;
  assign n26164 = pi15 ? n17039 : n16973;
  assign n26165 = pi14 ? n26163 : n26164;
  assign n26166 = pi13 ? n26162 : n26165;
  assign n26167 = pi14 ? n25138 : n25640;
  assign n26168 = pi14 ? n16520 : n24890;
  assign n26169 = pi13 ? n26167 : n26168;
  assign n26170 = pi12 ? n26166 : n26169;
  assign n26171 = pi15 ? n24712 : n24289;
  assign n26172 = pi14 ? n26171 : n16105;
  assign n26173 = pi13 ? n26172 : n26084;
  assign n26174 = pi15 ? n23094 : n14967;
  assign n26175 = pi14 ? n25001 : n26174;
  assign n26176 = pi13 ? n26087 : n26175;
  assign n26177 = pi12 ? n26173 : n26176;
  assign n26178 = pi11 ? n26170 : n26177;
  assign n26179 = pi10 ? n26160 : n26178;
  assign n26180 = pi09 ? n32 : n26179;
  assign n26181 = pi18 ? n32 : n18058;
  assign n26182 = pi17 ? n32 : n26181;
  assign n26183 = pi16 ? n32 : n26182;
  assign n26184 = pi15 ? n32 : n26183;
  assign n26185 = pi14 ? n32 : n26184;
  assign n26186 = pi13 ? n32 : n26185;
  assign n26187 = pi18 ? n32 : n18219;
  assign n26188 = pi17 ? n32 : n26187;
  assign n26189 = pi16 ? n32 : n26188;
  assign n26190 = pi15 ? n26189 : n26183;
  assign n26191 = pi15 ? n26183 : n25904;
  assign n26192 = pi14 ? n26190 : n26191;
  assign n26193 = pi13 ? n26192 : n26141;
  assign n26194 = pi12 ? n26186 : n26193;
  assign n26195 = pi15 ? n25988 : n17216;
  assign n26196 = pi14 ? n26195 : n17216;
  assign n26197 = pi13 ? n26146 : n26196;
  assign n26198 = pi19 ? n32 : n21561;
  assign n26199 = pi18 ? n32 : n26198;
  assign n26200 = pi17 ? n32 : n26199;
  assign n26201 = pi16 ? n32 : n26200;
  assign n26202 = pi15 ? n17298 : n26201;
  assign n26203 = pi14 ? n26155 : n26202;
  assign n26204 = pi13 ? n26203 : n32;
  assign n26205 = pi12 ? n26197 : n26204;
  assign n26206 = pi11 ? n26194 : n26205;
  assign n26207 = pi15 ? n26111 : n25814;
  assign n26208 = pi14 ? n25911 : n26207;
  assign n26209 = pi13 ? n26208 : n26165;
  assign n26210 = pi12 ? n26209 : n26169;
  assign n26211 = pi11 ? n26210 : n26177;
  assign n26212 = pi10 ? n26206 : n26211;
  assign n26213 = pi09 ? n32 : n26212;
  assign n26214 = pi08 ? n26180 : n26213;
  assign n26215 = pi07 ? n26132 : n26214;
  assign n26216 = pi06 ? n26030 : n26215;
  assign n26217 = pi05 ? n25860 : n26216;
  assign n26218 = pi04 ? n25373 : n26217;
  assign n26219 = pi03 ? n24156 : n26218;
  assign n26220 = pi02 ? n21540 : n26219;
  assign n26221 = pi01 ? n32 : n26220;
  assign n26222 = pi19 ? n32 : n2277;
  assign n26223 = pi18 ? n32 : n26222;
  assign n26224 = pi17 ? n32 : n26223;
  assign n26225 = pi16 ? n32 : n26224;
  assign n26226 = pi15 ? n32 : n26225;
  assign n26227 = pi14 ? n32 : n26226;
  assign n26228 = pi13 ? n32 : n26227;
  assign n26229 = pi15 ? n26225 : n17348;
  assign n26230 = pi14 ? n26225 : n26229;
  assign n26231 = pi15 ? n17348 : n26183;
  assign n26232 = pi14 ? n26231 : n26183;
  assign n26233 = pi13 ? n26230 : n26232;
  assign n26234 = pi12 ? n26228 : n26233;
  assign n26235 = pi15 ? n26183 : n17348;
  assign n26236 = pi14 ? n26235 : n32;
  assign n26237 = pi15 ? n17216 : n17056;
  assign n26238 = pi14 ? n26195 : n26237;
  assign n26239 = pi13 ? n26236 : n26238;
  assign n26240 = pi15 ? n25948 : n17061;
  assign n26241 = pi14 ? n26240 : n26201;
  assign n26242 = pi13 ? n26241 : n25755;
  assign n26243 = pi12 ? n26239 : n26242;
  assign n26244 = pi11 ? n26234 : n26243;
  assign n26245 = pi15 ? n17121 : n25556;
  assign n26246 = pi14 ? n26245 : n25563;
  assign n26247 = pi15 ? n16984 : n25763;
  assign n26248 = pi14 ? n26247 : n25633;
  assign n26249 = pi13 ? n26246 : n26248;
  assign n26250 = pi15 ? n16392 : n16837;
  assign n26251 = pi14 ? n26250 : n25640;
  assign n26252 = pi13 ? n26251 : n26168;
  assign n26253 = pi12 ? n26249 : n26252;
  assign n26254 = pi15 ? n24572 : n24289;
  assign n26255 = pi14 ? n26254 : n16105;
  assign n26256 = pi13 ? n26255 : n26084;
  assign n26257 = pi15 ? n23749 : n15518;
  assign n26258 = pi15 ? n22923 : n23340;
  assign n26259 = pi14 ? n26257 : n26258;
  assign n26260 = pi15 ? n25676 : n14967;
  assign n26261 = pi14 ? n23011 : n26260;
  assign n26262 = pi13 ? n26259 : n26261;
  assign n26263 = pi12 ? n26256 : n26262;
  assign n26264 = pi11 ? n26253 : n26263;
  assign n26265 = pi10 ? n26244 : n26264;
  assign n26266 = pi09 ? n32 : n26265;
  assign n26267 = pi18 ? n32 : n1819;
  assign n26268 = pi17 ? n32 : n26267;
  assign n26269 = pi16 ? n32 : n26268;
  assign n26270 = pi18 ? n32 : n17733;
  assign n26271 = pi17 ? n32 : n26270;
  assign n26272 = pi16 ? n32 : n26271;
  assign n26273 = pi15 ? n26269 : n26272;
  assign n26274 = pi14 ? n26269 : n26273;
  assign n26275 = pi14 ? n17348 : n26183;
  assign n26276 = pi13 ? n26274 : n26275;
  assign n26277 = pi12 ? n32 : n26276;
  assign n26278 = pi14 ? n26195 : n16852;
  assign n26279 = pi13 ? n26236 : n26278;
  assign n26280 = pi15 ? n16850 : n17056;
  assign n26281 = pi14 ? n26280 : n17056;
  assign n26282 = pi13 ? n26281 : n25755;
  assign n26283 = pi12 ? n26279 : n26282;
  assign n26284 = pi11 ? n26277 : n26283;
  assign n26285 = pi15 ? n23730 : n25331;
  assign n26286 = pi14 ? n26285 : n24170;
  assign n26287 = pi13 ? n26255 : n26286;
  assign n26288 = pi15 ? n22923 : n22728;
  assign n26289 = pi14 ? n26257 : n26288;
  assign n26290 = pi14 ? n24189 : n26260;
  assign n26291 = pi13 ? n26289 : n26290;
  assign n26292 = pi12 ? n26287 : n26291;
  assign n26293 = pi11 ? n26253 : n26292;
  assign n26294 = pi10 ? n26284 : n26293;
  assign n26295 = pi09 ? n32 : n26294;
  assign n26296 = pi08 ? n26266 : n26295;
  assign n26297 = pi15 ? n26269 : n17152;
  assign n26298 = pi14 ? n26269 : n26297;
  assign n26299 = pi15 ? n17152 : n26272;
  assign n26300 = pi14 ? n26299 : n26272;
  assign n26301 = pi13 ? n26298 : n26300;
  assign n26302 = pi12 ? n32 : n26301;
  assign n26303 = pi15 ? n26272 : n17348;
  assign n26304 = pi14 ? n26303 : n32;
  assign n26305 = pi14 ? n16851 : n16850;
  assign n26306 = pi13 ? n26304 : n26305;
  assign n26307 = pi19 ? n32 : n11145;
  assign n26308 = pi18 ? n32 : n26307;
  assign n26309 = pi17 ? n32 : n26308;
  assign n26310 = pi16 ? n32 : n26309;
  assign n26311 = pi15 ? n26310 : n17121;
  assign n26312 = pi19 ? n32 : n21699;
  assign n26313 = pi18 ? n32 : n26312;
  assign n26314 = pi17 ? n32 : n26313;
  assign n26315 = pi16 ? n32 : n26314;
  assign n26316 = pi15 ? n26315 : n25984;
  assign n26317 = pi14 ? n26311 : n26316;
  assign n26318 = pi15 ? n25904 : n25948;
  assign n26319 = pi19 ? n32 : n21637;
  assign n26320 = pi18 ? n32 : n26319;
  assign n26321 = pi17 ? n32 : n26320;
  assign n26322 = pi16 ? n32 : n26321;
  assign n26323 = pi15 ? n26322 : n25997;
  assign n26324 = pi14 ? n26318 : n26323;
  assign n26325 = pi13 ? n26317 : n26324;
  assign n26326 = pi12 ? n26306 : n26325;
  assign n26327 = pi11 ? n26302 : n26326;
  assign n26328 = pi15 ? n26201 : n25997;
  assign n26329 = pi14 ? n26328 : n25867;
  assign n26330 = pi15 ? n25763 : n16392;
  assign n26331 = pi14 ? n26247 : n26330;
  assign n26332 = pi13 ? n26329 : n26331;
  assign n26333 = pi14 ? n16392 : n25640;
  assign n26334 = pi13 ? n26333 : n26168;
  assign n26335 = pi12 ? n26332 : n26334;
  assign n26336 = pi15 ? n24572 : n16314;
  assign n26337 = pi14 ? n26336 : n24578;
  assign n26338 = pi15 ? n24256 : n23749;
  assign n26339 = pi14 ? n25331 : n26338;
  assign n26340 = pi13 ? n26337 : n26339;
  assign n26341 = pi15 ? n22923 : n23011;
  assign n26342 = pi14 ? n26257 : n26341;
  assign n26343 = pi14 ? n24189 : n26174;
  assign n26344 = pi13 ? n26342 : n26343;
  assign n26345 = pi12 ? n26340 : n26344;
  assign n26346 = pi11 ? n26335 : n26345;
  assign n26347 = pi10 ? n26327 : n26346;
  assign n26348 = pi09 ? n32 : n26347;
  assign n26349 = pi15 ? n32 : n17531;
  assign n26350 = pi14 ? n32 : n26349;
  assign n26351 = pi13 ? n32 : n26350;
  assign n26352 = pi18 ? n32 : n17714;
  assign n26353 = pi17 ? n32 : n26352;
  assign n26354 = pi16 ? n32 : n26353;
  assign n26355 = pi14 ? n26354 : n26297;
  assign n26356 = pi13 ? n26355 : n26300;
  assign n26357 = pi12 ? n26351 : n26356;
  assign n26358 = pi13 ? n26236 : n26305;
  assign n26359 = pi14 ? n26318 : n26328;
  assign n26360 = pi13 ? n26317 : n26359;
  assign n26361 = pi12 ? n26358 : n26360;
  assign n26362 = pi11 ? n26357 : n26361;
  assign n26363 = pi15 ? n26201 : n25814;
  assign n26364 = pi14 ? n26363 : n25867;
  assign n26365 = pi13 ? n26364 : n26248;
  assign n26366 = pi12 ? n26365 : n26252;
  assign n26367 = pi15 ? n16319 : n23730;
  assign n26368 = pi14 ? n26336 : n26367;
  assign n26369 = pi15 ? n25331 : n24256;
  assign n26370 = pi14 ? n26369 : n26338;
  assign n26371 = pi13 ? n26368 : n26370;
  assign n26372 = pi14 ? n15518 : n26341;
  assign n26373 = pi15 ? n23094 : n21928;
  assign n26374 = pi14 ? n24189 : n26373;
  assign n26375 = pi13 ? n26372 : n26374;
  assign n26376 = pi12 ? n26371 : n26375;
  assign n26377 = pi11 ? n26366 : n26376;
  assign n26378 = pi10 ? n26362 : n26377;
  assign n26379 = pi09 ? n32 : n26378;
  assign n26380 = pi08 ? n26348 : n26379;
  assign n26381 = pi07 ? n26296 : n26380;
  assign n26382 = pi15 ? n32 : n17514;
  assign n26383 = pi14 ? n32 : n26382;
  assign n26384 = pi13 ? n32 : n26383;
  assign n26385 = pi14 ? n17514 : n17348;
  assign n26386 = pi20 ? n32 : n20353;
  assign n26387 = pi19 ? n32 : n26386;
  assign n26388 = pi18 ? n32 : n26387;
  assign n26389 = pi17 ? n32 : n26388;
  assign n26390 = pi16 ? n32 : n26389;
  assign n26391 = pi13 ? n26385 : n26390;
  assign n26392 = pi12 ? n26384 : n26391;
  assign n26393 = pi15 ? n26390 : n17152;
  assign n26394 = pi15 ? n17152 : n17205;
  assign n26395 = pi14 ? n26393 : n26394;
  assign n26396 = pi15 ? n17205 : n17286;
  assign n26397 = pi19 ? n32 : n7795;
  assign n26398 = pi18 ? n32 : n26397;
  assign n26399 = pi17 ? n32 : n26398;
  assign n26400 = pi16 ? n32 : n26399;
  assign n26401 = pi15 ? n17286 : n26400;
  assign n26402 = pi14 ? n26396 : n26401;
  assign n26403 = pi13 ? n26395 : n26402;
  assign n26404 = pi15 ? n26315 : n25988;
  assign n26405 = pi14 ? n26400 : n26404;
  assign n26406 = pi14 ? n25904 : n26323;
  assign n26407 = pi13 ? n26405 : n26406;
  assign n26408 = pi12 ? n26403 : n26407;
  assign n26409 = pi11 ? n26392 : n26408;
  assign n26410 = pi15 ? n24572 : n24382;
  assign n26411 = pi15 ? n24247 : n25331;
  assign n26412 = pi14 ? n26410 : n26411;
  assign n26413 = pi15 ? n24097 : n24256;
  assign n26414 = pi14 ? n26413 : n24170;
  assign n26415 = pi13 ? n26412 : n26414;
  assign n26416 = pi14 ? n15255 : n23011;
  assign n26417 = pi14 ? n23443 : n21853;
  assign n26418 = pi13 ? n26416 : n26417;
  assign n26419 = pi12 ? n26415 : n26418;
  assign n26420 = pi11 ? n26335 : n26419;
  assign n26421 = pi10 ? n26409 : n26420;
  assign n26422 = pi09 ? n32 : n26421;
  assign n26423 = pi18 ? n32 : n17848;
  assign n26424 = pi17 ? n32 : n26423;
  assign n26425 = pi16 ? n32 : n26424;
  assign n26426 = pi18 ? n32 : n312;
  assign n26427 = pi17 ? n32 : n26426;
  assign n26428 = pi16 ? n32 : n26427;
  assign n26429 = pi15 ? n26425 : n26428;
  assign n26430 = pi14 ? n32 : n26429;
  assign n26431 = pi13 ? n32 : n26430;
  assign n26432 = pi15 ? n26428 : n17348;
  assign n26433 = pi14 ? n26432 : n17348;
  assign n26434 = pi15 ? n17152 : n26390;
  assign n26435 = pi14 ? n17152 : n26434;
  assign n26436 = pi13 ? n26433 : n26435;
  assign n26437 = pi12 ? n26431 : n26436;
  assign n26438 = pi14 ? n26393 : n17152;
  assign n26439 = pi15 ? n17152 : n17286;
  assign n26440 = pi14 ? n26439 : n26401;
  assign n26441 = pi13 ? n26438 : n26440;
  assign n26442 = pi12 ? n26441 : n26407;
  assign n26443 = pi11 ? n26437 : n26442;
  assign n26444 = pi13 ? n26329 : n26248;
  assign n26445 = pi15 ? n16837 : n16520;
  assign n26446 = pi14 ? n26250 : n26445;
  assign n26447 = pi15 ? n16520 : n16452;
  assign n26448 = pi14 ? n26447 : n24890;
  assign n26449 = pi13 ? n26446 : n26448;
  assign n26450 = pi12 ? n26444 : n26449;
  assign n26451 = pi15 ? n16377 : n24382;
  assign n26452 = pi14 ? n26451 : n26411;
  assign n26453 = pi15 ? n23933 : n15518;
  assign n26454 = pi14 ? n26413 : n26453;
  assign n26455 = pi13 ? n26452 : n26454;
  assign n26456 = pi12 ? n26455 : n26418;
  assign n26457 = pi11 ? n26450 : n26456;
  assign n26458 = pi10 ? n26443 : n26457;
  assign n26459 = pi09 ? n32 : n26458;
  assign n26460 = pi08 ? n26422 : n26459;
  assign n26461 = pi17 ? n32 : n23052;
  assign n26462 = pi16 ? n32 : n26461;
  assign n26463 = pi15 ? n26462 : n17465;
  assign n26464 = pi14 ? n32 : n26463;
  assign n26465 = pi13 ? n32 : n26464;
  assign n26466 = pi15 ? n17465 : n17152;
  assign n26467 = pi14 ? n26466 : n17152;
  assign n26468 = pi13 ? n26467 : n26435;
  assign n26469 = pi12 ? n26465 : n26468;
  assign n26470 = pi15 ? n17152 : n17348;
  assign n26471 = pi14 ? n26393 : n26470;
  assign n26472 = pi15 ? n26272 : n17286;
  assign n26473 = pi14 ? n26472 : n17286;
  assign n26474 = pi13 ? n26471 : n26473;
  assign n26475 = pi15 ? n26400 : n25984;
  assign n26476 = pi14 ? n26400 : n26475;
  assign n26477 = pi18 ? n32 : n19209;
  assign n26478 = pi17 ? n32 : n26477;
  assign n26479 = pi16 ? n32 : n26478;
  assign n26480 = pi15 ? n26322 : n26479;
  assign n26481 = pi14 ? n25904 : n26480;
  assign n26482 = pi13 ? n26476 : n26481;
  assign n26483 = pi12 ? n26474 : n26482;
  assign n26484 = pi11 ? n26469 : n26483;
  assign n26485 = pi14 ? n25997 : n25563;
  assign n26486 = pi13 ? n26485 : n26248;
  assign n26487 = pi12 ? n26486 : n26449;
  assign n26488 = pi15 ? n24289 : n24382;
  assign n26489 = pi14 ? n26488 : n24097;
  assign n26490 = pi15 ? n23933 : n24256;
  assign n26491 = pi14 ? n26490 : n15518;
  assign n26492 = pi13 ? n26489 : n26491;
  assign n26493 = pi15 ? n15255 : n15119;
  assign n26494 = pi14 ? n26493 : n22817;
  assign n26495 = pi15 ? n23443 : n14790;
  assign n26496 = pi18 ? n32 : n25116;
  assign n26497 = pi17 ? n32 : n26496;
  assign n26498 = pi16 ? n32 : n26497;
  assign n26499 = pi15 ? n21853 : n26498;
  assign n26500 = pi14 ? n26495 : n26499;
  assign n26501 = pi13 ? n26494 : n26500;
  assign n26502 = pi12 ? n26492 : n26501;
  assign n26503 = pi11 ? n26487 : n26502;
  assign n26504 = pi10 ? n26484 : n26503;
  assign n26505 = pi09 ? n32 : n26504;
  assign n26506 = pi15 ? n26462 : n17618;
  assign n26507 = pi14 ? n32 : n26506;
  assign n26508 = pi13 ? n32 : n26507;
  assign n26509 = pi15 ? n17618 : n17278;
  assign n26510 = pi14 ? n26509 : n17278;
  assign n26511 = pi13 ? n26510 : n17278;
  assign n26512 = pi12 ? n26508 : n26511;
  assign n26513 = pi18 ? n32 : n728;
  assign n26514 = pi17 ? n32 : n26513;
  assign n26515 = pi16 ? n32 : n26514;
  assign n26516 = pi15 ? n26515 : n17348;
  assign n26517 = pi14 ? n26515 : n26516;
  assign n26518 = pi13 ? n26517 : n26473;
  assign n26519 = pi13 ? n26476 : n26406;
  assign n26520 = pi12 ? n26518 : n26519;
  assign n26521 = pi11 ? n26512 : n26520;
  assign n26522 = pi14 ? n26447 : n16457;
  assign n26523 = pi13 ? n26446 : n26522;
  assign n26524 = pi12 ? n26486 : n26523;
  assign n26525 = pi14 ? n23679 : n26499;
  assign n26526 = pi13 ? n26494 : n26525;
  assign n26527 = pi12 ? n26492 : n26526;
  assign n26528 = pi11 ? n26524 : n26527;
  assign n26529 = pi10 ? n26521 : n26528;
  assign n26530 = pi09 ? n32 : n26529;
  assign n26531 = pi08 ? n26505 : n26530;
  assign n26532 = pi07 ? n26460 : n26531;
  assign n26533 = pi06 ? n26381 : n26532;
  assign n26534 = pi14 ? n32 : n17619;
  assign n26535 = pi13 ? n32 : n26534;
  assign n26536 = pi12 ? n32 : n26535;
  assign n26537 = pi15 ? n26515 : n32;
  assign n26538 = pi14 ? n26515 : n26537;
  assign n26539 = pi14 ? n26269 : n17286;
  assign n26540 = pi13 ? n26538 : n26539;
  assign n26541 = pi14 ? n26400 : n26145;
  assign n26542 = pi14 ? n25904 : n26328;
  assign n26543 = pi13 ? n26541 : n26542;
  assign n26544 = pi12 ? n26540 : n26543;
  assign n26545 = pi11 ? n26536 : n26544;
  assign n26546 = pi15 ? n25997 : n25556;
  assign n26547 = pi14 ? n26546 : n25630;
  assign n26548 = pi15 ? n25708 : n16485;
  assign n26549 = pi14 ? n26548 : n25633;
  assign n26550 = pi13 ? n26547 : n26549;
  assign n26551 = pi14 ? n16837 : n24880;
  assign n26552 = pi14 ? n16452 : n26451;
  assign n26553 = pi13 ? n26551 : n26552;
  assign n26554 = pi12 ? n26550 : n26553;
  assign n26555 = pi15 ? n24289 : n24247;
  assign n26556 = pi14 ? n26555 : n23933;
  assign n26557 = pi15 ? n23933 : n23160;
  assign n26558 = pi14 ? n26557 : n23761;
  assign n26559 = pi13 ? n26556 : n26558;
  assign n26560 = pi14 ? n24747 : n22931;
  assign n26561 = pi15 ? n14790 : n22958;
  assign n26562 = pi14 ? n26561 : n14389;
  assign n26563 = pi13 ? n26560 : n26562;
  assign n26564 = pi12 ? n26559 : n26563;
  assign n26565 = pi11 ? n26554 : n26564;
  assign n26566 = pi10 ? n26545 : n26565;
  assign n26567 = pi09 ? n32 : n26566;
  assign n26568 = pi14 ? n32 : n17443;
  assign n26569 = pi13 ? n32 : n26568;
  assign n26570 = pi12 ? n32 : n26569;
  assign n26571 = pi15 ? n17278 : n26515;
  assign n26572 = pi14 ? n26571 : n26537;
  assign n26573 = pi13 ? n26572 : n26539;
  assign n26574 = pi12 ? n26573 : n26543;
  assign n26575 = pi11 ? n26570 : n26574;
  assign n26576 = pi15 ? n23484 : n23160;
  assign n26577 = pi14 ? n26576 : n23761;
  assign n26578 = pi13 ? n26556 : n26577;
  assign n26579 = pi15 ? n14606 : n22958;
  assign n26580 = pi15 ? n14389 : n14394;
  assign n26581 = pi14 ? n26579 : n26580;
  assign n26582 = pi13 ? n26560 : n26581;
  assign n26583 = pi12 ? n26578 : n26582;
  assign n26584 = pi11 ? n26554 : n26583;
  assign n26585 = pi10 ? n26575 : n26584;
  assign n26586 = pi09 ? n32 : n26585;
  assign n26587 = pi08 ? n26567 : n26586;
  assign n26588 = pi18 ? n32 : n17843;
  assign n26589 = pi17 ? n32 : n26588;
  assign n26590 = pi16 ? n32 : n26589;
  assign n26591 = pi15 ? n32 : n26590;
  assign n26592 = pi14 ? n32 : n26591;
  assign n26593 = pi13 ? n32 : n26592;
  assign n26594 = pi12 ? n32 : n26593;
  assign n26595 = pi14 ? n26269 : n26401;
  assign n26596 = pi13 ? n26572 : n26595;
  assign n26597 = pi14 ? n25904 : n26201;
  assign n26598 = pi13 ? n26541 : n26597;
  assign n26599 = pi12 ? n26596 : n26598;
  assign n26600 = pi11 ? n26594 : n26599;
  assign n26601 = pi14 ? n26548 : n16838;
  assign n26602 = pi13 ? n26547 : n26601;
  assign n26603 = pi13 ? n25919 : n26552;
  assign n26604 = pi12 ? n26602 : n26603;
  assign n26605 = pi15 ? n16314 : n24247;
  assign n26606 = pi14 ? n26605 : n23933;
  assign n26607 = pi14 ? n24840 : n23761;
  assign n26608 = pi13 ? n26606 : n26607;
  assign n26609 = pi14 ? n24189 : n15123;
  assign n26610 = pi15 ? n14973 : n22958;
  assign n26611 = pi14 ? n26610 : n26580;
  assign n26612 = pi13 ? n26609 : n26611;
  assign n26613 = pi12 ? n26608 : n26612;
  assign n26614 = pi11 ? n26604 : n26613;
  assign n26615 = pi10 ? n26600 : n26614;
  assign n26616 = pi09 ? n32 : n26615;
  assign n26617 = pi14 ? n25521 : n26451;
  assign n26618 = pi13 ? n25919 : n26617;
  assign n26619 = pi12 ? n26602 : n26618;
  assign n26620 = pi19 ? n594 : ~n813;
  assign n26621 = pi18 ? n32 : n26620;
  assign n26622 = pi17 ? n32 : n26621;
  assign n26623 = pi16 ? n32 : n26622;
  assign n26624 = pi15 ? n23933 : n26623;
  assign n26625 = pi14 ? n26605 : n26624;
  assign n26626 = pi13 ? n26625 : n26607;
  assign n26627 = pi14 ? n24189 : n22635;
  assign n26628 = pi14 ? n26610 : n14394;
  assign n26629 = pi13 ? n26627 : n26628;
  assign n26630 = pi12 ? n26626 : n26629;
  assign n26631 = pi11 ? n26619 : n26630;
  assign n26632 = pi10 ? n26600 : n26631;
  assign n26633 = pi09 ? n32 : n26632;
  assign n26634 = pi08 ? n26616 : n26633;
  assign n26635 = pi07 ? n26587 : n26634;
  assign n26636 = pi15 ? n26515 : n26269;
  assign n26637 = pi14 ? n26571 : n26636;
  assign n26638 = pi13 ? n26637 : n26595;
  assign n26639 = pi14 ? n26400 : n25984;
  assign n26640 = pi15 ? n25948 : n26322;
  assign n26641 = pi14 ? n26640 : n26201;
  assign n26642 = pi13 ? n26639 : n26641;
  assign n26643 = pi12 ? n26638 : n26642;
  assign n26644 = pi11 ? n26536 : n26643;
  assign n26645 = pi15 ? n25997 : n25563;
  assign n26646 = pi14 ? n26645 : n25815;
  assign n26647 = pi14 ? n25816 : n16838;
  assign n26648 = pi13 ? n26646 : n26647;
  assign n26649 = pi15 ? n16837 : n26009;
  assign n26650 = pi14 ? n26649 : n26447;
  assign n26651 = pi15 ? n16452 : n16308;
  assign n26652 = pi14 ? n26651 : n16314;
  assign n26653 = pi13 ? n26650 : n26652;
  assign n26654 = pi12 ? n26648 : n26653;
  assign n26655 = pi15 ? n24289 : n24097;
  assign n26656 = pi15 ? n23933 : n23484;
  assign n26657 = pi14 ? n26655 : n26656;
  assign n26658 = pi14 ? n24840 : n15255;
  assign n26659 = pi13 ? n26657 : n26658;
  assign n26660 = pi19 ? n519 : n32;
  assign n26661 = pi18 ? n32 : n26660;
  assign n26662 = pi17 ? n32 : n26661;
  assign n26663 = pi16 ? n32 : n26662;
  assign n26664 = pi15 ? n23011 : n26663;
  assign n26665 = pi15 ? n14967 : n25850;
  assign n26666 = pi14 ? n26664 : n26665;
  assign n26667 = pi21 ? n100 : ~n1939;
  assign n26668 = pi20 ? n32 : n26667;
  assign n26669 = pi19 ? n26668 : n32;
  assign n26670 = pi18 ? n32 : n26669;
  assign n26671 = pi17 ? n32 : n26670;
  assign n26672 = pi16 ? n32 : n26671;
  assign n26673 = pi15 ? n14152 : n14394;
  assign n26674 = pi14 ? n26672 : n26673;
  assign n26675 = pi13 ? n26666 : n26674;
  assign n26676 = pi12 ? n26659 : n26675;
  assign n26677 = pi11 ? n26654 : n26676;
  assign n26678 = pi10 ? n26644 : n26677;
  assign n26679 = pi09 ? n32 : n26678;
  assign n26680 = pi14 ? n26515 : n26636;
  assign n26681 = pi13 ? n26680 : n26595;
  assign n26682 = pi12 ? n26681 : n26642;
  assign n26683 = pi11 ? n26570 : n26682;
  assign n26684 = pi15 ? n25814 : n25563;
  assign n26685 = pi14 ? n26684 : n25815;
  assign n26686 = pi14 ? n16832 : n16838;
  assign n26687 = pi13 ? n26685 : n26686;
  assign n26688 = pi12 ? n26687 : n26653;
  assign n26689 = pi15 ? n15255 : n23011;
  assign n26690 = pi14 ? n24840 : n26689;
  assign n26691 = pi13 ? n26657 : n26690;
  assign n26692 = pi15 ? n23011 : n14967;
  assign n26693 = pi14 ? n26692 : n26665;
  assign n26694 = pi15 ? n14790 : n14606;
  assign n26695 = pi15 ? n14152 : n14397;
  assign n26696 = pi14 ? n26694 : n26695;
  assign n26697 = pi13 ? n26693 : n26696;
  assign n26698 = pi12 ? n26691 : n26697;
  assign n26699 = pi11 ? n26688 : n26698;
  assign n26700 = pi10 ? n26683 : n26699;
  assign n26701 = pi09 ? n32 : n26700;
  assign n26702 = pi08 ? n26679 : n26701;
  assign n26703 = pi14 ? n26322 : n26201;
  assign n26704 = pi13 ? n26639 : n26703;
  assign n26705 = pi12 ? n26681 : n26704;
  assign n26706 = pi11 ? n26570 : n26705;
  assign n26707 = pi14 ? n16832 : n25138;
  assign n26708 = pi13 ? n26685 : n26707;
  assign n26709 = pi14 ? n26009 : n16452;
  assign n26710 = pi15 ? n16314 : n24289;
  assign n26711 = pi14 ? n16308 : n26710;
  assign n26712 = pi13 ? n26709 : n26711;
  assign n26713 = pi12 ? n26708 : n26712;
  assign n26714 = pi19 ? n594 : ~n1812;
  assign n26715 = pi18 ? n32 : n26714;
  assign n26716 = pi17 ? n32 : n26715;
  assign n26717 = pi16 ? n32 : n26716;
  assign n26718 = pi15 ? n24289 : n26717;
  assign n26719 = pi15 ? n26623 : n25888;
  assign n26720 = pi14 ? n26718 : n26719;
  assign n26721 = pi15 ? n25888 : n15260;
  assign n26722 = pi19 ? n2141 : ~n1105;
  assign n26723 = pi18 ? n32 : n26722;
  assign n26724 = pi17 ? n32 : n26723;
  assign n26725 = pi16 ? n32 : n26724;
  assign n26726 = pi15 ? n15386 : n26725;
  assign n26727 = pi14 ? n26721 : n26726;
  assign n26728 = pi13 ? n26720 : n26727;
  assign n26729 = pi14 ? n26692 : n22437;
  assign n26730 = pi15 ? n22958 : n22006;
  assign n26731 = pi15 ? n14156 : n21954;
  assign n26732 = pi14 ? n26730 : n26731;
  assign n26733 = pi13 ? n26729 : n26732;
  assign n26734 = pi12 ? n26728 : n26733;
  assign n26735 = pi11 ? n26713 : n26734;
  assign n26736 = pi10 ? n26706 : n26735;
  assign n26737 = pi09 ? n32 : n26736;
  assign n26738 = pi14 ? n16308 : n24289;
  assign n26739 = pi13 ? n26709 : n26738;
  assign n26740 = pi12 ? n26708 : n26739;
  assign n26741 = pi15 ? n23730 : n26717;
  assign n26742 = pi14 ? n26741 : n25888;
  assign n26743 = pi15 ? n25888 : n15386;
  assign n26744 = pi15 ? n15386 : n22728;
  assign n26745 = pi14 ? n26743 : n26744;
  assign n26746 = pi13 ? n26742 : n26745;
  assign n26747 = pi15 ? n22347 : n14967;
  assign n26748 = pi14 ? n26747 : n22437;
  assign n26749 = pi13 ? n26748 : n26732;
  assign n26750 = pi12 ? n26746 : n26749;
  assign n26751 = pi11 ? n26740 : n26750;
  assign n26752 = pi10 ? n26706 : n26751;
  assign n26753 = pi09 ? n32 : n26752;
  assign n26754 = pi08 ? n26737 : n26753;
  assign n26755 = pi07 ? n26702 : n26754;
  assign n26756 = pi06 ? n26635 : n26755;
  assign n26757 = pi05 ? n26533 : n26756;
  assign n26758 = pi14 ? n17286 : n26401;
  assign n26759 = pi13 ? n26680 : n26758;
  assign n26760 = pi15 ? n26400 : n25988;
  assign n26761 = pi15 ? n25984 : n17216;
  assign n26762 = pi14 ? n26760 : n26761;
  assign n26763 = pi15 ? n26322 : n26201;
  assign n26764 = pi14 ? n26763 : n26201;
  assign n26765 = pi13 ? n26762 : n26764;
  assign n26766 = pi12 ? n26759 : n26765;
  assign n26767 = pi11 ? n26570 : n26766;
  assign n26768 = pi15 ? n25563 : n25814;
  assign n26769 = pi14 ? n26768 : n25815;
  assign n26770 = pi15 ? n16899 : n24874;
  assign n26771 = pi14 ? n16832 : n26770;
  assign n26772 = pi13 ? n26769 : n26771;
  assign n26773 = pi14 ? n24504 : n24289;
  assign n26774 = pi13 ? n26709 : n26773;
  assign n26775 = pi12 ? n26772 : n26774;
  assign n26776 = pi21 ? n20130 : n32;
  assign n26777 = pi20 ? n26776 : n32;
  assign n26778 = pi19 ? n507 : n26777;
  assign n26779 = pi18 ? n32 : n26778;
  assign n26780 = pi17 ? n32 : n26779;
  assign n26781 = pi16 ? n32 : n26780;
  assign n26782 = pi15 ? n23730 : n26781;
  assign n26783 = pi15 ? n23484 : n25888;
  assign n26784 = pi14 ? n26782 : n26783;
  assign n26785 = pi14 ? n26743 : n23174;
  assign n26786 = pi13 ? n26784 : n26785;
  assign n26787 = pi15 ? n25676 : n22437;
  assign n26788 = pi15 ? n22437 : n21853;
  assign n26789 = pi14 ? n26787 : n26788;
  assign n26790 = pi14 ? n21801 : n14156;
  assign n26791 = pi13 ? n26789 : n26790;
  assign n26792 = pi12 ? n26786 : n26791;
  assign n26793 = pi11 ? n26775 : n26792;
  assign n26794 = pi10 ? n26767 : n26793;
  assign n26795 = pi09 ? n32 : n26794;
  assign n26796 = pi15 ? n26201 : n26111;
  assign n26797 = pi14 ? n26763 : n26796;
  assign n26798 = pi13 ? n26762 : n26797;
  assign n26799 = pi12 ? n26759 : n26798;
  assign n26800 = pi11 ? n26570 : n26799;
  assign n26801 = pi15 ? n25814 : n16832;
  assign n26802 = pi14 ? n26768 : n26801;
  assign n26803 = pi15 ? n16832 : n16899;
  assign n26804 = pi14 ? n26803 : n26770;
  assign n26805 = pi13 ? n26802 : n26804;
  assign n26806 = pi15 ? n26009 : n16606;
  assign n26807 = pi14 ? n26806 : n25521;
  assign n26808 = pi13 ? n26807 : n26773;
  assign n26809 = pi12 ? n26805 : n26808;
  assign n26810 = pi19 ? n507 : n7502;
  assign n26811 = pi18 ? n32 : n26810;
  assign n26812 = pi17 ? n32 : n26811;
  assign n26813 = pi16 ? n32 : n26812;
  assign n26814 = pi15 ? n23730 : n26813;
  assign n26815 = pi14 ? n26814 : n26783;
  assign n26816 = pi13 ? n26815 : n26785;
  assign n26817 = pi14 ? n25974 : n26788;
  assign n26818 = pi13 ? n26817 : n26790;
  assign n26819 = pi12 ? n26816 : n26818;
  assign n26820 = pi11 ? n26809 : n26819;
  assign n26821 = pi10 ? n26800 : n26820;
  assign n26822 = pi09 ? n32 : n26821;
  assign n26823 = pi08 ? n26795 : n26822;
  assign n26824 = pi15 ? n25984 : n17056;
  assign n26825 = pi14 ? n26760 : n26824;
  assign n26826 = pi15 ? n26201 : n25563;
  assign n26827 = pi14 ? n26763 : n26826;
  assign n26828 = pi13 ? n26825 : n26827;
  assign n26829 = pi12 ? n26759 : n26828;
  assign n26830 = pi11 ? n26570 : n26829;
  assign n26831 = pi15 ? n24874 : n16452;
  assign n26832 = pi21 ? n1939 : ~n259;
  assign n26833 = pi20 ? n26832 : n32;
  assign n26834 = pi19 ? n32 : n26833;
  assign n26835 = pi18 ? n32 : n26834;
  assign n26836 = pi17 ? n32 : n26835;
  assign n26837 = pi16 ? n32 : n26836;
  assign n26838 = pi15 ? n16452 : n26837;
  assign n26839 = pi14 ? n26831 : n26838;
  assign n26840 = pi15 ? n24289 : n23730;
  assign n26841 = pi14 ? n26837 : n26840;
  assign n26842 = pi13 ? n26839 : n26841;
  assign n26843 = pi12 ? n26805 : n26842;
  assign n26844 = pi19 ? n18741 : ~n236;
  assign n26845 = pi18 ? n32 : n26844;
  assign n26846 = pi17 ? n32 : n26845;
  assign n26847 = pi16 ? n32 : n26846;
  assign n26848 = pi15 ? n24742 : n26847;
  assign n26849 = pi14 ? n25783 : n26848;
  assign n26850 = pi19 ? n1165 : ~n617;
  assign n26851 = pi18 ? n32 : n26850;
  assign n26852 = pi17 ? n32 : n26851;
  assign n26853 = pi16 ? n32 : n26852;
  assign n26854 = pi15 ? n26853 : n15389;
  assign n26855 = pi14 ? n26854 : n23094;
  assign n26856 = pi13 ? n26849 : n26855;
  assign n26857 = pi20 ? n32 : ~n9367;
  assign n26858 = pi19 ? n26857 : n32;
  assign n26859 = pi18 ? n32 : n26858;
  assign n26860 = pi17 ? n32 : n26859;
  assign n26861 = pi16 ? n32 : n26860;
  assign n26862 = pi15 ? n21853 : n26861;
  assign n26863 = pi14 ? n25974 : n26862;
  assign n26864 = pi15 ? n14156 : n14168;
  assign n26865 = pi14 ? n21801 : n26864;
  assign n26866 = pi13 ? n26863 : n26865;
  assign n26867 = pi12 ? n26856 : n26866;
  assign n26868 = pi11 ? n26843 : n26867;
  assign n26869 = pi10 ? n26830 : n26868;
  assign n26870 = pi09 ? n32 : n26869;
  assign n26871 = pi15 ? n17152 : n26269;
  assign n26872 = pi14 ? n26515 : n26871;
  assign n26873 = pi14 ? n17286 : n26400;
  assign n26874 = pi13 ? n26872 : n26873;
  assign n26875 = pi12 ? n26874 : n26828;
  assign n26876 = pi11 ? n26570 : n26875;
  assign n26877 = pi19 ? n32 : n10879;
  assign n26878 = pi18 ? n32 : n26877;
  assign n26879 = pi17 ? n32 : n26878;
  assign n26880 = pi16 ? n32 : n26879;
  assign n26881 = pi15 ? n26880 : n16293;
  assign n26882 = pi19 ? n32 : n5597;
  assign n26883 = pi18 ? n32 : n26882;
  assign n26884 = pi17 ? n32 : n26883;
  assign n26885 = pi16 ? n32 : n26884;
  assign n26886 = pi15 ? n26885 : n16308;
  assign n26887 = pi14 ? n26881 : n26886;
  assign n26888 = pi14 ? n24504 : n26840;
  assign n26889 = pi13 ? n26887 : n26888;
  assign n26890 = pi12 ? n26805 : n26889;
  assign n26891 = pi15 ? n26853 : n22347;
  assign n26892 = pi14 ? n26891 : n23094;
  assign n26893 = pi13 ? n26849 : n26892;
  assign n26894 = pi15 ? n23094 : n14790;
  assign n26895 = pi15 ? n32 : n26861;
  assign n26896 = pi14 ? n26894 : n26895;
  assign n26897 = pi13 ? n26896 : n26865;
  assign n26898 = pi12 ? n26893 : n26897;
  assign n26899 = pi11 ? n26890 : n26898;
  assign n26900 = pi10 ? n26876 : n26899;
  assign n26901 = pi09 ? n32 : n26900;
  assign n26902 = pi08 ? n26870 : n26901;
  assign n26903 = pi07 ? n26823 : n26902;
  assign n26904 = pi15 ? n32 : n26269;
  assign n26905 = pi14 ? n26515 : n26904;
  assign n26906 = pi13 ? n26905 : n26873;
  assign n26907 = pi14 ? n26031 : n26824;
  assign n26908 = pi15 ? n32 : n25563;
  assign n26909 = pi14 ? n26201 : n26908;
  assign n26910 = pi13 ? n26907 : n26909;
  assign n26911 = pi12 ? n26906 : n26910;
  assign n26912 = pi11 ? n26570 : n26911;
  assign n26913 = pi14 ? n26768 : n16832;
  assign n26914 = pi15 ? n32 : n25384;
  assign n26915 = pi15 ? n25384 : n24874;
  assign n26916 = pi14 ? n26914 : n26915;
  assign n26917 = pi13 ? n26913 : n26916;
  assign n26918 = pi14 ? n24498 : n24504;
  assign n26919 = pi15 ? n24504 : n16105;
  assign n26920 = pi14 ? n26919 : n22818;
  assign n26921 = pi13 ? n26918 : n26920;
  assign n26922 = pi12 ? n26917 : n26921;
  assign n26923 = pi19 ? n11183 : ~n236;
  assign n26924 = pi18 ? n32 : n26923;
  assign n26925 = pi17 ? n32 : n26924;
  assign n26926 = pi16 ? n32 : n26925;
  assign n26927 = pi19 ? n11183 : ~n617;
  assign n26928 = pi18 ? n32 : n26927;
  assign n26929 = pi17 ? n32 : n26928;
  assign n26930 = pi16 ? n32 : n26929;
  assign n26931 = pi15 ? n26926 : n26930;
  assign n26932 = pi14 ? n25783 : n26931;
  assign n26933 = pi15 ? n14967 : n22347;
  assign n26934 = pi21 ? n32 : n17044;
  assign n26935 = pi20 ? n32 : n26934;
  assign n26936 = pi19 ? n26935 : n32;
  assign n26937 = pi18 ? n32 : n26936;
  assign n26938 = pi17 ? n32 : n26937;
  assign n26939 = pi16 ? n32 : n26938;
  assign n26940 = pi14 ? n26933 : n26939;
  assign n26941 = pi13 ? n26932 : n26940;
  assign n26942 = pi15 ? n14156 : n26861;
  assign n26943 = pi14 ? n14799 : n26942;
  assign n26944 = pi13 ? n26943 : n26865;
  assign n26945 = pi12 ? n26941 : n26944;
  assign n26946 = pi11 ? n26922 : n26945;
  assign n26947 = pi10 ? n26912 : n26946;
  assign n26948 = pi09 ? n32 : n26947;
  assign n26949 = pi18 ? n32 : n17834;
  assign n26950 = pi17 ? n32 : n26949;
  assign n26951 = pi16 ? n32 : n26950;
  assign n26952 = pi15 ? n26951 : n17278;
  assign n26953 = pi14 ? n32 : n26952;
  assign n26954 = pi13 ? n32 : n26953;
  assign n26955 = pi12 ? n32 : n26954;
  assign n26956 = pi11 ? n26955 : n26911;
  assign n26957 = pi19 ? n507 : n53;
  assign n26958 = pi18 ? n32 : n26957;
  assign n26959 = pi17 ? n32 : n26958;
  assign n26960 = pi16 ? n32 : n26959;
  assign n26961 = pi15 ? n32 : n26960;
  assign n26962 = pi14 ? n26919 : n26961;
  assign n26963 = pi13 ? n26918 : n26962;
  assign n26964 = pi12 ? n26917 : n26963;
  assign n26965 = pi15 ? n15255 : n15123;
  assign n26966 = pi14 ? n25783 : n26965;
  assign n26967 = pi15 ? n14967 : n24406;
  assign n26968 = pi14 ? n26967 : n23094;
  assign n26969 = pi13 ? n26966 : n26968;
  assign n26970 = pi15 ? n14790 : n32;
  assign n26971 = pi14 ? n26970 : n21801;
  assign n26972 = pi15 ? n21801 : n14156;
  assign n26973 = pi14 ? n26972 : n21558;
  assign n26974 = pi13 ? n26971 : n26973;
  assign n26975 = pi12 ? n26969 : n26974;
  assign n26976 = pi11 ? n26964 : n26975;
  assign n26977 = pi10 ? n26956 : n26976;
  assign n26978 = pi09 ? n32 : n26977;
  assign n26979 = pi08 ? n26948 : n26978;
  assign n26980 = pi20 ? n23122 : ~n141;
  assign n26981 = pi19 ? n32 : n26980;
  assign n26982 = pi18 ? n32 : n26981;
  assign n26983 = pi17 ? n32 : n26982;
  assign n26984 = pi16 ? n32 : n26983;
  assign n26985 = pi15 ? n26984 : n32;
  assign n26986 = pi14 ? n26207 : n26985;
  assign n26987 = pi19 ? n32 : n19852;
  assign n26988 = pi18 ? n32 : n26987;
  assign n26989 = pi17 ? n32 : n26988;
  assign n26990 = pi16 ? n32 : n26989;
  assign n26991 = pi15 ? n26990 : n16601;
  assign n26992 = pi14 ? n26914 : n26991;
  assign n26993 = pi13 ? n26986 : n26992;
  assign n26994 = pi15 ? n32 : n24237;
  assign n26995 = pi14 ? n26994 : n24504;
  assign n26996 = pi13 ? n26995 : n26962;
  assign n26997 = pi12 ? n26993 : n26996;
  assign n26998 = pi15 ? n24612 : n32;
  assign n26999 = pi14 ? n25783 : n26998;
  assign n27000 = pi22 ? n173 : n13584;
  assign n27001 = pi21 ? n32 : n27000;
  assign n27002 = pi20 ? n32 : n27001;
  assign n27003 = pi19 ? n27002 : n32;
  assign n27004 = pi18 ? n32 : n27003;
  assign n27005 = pi17 ? n32 : n27004;
  assign n27006 = pi16 ? n32 : n27005;
  assign n27007 = pi15 ? n21853 : n27006;
  assign n27008 = pi14 ? n27007 : n23094;
  assign n27009 = pi13 ? n26999 : n27008;
  assign n27010 = pi15 ? n14790 : n14397;
  assign n27011 = pi14 ? n27010 : n21801;
  assign n27012 = pi15 ? n20660 : n19972;
  assign n27013 = pi14 ? n26972 : n27012;
  assign n27014 = pi13 ? n27011 : n27013;
  assign n27015 = pi12 ? n27009 : n27014;
  assign n27016 = pi11 ? n26997 : n27015;
  assign n27017 = pi10 ? n26956 : n27016;
  assign n27018 = pi09 ? n32 : n27017;
  assign n27019 = pi15 ? n16953 : n32;
  assign n27020 = pi14 ? n26055 : n27019;
  assign n27021 = pi15 ? n16973 : n25384;
  assign n27022 = pi14 ? n27021 : n26991;
  assign n27023 = pi13 ? n27020 : n27022;
  assign n27024 = pi15 ? n24289 : n32;
  assign n27025 = pi14 ? n27024 : n26961;
  assign n27026 = pi13 ? n26995 : n27025;
  assign n27027 = pi12 ? n27023 : n27026;
  assign n27028 = pi15 ? n24659 : n32;
  assign n27029 = pi14 ? n25783 : n27028;
  assign n27030 = pi21 ? n32 : ~n9326;
  assign n27031 = pi20 ? n32 : n27030;
  assign n27032 = pi19 ? n27031 : n32;
  assign n27033 = pi18 ? n32 : n27032;
  assign n27034 = pi17 ? n32 : n27033;
  assign n27035 = pi16 ? n32 : n27034;
  assign n27036 = pi15 ? n27035 : n25676;
  assign n27037 = pi14 ? n27036 : n25974;
  assign n27038 = pi13 ? n27029 : n27037;
  assign n27039 = pi15 ? n21686 : n14397;
  assign n27040 = pi14 ? n27039 : n21801;
  assign n27041 = pi15 ? n21801 : n13943;
  assign n27042 = pi15 ? n20660 : n13671;
  assign n27043 = pi14 ? n27041 : n27042;
  assign n27044 = pi13 ? n27040 : n27043;
  assign n27045 = pi12 ? n27038 : n27044;
  assign n27046 = pi11 ? n27027 : n27045;
  assign n27047 = pi10 ? n26956 : n27046;
  assign n27048 = pi09 ? n32 : n27047;
  assign n27049 = pi08 ? n27018 : n27048;
  assign n27050 = pi07 ? n26979 : n27049;
  assign n27051 = pi06 ? n26903 : n27050;
  assign n27052 = pi14 ? n32 : n26509;
  assign n27053 = pi13 ? n32 : n27052;
  assign n27054 = pi12 ? n32 : n27053;
  assign n27055 = pi14 ? n26515 : n26269;
  assign n27056 = pi13 ? n27055 : n26873;
  assign n27057 = pi15 ? n32 : n26315;
  assign n27058 = pi14 ? n27057 : n17056;
  assign n27059 = pi15 ? n16984 : n25563;
  assign n27060 = pi14 ? n26201 : n27059;
  assign n27061 = pi13 ? n27058 : n27060;
  assign n27062 = pi12 ? n27056 : n27061;
  assign n27063 = pi11 ? n27054 : n27062;
  assign n27064 = pi15 ? n16953 : n16452;
  assign n27065 = pi14 ? n25814 : n27064;
  assign n27066 = pi20 ? n27030 : n32;
  assign n27067 = pi19 ? n32 : n27066;
  assign n27068 = pi18 ? n32 : n27067;
  assign n27069 = pi17 ? n32 : n27068;
  assign n27070 = pi16 ? n32 : n27069;
  assign n27071 = pi15 ? n27070 : n25384;
  assign n27072 = pi15 ? n25384 : n16601;
  assign n27073 = pi14 ? n27071 : n27072;
  assign n27074 = pi13 ? n27065 : n27073;
  assign n27075 = pi15 ? n26837 : n24504;
  assign n27076 = pi14 ? n26994 : n27075;
  assign n27077 = pi15 ? n24382 : n23250;
  assign n27078 = pi19 ? n507 : ~n10447;
  assign n27079 = pi18 ? n32 : n27078;
  assign n27080 = pi17 ? n32 : n27079;
  assign n27081 = pi16 ? n32 : n27080;
  assign n27082 = pi15 ? n23484 : n27081;
  assign n27083 = pi14 ? n27077 : n27082;
  assign n27084 = pi13 ? n27076 : n27083;
  assign n27085 = pi12 ? n27074 : n27084;
  assign n27086 = pi15 ? n24838 : n25466;
  assign n27087 = pi15 ? n24742 : n21928;
  assign n27088 = pi14 ? n27086 : n27087;
  assign n27089 = pi14 ? n25676 : n25974;
  assign n27090 = pi13 ? n27088 : n27089;
  assign n27091 = pi15 ? n21686 : n21695;
  assign n27092 = pi15 ? n21695 : n21801;
  assign n27093 = pi14 ? n27091 : n27092;
  assign n27094 = pi15 ? n14168 : n21232;
  assign n27095 = pi15 ? n21571 : n20301;
  assign n27096 = pi14 ? n27094 : n27095;
  assign n27097 = pi13 ? n27093 : n27096;
  assign n27098 = pi12 ? n27090 : n27097;
  assign n27099 = pi11 ? n27085 : n27098;
  assign n27100 = pi10 ? n27063 : n27099;
  assign n27101 = pi09 ? n32 : n27100;
  assign n27102 = pi14 ? n32 : n17278;
  assign n27103 = pi13 ? n32 : n27102;
  assign n27104 = pi12 ? n32 : n27103;
  assign n27105 = pi15 ? n25988 : n26315;
  assign n27106 = pi15 ? n17056 : n17255;
  assign n27107 = pi14 ? n27105 : n27106;
  assign n27108 = pi15 ? n26201 : n16984;
  assign n27109 = pi14 ? n27108 : n25563;
  assign n27110 = pi13 ? n27107 : n27109;
  assign n27111 = pi12 ? n27056 : n27110;
  assign n27112 = pi11 ? n27104 : n27111;
  assign n27113 = pi14 ? n25815 : n24691;
  assign n27114 = pi14 ? n27071 : n25504;
  assign n27115 = pi13 ? n27113 : n27114;
  assign n27116 = pi15 ? n24382 : n23631;
  assign n27117 = pi14 ? n27116 : n25783;
  assign n27118 = pi13 ? n27076 : n27117;
  assign n27119 = pi12 ? n27115 : n27118;
  assign n27120 = pi15 ? n24838 : n24659;
  assign n27121 = pi19 ? n11183 : ~n1105;
  assign n27122 = pi18 ? n32 : n27121;
  assign n27123 = pi17 ? n32 : n27122;
  assign n27124 = pi16 ? n32 : n27123;
  assign n27125 = pi15 ? n27124 : n21928;
  assign n27126 = pi14 ? n27120 : n27125;
  assign n27127 = pi15 ? n26939 : n25676;
  assign n27128 = pi15 ? n26939 : n21853;
  assign n27129 = pi14 ? n27127 : n27128;
  assign n27130 = pi13 ? n27126 : n27129;
  assign n27131 = pi20 ? n101 : ~n1839;
  assign n27132 = pi19 ? n27131 : n32;
  assign n27133 = pi18 ? n32 : n27132;
  assign n27134 = pi17 ? n32 : n27133;
  assign n27135 = pi16 ? n32 : n27134;
  assign n27136 = pi15 ? n21695 : n27135;
  assign n27137 = pi14 ? n27091 : n27136;
  assign n27138 = pi19 ? n17224 : n32;
  assign n27139 = pi18 ? n32 : n27138;
  assign n27140 = pi17 ? n32 : n27139;
  assign n27141 = pi16 ? n32 : n27140;
  assign n27142 = pi15 ? n14168 : n27141;
  assign n27143 = pi15 ? n21571 : n13684;
  assign n27144 = pi14 ? n27142 : n27143;
  assign n27145 = pi13 ? n27137 : n27144;
  assign n27146 = pi12 ? n27130 : n27145;
  assign n27147 = pi11 ? n27119 : n27146;
  assign n27148 = pi10 ? n27112 : n27147;
  assign n27149 = pi09 ? n32 : n27148;
  assign n27150 = pi08 ? n27101 : n27149;
  assign n27151 = pi15 ? n25988 : n17056;
  assign n27152 = pi14 ? n27151 : n17056;
  assign n27153 = pi15 ? n26201 : n25556;
  assign n27154 = pi14 ? n27153 : n26207;
  assign n27155 = pi13 ? n27152 : n27154;
  assign n27156 = pi12 ? n27056 : n27155;
  assign n27157 = pi11 ? n27104 : n27156;
  assign n27158 = pi14 ? n25815 : n27021;
  assign n27159 = pi15 ? n24874 : n24504;
  assign n27160 = pi14 ? n25384 : n27159;
  assign n27161 = pi13 ? n27158 : n27160;
  assign n27162 = pi15 ? n24289 : n23631;
  assign n27163 = pi14 ? n27162 : n23749;
  assign n27164 = pi13 ? n24504 : n27163;
  assign n27165 = pi12 ? n27161 : n27164;
  assign n27166 = pi15 ? n23749 : n24659;
  assign n27167 = pi15 ? n23011 : n23094;
  assign n27168 = pi14 ? n27166 : n27167;
  assign n27169 = pi15 ? n26498 : n22006;
  assign n27170 = pi14 ? n23094 : n27169;
  assign n27171 = pi13 ? n27168 : n27170;
  assign n27172 = pi15 ? n22006 : n21695;
  assign n27173 = pi14 ? n27172 : n14168;
  assign n27174 = pi15 ? n21490 : n21346;
  assign n27175 = pi15 ? n19972 : n19856;
  assign n27176 = pi14 ? n27174 : n27175;
  assign n27177 = pi13 ? n27173 : n27176;
  assign n27178 = pi12 ? n27171 : n27177;
  assign n27179 = pi11 ? n27165 : n27178;
  assign n27180 = pi10 ? n27157 : n27179;
  assign n27181 = pi09 ? n32 : n27180;
  assign n27182 = pi14 ? n24504 : n25590;
  assign n27183 = pi14 ? n25333 : n23749;
  assign n27184 = pi13 ? n27182 : n27183;
  assign n27185 = pi12 ? n27161 : n27184;
  assign n27186 = pi15 ? n23749 : n25247;
  assign n27187 = pi14 ? n27186 : n27167;
  assign n27188 = pi13 ? n27187 : n27170;
  assign n27189 = pi15 ? n22006 : n14397;
  assign n27190 = pi14 ? n27189 : n13943;
  assign n27191 = pi13 ? n27190 : n27176;
  assign n27192 = pi12 ? n27188 : n27191;
  assign n27193 = pi11 ? n27185 : n27192;
  assign n27194 = pi10 ? n27157 : n27193;
  assign n27195 = pi09 ? n32 : n27194;
  assign n27196 = pi08 ? n27181 : n27195;
  assign n27197 = pi07 ? n27150 : n27196;
  assign n27198 = pi15 ? n26269 : n17286;
  assign n27199 = pi14 ? n26515 : n27198;
  assign n27200 = pi15 ? n26400 : n32;
  assign n27201 = pi14 ? n17286 : n27200;
  assign n27202 = pi13 ? n27199 : n27201;
  assign n27203 = pi15 ? n17216 : n26322;
  assign n27204 = pi14 ? n26237 : n27203;
  assign n27205 = pi15 ? n32 : n26111;
  assign n27206 = pi14 ? n27205 : n26111;
  assign n27207 = pi13 ? n27204 : n27206;
  assign n27208 = pi12 ? n27202 : n27207;
  assign n27209 = pi11 ? n27104 : n27208;
  assign n27210 = pi19 ? n32 : ~n9321;
  assign n27211 = pi18 ? n32 : n27210;
  assign n27212 = pi17 ? n32 : n27211;
  assign n27213 = pi16 ? n32 : n27212;
  assign n27214 = pi15 ? n27213 : n32;
  assign n27215 = pi14 ? n27214 : n27021;
  assign n27216 = pi15 ? n26990 : n25384;
  assign n27217 = pi19 ? n32 : n20326;
  assign n27218 = pi18 ? n32 : n27217;
  assign n27219 = pi17 ? n32 : n27218;
  assign n27220 = pi16 ? n32 : n27219;
  assign n27221 = pi15 ? n27220 : n24504;
  assign n27222 = pi14 ? n27216 : n27221;
  assign n27223 = pi13 ? n27215 : n27222;
  assign n27224 = pi15 ? n24504 : n24382;
  assign n27225 = pi14 ? n24504 : n27224;
  assign n27226 = pi19 ? n1464 : ~n1941;
  assign n27227 = pi18 ? n32 : n27226;
  assign n27228 = pi17 ? n32 : n27227;
  assign n27229 = pi16 ? n32 : n27228;
  assign n27230 = pi15 ? n23749 : n27229;
  assign n27231 = pi14 ? n24170 : n27230;
  assign n27232 = pi13 ? n27225 : n27231;
  assign n27233 = pi12 ? n27223 : n27232;
  assign n27234 = pi15 ? n14580 : n25251;
  assign n27235 = pi21 ? n405 : ~n100;
  assign n27236 = pi20 ? n32 : n27235;
  assign n27237 = pi19 ? n27236 : n32;
  assign n27238 = pi18 ? n32 : n27237;
  assign n27239 = pi17 ? n32 : n27238;
  assign n27240 = pi16 ? n32 : n27239;
  assign n27241 = pi15 ? n25251 : n27240;
  assign n27242 = pi14 ? n27234 : n27241;
  assign n27243 = pi15 ? n22376 : n14394;
  assign n27244 = pi14 ? n26499 : n27243;
  assign n27245 = pi13 ? n27242 : n27244;
  assign n27246 = pi19 ? n633 : n32;
  assign n27247 = pi18 ? n32 : n27246;
  assign n27248 = pi17 ? n32 : n27247;
  assign n27249 = pi16 ? n32 : n27248;
  assign n27250 = pi15 ? n14164 : n27249;
  assign n27251 = pi14 ? n27250 : n22236;
  assign n27252 = pi15 ? n21571 : n20779;
  assign n27253 = pi15 ? n20618 : n19856;
  assign n27254 = pi14 ? n27252 : n27253;
  assign n27255 = pi13 ? n27251 : n27254;
  assign n27256 = pi12 ? n27245 : n27255;
  assign n27257 = pi11 ? n27233 : n27256;
  assign n27258 = pi10 ? n27209 : n27257;
  assign n27259 = pi09 ? n32 : n27258;
  assign n27260 = pi14 ? n17286 : n26760;
  assign n27261 = pi13 ? n27199 : n27260;
  assign n27262 = pi15 ? n25556 : n26111;
  assign n27263 = pi14 ? n27262 : n26111;
  assign n27264 = pi13 ? n27204 : n27263;
  assign n27265 = pi12 ? n27261 : n27264;
  assign n27266 = pi11 ? n27104 : n27265;
  assign n27267 = pi15 ? n26990 : n24874;
  assign n27268 = pi15 ? n25155 : n24504;
  assign n27269 = pi14 ? n27267 : n27268;
  assign n27270 = pi13 ? n27215 : n27269;
  assign n27271 = pi15 ? n24504 : n24097;
  assign n27272 = pi14 ? n24504 : n27271;
  assign n27273 = pi19 ? n1325 : ~n1941;
  assign n27274 = pi18 ? n32 : n27273;
  assign n27275 = pi17 ? n32 : n27274;
  assign n27276 = pi16 ? n32 : n27275;
  assign n27277 = pi15 ? n23749 : n27276;
  assign n27278 = pi14 ? n24170 : n27277;
  assign n27279 = pi13 ? n27272 : n27278;
  assign n27280 = pi12 ? n27270 : n27279;
  assign n27281 = pi15 ? n25251 : n25850;
  assign n27282 = pi14 ? n27234 : n27281;
  assign n27283 = pi15 ? n22376 : n21863;
  assign n27284 = pi14 ? n26498 : n27283;
  assign n27285 = pi13 ? n27282 : n27284;
  assign n27286 = pi15 ? n27249 : n13948;
  assign n27287 = pi14 ? n21552 : n27286;
  assign n27288 = pi19 ? n16625 : n32;
  assign n27289 = pi18 ? n32 : n27288;
  assign n27290 = pi17 ? n32 : n27289;
  assign n27291 = pi16 ? n32 : n27290;
  assign n27292 = pi15 ? n13671 : n27291;
  assign n27293 = pi14 ? n27292 : n13393;
  assign n27294 = pi13 ? n27287 : n27293;
  assign n27295 = pi12 ? n27285 : n27294;
  assign n27296 = pi11 ? n27280 : n27295;
  assign n27297 = pi10 ? n27266 : n27296;
  assign n27298 = pi09 ? n32 : n27297;
  assign n27299 = pi08 ? n27259 : n27298;
  assign n27300 = pi15 ? n27213 : n16973;
  assign n27301 = pi19 ? n32 : n13085;
  assign n27302 = pi18 ? n32 : n27301;
  assign n27303 = pi17 ? n32 : n27302;
  assign n27304 = pi16 ? n32 : n27303;
  assign n27305 = pi15 ? n26990 : n27304;
  assign n27306 = pi14 ? n27300 : n27305;
  assign n27307 = pi15 ? n27304 : n24874;
  assign n27308 = pi15 ? n24712 : n24504;
  assign n27309 = pi14 ? n27307 : n27308;
  assign n27310 = pi13 ? n27306 : n27309;
  assign n27311 = pi15 ? n25331 : n23933;
  assign n27312 = pi14 ? n25724 : n27311;
  assign n27313 = pi15 ? n23933 : n24838;
  assign n27314 = pi19 ? n2141 : ~n617;
  assign n27315 = pi18 ? n32 : n27314;
  assign n27316 = pi17 ? n32 : n27315;
  assign n27317 = pi16 ? n32 : n27316;
  assign n27318 = pi15 ? n27317 : n25247;
  assign n27319 = pi14 ? n27313 : n27318;
  assign n27320 = pi13 ? n27312 : n27319;
  assign n27321 = pi12 ? n27310 : n27320;
  assign n27322 = pi15 ? n25251 : n23443;
  assign n27323 = pi15 ? n22958 : n26498;
  assign n27324 = pi14 ? n27322 : n27323;
  assign n27325 = pi19 ? n624 : n32;
  assign n27326 = pi18 ? n32 : n27325;
  assign n27327 = pi17 ? n32 : n27326;
  assign n27328 = pi16 ? n32 : n27327;
  assign n27329 = pi15 ? n27328 : n21551;
  assign n27330 = pi14 ? n27169 : n27329;
  assign n27331 = pi13 ? n27324 : n27330;
  assign n27332 = pi14 ? n21552 : n13953;
  assign n27333 = pi14 ? n13684 : n32;
  assign n27334 = pi13 ? n27332 : n27333;
  assign n27335 = pi12 ? n27331 : n27334;
  assign n27336 = pi11 ? n27321 : n27335;
  assign n27337 = pi10 ? n27266 : n27336;
  assign n27338 = pi09 ? n32 : n27337;
  assign n27339 = pi15 ? n26515 : n17152;
  assign n27340 = pi14 ? n27339 : n27198;
  assign n27341 = pi15 ? n25948 : n25988;
  assign n27342 = pi14 ? n26401 : n27341;
  assign n27343 = pi13 ? n27340 : n27342;
  assign n27344 = pi15 ? n25948 : n17066;
  assign n27345 = pi14 ? n26237 : n27344;
  assign n27346 = pi13 ? n27345 : n27263;
  assign n27347 = pi12 ? n27343 : n27346;
  assign n27348 = pi11 ? n27104 : n27347;
  assign n27349 = pi15 ? n27304 : n16452;
  assign n27350 = pi14 ? n27349 : n27308;
  assign n27351 = pi13 ? n27306 : n27350;
  assign n27352 = pi19 ? n857 : ~n813;
  assign n27353 = pi18 ? n32 : n27352;
  assign n27354 = pi17 ? n32 : n27353;
  assign n27355 = pi16 ? n32 : n27354;
  assign n27356 = pi15 ? n27355 : n24742;
  assign n27357 = pi15 ? n15119 : n25247;
  assign n27358 = pi14 ? n27356 : n27357;
  assign n27359 = pi13 ? n27312 : n27358;
  assign n27360 = pi12 ? n27351 : n27359;
  assign n27361 = pi15 ? n21954 : n21551;
  assign n27362 = pi14 ? n26580 : n27361;
  assign n27363 = pi13 ? n27324 : n27362;
  assign n27364 = pi12 ? n27363 : n13955;
  assign n27365 = pi11 ? n27360 : n27364;
  assign n27366 = pi10 ? n27348 : n27365;
  assign n27367 = pi09 ? n32 : n27366;
  assign n27368 = pi08 ? n27338 : n27367;
  assign n27369 = pi07 ? n27299 : n27368;
  assign n27370 = pi06 ? n27197 : n27369;
  assign n27371 = pi05 ? n27051 : n27370;
  assign n27372 = pi04 ? n26757 : n27371;
  assign n27373 = pi14 ? n26537 : n27198;
  assign n27374 = pi14 ? n26401 : n26031;
  assign n27375 = pi13 ? n27373 : n27374;
  assign n27376 = pi15 ? n25948 : n32;
  assign n27377 = pi14 ? n26237 : n27376;
  assign n27378 = pi15 ? n26111 : n17066;
  assign n27379 = pi14 ? n27262 : n27378;
  assign n27380 = pi13 ? n27377 : n27379;
  assign n27381 = pi12 ? n27375 : n27380;
  assign n27382 = pi11 ? n27104 : n27381;
  assign n27383 = pi15 ? n24237 : n16899;
  assign n27384 = pi14 ? n27383 : n27216;
  assign n27385 = pi19 ? n32 : ~n7206;
  assign n27386 = pi18 ? n32 : n27385;
  assign n27387 = pi17 ? n32 : n27386;
  assign n27388 = pi16 ? n32 : n27387;
  assign n27389 = pi15 ? n27388 : n24640;
  assign n27390 = pi14 ? n27389 : n27308;
  assign n27391 = pi13 ? n27384 : n27390;
  assign n27392 = pi14 ? n26285 : n26338;
  assign n27393 = pi15 ? n25247 : n25001;
  assign n27394 = pi14 ? n26258 : n27393;
  assign n27395 = pi13 ? n27392 : n27394;
  assign n27396 = pi12 ? n27391 : n27395;
  assign n27397 = pi15 ? n23443 : n22958;
  assign n27398 = pi15 ? n22958 : n14389;
  assign n27399 = pi14 ? n27397 : n27398;
  assign n27400 = pi15 ? n14394 : n21954;
  assign n27401 = pi14 ? n27400 : n14164;
  assign n27402 = pi13 ? n27399 : n27401;
  assign n27403 = pi12 ? n27402 : n32;
  assign n27404 = pi11 ? n27396 : n27403;
  assign n27405 = pi10 ? n27382 : n27404;
  assign n27406 = pi09 ? n32 : n27405;
  assign n27407 = pi19 ? n32 : n20132;
  assign n27408 = pi18 ? n32 : n27407;
  assign n27409 = pi17 ? n32 : n27408;
  assign n27410 = pi16 ? n32 : n27409;
  assign n27411 = pi15 ? n27410 : n25384;
  assign n27412 = pi14 ? n27383 : n27411;
  assign n27413 = pi21 ? n1392 : ~n140;
  assign n27414 = pi20 ? n27413 : n32;
  assign n27415 = pi19 ? n32 : n27414;
  assign n27416 = pi18 ? n32 : n27415;
  assign n27417 = pi17 ? n32 : n27416;
  assign n27418 = pi16 ? n32 : n27417;
  assign n27419 = pi15 ? n24712 : n27418;
  assign n27420 = pi14 ? n27389 : n27419;
  assign n27421 = pi13 ? n27412 : n27420;
  assign n27422 = pi22 ? n65 : ~n34;
  assign n27423 = pi21 ? n27422 : n32;
  assign n27424 = pi20 ? n27423 : n32;
  assign n27425 = pi19 ? n32 : n27424;
  assign n27426 = pi18 ? n32 : n27425;
  assign n27427 = pi17 ? n32 : n27426;
  assign n27428 = pi16 ? n32 : n27427;
  assign n27429 = pi15 ? n27428 : n25331;
  assign n27430 = pi14 ? n27429 : n26338;
  assign n27431 = pi15 ? n25247 : n23443;
  assign n27432 = pi14 ? n26258 : n27431;
  assign n27433 = pi13 ? n27430 : n27432;
  assign n27434 = pi12 ? n27421 : n27433;
  assign n27435 = pi15 ? n22437 : n22958;
  assign n27436 = pi14 ? n27435 : n27398;
  assign n27437 = pi13 ? n27436 : n14406;
  assign n27438 = pi12 ? n27437 : n32;
  assign n27439 = pi11 ? n27434 : n27438;
  assign n27440 = pi10 ? n27382 : n27439;
  assign n27441 = pi09 ? n32 : n27440;
  assign n27442 = pi08 ? n27406 : n27441;
  assign n27443 = pi15 ? n26479 : n32;
  assign n27444 = pi14 ? n17216 : n27443;
  assign n27445 = pi15 ? n26111 : n17039;
  assign n27446 = pi14 ? n26111 : n27445;
  assign n27447 = pi13 ? n27444 : n27446;
  assign n27448 = pi12 ? n27375 : n27447;
  assign n27449 = pi11 ? n27104 : n27448;
  assign n27450 = pi15 ? n16837 : n16899;
  assign n27451 = pi15 ? n27410 : n16606;
  assign n27452 = pi14 ? n27450 : n27451;
  assign n27453 = pi15 ? n24700 : n24640;
  assign n27454 = pi15 ? n16308 : n23730;
  assign n27455 = pi14 ? n27453 : n27454;
  assign n27456 = pi13 ? n27452 : n27455;
  assign n27457 = pi15 ? n24097 : n25331;
  assign n27458 = pi14 ? n27457 : n26019;
  assign n27459 = pi19 ? n1818 : ~n617;
  assign n27460 = pi18 ? n32 : n27459;
  assign n27461 = pi17 ? n32 : n27460;
  assign n27462 = pi16 ? n32 : n27461;
  assign n27463 = pi19 ? n1325 : ~n617;
  assign n27464 = pi18 ? n32 : n27463;
  assign n27465 = pi17 ? n32 : n27464;
  assign n27466 = pi16 ? n32 : n27465;
  assign n27467 = pi15 ? n27462 : n27466;
  assign n27468 = pi19 ? n750 : n32;
  assign n27469 = pi18 ? n32 : n27468;
  assign n27470 = pi17 ? n32 : n27469;
  assign n27471 = pi16 ? n32 : n27470;
  assign n27472 = pi15 ? n25247 : n27471;
  assign n27473 = pi14 ? n27467 : n27472;
  assign n27474 = pi13 ? n27458 : n27473;
  assign n27475 = pi12 ? n27456 : n27474;
  assign n27476 = pi15 ? n22437 : n14606;
  assign n27477 = pi15 ? n14790 : n658;
  assign n27478 = pi14 ? n27476 : n27477;
  assign n27479 = pi13 ? n27478 : n14614;
  assign n27480 = pi12 ? n27479 : n32;
  assign n27481 = pi11 ? n27475 : n27480;
  assign n27482 = pi10 ? n27449 : n27481;
  assign n27483 = pi09 ? n32 : n27482;
  assign n27484 = pi14 ? n16899 : n27451;
  assign n27485 = pi13 ? n27484 : n27455;
  assign n27486 = pi15 ? n23631 : n23160;
  assign n27487 = pi14 ? n27457 : n27486;
  assign n27488 = pi20 ? n32 : n7229;
  assign n27489 = pi19 ? n27488 : ~n617;
  assign n27490 = pi18 ? n32 : n27489;
  assign n27491 = pi17 ? n32 : n27490;
  assign n27492 = pi16 ? n32 : n27491;
  assign n27493 = pi21 ? n100 : ~n51;
  assign n27494 = pi20 ? n32 : n27493;
  assign n27495 = pi19 ? n27494 : n32;
  assign n27496 = pi18 ? n32 : n27495;
  assign n27497 = pi17 ? n32 : n27496;
  assign n27498 = pi16 ? n32 : n27497;
  assign n27499 = pi15 ? n27492 : n27498;
  assign n27500 = pi14 ? n27467 : n27499;
  assign n27501 = pi13 ? n27487 : n27500;
  assign n27502 = pi12 ? n27485 : n27501;
  assign n27503 = pi14 ? n23679 : n14799;
  assign n27504 = pi13 ? n27503 : n32;
  assign n27505 = pi12 ? n27504 : n32;
  assign n27506 = pi11 ? n27502 : n27505;
  assign n27507 = pi10 ? n27449 : n27506;
  assign n27508 = pi09 ? n32 : n27507;
  assign n27509 = pi08 ? n27483 : n27508;
  assign n27510 = pi07 ? n27442 : n27509;
  assign n27511 = pi14 ? n17421 : n17278;
  assign n27512 = pi13 ? n32 : n27511;
  assign n27513 = pi12 ? n32 : n27512;
  assign n27514 = pi14 ? n26636 : n26439;
  assign n27515 = pi15 ? n17121 : n26315;
  assign n27516 = pi14 ? n26401 : n27515;
  assign n27517 = pi13 ? n27514 : n27516;
  assign n27518 = pi15 ? n26479 : n16392;
  assign n27519 = pi14 ? n17216 : n27518;
  assign n27520 = pi15 ? n25814 : n26111;
  assign n27521 = pi14 ? n27520 : n27445;
  assign n27522 = pi13 ? n27519 : n27521;
  assign n27523 = pi12 ? n27517 : n27522;
  assign n27524 = pi11 ? n27513 : n27523;
  assign n27525 = pi19 ? n32 : ~n429;
  assign n27526 = pi18 ? n32 : n27525;
  assign n27527 = pi17 ? n32 : n27526;
  assign n27528 = pi16 ? n32 : n27527;
  assign n27529 = pi15 ? n27528 : n16452;
  assign n27530 = pi14 ? n16899 : n27529;
  assign n27531 = pi15 ? n16452 : n24640;
  assign n27532 = pi15 ? n16308 : n26717;
  assign n27533 = pi14 ? n27531 : n27532;
  assign n27534 = pi13 ? n27530 : n27533;
  assign n27535 = pi15 ? n24097 : n26717;
  assign n27536 = pi15 ? n23631 : n15260;
  assign n27537 = pi14 ? n27535 : n27536;
  assign n27538 = pi15 ? n26930 : n15119;
  assign n27539 = pi21 ? n32 : n454;
  assign n27540 = pi20 ? n32 : n27539;
  assign n27541 = pi19 ? n27540 : n32;
  assign n27542 = pi18 ? n32 : n27541;
  assign n27543 = pi17 ? n32 : n27542;
  assign n27544 = pi16 ? n32 : n27543;
  assign n27545 = pi15 ? n27544 : n15263;
  assign n27546 = pi14 ? n27538 : n27545;
  assign n27547 = pi13 ? n27537 : n27546;
  assign n27548 = pi12 ? n27534 : n27547;
  assign n27549 = pi11 ? n27548 : n14978;
  assign n27550 = pi10 ? n27524 : n27549;
  assign n27551 = pi09 ? n32 : n27550;
  assign n27552 = pi14 ? n17443 : n17278;
  assign n27553 = pi13 ? n32 : n27552;
  assign n27554 = pi12 ? n32 : n27553;
  assign n27555 = pi14 ? n26636 : n26396;
  assign n27556 = pi13 ? n27555 : n27516;
  assign n27557 = pi15 ? n16804 : n16392;
  assign n27558 = pi14 ? n17216 : n27557;
  assign n27559 = pi14 ? n27520 : n17039;
  assign n27560 = pi13 ? n27558 : n27559;
  assign n27561 = pi12 ? n27556 : n27560;
  assign n27562 = pi11 ? n27554 : n27561;
  assign n27563 = pi15 ? n24700 : n16452;
  assign n27564 = pi14 ? n25138 : n27563;
  assign n27565 = pi15 ? n16452 : n24511;
  assign n27566 = pi15 ? n16319 : n26717;
  assign n27567 = pi14 ? n27565 : n27566;
  assign n27568 = pi13 ? n27564 : n27567;
  assign n27569 = pi15 ? n23631 : n15386;
  assign n27570 = pi14 ? n27535 : n27569;
  assign n27571 = pi13 ? n27570 : n15124;
  assign n27572 = pi12 ? n27568 : n27571;
  assign n27573 = pi11 ? n27572 : n15130;
  assign n27574 = pi10 ? n27562 : n27573;
  assign n27575 = pi09 ? n32 : n27574;
  assign n27576 = pi08 ? n27551 : n27575;
  assign n27577 = pi14 ? n26401 : n17216;
  assign n27578 = pi13 ? n27555 : n27577;
  assign n27579 = pi14 ? n17216 : n25911;
  assign n27580 = pi14 ? n25814 : n16392;
  assign n27581 = pi13 ? n27579 : n27580;
  assign n27582 = pi12 ? n27578 : n27581;
  assign n27583 = pi11 ? n27554 : n27582;
  assign n27584 = pi14 ? n26010 : n27563;
  assign n27585 = pi15 ? n16452 : n15357;
  assign n27586 = pi15 ? n15362 : n26717;
  assign n27587 = pi14 ? n27585 : n27586;
  assign n27588 = pi13 ? n27584 : n27587;
  assign n27589 = pi15 ? n24097 : n15518;
  assign n27590 = pi15 ? n15386 : n15255;
  assign n27591 = pi14 ? n27589 : n27590;
  assign n27592 = pi13 ? n27591 : n15264;
  assign n27593 = pi12 ? n27588 : n27592;
  assign n27594 = pi11 ? n27593 : n15270;
  assign n27595 = pi10 ? n27583 : n27594;
  assign n27596 = pi09 ? n32 : n27595;
  assign n27597 = pi14 ? n25815 : n16392;
  assign n27598 = pi13 ? n27579 : n27597;
  assign n27599 = pi12 ? n27578 : n27598;
  assign n27600 = pi11 ? n27554 : n27599;
  assign n27601 = pi15 ? n15511 : n15382;
  assign n27602 = pi14 ? n27601 : n15387;
  assign n27603 = pi13 ? n27602 : n15391;
  assign n27604 = pi12 ? n27588 : n27603;
  assign n27605 = pi11 ? n27604 : n32;
  assign n27606 = pi10 ? n27600 : n27605;
  assign n27607 = pi09 ? n32 : n27606;
  assign n27608 = pi08 ? n27596 : n27607;
  assign n27609 = pi07 ? n27576 : n27608;
  assign n27610 = pi06 ? n27510 : n27609;
  assign n27611 = pi15 ? n26515 : n17205;
  assign n27612 = pi14 ? n27611 : n17205;
  assign n27613 = pi15 ? n17286 : n25948;
  assign n27614 = pi14 ? n27613 : n17216;
  assign n27615 = pi13 ? n27612 : n27614;
  assign n27616 = pi15 ? n17216 : n16804;
  assign n27617 = pi14 ? n27616 : n25911;
  assign n27618 = pi14 ? n26330 : n16392;
  assign n27619 = pi13 ? n27617 : n27618;
  assign n27620 = pi12 ? n27615 : n27619;
  assign n27621 = pi11 ? n27554 : n27620;
  assign n27622 = pi14 ? n26806 : n25051;
  assign n27623 = pi19 ? n1574 : n1885;
  assign n27624 = pi18 ? n32 : n27623;
  assign n27625 = pi17 ? n32 : n27624;
  assign n27626 = pi16 ? n32 : n27625;
  assign n27627 = pi15 ? n15834 : n27626;
  assign n27628 = pi19 ? n1574 : n19892;
  assign n27629 = pi18 ? n32 : n27628;
  assign n27630 = pi17 ? n32 : n27629;
  assign n27631 = pi16 ? n32 : n27630;
  assign n27632 = pi15 ? n27626 : n27631;
  assign n27633 = pi14 ? n27627 : n27632;
  assign n27634 = pi13 ? n27622 : n27633;
  assign n27635 = pi12 ? n27634 : n15522;
  assign n27636 = pi11 ? n27635 : n32;
  assign n27637 = pi10 ? n27621 : n27636;
  assign n27638 = pi09 ? n32 : n27637;
  assign n27639 = pi15 ? n17286 : n17216;
  assign n27640 = pi14 ? n27639 : n17216;
  assign n27641 = pi13 ? n27612 : n27640;
  assign n27642 = pi12 ? n27641 : n27619;
  assign n27643 = pi11 ? n27554 : n27642;
  assign n27644 = pi14 ? n26831 : n25051;
  assign n27645 = pi14 ? n15834 : n15837;
  assign n27646 = pi13 ? n27644 : n27645;
  assign n27647 = pi12 ? n27646 : n15668;
  assign n27648 = pi11 ? n27647 : n32;
  assign n27649 = pi10 ? n27643 : n27648;
  assign n27650 = pi09 ? n32 : n27649;
  assign n27651 = pi08 ? n27638 : n27650;
  assign n27652 = pi15 ? n25948 : n16804;
  assign n27653 = pi14 ? n27652 : n25911;
  assign n27654 = pi15 ? n17066 : n16392;
  assign n27655 = pi14 ? n27654 : n25502;
  assign n27656 = pi13 ? n27653 : n27655;
  assign n27657 = pi12 ? n27641 : n27656;
  assign n27658 = pi11 ? n27554 : n27657;
  assign n27659 = pi19 ? n32 : n22410;
  assign n27660 = pi18 ? n32 : n27659;
  assign n27661 = pi17 ? n32 : n27660;
  assign n27662 = pi16 ? n32 : n27661;
  assign n27663 = pi15 ? n27662 : n16452;
  assign n27664 = pi15 ? n16452 : n15829;
  assign n27665 = pi14 ? n27663 : n27664;
  assign n27666 = pi13 ? n27665 : n15838;
  assign n27667 = pi12 ? n27666 : n32;
  assign n27668 = pi11 ? n27667 : n32;
  assign n27669 = pi10 ? n27658 : n27668;
  assign n27670 = pi09 ? n32 : n27669;
  assign n27671 = pi14 ? n26394 : n17205;
  assign n27672 = pi15 ? n17216 : n25948;
  assign n27673 = pi14 ? n17216 : n27672;
  assign n27674 = pi13 ? n27671 : n27673;
  assign n27675 = pi15 ? n17121 : n16804;
  assign n27676 = pi15 ? n16804 : n25763;
  assign n27677 = pi14 ? n27675 : n27676;
  assign n27678 = pi15 ? n16392 : n16452;
  assign n27679 = pi14 ? n25378 : n27678;
  assign n27680 = pi13 ? n27677 : n27679;
  assign n27681 = pi12 ? n27674 : n27680;
  assign n27682 = pi11 ? n27554 : n27681;
  assign n27683 = pi19 ? n32 : n5855;
  assign n27684 = pi18 ? n32 : n27683;
  assign n27685 = pi17 ? n32 : n27684;
  assign n27686 = pi16 ? n32 : n27685;
  assign n27687 = pi15 ? n27686 : n16452;
  assign n27688 = pi15 ? n16377 : n15700;
  assign n27689 = pi14 ? n27687 : n27688;
  assign n27690 = pi15 ? n16105 : n15966;
  assign n27691 = pi14 ? n27690 : n15968;
  assign n27692 = pi13 ? n27689 : n27691;
  assign n27693 = pi12 ? n27692 : n32;
  assign n27694 = pi11 ? n27693 : n32;
  assign n27695 = pi10 ? n27682 : n27694;
  assign n27696 = pi09 ? n32 : n27695;
  assign n27697 = pi08 ? n27670 : n27696;
  assign n27698 = pi07 ? n27651 : n27697;
  assign n27699 = pi15 ? n26269 : n17205;
  assign n27700 = pi14 ? n27699 : n17205;
  assign n27701 = pi14 ? n26195 : n27672;
  assign n27702 = pi13 ? n27700 : n27701;
  assign n27703 = pi15 ? n17121 : n16237;
  assign n27704 = pi15 ? n16804 : n17066;
  assign n27705 = pi14 ? n27703 : n27704;
  assign n27706 = pi14 ? n16392 : n27678;
  assign n27707 = pi13 ? n27705 : n27706;
  assign n27708 = pi12 ? n27702 : n27707;
  assign n27709 = pi11 ? n27554 : n27708;
  assign n27710 = pi14 ? n27687 : n16216;
  assign n27711 = pi13 ? n27710 : n16111;
  assign n27712 = pi12 ? n27711 : n32;
  assign n27713 = pi11 ? n27712 : n32;
  assign n27714 = pi10 ? n27709 : n27713;
  assign n27715 = pi09 ? n32 : n27714;
  assign n27716 = pi20 ? n32 : n16570;
  assign n27717 = pi19 ? n32 : n27716;
  assign n27718 = pi18 ? n32 : n27717;
  assign n27719 = pi17 ? n32 : n27718;
  assign n27720 = pi16 ? n32 : n27719;
  assign n27721 = pi15 ? n17205 : n27720;
  assign n27722 = pi14 ? n27699 : n27721;
  assign n27723 = pi13 ? n27722 : n27701;
  assign n27724 = pi12 ? n27723 : n27707;
  assign n27725 = pi11 ? n27554 : n27724;
  assign n27726 = pi14 ? n16452 : n16216;
  assign n27727 = pi13 ? n27726 : n16219;
  assign n27728 = pi12 ? n27727 : n32;
  assign n27729 = pi11 ? n27728 : n32;
  assign n27730 = pi10 ? n27725 : n27729;
  assign n27731 = pi09 ? n32 : n27730;
  assign n27732 = pi08 ? n27715 : n27731;
  assign n27733 = pi15 ? n16804 : n16237;
  assign n27734 = pi15 ? n17061 : n16392;
  assign n27735 = pi14 ? n27733 : n27734;
  assign n27736 = pi14 ? n16392 : n25918;
  assign n27737 = pi13 ? n27735 : n27736;
  assign n27738 = pi12 ? n27723 : n27737;
  assign n27739 = pi11 ? n27554 : n27738;
  assign n27740 = pi15 ? n16314 : n16319;
  assign n27741 = pi14 ? n16457 : n27740;
  assign n27742 = pi13 ? n27741 : n16322;
  assign n27743 = pi12 ? n27742 : n32;
  assign n27744 = pi11 ? n27743 : n32;
  assign n27745 = pi10 ? n27739 : n27744;
  assign n27746 = pi09 ? n32 : n27745;
  assign n27747 = pi15 ? n17128 : n16392;
  assign n27748 = pi14 ? n27733 : n27747;
  assign n27749 = pi20 ? n14793 : n32;
  assign n27750 = pi19 ? n32 : n27749;
  assign n27751 = pi18 ? n32 : n27750;
  assign n27752 = pi17 ? n32 : n27751;
  assign n27753 = pi16 ? n32 : n27752;
  assign n27754 = pi15 ? n27753 : n16515;
  assign n27755 = pi14 ? n16392 : n27754;
  assign n27756 = pi13 ? n27748 : n27755;
  assign n27757 = pi12 ? n27723 : n27756;
  assign n27758 = pi11 ? n27554 : n27757;
  assign n27759 = pi15 ? n16293 : n16377;
  assign n27760 = pi14 ? n27759 : n16378;
  assign n27761 = pi13 ? n27760 : n32;
  assign n27762 = pi12 ? n27761 : n32;
  assign n27763 = pi11 ? n27762 : n32;
  assign n27764 = pi10 ? n27758 : n27763;
  assign n27765 = pi09 ? n32 : n27764;
  assign n27766 = pi08 ? n27746 : n27765;
  assign n27767 = pi07 ? n27732 : n27766;
  assign n27768 = pi06 ? n27698 : n27767;
  assign n27769 = pi05 ? n27610 : n27768;
  assign n27770 = pi15 ? n17465 : n17278;
  assign n27771 = pi14 ? n27770 : n26571;
  assign n27772 = pi13 ? n32 : n27771;
  assign n27773 = pi12 ? n32 : n27772;
  assign n27774 = pi15 ? n26272 : n17205;
  assign n27775 = pi14 ? n27774 : n27721;
  assign n27776 = pi15 ? n26315 : n17216;
  assign n27777 = pi14 ? n27776 : n27672;
  assign n27778 = pi13 ? n27775 : n27777;
  assign n27779 = pi14 ? n16804 : n27557;
  assign n27780 = pi13 ? n27779 : n27755;
  assign n27781 = pi12 ? n27778 : n27780;
  assign n27782 = pi11 ? n27773 : n27781;
  assign n27783 = pi10 ? n27782 : n16461;
  assign n27784 = pi09 ? n32 : n27783;
  assign n27785 = pi15 ? n17216 : n17121;
  assign n27786 = pi14 ? n27776 : n27785;
  assign n27787 = pi13 ? n27775 : n27786;
  assign n27788 = pi14 ? n16804 : n25633;
  assign n27789 = pi15 ? n16392 : n16786;
  assign n27790 = pi15 ? n27753 : n16526;
  assign n27791 = pi14 ? n27789 : n27790;
  assign n27792 = pi13 ? n27788 : n27791;
  assign n27793 = pi12 ? n27787 : n27792;
  assign n27794 = pi11 ? n27773 : n27793;
  assign n27795 = pi10 ? n27794 : n32;
  assign n27796 = pi09 ? n32 : n27795;
  assign n27797 = pi08 ? n27784 : n27796;
  assign n27798 = pi14 ? n17278 : n26571;
  assign n27799 = pi13 ? n32 : n27798;
  assign n27800 = pi12 ? n32 : n27799;
  assign n27801 = pi15 ? n17205 : n26400;
  assign n27802 = pi14 ? n17205 : n27801;
  assign n27803 = pi15 ? n17216 : n17061;
  assign n27804 = pi14 ? n17216 : n27803;
  assign n27805 = pi13 ? n27802 : n27804;
  assign n27806 = pi13 ? n27788 : n16608;
  assign n27807 = pi12 ? n27805 : n27806;
  assign n27808 = pi11 ? n27800 : n27807;
  assign n27809 = pi10 ? n27808 : n32;
  assign n27810 = pi09 ? n32 : n27809;
  assign n27811 = pi13 ? n27788 : n16657;
  assign n27812 = pi12 ? n27805 : n27811;
  assign n27813 = pi11 ? n27800 : n27812;
  assign n27814 = pi10 ? n27813 : n32;
  assign n27815 = pi09 ? n32 : n27814;
  assign n27816 = pi08 ? n27810 : n27815;
  assign n27817 = pi07 ? n27797 : n27816;
  assign n27818 = pi15 ? n17205 : n17216;
  assign n27819 = pi14 ? n17205 : n27818;
  assign n27820 = pi14 ? n17216 : n17121;
  assign n27821 = pi13 ? n27819 : n27820;
  assign n27822 = pi15 ? n17061 : n16832;
  assign n27823 = pi15 ? n16832 : n16467;
  assign n27824 = pi14 ? n27822 : n27823;
  assign n27825 = pi13 ? n27824 : n16727;
  assign n27826 = pi12 ? n27821 : n27825;
  assign n27827 = pi11 ? n27800 : n27826;
  assign n27828 = pi10 ? n27827 : n32;
  assign n27829 = pi09 ? n32 : n27828;
  assign n27830 = pi14 ? n27822 : n16725;
  assign n27831 = pi13 ? n27830 : n16787;
  assign n27832 = pi12 ? n27821 : n27831;
  assign n27833 = pi11 ? n27800 : n27832;
  assign n27834 = pi10 ? n27833 : n32;
  assign n27835 = pi09 ? n32 : n27834;
  assign n27836 = pi08 ? n27829 : n27835;
  assign n27837 = pi15 ? n17121 : n17061;
  assign n27838 = pi14 ? n17216 : n27837;
  assign n27839 = pi13 ? n27819 : n27838;
  assign n27840 = pi12 ? n27839 : n16842;
  assign n27841 = pi11 ? n27800 : n27840;
  assign n27842 = pi10 ? n27841 : n32;
  assign n27843 = pi09 ? n32 : n27842;
  assign n27844 = pi14 ? n17278 : n17494;
  assign n27845 = pi13 ? n32 : n27844;
  assign n27846 = pi12 ? n32 : n27845;
  assign n27847 = pi15 ? n17331 : n17216;
  assign n27848 = pi14 ? n17205 : n27847;
  assign n27849 = pi14 ? n27785 : n27837;
  assign n27850 = pi13 ? n27848 : n27849;
  assign n27851 = pi12 ? n27850 : n16902;
  assign n27852 = pi11 ? n27846 : n27851;
  assign n27853 = pi10 ? n27852 : n32;
  assign n27854 = pi09 ? n32 : n27853;
  assign n27855 = pi08 ? n27843 : n27854;
  assign n27856 = pi07 ? n27836 : n27855;
  assign n27857 = pi06 ? n27817 : n27856;
  assign n27858 = pi15 ? n17036 : n16953;
  assign n27859 = pi14 ? n27858 : n16974;
  assign n27860 = pi13 ? n27859 : n32;
  assign n27861 = pi12 ? n27850 : n27860;
  assign n27862 = pi11 ? n27846 : n27861;
  assign n27863 = pi10 ? n27862 : n32;
  assign n27864 = pi09 ? n32 : n27863;
  assign n27865 = pi15 ? n17121 : n17013;
  assign n27866 = pi14 ? n27785 : n27865;
  assign n27867 = pi13 ? n27848 : n27866;
  assign n27868 = pi12 ? n27867 : n17019;
  assign n27869 = pi11 ? n27846 : n27868;
  assign n27870 = pi10 ? n27869 : n32;
  assign n27871 = pi09 ? n32 : n27870;
  assign n27872 = pi08 ? n27864 : n27871;
  assign n27873 = pi14 ? n17205 : n17331;
  assign n27874 = pi14 ? n27785 : n17067;
  assign n27875 = pi13 ? n27873 : n27874;
  assign n27876 = pi12 ? n27875 : n17072;
  assign n27877 = pi11 ? n27846 : n27876;
  assign n27878 = pi10 ? n27877 : n32;
  assign n27879 = pi09 ? n32 : n27878;
  assign n27880 = pi15 ? n17061 : n17170;
  assign n27881 = pi14 ? n27785 : n27880;
  assign n27882 = pi13 ? n27873 : n27881;
  assign n27883 = pi12 ? n27882 : n17102;
  assign n27884 = pi11 ? n27846 : n27883;
  assign n27885 = pi10 ? n27884 : n32;
  assign n27886 = pi09 ? n32 : n27885;
  assign n27887 = pi08 ? n27879 : n27886;
  assign n27888 = pi07 ? n27872 : n27887;
  assign n27889 = pi14 ? n17262 : n26121;
  assign n27890 = pi13 ? n27873 : n27889;
  assign n27891 = pi12 ? n27890 : n32;
  assign n27892 = pi11 ? n27846 : n27891;
  assign n27893 = pi10 ? n27892 : n32;
  assign n27894 = pi09 ? n32 : n27893;
  assign n27895 = pi15 ? n17261 : n17128;
  assign n27896 = pi14 ? n27895 : n17230;
  assign n27897 = pi13 ? n27848 : n27896;
  assign n27898 = pi12 ? n27897 : n32;
  assign n27899 = pi11 ? n27846 : n27898;
  assign n27900 = pi10 ? n27899 : n32;
  assign n27901 = pi09 ? n32 : n27900;
  assign n27902 = pi08 ? n27894 : n27901;
  assign n27903 = pi13 ? n27848 : n17263;
  assign n27904 = pi12 ? n27903 : n32;
  assign n27905 = pi11 ? n27846 : n27904;
  assign n27906 = pi10 ? n27905 : n32;
  assign n27907 = pi09 ? n32 : n27906;
  assign n27908 = pi15 ? n17205 : n17363;
  assign n27909 = pi15 ? n17331 : n17261;
  assign n27910 = pi14 ? n27908 : n27909;
  assign n27911 = pi13 ? n27910 : n17301;
  assign n27912 = pi12 ? n27911 : n32;
  assign n27913 = pi11 ? n27846 : n27912;
  assign n27914 = pi10 ? n27913 : n32;
  assign n27915 = pi09 ? n32 : n27914;
  assign n27916 = pi08 ? n27907 : n27915;
  assign n27917 = pi07 ? n27902 : n27916;
  assign n27918 = pi06 ? n27888 : n27917;
  assign n27919 = pi05 ? n27857 : n27918;
  assign n27920 = pi04 ? n27769 : n27919;
  assign n27921 = pi03 ? n27372 : n27920;
  assign n27922 = pi21 ? n140 : ~n242;
  assign n27923 = pi20 ? n32 : n27922;
  assign n27924 = pi19 ? n32 : n27923;
  assign n27925 = pi18 ? n32 : n27924;
  assign n27926 = pi17 ? n32 : n27925;
  assign n27927 = pi16 ? n32 : n27926;
  assign n27928 = pi15 ? n27927 : n17205;
  assign n27929 = pi14 ? n17278 : n27928;
  assign n27930 = pi13 ? n32 : n27929;
  assign n27931 = pi12 ? n32 : n27930;
  assign n27932 = pi15 ? n17454 : n17121;
  assign n27933 = pi14 ? n17448 : n27932;
  assign n27934 = pi15 ? n16984 : n17188;
  assign n27935 = pi14 ? n27934 : n32;
  assign n27936 = pi13 ? n27933 : n27935;
  assign n27937 = pi12 ? n27936 : n32;
  assign n27938 = pi11 ? n27931 : n27937;
  assign n27939 = pi10 ? n27938 : n32;
  assign n27940 = pi09 ? n32 : n27939;
  assign n27941 = pi07 ? n27915 : n27940;
  assign n27942 = pi13 ? n27933 : n17413;
  assign n27943 = pi12 ? n27942 : n32;
  assign n27944 = pi11 ? n27931 : n27943;
  assign n27945 = pi10 ? n27944 : n32;
  assign n27946 = pi09 ? n32 : n27945;
  assign n27947 = pi08 ? n27940 : n27946;
  assign n27948 = pi14 ? n17448 : n17262;
  assign n27949 = pi13 ? n27948 : n17413;
  assign n27950 = pi12 ? n27949 : n32;
  assign n27951 = pi11 ? n27931 : n27950;
  assign n27952 = pi10 ? n27951 : n32;
  assign n27953 = pi09 ? n32 : n27952;
  assign n27954 = pi08 ? n27953 : n27946;
  assign n27955 = pi07 ? n27947 : n27954;
  assign n27956 = pi06 ? n27941 : n27955;
  assign n27957 = pi11 ? n27931 : n17458;
  assign n27958 = pi10 ? n27957 : n32;
  assign n27959 = pi09 ? n32 : n27958;
  assign n27960 = pi11 ? n27931 : n17473;
  assign n27961 = pi10 ? n27960 : n32;
  assign n27962 = pi09 ? n32 : n27961;
  assign n27963 = pi11 ? n27931 : n17480;
  assign n27964 = pi10 ? n27963 : n32;
  assign n27965 = pi09 ? n32 : n27964;
  assign n27966 = pi08 ? n27962 : n27965;
  assign n27967 = pi07 ? n27959 : n27966;
  assign n27968 = pi14 ? n17443 : n17494;
  assign n27969 = pi13 ? n32 : n27968;
  assign n27970 = pi12 ? n32 : n27969;
  assign n27971 = pi11 ? n27970 : n17480;
  assign n27972 = pi10 ? n27971 : n32;
  assign n27973 = pi09 ? n32 : n27972;
  assign n27974 = pi11 ? n27970 : n17504;
  assign n27975 = pi10 ? n27974 : n32;
  assign n27976 = pi09 ? n32 : n27975;
  assign n27977 = pi08 ? n27973 : n27976;
  assign n27978 = pi15 ? n27927 : n17363;
  assign n27979 = pi14 ? n17443 : n27978;
  assign n27980 = pi13 ? n32 : n27979;
  assign n27981 = pi12 ? n32 : n27980;
  assign n27982 = pi11 ? n27981 : n17521;
  assign n27983 = pi10 ? n27982 : n32;
  assign n27984 = pi09 ? n32 : n27983;
  assign n27985 = pi07 ? n27977 : n27984;
  assign n27986 = pi06 ? n27967 : n27985;
  assign n27987 = pi05 ? n27956 : n27986;
  assign n27988 = pi15 ? n27927 : n17331;
  assign n27989 = pi14 ? n17443 : n27988;
  assign n27990 = pi13 ? n32 : n27989;
  assign n27991 = pi12 ? n32 : n27990;
  assign n27992 = pi11 ? n27991 : n32;
  assign n27993 = pi10 ? n27992 : n32;
  assign n27994 = pi09 ? n32 : n27993;
  assign n27995 = pi08 ? n27994 : n17554;
  assign n27996 = pi07 ? n27994 : n27995;
  assign n27997 = pi06 ? n27996 : n17561;
  assign n27998 = pi05 ? n27997 : n17565;
  assign n27999 = pi04 ? n27987 : n27998;
  assign n28000 = pi03 ? n27999 : n32;
  assign n28001 = pi02 ? n27921 : n28000;
  assign n28002 = pi06 ? n17586 : n17568;
  assign n28003 = pi05 ? n28002 : n17568;
  assign n28004 = pi08 ? n17568 : n32;
  assign n28005 = pi07 ? n28004 : n32;
  assign n28006 = pi06 ? n17568 : n28005;
  assign n28007 = pi05 ? n28006 : n32;
  assign n28008 = pi04 ? n28003 : n28007;
  assign n28009 = pi03 ? n32 : n28008;
  assign n28010 = pi02 ? n28009 : n32;
  assign n28011 = pi01 ? n28001 : n28010;
  assign n28012 = pi00 ? n26221 : n28011;
  assign n28013 = pi20 ? n357 : n67;
  assign n28014 = pi19 ? n857 : n28013;
  assign n28015 = pi18 ? n28014 : n32;
  assign n28016 = pi17 ? n21317 : n28015;
  assign n28017 = pi16 ? n32 : n28016;
  assign n28018 = pi15 ? n32 : n28017;
  assign n28019 = pi19 ? n32 : n1785;
  assign n28020 = pi18 ? n28019 : n32;
  assign n28021 = pi17 ? n32 : n28020;
  assign n28022 = pi16 ? n32 : n28021;
  assign n28023 = pi15 ? n28017 : n28022;
  assign n28024 = pi14 ? n28018 : n28023;
  assign n28025 = pi13 ? n32 : n28024;
  assign n28026 = pi12 ? n32 : n28025;
  assign n28027 = pi16 ? n17884 : n28021;
  assign n28028 = pi15 ? n28022 : n28027;
  assign n28029 = pi18 ? n863 : n237;
  assign n28030 = pi17 ? n32 : n28029;
  assign n28031 = pi18 ? n17118 : n20172;
  assign n28032 = pi19 ? n9007 : n342;
  assign n28033 = pi18 ? n28032 : ~n32;
  assign n28034 = pi17 ? n28031 : n28033;
  assign n28035 = pi16 ? n28030 : ~n28034;
  assign n28036 = pi20 ? n206 : ~n246;
  assign n28037 = pi19 ? n28036 : ~n4670;
  assign n28038 = pi18 ? n863 : n28037;
  assign n28039 = pi17 ? n32 : n28038;
  assign n28040 = pi19 ? n18502 : ~n9007;
  assign n28041 = pi20 ? n206 : ~n266;
  assign n28042 = pi19 ? n266 : ~n28041;
  assign n28043 = pi18 ? n28040 : ~n28042;
  assign n28044 = pi19 ? n11879 : ~n6308;
  assign n28045 = pi18 ? n28044 : ~n32;
  assign n28046 = pi17 ? n28043 : ~n28045;
  assign n28047 = pi16 ? n28039 : n28046;
  assign n28048 = pi15 ? n28035 : n28047;
  assign n28049 = pi14 ? n28028 : n28048;
  assign n28050 = pi13 ? n28049 : n32;
  assign n28051 = pi15 ? n17637 : n32;
  assign n28052 = pi14 ? n17852 : n28051;
  assign n28053 = pi19 ? n32 : n19141;
  assign n28054 = pi20 ? n18281 : n18253;
  assign n28055 = pi19 ? n28054 : n18409;
  assign n28056 = pi18 ? n28053 : ~n28055;
  assign n28057 = pi17 ? n32 : n28056;
  assign n28058 = pi20 ? n9194 : n9488;
  assign n28059 = pi20 ? n17652 : n18415;
  assign n28060 = pi19 ? n28058 : ~n28059;
  assign n28061 = pi20 ? n18415 : ~n18129;
  assign n28062 = pi19 ? n28061 : n18281;
  assign n28063 = pi18 ? n28060 : ~n28062;
  assign n28064 = pi20 ? n18415 : ~n17665;
  assign n28065 = pi20 ? n18073 : n12884;
  assign n28066 = pi19 ? n28064 : ~n28065;
  assign n28067 = pi18 ? n28066 : ~n32;
  assign n28068 = pi17 ? n28063 : ~n28067;
  assign n28069 = pi16 ? n28057 : n28068;
  assign n28070 = pi20 ? n32 : n3843;
  assign n28071 = pi19 ? n32 : n28070;
  assign n28072 = pi20 ? n18832 : n18408;
  assign n28073 = pi19 ? n28072 : ~n18782;
  assign n28074 = pi18 ? n28071 : ~n28073;
  assign n28075 = pi17 ? n32 : n28074;
  assign n28076 = pi20 ? n18253 : n9491;
  assign n28077 = pi19 ? n18404 : ~n28076;
  assign n28078 = pi20 ? n18073 : n2180;
  assign n28079 = pi19 ? n28078 : n18832;
  assign n28080 = pi18 ? n28077 : ~n28079;
  assign n28081 = pi20 ? n18073 : n333;
  assign n28082 = pi21 ? n173 : ~n10445;
  assign n28083 = pi20 ? n18832 : n28082;
  assign n28084 = pi19 ? n28081 : ~n28083;
  assign n28085 = pi18 ? n28084 : ~n32;
  assign n28086 = pi17 ? n28080 : ~n28085;
  assign n28087 = pi16 ? n28075 : n28086;
  assign n28088 = pi15 ? n28069 : n28087;
  assign n28089 = pi20 ? n9491 : n18253;
  assign n28090 = pi19 ? n28089 : n18832;
  assign n28091 = pi18 ? n28077 : ~n28090;
  assign n28092 = pi20 ? n9491 : n17652;
  assign n28093 = pi20 ? n9488 : n28082;
  assign n28094 = pi19 ? n28092 : ~n28093;
  assign n28095 = pi18 ? n28094 : ~n32;
  assign n28096 = pi17 ? n28091 : ~n28095;
  assign n28097 = pi16 ? n28075 : n28096;
  assign n28098 = pi16 ? n18561 : n32;
  assign n28099 = pi15 ? n28097 : n28098;
  assign n28100 = pi14 ? n28088 : n28099;
  assign n28101 = pi13 ? n28052 : n28100;
  assign n28102 = pi12 ? n28050 : n28101;
  assign n28103 = pi11 ? n28026 : n28102;
  assign n28104 = pi15 ? n32 : n17837;
  assign n28105 = pi14 ? n28104 : n17702;
  assign n28106 = pi15 ? n17702 : n17825;
  assign n28107 = pi14 ? n28106 : n17702;
  assign n28108 = pi13 ? n28105 : n28107;
  assign n28109 = pi14 ? n17702 : n17708;
  assign n28110 = pi15 ? n17707 : n17736;
  assign n28111 = pi15 ? n17856 : n17717;
  assign n28112 = pi14 ? n28110 : n28111;
  assign n28113 = pi13 ? n28109 : n28112;
  assign n28114 = pi12 ? n28108 : n28113;
  assign n28115 = pi20 ? n246 : n7388;
  assign n28116 = pi19 ? n32 : n28115;
  assign n28117 = pi18 ? n28116 : n32;
  assign n28118 = pi17 ? n32 : n28117;
  assign n28119 = pi16 ? n32 : n28118;
  assign n28120 = pi19 ? n32 : n23699;
  assign n28121 = pi18 ? n28120 : n32;
  assign n28122 = pi17 ? n32 : n28121;
  assign n28123 = pi16 ? n32 : n28122;
  assign n28124 = pi15 ? n28119 : n28123;
  assign n28125 = pi14 ? n32 : n28124;
  assign n28126 = pi19 ? n32 : n17752;
  assign n28127 = pi18 ? n28126 : n32;
  assign n28128 = pi17 ? n17768 : n28127;
  assign n28129 = pi16 ? n32 : n28128;
  assign n28130 = pi20 ? n7839 : n266;
  assign n28131 = pi19 ? n28130 : n4670;
  assign n28132 = pi18 ? n32 : n28131;
  assign n28133 = pi17 ? n32 : n28132;
  assign n28134 = pi20 ? n207 : ~n220;
  assign n28135 = pi19 ? n28134 : n32;
  assign n28136 = pi18 ? n28135 : n15984;
  assign n28137 = pi17 ? n28136 : n1842;
  assign n28138 = pi16 ? n28133 : ~n28137;
  assign n28139 = pi15 ? n28129 : n28138;
  assign n28140 = pi20 ? n220 : ~n17669;
  assign n28141 = pi19 ? n28140 : n19129;
  assign n28142 = pi18 ? n1819 : n28141;
  assign n28143 = pi17 ? n32 : n28142;
  assign n28144 = pi20 ? n6050 : n310;
  assign n28145 = pi19 ? n28144 : ~n236;
  assign n28146 = pi19 ? n247 : ~n23644;
  assign n28147 = pi18 ? n28145 : n28146;
  assign n28148 = pi19 ? n9037 : ~n18211;
  assign n28149 = pi18 ? n28148 : ~n32;
  assign n28150 = pi17 ? n28147 : n28149;
  assign n28151 = pi16 ? n28143 : ~n28150;
  assign n28152 = pi20 ? n266 : ~n2358;
  assign n28153 = pi19 ? n9037 : ~n28152;
  assign n28154 = pi18 ? n28153 : ~n32;
  assign n28155 = pi17 ? n28147 : n28154;
  assign n28156 = pi16 ? n28143 : ~n28155;
  assign n28157 = pi15 ? n28151 : n28156;
  assign n28158 = pi14 ? n28139 : n28157;
  assign n28159 = pi13 ? n28125 : n28158;
  assign n28160 = pi19 ? n32 : n206;
  assign n28161 = pi20 ? n274 : ~n207;
  assign n28162 = pi19 ? n28161 : n32;
  assign n28163 = pi18 ? n28160 : n28162;
  assign n28164 = pi19 ? n9007 : n1757;
  assign n28165 = pi18 ? n28164 : n32;
  assign n28166 = pi17 ? n28163 : n28165;
  assign n28167 = pi16 ? n32 : n28166;
  assign n28168 = pi16 ? n32 : n270;
  assign n28169 = pi15 ? n28167 : n28168;
  assign n28170 = pi14 ? n28169 : n32;
  assign n28171 = pi18 ? n6600 : n32;
  assign n28172 = pi19 ? n7089 : n9007;
  assign n28173 = pi18 ? n28172 : n32;
  assign n28174 = pi17 ? n28171 : n28173;
  assign n28175 = pi16 ? n32 : n28174;
  assign n28176 = pi15 ? n32 : n28175;
  assign n28177 = pi20 ? n32 : n287;
  assign n28178 = pi19 ? n32 : n28177;
  assign n28179 = pi20 ? n206 : ~n207;
  assign n28180 = pi19 ? n21349 : n28179;
  assign n28181 = pi18 ? n28178 : ~n28180;
  assign n28182 = pi17 ? n32 : n28181;
  assign n28183 = pi19 ? n4391 : ~n17766;
  assign n28184 = pi20 ? n206 : ~n206;
  assign n28185 = pi19 ? n507 : n28184;
  assign n28186 = pi18 ? n28183 : ~n28185;
  assign n28187 = pi19 ? n267 : n24218;
  assign n28188 = pi18 ? n28187 : ~n32;
  assign n28189 = pi17 ? n28186 : ~n28188;
  assign n28190 = pi16 ? n28182 : n28189;
  assign n28191 = pi20 ? n246 : ~n246;
  assign n28192 = pi19 ? n322 : ~n28191;
  assign n28193 = pi19 ? n1248 : ~n32;
  assign n28194 = pi18 ? n28192 : ~n28193;
  assign n28195 = pi19 ? n1757 : n208;
  assign n28196 = pi18 ? n28195 : ~n32;
  assign n28197 = pi17 ? n28194 : ~n28196;
  assign n28198 = pi16 ? n18813 : n28197;
  assign n28199 = pi15 ? n28190 : n28198;
  assign n28200 = pi14 ? n28176 : n28199;
  assign n28201 = pi13 ? n28170 : n28200;
  assign n28202 = pi12 ? n28159 : n28201;
  assign n28203 = pi11 ? n28114 : n28202;
  assign n28204 = pi10 ? n28103 : n28203;
  assign n28205 = pi09 ? n32 : n28204;
  assign n28206 = pi20 ? n357 : n2077;
  assign n28207 = pi19 ? n857 : n28206;
  assign n28208 = pi18 ? n28207 : n32;
  assign n28209 = pi17 ? n21317 : n28208;
  assign n28210 = pi16 ? n32 : n28209;
  assign n28211 = pi15 ? n32 : n28210;
  assign n28212 = pi20 ? n357 : n13387;
  assign n28213 = pi19 ? n857 : n28212;
  assign n28214 = pi18 ? n28213 : n32;
  assign n28215 = pi17 ? n21317 : n28214;
  assign n28216 = pi16 ? n32 : n28215;
  assign n28217 = pi15 ? n28216 : n17813;
  assign n28218 = pi14 ? n28211 : n28217;
  assign n28219 = pi13 ? n32 : n28218;
  assign n28220 = pi12 ? n32 : n28219;
  assign n28221 = pi16 ? n17884 : n17812;
  assign n28222 = pi15 ? n17813 : n28221;
  assign n28223 = pi20 ? n342 : n12019;
  assign n28224 = pi19 ? n9007 : n28223;
  assign n28225 = pi18 ? n28224 : ~n32;
  assign n28226 = pi17 ? n28031 : n28225;
  assign n28227 = pi16 ? n28030 : ~n28226;
  assign n28228 = pi20 ? n220 : ~n12019;
  assign n28229 = pi19 ? n11879 : ~n28228;
  assign n28230 = pi18 ? n28229 : ~n32;
  assign n28231 = pi17 ? n28043 : ~n28230;
  assign n28232 = pi16 ? n28039 : n28231;
  assign n28233 = pi15 ? n28227 : n28232;
  assign n28234 = pi14 ? n28222 : n28233;
  assign n28235 = pi13 ? n28234 : n17813;
  assign n28236 = pi15 ? n17851 : n17813;
  assign n28237 = pi14 ? n28236 : n17813;
  assign n28238 = pi20 ? n18073 : n17665;
  assign n28239 = pi19 ? n28064 : ~n28238;
  assign n28240 = pi18 ? n28239 : ~n32;
  assign n28241 = pi17 ? n28063 : ~n28240;
  assign n28242 = pi16 ? n28057 : n28241;
  assign n28243 = pi20 ? n17671 : n1817;
  assign n28244 = pi19 ? n18173 : ~n28243;
  assign n28245 = pi18 ? n19082 : ~n28244;
  assign n28246 = pi17 ? n32 : n28245;
  assign n28247 = pi20 ? n314 : n18253;
  assign n28248 = pi19 ? n18567 : ~n28247;
  assign n28249 = pi20 ? n18281 : n501;
  assign n28250 = pi19 ? n28249 : n18173;
  assign n28251 = pi18 ? n28248 : ~n28250;
  assign n28252 = pi20 ? n9491 : n17665;
  assign n28253 = pi19 ? n18621 : ~n28252;
  assign n28254 = pi18 ? n28253 : ~n32;
  assign n28255 = pi17 ? n28251 : ~n28254;
  assign n28256 = pi16 ? n28246 : n28255;
  assign n28257 = pi15 ? n28242 : n28256;
  assign n28258 = pi20 ? n9488 : n2019;
  assign n28259 = pi19 ? n28092 : ~n28258;
  assign n28260 = pi18 ? n28259 : ~n32;
  assign n28261 = pi17 ? n28091 : ~n28260;
  assign n28262 = pi16 ? n28075 : n28261;
  assign n28263 = pi15 ? n28262 : n28098;
  assign n28264 = pi14 ? n28257 : n28263;
  assign n28265 = pi13 ? n28237 : n28264;
  assign n28266 = pi12 ? n28235 : n28265;
  assign n28267 = pi11 ? n28220 : n28266;
  assign n28268 = pi14 ? n32 : n17825;
  assign n28269 = pi15 ? n17825 : n17915;
  assign n28270 = pi14 ? n28269 : n17825;
  assign n28271 = pi13 ? n28268 : n28270;
  assign n28272 = pi14 ? n18327 : n17708;
  assign n28273 = pi19 ? n32 : n383;
  assign n28274 = pi18 ? n28273 : n32;
  assign n28275 = pi17 ? n32 : n28274;
  assign n28276 = pi16 ? n32 : n28275;
  assign n28277 = pi15 ? n28276 : n17736;
  assign n28278 = pi14 ? n28277 : n19012;
  assign n28279 = pi13 ? n28272 : n28278;
  assign n28280 = pi12 ? n28271 : n28279;
  assign n28281 = pi20 ? n246 : n1685;
  assign n28282 = pi19 ? n32 : n28281;
  assign n28283 = pi18 ? n28282 : n32;
  assign n28284 = pi17 ? n32 : n28283;
  assign n28285 = pi16 ? n32 : n28284;
  assign n28286 = pi18 ? n16603 : n32;
  assign n28287 = pi19 ? n32 : n13340;
  assign n28288 = pi18 ? n28287 : n32;
  assign n28289 = pi17 ? n28286 : n28288;
  assign n28290 = pi16 ? n32 : n28289;
  assign n28291 = pi15 ? n28285 : n28290;
  assign n28292 = pi14 ? n32 : n28291;
  assign n28293 = pi20 ? n246 : ~n518;
  assign n28294 = pi19 ? n32 : n28293;
  assign n28295 = pi18 ? n28294 : n32;
  assign n28296 = pi17 ? n17768 : n28295;
  assign n28297 = pi16 ? n32 : n28296;
  assign n28298 = pi17 ? n28136 : n1593;
  assign n28299 = pi16 ? n28133 : ~n28298;
  assign n28300 = pi15 ? n28297 : n28299;
  assign n28301 = pi14 ? n28300 : n28157;
  assign n28302 = pi13 ? n28292 : n28301;
  assign n28303 = pi19 ? n1757 : n1969;
  assign n28304 = pi18 ? n28303 : ~n32;
  assign n28305 = pi17 ? n28194 : ~n28304;
  assign n28306 = pi16 ? n18813 : n28305;
  assign n28307 = pi15 ? n28190 : n28306;
  assign n28308 = pi14 ? n28176 : n28307;
  assign n28309 = pi13 ? n28170 : n28308;
  assign n28310 = pi12 ? n28302 : n28309;
  assign n28311 = pi11 ? n28280 : n28310;
  assign n28312 = pi10 ? n28267 : n28311;
  assign n28313 = pi09 ? n32 : n28312;
  assign n28314 = pi08 ? n28205 : n28313;
  assign n28315 = pi07 ? n32 : n28314;
  assign n28316 = pi06 ? n32 : n28315;
  assign n28317 = pi19 ? n857 : n358;
  assign n28318 = pi18 ? n28317 : n32;
  assign n28319 = pi17 ? n21317 : n28318;
  assign n28320 = pi16 ? n32 : n28319;
  assign n28321 = pi14 ? n28320 : n17885;
  assign n28322 = pi13 ? n32 : n28321;
  assign n28323 = pi12 ? n32 : n28322;
  assign n28324 = pi14 ? n32 : n17885;
  assign n28325 = pi13 ? n17897 : n28324;
  assign n28326 = pi18 ? n858 : ~n28055;
  assign n28327 = pi17 ? n32 : n28326;
  assign n28328 = pi20 ? n354 : n314;
  assign n28329 = pi19 ? n28058 : ~n28328;
  assign n28330 = pi19 ? n18333 : n18266;
  assign n28331 = pi18 ? n28329 : ~n28330;
  assign n28332 = pi20 ? n17665 : n17669;
  assign n28333 = pi19 ? n18789 : n28332;
  assign n28334 = pi18 ? n28333 : n32;
  assign n28335 = pi17 ? n28331 : n28334;
  assign n28336 = pi16 ? n28327 : n28335;
  assign n28337 = pi15 ? n32 : n28336;
  assign n28338 = pi20 ? n17665 : n18073;
  assign n28339 = pi19 ? n18789 : n28338;
  assign n28340 = pi18 ? n28339 : n32;
  assign n28341 = pi17 ? n28331 : n28340;
  assign n28342 = pi16 ? n28327 : n28341;
  assign n28343 = pi19 ? n5748 : n9007;
  assign n28344 = pi18 ? n24063 : n28343;
  assign n28345 = pi20 ? n342 : n428;
  assign n28346 = pi19 ? n267 : ~n28345;
  assign n28347 = pi18 ? n28346 : ~n32;
  assign n28348 = pi17 ? n28344 : ~n28347;
  assign n28349 = pi16 ? n20257 : n28348;
  assign n28350 = pi15 ? n28342 : n28349;
  assign n28351 = pi14 ? n28337 : n28350;
  assign n28352 = pi20 ? n1817 : n342;
  assign n28353 = pi19 ? n32 : n28352;
  assign n28354 = pi19 ? n17649 : n462;
  assign n28355 = pi18 ? n28353 : n28354;
  assign n28356 = pi20 ? n9491 : n17669;
  assign n28357 = pi20 ? n1324 : n27030;
  assign n28358 = pi19 ? n28356 : n28357;
  assign n28359 = pi18 ? n28358 : n32;
  assign n28360 = pi17 ? n28355 : n28359;
  assign n28361 = pi16 ? n17706 : n28360;
  assign n28362 = pi19 ? n207 : ~n23644;
  assign n28363 = pi18 ? n19082 : ~n28362;
  assign n28364 = pi17 ? n32 : n28363;
  assign n28365 = pi20 ? n501 : n17652;
  assign n28366 = pi19 ? n4670 : ~n28365;
  assign n28367 = pi20 ? n5854 : ~n357;
  assign n28368 = pi19 ? n28367 : n6050;
  assign n28369 = pi18 ? n28366 : ~n28368;
  assign n28370 = pi20 ? n1324 : n246;
  assign n28371 = pi19 ? n18133 : ~n28370;
  assign n28372 = pi18 ? n28371 : ~n32;
  assign n28373 = pi17 ? n28369 : ~n28372;
  assign n28374 = pi16 ? n28364 : n28373;
  assign n28375 = pi15 ? n28361 : n28374;
  assign n28376 = pi14 ? n28375 : n32;
  assign n28377 = pi13 ? n28351 : n28376;
  assign n28378 = pi12 ? n28325 : n28377;
  assign n28379 = pi11 ? n28323 : n28378;
  assign n28380 = pi16 ? n19804 : n17884;
  assign n28381 = pi15 ? n28380 : n17885;
  assign n28382 = pi19 ? n1757 : n507;
  assign n28383 = pi18 ? n28382 : n32;
  assign n28384 = pi17 ? n32 : n28383;
  assign n28385 = pi16 ? n32 : n28384;
  assign n28386 = pi15 ? n17903 : n28385;
  assign n28387 = pi14 ? n28381 : n28386;
  assign n28388 = pi19 ? n11374 : n17655;
  assign n28389 = pi18 ? n28388 : n32;
  assign n28390 = pi17 ? n3282 : n28389;
  assign n28391 = pi16 ? n32 : n28390;
  assign n28392 = pi15 ? n32 : n28391;
  assign n28393 = pi14 ? n17903 : n28392;
  assign n28394 = pi13 ? n28387 : n28393;
  assign n28395 = pi15 ? n17915 : n18326;
  assign n28396 = pi15 ? n18326 : n32;
  assign n28397 = pi14 ? n28395 : n28396;
  assign n28398 = pi14 ? n28396 : n32;
  assign n28399 = pi13 ? n28397 : n28398;
  assign n28400 = pi12 ? n28394 : n28399;
  assign n28401 = pi18 ? n16801 : n32;
  assign n28402 = pi20 ? n321 : n1817;
  assign n28403 = pi19 ? n507 : n28402;
  assign n28404 = pi18 ? n28403 : n32;
  assign n28405 = pi17 ? n28401 : n28404;
  assign n28406 = pi16 ? n32 : n28405;
  assign n28407 = pi18 ? n16389 : n32;
  assign n28408 = pi20 ? n207 : n1685;
  assign n28409 = pi19 ? n1464 : n28408;
  assign n28410 = pi18 ? n28409 : n32;
  assign n28411 = pi17 ? n28407 : n28410;
  assign n28412 = pi16 ? n32 : n28411;
  assign n28413 = pi15 ? n28406 : n28412;
  assign n28414 = pi14 ? n32 : n28413;
  assign n28415 = pi18 ? n15844 : n32;
  assign n28416 = pi20 ? n32 : ~n1685;
  assign n28417 = pi19 ? n1464 : ~n28416;
  assign n28418 = pi18 ? n28417 : n32;
  assign n28419 = pi17 ? n28415 : n28418;
  assign n28420 = pi16 ? n32 : n28419;
  assign n28421 = pi19 ? n4670 : ~n32;
  assign n28422 = pi18 ? n702 : ~n28421;
  assign n28423 = pi19 ? n343 : ~n519;
  assign n28424 = pi18 ? n28423 : n32;
  assign n28425 = pi17 ? n28422 : n28424;
  assign n28426 = pi16 ? n19804 : n28425;
  assign n28427 = pi15 ? n28420 : n28426;
  assign n28428 = pi18 ? n21888 : ~n237;
  assign n28429 = pi19 ? n208 : ~n11027;
  assign n28430 = pi18 ? n28429 : n32;
  assign n28431 = pi17 ? n28428 : n28430;
  assign n28432 = pi16 ? n32 : n28431;
  assign n28433 = pi19 ? n208 : ~n349;
  assign n28434 = pi18 ? n28433 : n32;
  assign n28435 = pi17 ? n28428 : n28434;
  assign n28436 = pi16 ? n32 : n28435;
  assign n28437 = pi15 ? n28432 : n28436;
  assign n28438 = pi14 ? n28427 : n28437;
  assign n28439 = pi13 ? n28414 : n28438;
  assign n28440 = pi18 ? n23440 : n32;
  assign n28441 = pi17 ? n32 : n28440;
  assign n28442 = pi16 ? n32 : n28441;
  assign n28443 = pi15 ? n28442 : n32;
  assign n28444 = pi14 ? n28443 : n32;
  assign n28445 = pi18 ? n5749 : n32;
  assign n28446 = pi17 ? n32 : n28445;
  assign n28447 = pi16 ? n32 : n28446;
  assign n28448 = pi15 ? n32 : n28447;
  assign n28449 = pi17 ? n32 : n6119;
  assign n28450 = pi18 ? n17975 : n4671;
  assign n28451 = pi20 ? n915 : n207;
  assign n28452 = pi19 ? n786 : n28451;
  assign n28453 = pi18 ? n28452 : ~n32;
  assign n28454 = pi17 ? n28450 : n28453;
  assign n28455 = pi16 ? n28449 : ~n28454;
  assign n28456 = pi20 ? n4279 : ~n1817;
  assign n28457 = pi19 ? n28456 : ~n208;
  assign n28458 = pi18 ? n28457 : n32;
  assign n28459 = pi17 ? n32 : n28458;
  assign n28460 = pi16 ? n32 : n28459;
  assign n28461 = pi15 ? n28455 : n28460;
  assign n28462 = pi14 ? n28448 : n28461;
  assign n28463 = pi13 ? n28444 : n28462;
  assign n28464 = pi12 ? n28439 : n28463;
  assign n28465 = pi11 ? n28400 : n28464;
  assign n28466 = pi10 ? n28379 : n28465;
  assign n28467 = pi09 ? n32 : n28466;
  assign n28468 = pi18 ? n28317 : ~n1676;
  assign n28469 = pi17 ? n21317 : n28468;
  assign n28470 = pi16 ? n32 : n28469;
  assign n28471 = pi15 ? n18972 : n17894;
  assign n28472 = pi14 ? n28470 : n28471;
  assign n28473 = pi13 ? n32 : n28472;
  assign n28474 = pi12 ? n32 : n28473;
  assign n28475 = pi14 ? n17894 : n19717;
  assign n28476 = pi13 ? n17894 : n28475;
  assign n28477 = pi20 ? n18129 : n1331;
  assign n28478 = pi19 ? n28477 : ~n18571;
  assign n28479 = pi18 ? n858 : n28478;
  assign n28480 = pi17 ? n32 : n28479;
  assign n28481 = pi20 ? n1817 : n6085;
  assign n28482 = pi19 ? n28481 : n20937;
  assign n28483 = pi20 ? n1331 : n175;
  assign n28484 = pi19 ? n28483 : n1331;
  assign n28485 = pi18 ? n28482 : n28484;
  assign n28486 = pi20 ? n1817 : n1324;
  assign n28487 = pi19 ? n18789 : n28486;
  assign n28488 = pi18 ? n28487 : ~n618;
  assign n28489 = pi17 ? n28485 : n28488;
  assign n28490 = pi16 ? n28480 : n28489;
  assign n28491 = pi15 ? n18008 : n28490;
  assign n28492 = pi20 ? n1817 : n9641;
  assign n28493 = pi19 ? n18789 : n28492;
  assign n28494 = pi18 ? n28493 : n32;
  assign n28495 = pi17 ? n28485 : n28494;
  assign n28496 = pi16 ? n28480 : n28495;
  assign n28497 = pi15 ? n28496 : n28349;
  assign n28498 = pi14 ? n28491 : n28497;
  assign n28499 = pi19 ? n28356 : n1324;
  assign n28500 = pi18 ? n28499 : n32;
  assign n28501 = pi17 ? n28355 : n28500;
  assign n28502 = pi16 ? n17706 : n28501;
  assign n28503 = pi18 ? n18134 : ~n32;
  assign n28504 = pi17 ? n28369 : ~n28503;
  assign n28505 = pi16 ? n28364 : n28504;
  assign n28506 = pi15 ? n28502 : n28505;
  assign n28507 = pi15 ? n17885 : n32;
  assign n28508 = pi14 ? n28506 : n28507;
  assign n28509 = pi13 ? n28498 : n28508;
  assign n28510 = pi12 ? n28476 : n28509;
  assign n28511 = pi11 ? n28474 : n28510;
  assign n28512 = pi16 ? n19804 : n18971;
  assign n28513 = pi15 ? n28512 : n18972;
  assign n28514 = pi18 ? n28382 : ~n1676;
  assign n28515 = pi17 ? n32 : n28514;
  assign n28516 = pi16 ? n32 : n28515;
  assign n28517 = pi15 ? n17891 : n28516;
  assign n28518 = pi14 ? n28513 : n28517;
  assign n28519 = pi19 ? n11374 : n322;
  assign n28520 = pi18 ? n28519 : n32;
  assign n28521 = pi17 ? n3282 : n28520;
  assign n28522 = pi16 ? n32 : n28521;
  assign n28523 = pi15 ? n32 : n28522;
  assign n28524 = pi14 ? n17891 : n28523;
  assign n28525 = pi13 ? n28518 : n28524;
  assign n28526 = pi15 ? n18019 : n18326;
  assign n28527 = pi14 ? n28526 : n28396;
  assign n28528 = pi13 ? n28527 : n28398;
  assign n28529 = pi12 ? n28525 : n28528;
  assign n28530 = pi19 ? n322 : n2092;
  assign n28531 = pi18 ? n28530 : n32;
  assign n28532 = pi17 ? n32 : n28531;
  assign n28533 = pi16 ? n32 : n28532;
  assign n28534 = pi15 ? n28533 : n17856;
  assign n28535 = pi14 ? n28534 : n32;
  assign n28536 = pi20 ? n20944 : n354;
  assign n28537 = pi19 ? n20006 : ~n28536;
  assign n28538 = pi20 ? n333 : n428;
  assign n28539 = pi20 ? n3523 : n428;
  assign n28540 = pi19 ? n28538 : n28539;
  assign n28541 = pi18 ? n28537 : n28540;
  assign n28542 = pi20 ? n19554 : n207;
  assign n28543 = pi19 ? n28542 : ~n32;
  assign n28544 = pi18 ? n28543 : ~n32;
  assign n28545 = pi17 ? n28541 : ~n28544;
  assign n28546 = pi16 ? n278 : n28545;
  assign n28547 = pi15 ? n32 : n28546;
  assign n28548 = pi18 ? n23571 : n4671;
  assign n28549 = pi19 ? n4126 : n28451;
  assign n28550 = pi18 ? n28549 : ~n32;
  assign n28551 = pi17 ? n28548 : n28550;
  assign n28552 = pi16 ? n28449 : ~n28551;
  assign n28553 = pi21 ? n313 : n173;
  assign n28554 = pi20 ? n32 : n28553;
  assign n28555 = pi19 ? n32 : n28554;
  assign n28556 = pi20 ? n9491 : ~n18624;
  assign n28557 = pi19 ? n28556 : n18761;
  assign n28558 = pi18 ? n28555 : ~n28557;
  assign n28559 = pi17 ? n32 : n28558;
  assign n28560 = pi20 ? n18073 : ~n174;
  assign n28561 = pi20 ? n19554 : n18073;
  assign n28562 = pi19 ? n28560 : ~n28561;
  assign n28563 = pi20 ? n13171 : ~n13171;
  assign n28564 = pi18 ? n28562 : n28563;
  assign n28565 = pi20 ? n309 : n32;
  assign n28566 = pi19 ? n28565 : n208;
  assign n28567 = pi18 ? n28566 : ~n32;
  assign n28568 = pi17 ? n28564 : ~n28567;
  assign n28569 = pi16 ? n28559 : n28568;
  assign n28570 = pi15 ? n28552 : n28569;
  assign n28571 = pi14 ? n28547 : n28570;
  assign n28572 = pi13 ? n28535 : n28571;
  assign n28573 = pi12 ? n28439 : n28572;
  assign n28574 = pi11 ? n28529 : n28573;
  assign n28575 = pi10 ? n28511 : n28574;
  assign n28576 = pi09 ? n32 : n28575;
  assign n28577 = pi08 ? n28467 : n28576;
  assign n28578 = pi20 ? n3523 : ~n339;
  assign n28579 = pi19 ? n32 : n28578;
  assign n28580 = pi20 ? n2358 : n9491;
  assign n28581 = pi19 ? n28580 : ~n311;
  assign n28582 = pi18 ? n28579 : ~n28581;
  assign n28583 = pi20 ? n310 : ~n18073;
  assign n28584 = pi19 ? n28583 : ~n501;
  assign n28585 = pi18 ? n28584 : n32;
  assign n28586 = pi17 ? n28582 : n28585;
  assign n28587 = pi16 ? n32 : n28586;
  assign n28588 = pi15 ? n32 : n28587;
  assign n28589 = pi14 ? n32 : n28588;
  assign n28590 = pi13 ? n28589 : n32;
  assign n28591 = pi12 ? n32 : n28590;
  assign n28592 = pi15 ? n18008 : n17997;
  assign n28593 = pi14 ? n32 : n28592;
  assign n28594 = pi14 ? n17997 : n19913;
  assign n28595 = pi13 ? n28593 : n28594;
  assign n28596 = pi18 ? n4380 : n18242;
  assign n28597 = pi17 ? n32 : n28596;
  assign n28598 = pi18 ? n18249 : n32;
  assign n28599 = pi17 ? n18248 : ~n28598;
  assign n28600 = pi16 ? n28597 : ~n28599;
  assign n28601 = pi15 ? n28600 : n32;
  assign n28602 = pi19 ? n18390 : n32;
  assign n28603 = pi18 ? n28602 : ~n3350;
  assign n28604 = pi17 ? n32 : n28603;
  assign n28605 = pi16 ? n32 : n28604;
  assign n28606 = pi15 ? n32 : n28605;
  assign n28607 = pi14 ? n28601 : n28606;
  assign n28608 = pi18 ? n18397 : ~n618;
  assign n28609 = pi17 ? n18395 : n28608;
  assign n28610 = pi16 ? n32 : n28609;
  assign n28611 = pi15 ? n28610 : n18008;
  assign n28612 = pi15 ? n18008 : n32;
  assign n28613 = pi14 ? n28611 : n28612;
  assign n28614 = pi13 ? n28607 : n28613;
  assign n28615 = pi12 ? n28595 : n28614;
  assign n28616 = pi11 ? n28591 : n28615;
  assign n28617 = pi19 ? n19601 : ~n342;
  assign n28618 = pi18 ? n28617 : n1676;
  assign n28619 = pi17 ? n16982 : ~n28618;
  assign n28620 = pi16 ? n32 : n28619;
  assign n28621 = pi15 ? n17891 : n28620;
  assign n28622 = pi14 ? n32 : n28621;
  assign n28623 = pi20 ? n342 : n206;
  assign n28624 = pi19 ? n32 : n28623;
  assign n28625 = pi18 ? n28624 : n32;
  assign n28626 = pi17 ? n32 : n28625;
  assign n28627 = pi16 ? n32 : n28626;
  assign n28628 = pi15 ? n28627 : n17903;
  assign n28629 = pi14 ? n17891 : n28628;
  assign n28630 = pi13 ? n28622 : n28629;
  assign n28631 = pi14 ? n32 : n28396;
  assign n28632 = pi16 ? n32 : n224;
  assign n28633 = pi15 ? n28632 : n32;
  assign n28634 = pi15 ? n32 : n17851;
  assign n28635 = pi14 ? n28633 : n28634;
  assign n28636 = pi13 ? n28631 : n28635;
  assign n28637 = pi12 ? n28630 : n28636;
  assign n28638 = pi18 ? n16981 : n32;
  assign n28639 = pi20 ? n749 : ~n339;
  assign n28640 = pi19 ? n32 : n28639;
  assign n28641 = pi18 ? n28640 : n32;
  assign n28642 = pi17 ? n28638 : n28641;
  assign n28643 = pi16 ? n32 : n28642;
  assign n28644 = pi18 ? n15400 : n32;
  assign n28645 = pi17 ? n32 : n28644;
  assign n28646 = pi16 ? n32 : n28645;
  assign n28647 = pi15 ? n28643 : n28646;
  assign n28648 = pi14 ? n32 : n28647;
  assign n28649 = pi19 ? n507 : ~n1248;
  assign n28650 = pi18 ? n28649 : n32;
  assign n28651 = pi17 ? n32 : n28650;
  assign n28652 = pi16 ? n32 : n28651;
  assign n28653 = pi19 ? n208 : ~n519;
  assign n28654 = pi18 ? n28653 : n32;
  assign n28655 = pi17 ? n32 : n28654;
  assign n28656 = pi16 ? n32 : n28655;
  assign n28657 = pi15 ? n28652 : n28656;
  assign n28658 = pi19 ? n208 : ~n208;
  assign n28659 = pi18 ? n28658 : n32;
  assign n28660 = pi17 ? n32 : n28659;
  assign n28661 = pi16 ? n32 : n28660;
  assign n28662 = pi17 ? n32 : n28434;
  assign n28663 = pi16 ? n32 : n28662;
  assign n28664 = pi15 ? n28661 : n28663;
  assign n28665 = pi14 ? n28657 : n28664;
  assign n28666 = pi13 ? n28648 : n28665;
  assign n28667 = pi19 ? n208 : n358;
  assign n28668 = pi18 ? n28667 : n32;
  assign n28669 = pi17 ? n32 : n28668;
  assign n28670 = pi16 ? n32 : n28669;
  assign n28671 = pi15 ? n28670 : n32;
  assign n28672 = pi14 ? n28671 : n32;
  assign n28673 = pi21 ? n1392 : ~n206;
  assign n28674 = pi20 ? n32 : n28673;
  assign n28675 = pi19 ? n32 : n28674;
  assign n28676 = pi18 ? n28675 : ~n32;
  assign n28677 = pi17 ? n32 : n28676;
  assign n28678 = pi19 ? n236 : ~n5004;
  assign n28679 = pi18 ? n28678 : ~n32;
  assign n28680 = pi17 ? n18213 : n28679;
  assign n28681 = pi16 ? n28677 : ~n28680;
  assign n28682 = pi19 ? n23895 : ~n207;
  assign n28683 = pi18 ? n18199 : ~n28682;
  assign n28684 = pi17 ? n32 : n28683;
  assign n28685 = pi20 ? n220 : ~n206;
  assign n28686 = pi20 ? n206 : n266;
  assign n28687 = pi19 ? n28685 : ~n28686;
  assign n28688 = pi18 ? n28687 : n28041;
  assign n28689 = pi19 ? n22185 : ~n750;
  assign n28690 = pi18 ? n28689 : n32;
  assign n28691 = pi17 ? n28688 : n28690;
  assign n28692 = pi16 ? n28684 : n28691;
  assign n28693 = pi15 ? n28681 : n28692;
  assign n28694 = pi14 ? n32 : n28693;
  assign n28695 = pi13 ? n28672 : n28694;
  assign n28696 = pi12 ? n28666 : n28695;
  assign n28697 = pi11 ? n28637 : n28696;
  assign n28698 = pi10 ? n28616 : n28697;
  assign n28699 = pi09 ? n32 : n28698;
  assign n28700 = pi18 ? n28584 : n18076;
  assign n28701 = pi17 ? n28582 : n28700;
  assign n28702 = pi16 ? n32 : n28701;
  assign n28703 = pi15 ? n32 : n28702;
  assign n28704 = pi14 ? n32 : n28703;
  assign n28705 = pi14 ? n32 : n18585;
  assign n28706 = pi13 ? n28704 : n28705;
  assign n28707 = pi12 ? n32 : n28706;
  assign n28708 = pi15 ? n19172 : n18294;
  assign n28709 = pi14 ? n18585 : n28708;
  assign n28710 = pi15 ? n18294 : n18008;
  assign n28711 = pi14 ? n18294 : n28710;
  assign n28712 = pi13 ? n28709 : n28711;
  assign n28713 = pi18 ? n28602 : ~n237;
  assign n28714 = pi17 ? n32 : n28713;
  assign n28715 = pi16 ? n32 : n28714;
  assign n28716 = pi15 ? n32 : n28715;
  assign n28717 = pi14 ? n28601 : n28716;
  assign n28718 = pi16 ? n18561 : n28609;
  assign n28719 = pi15 ? n28718 : n18008;
  assign n28720 = pi15 ? n18297 : n32;
  assign n28721 = pi14 ? n28719 : n28720;
  assign n28722 = pi13 ? n28717 : n28721;
  assign n28723 = pi12 ? n28712 : n28722;
  assign n28724 = pi11 ? n28707 : n28723;
  assign n28725 = pi18 ? n28617 : n618;
  assign n28726 = pi17 ? n16982 : ~n28725;
  assign n28727 = pi16 ? n32 : n28726;
  assign n28728 = pi15 ? n18439 : n28727;
  assign n28729 = pi14 ? n18143 : n28728;
  assign n28730 = pi18 ? n28624 : ~n1676;
  assign n28731 = pi17 ? n32 : n28730;
  assign n28732 = pi16 ? n32 : n28731;
  assign n28733 = pi15 ? n28732 : n17891;
  assign n28734 = pi14 ? n18439 : n28733;
  assign n28735 = pi13 ? n28729 : n28734;
  assign n28736 = pi12 ? n28735 : n28636;
  assign n28737 = pi17 ? n32 : n28641;
  assign n28738 = pi16 ? n32 : n28737;
  assign n28739 = pi20 ? n207 : n111;
  assign n28740 = pi19 ? n32 : n28739;
  assign n28741 = pi18 ? n28740 : n32;
  assign n28742 = pi17 ? n32 : n28741;
  assign n28743 = pi16 ? n32 : n28742;
  assign n28744 = pi15 ? n28738 : n28743;
  assign n28745 = pi14 ? n32 : n28744;
  assign n28746 = pi21 ? n8275 : n206;
  assign n28747 = pi20 ? n32 : n28746;
  assign n28748 = pi19 ? n32 : n28747;
  assign n28749 = pi20 ? n18073 : n17671;
  assign n28750 = pi20 ? n6822 : n333;
  assign n28751 = pi19 ? n28749 : n28750;
  assign n28752 = pi18 ? n28748 : n28751;
  assign n28753 = pi17 ? n32 : n28752;
  assign n28754 = pi20 ? n18073 : n4279;
  assign n28755 = pi20 ? n6621 : n313;
  assign n28756 = pi19 ? n28754 : n28755;
  assign n28757 = pi20 ? n18624 : n18415;
  assign n28758 = pi20 ? n17669 : ~n18415;
  assign n28759 = pi19 ? n28757 : ~n28758;
  assign n28760 = pi18 ? n28756 : ~n28759;
  assign n28761 = pi21 ? n309 : n313;
  assign n28762 = pi20 ? n28761 : n357;
  assign n28763 = pi19 ? n28762 : n519;
  assign n28764 = pi18 ? n28763 : ~n32;
  assign n28765 = pi17 ? n28760 : n28764;
  assign n28766 = pi16 ? n28753 : ~n28765;
  assign n28767 = pi15 ? n28652 : n28766;
  assign n28768 = pi21 ? n124 : n174;
  assign n28769 = pi20 ? n32 : n28768;
  assign n28770 = pi19 ? n32 : n28769;
  assign n28771 = pi19 ? n18574 : n21107;
  assign n28772 = pi18 ? n28770 : n28771;
  assign n28773 = pi17 ? n32 : n28772;
  assign n28774 = pi20 ? n333 : ~n18834;
  assign n28775 = pi20 ? n18624 : n313;
  assign n28776 = pi19 ? n28774 : ~n28775;
  assign n28777 = pi20 ? n18337 : n18073;
  assign n28778 = pi20 ? n6621 : n18073;
  assign n28779 = pi19 ? n28777 : n28778;
  assign n28780 = pi18 ? n28776 : n28779;
  assign n28781 = pi20 ? n18256 : ~n357;
  assign n28782 = pi19 ? n28781 : ~n208;
  assign n28783 = pi18 ? n28782 : n32;
  assign n28784 = pi17 ? n28780 : n28783;
  assign n28785 = pi16 ? n28773 : n28784;
  assign n28786 = pi20 ? n11107 : n207;
  assign n28787 = pi19 ? n28786 : ~n349;
  assign n28788 = pi18 ? n28787 : n32;
  assign n28789 = pi17 ? n28780 : n28788;
  assign n28790 = pi16 ? n28773 : n28789;
  assign n28791 = pi15 ? n28785 : n28790;
  assign n28792 = pi14 ? n28767 : n28791;
  assign n28793 = pi13 ? n28745 : n28792;
  assign n28794 = pi19 ? n18919 : n21107;
  assign n28795 = pi18 ? n28770 : n28794;
  assign n28796 = pi17 ? n32 : n28795;
  assign n28797 = pi19 ? n28786 : n358;
  assign n28798 = pi18 ? n28797 : n32;
  assign n28799 = pi17 ? n28780 : n28798;
  assign n28800 = pi16 ? n28796 : n28799;
  assign n28801 = pi15 ? n28800 : n32;
  assign n28802 = pi14 ? n28801 : n32;
  assign n28803 = pi18 ? n222 : ~n32;
  assign n28804 = pi17 ? n32 : n28803;
  assign n28805 = pi16 ? n28804 : ~n28680;
  assign n28806 = pi18 ? n4127 : ~n28682;
  assign n28807 = pi17 ? n32 : n28806;
  assign n28808 = pi16 ? n28807 : n28691;
  assign n28809 = pi15 ? n28805 : n28808;
  assign n28810 = pi14 ? n32 : n28809;
  assign n28811 = pi13 ? n28802 : n28810;
  assign n28812 = pi12 ? n28793 : n28811;
  assign n28813 = pi11 ? n28736 : n28812;
  assign n28814 = pi10 ? n28724 : n28813;
  assign n28815 = pi09 ? n32 : n28814;
  assign n28816 = pi08 ? n28699 : n28815;
  assign n28817 = pi07 ? n28577 : n28816;
  assign n28818 = pi18 ? n32 : n21194;
  assign n28819 = pi17 ? n32 : n28818;
  assign n28820 = pi20 ? n32 : n9194;
  assign n28821 = pi19 ? n32 : n28820;
  assign n28822 = pi20 ? n1368 : n428;
  assign n28823 = pi20 ? n9194 : n6085;
  assign n28824 = pi19 ? n28822 : n28823;
  assign n28825 = pi18 ? n28821 : n28824;
  assign n28826 = pi20 ? n6085 : n357;
  assign n28827 = pi19 ? n28826 : n4491;
  assign n28828 = pi18 ? n28827 : n32;
  assign n28829 = pi17 ? n28825 : n28828;
  assign n28830 = pi16 ? n28819 : n28829;
  assign n28831 = pi15 ? n28830 : n32;
  assign n28832 = pi14 ? n28831 : n32;
  assign n28833 = pi20 ? n175 : n357;
  assign n28834 = pi19 ? n28833 : n4491;
  assign n28835 = pi18 ? n28834 : n32;
  assign n28836 = pi17 ? n17661 : n28835;
  assign n28837 = pi16 ? n32 : n28836;
  assign n28838 = pi15 ? n32 : n28837;
  assign n28839 = pi14 ? n32 : n28838;
  assign n28840 = pi13 ? n28832 : n28839;
  assign n28841 = pi12 ? n32 : n28840;
  assign n28842 = pi20 ? n18253 : n18255;
  assign n28843 = pi19 ? n18261 : ~n28842;
  assign n28844 = pi18 ? n4519 : n28843;
  assign n28845 = pi17 ? n32 : n28844;
  assign n28846 = pi20 ? n18256 : n3695;
  assign n28847 = pi20 ? n3695 : n820;
  assign n28848 = pi19 ? n28846 : n28847;
  assign n28849 = pi20 ? n820 : n1385;
  assign n28850 = pi20 ? n18261 : ~n5854;
  assign n28851 = pi19 ? n28849 : n28850;
  assign n28852 = pi18 ? n28848 : n28851;
  assign n28853 = pi20 ? n274 : n206;
  assign n28854 = pi20 ? n785 : n1685;
  assign n28855 = pi19 ? n28853 : ~n28854;
  assign n28856 = pi18 ? n28855 : ~n54;
  assign n28857 = pi17 ? n28852 : ~n28856;
  assign n28858 = pi16 ? n28845 : n28857;
  assign n28859 = pi15 ? n32 : n28858;
  assign n28860 = pi20 ? n3695 : n448;
  assign n28861 = pi19 ? n28846 : n28860;
  assign n28862 = pi20 ? n18261 : n2385;
  assign n28863 = pi19 ? n18785 : n28862;
  assign n28864 = pi18 ? n28861 : n28863;
  assign n28865 = pi19 ? n18116 : n1685;
  assign n28866 = pi18 ? n28865 : n54;
  assign n28867 = pi17 ? n28864 : n28866;
  assign n28868 = pi16 ? n28845 : n28867;
  assign n28869 = pi18 ? n858 : n28843;
  assign n28870 = pi17 ? n32 : n28869;
  assign n28871 = pi20 ? n357 : n448;
  assign n28872 = pi19 ? n28846 : n28871;
  assign n28873 = pi20 ? n18261 : n342;
  assign n28874 = pi19 ? n28483 : n28873;
  assign n28875 = pi18 ? n28872 : n28874;
  assign n28876 = pi19 ? n32 : n1817;
  assign n28877 = pi18 ? n28876 : n54;
  assign n28878 = pi17 ? n28875 : n28877;
  assign n28879 = pi16 ? n28870 : n28878;
  assign n28880 = pi15 ? n28868 : n28879;
  assign n28881 = pi14 ? n28859 : n28880;
  assign n28882 = pi15 ? n57 : n19166;
  assign n28883 = pi14 ? n28882 : n57;
  assign n28884 = pi13 ? n28881 : n28883;
  assign n28885 = pi14 ? n57 : n28882;
  assign n28886 = pi19 ? n18403 : ~n18678;
  assign n28887 = pi18 ? n18908 : n28886;
  assign n28888 = pi17 ? n32 : n28887;
  assign n28889 = pi20 ? n266 : n310;
  assign n28890 = pi19 ? n9007 : n28889;
  assign n28891 = pi19 ? n6314 : n28152;
  assign n28892 = pi18 ? n28890 : n28891;
  assign n28893 = pi20 ? n2358 : n339;
  assign n28894 = pi19 ? n28893 : ~n175;
  assign n28895 = pi18 ? n28894 : ~n237;
  assign n28896 = pi17 ? n28892 : ~n28895;
  assign n28897 = pi16 ? n28888 : ~n28896;
  assign n28898 = pi20 ? n9488 : ~n2180;
  assign n28899 = pi19 ? n28898 : ~n9491;
  assign n28900 = pi20 ? n9491 : ~n3843;
  assign n28901 = pi19 ? n28900 : n9491;
  assign n28902 = pi18 ? n28899 : ~n28901;
  assign n28903 = pi20 ? n9491 : n339;
  assign n28904 = pi19 ? n28903 : ~n9488;
  assign n28905 = pi18 ? n28904 : ~n3350;
  assign n28906 = pi17 ? n28902 : ~n28905;
  assign n28907 = pi16 ? n18938 : ~n28906;
  assign n28908 = pi15 ? n28897 : n28907;
  assign n28909 = pi14 ? n28908 : n18304;
  assign n28910 = pi13 ? n28885 : n28909;
  assign n28911 = pi12 ? n28884 : n28910;
  assign n28912 = pi11 ? n28841 : n28911;
  assign n28913 = pi19 ? n349 : ~n342;
  assign n28914 = pi18 ? n28913 : ~n32;
  assign n28915 = pi17 ? n32 : ~n28914;
  assign n28916 = pi16 ? n32 : n28915;
  assign n28917 = pi15 ? n32 : n28916;
  assign n28918 = pi20 ? n3523 : ~n342;
  assign n28919 = pi19 ? n32 : n28918;
  assign n28920 = pi18 ? n32 : n28919;
  assign n28921 = pi18 ? n5657 : n618;
  assign n28922 = pi17 ? n28920 : ~n28921;
  assign n28923 = pi16 ? n32 : n28922;
  assign n28924 = pi15 ? n28923 : n18439;
  assign n28925 = pi14 ? n28917 : n28924;
  assign n28926 = pi20 ? n428 : n342;
  assign n28927 = pi19 ? n32 : n28926;
  assign n28928 = pi18 ? n28927 : ~n618;
  assign n28929 = pi17 ? n32 : n28928;
  assign n28930 = pi16 ? n32 : n28929;
  assign n28931 = pi15 ? n28930 : n18594;
  assign n28932 = pi14 ? n28931 : n18005;
  assign n28933 = pi13 ? n28925 : n28932;
  assign n28934 = pi15 ? n17903 : n18326;
  assign n28935 = pi14 ? n18827 : n28934;
  assign n28936 = pi14 ? n32 : n28634;
  assign n28937 = pi13 ? n28935 : n28936;
  assign n28938 = pi12 ? n28933 : n28937;
  assign n28939 = pi17 ? n32 : n28415;
  assign n28940 = pi16 ? n32 : n28939;
  assign n28941 = pi19 ? n507 : ~n4721;
  assign n28942 = pi18 ? n28941 : n32;
  assign n28943 = pi17 ? n32 : n28942;
  assign n28944 = pi16 ? n32 : n28943;
  assign n28945 = pi15 ? n28940 : n28944;
  assign n28946 = pi14 ? n17852 : n28945;
  assign n28947 = pi16 ? n1135 : ~n1581;
  assign n28948 = pi18 ? n341 : ~n6145;
  assign n28949 = pi17 ? n32 : n28948;
  assign n28950 = pi16 ? n28949 : ~n1471;
  assign n28951 = pi15 ? n28947 : n28950;
  assign n28952 = pi20 ? n206 : n321;
  assign n28953 = pi19 ? n28952 : n6997;
  assign n28954 = pi18 ? n4127 : ~n28953;
  assign n28955 = pi17 ? n32 : n28954;
  assign n28956 = pi19 ? n4391 : ~n4126;
  assign n28957 = pi20 ? n266 : ~n206;
  assign n28958 = pi19 ? n20006 : n28957;
  assign n28959 = pi18 ? n28956 : ~n28958;
  assign n28960 = pi19 ? n28686 : n343;
  assign n28961 = pi18 ? n28960 : ~n32;
  assign n28962 = pi17 ? n28959 : ~n28961;
  assign n28963 = pi16 ? n28955 : n28962;
  assign n28964 = pi20 ? n18173 : n2358;
  assign n28965 = pi20 ? n2358 : ~n18129;
  assign n28966 = pi19 ? n28964 : n28965;
  assign n28967 = pi18 ? n18331 : ~n28966;
  assign n28968 = pi17 ? n32 : n28967;
  assign n28969 = pi20 ? n1076 : n21111;
  assign n28970 = pi20 ? n405 : n206;
  assign n28971 = pi19 ? n28969 : ~n28970;
  assign n28972 = pi20 ? n309 : ~n6621;
  assign n28973 = pi20 ? n310 : ~n6621;
  assign n28974 = pi19 ? n28972 : n28973;
  assign n28975 = pi18 ? n28971 : ~n28974;
  assign n28976 = pi20 ? n206 : n915;
  assign n28977 = pi19 ? n28976 : ~n5614;
  assign n28978 = pi18 ? n28977 : ~n32;
  assign n28979 = pi17 ? n28975 : ~n28978;
  assign n28980 = pi16 ? n28968 : n28979;
  assign n28981 = pi15 ? n28963 : n28980;
  assign n28982 = pi14 ? n28951 : n28981;
  assign n28983 = pi13 ? n28946 : n28982;
  assign n28984 = pi18 ? n32 : n28032;
  assign n28985 = pi17 ? n32 : n28984;
  assign n28986 = pi18 ? n4380 : ~n18503;
  assign n28987 = pi19 ? n32 : n7642;
  assign n28988 = pi18 ? n28987 : n32;
  assign n28989 = pi17 ? n28986 : n28988;
  assign n28990 = pi16 ? n28985 : n28989;
  assign n28991 = pi15 ? n32 : n28990;
  assign n28992 = pi16 ? n1214 : ~n1471;
  assign n28993 = pi17 ? n32 : n5699;
  assign n28994 = pi16 ? n28993 : ~n1471;
  assign n28995 = pi15 ? n28992 : n28994;
  assign n28996 = pi14 ? n28991 : n28995;
  assign n28997 = pi13 ? n32 : n28996;
  assign n28998 = pi12 ? n28983 : n28997;
  assign n28999 = pi11 ? n28938 : n28998;
  assign n29000 = pi10 ? n28912 : n28999;
  assign n29001 = pi09 ? n32 : n29000;
  assign n29002 = pi20 ? n1817 : n428;
  assign n29003 = pi20 ? n1817 : n357;
  assign n29004 = pi19 ? n29002 : n29003;
  assign n29005 = pi18 ? n1819 : n29004;
  assign n29006 = pi17 ? n29005 : n1124;
  assign n29007 = pi16 ? n32 : n29006;
  assign n29008 = pi15 ? n29007 : n32;
  assign n29009 = pi14 ? n29008 : n32;
  assign n29010 = pi18 ? n18520 : ~n18532;
  assign n29011 = pi17 ? n18518 : ~n29010;
  assign n29012 = pi16 ? n32 : n29011;
  assign n29013 = pi15 ? n32 : n29012;
  assign n29014 = pi14 ? n32 : n29013;
  assign n29015 = pi13 ? n29009 : n29014;
  assign n29016 = pi12 ? n32 : n29015;
  assign n29017 = pi19 ? n1611 : n18095;
  assign n29018 = pi18 ? n4380 : n29017;
  assign n29019 = pi17 ? n32 : n29018;
  assign n29020 = pi20 ? n12884 : n2358;
  assign n29021 = pi19 ? n18099 : n29020;
  assign n29022 = pi20 ? n2358 : n246;
  assign n29023 = pi20 ? n1611 : ~n220;
  assign n29024 = pi19 ? n29022 : n29023;
  assign n29025 = pi18 ? n29021 : n29024;
  assign n29026 = pi19 ? n17757 : ~n28686;
  assign n29027 = pi18 ? n29026 : ~n32;
  assign n29028 = pi17 ? n29025 : ~n29027;
  assign n29029 = pi16 ? n29019 : n29028;
  assign n29030 = pi15 ? n32 : n29029;
  assign n29031 = pi20 ? n12884 : n357;
  assign n29032 = pi19 ? n18099 : n29031;
  assign n29033 = pi20 ? n1611 : n342;
  assign n29034 = pi19 ? n18665 : n29033;
  assign n29035 = pi18 ? n29032 : n29034;
  assign n29036 = pi19 ? n4670 : n266;
  assign n29037 = pi18 ? n29036 : n32;
  assign n29038 = pi17 ? n29035 : n29037;
  assign n29039 = pi16 ? n29019 : n29038;
  assign n29040 = pi18 ? n32 : n29017;
  assign n29041 = pi17 ? n32 : n29040;
  assign n29042 = pi19 ? n18099 : n357;
  assign n29043 = pi19 ? n32 : n29033;
  assign n29044 = pi18 ? n29042 : n29043;
  assign n29045 = pi17 ? n29044 : n32;
  assign n29046 = pi16 ? n29041 : n29045;
  assign n29047 = pi15 ? n29039 : n29046;
  assign n29048 = pi14 ? n29030 : n29047;
  assign n29049 = pi15 ? n32 : n19166;
  assign n29050 = pi15 ? n57 : n32;
  assign n29051 = pi14 ? n29049 : n29050;
  assign n29052 = pi13 ? n29048 : n29051;
  assign n29053 = pi16 ? n18561 : n18687;
  assign n29054 = pi16 ? n18561 : n19165;
  assign n29055 = pi15 ? n29053 : n29054;
  assign n29056 = pi14 ? n32 : n29055;
  assign n29057 = pi20 ? n17665 : n9194;
  assign n29058 = pi19 ? n29057 : ~n18678;
  assign n29059 = pi18 ? n32 : n29058;
  assign n29060 = pi17 ? n32 : n29059;
  assign n29061 = pi16 ? n29060 : ~n28896;
  assign n29062 = pi18 ? n28904 : ~n237;
  assign n29063 = pi17 ? n28902 : ~n29062;
  assign n29064 = pi16 ? n19048 : ~n29063;
  assign n29065 = pi15 ? n29061 : n29064;
  assign n29066 = pi14 ? n29065 : n18590;
  assign n29067 = pi13 ? n29056 : n29066;
  assign n29068 = pi12 ? n29052 : n29067;
  assign n29069 = pi11 ? n29016 : n29068;
  assign n29070 = pi18 ? n28913 : ~n18076;
  assign n29071 = pi17 ? n32 : ~n29070;
  assign n29072 = pi16 ? n32 : n29071;
  assign n29073 = pi15 ? n18142 : n29072;
  assign n29074 = pi15 ? n28923 : n18594;
  assign n29075 = pi14 ? n29073 : n29074;
  assign n29076 = pi18 ? n28927 : ~n3350;
  assign n29077 = pi17 ? n32 : n29076;
  assign n29078 = pi16 ? n32 : n29077;
  assign n29079 = pi15 ? n29078 : n18594;
  assign n29080 = pi14 ? n29079 : n18005;
  assign n29081 = pi13 ? n29075 : n29080;
  assign n29082 = pi14 ? n18019 : n28934;
  assign n29083 = pi13 ? n29082 : n28936;
  assign n29084 = pi12 ? n29081 : n29083;
  assign n29085 = pi20 ? n32 : n18408;
  assign n29086 = pi19 ? n32 : n29085;
  assign n29087 = pi20 ? n333 : ~n18832;
  assign n29088 = pi19 ? n18621 : n29087;
  assign n29089 = pi18 ? n29086 : n29088;
  assign n29090 = pi17 ? n32 : n29089;
  assign n29091 = pi19 ? n18621 : n18339;
  assign n29092 = pi20 ? n18337 : ~n6621;
  assign n29093 = pi20 ? n18073 : ~n17669;
  assign n29094 = pi19 ? n29092 : ~n29093;
  assign n29095 = pi18 ? n29091 : ~n29094;
  assign n29096 = pi20 ? n17665 : ~n4279;
  assign n29097 = pi19 ? n29096 : n4721;
  assign n29098 = pi18 ? n29097 : ~n32;
  assign n29099 = pi17 ? n29095 : n29098;
  assign n29100 = pi16 ? n29090 : ~n29099;
  assign n29101 = pi15 ? n28940 : n29100;
  assign n29102 = pi14 ? n17852 : n29101;
  assign n29103 = pi20 ? n3523 : ~n2358;
  assign n29104 = pi19 ? n29103 : ~n28965;
  assign n29105 = pi18 ? n18331 : n29104;
  assign n29106 = pi17 ? n32 : n29105;
  assign n29107 = pi20 ? n206 : n287;
  assign n29108 = pi19 ? n17644 : ~n29107;
  assign n29109 = pi20 ? n12884 : ~n174;
  assign n29110 = pi20 ? n310 : ~n174;
  assign n29111 = pi19 ? n29109 : n29110;
  assign n29112 = pi18 ? n29108 : ~n29111;
  assign n29113 = pi20 ? n287 : n623;
  assign n29114 = pi19 ? n29113 : ~n5614;
  assign n29115 = pi18 ? n29114 : ~n32;
  assign n29116 = pi17 ? n29112 : ~n29115;
  assign n29117 = pi16 ? n29106 : n29116;
  assign n29118 = pi15 ? n28963 : n29117;
  assign n29119 = pi14 ? n28951 : n29118;
  assign n29120 = pi13 ? n29102 : n29119;
  assign n29121 = pi14 ? n17852 : n32;
  assign n29122 = pi13 ? n29121 : n28996;
  assign n29123 = pi12 ? n29120 : n29122;
  assign n29124 = pi11 ? n29084 : n29123;
  assign n29125 = pi10 ? n29069 : n29124;
  assign n29126 = pi09 ? n32 : n29125;
  assign n29127 = pi08 ? n29001 : n29126;
  assign n29128 = pi14 ? n32 : n18661;
  assign n29129 = pi13 ? n32 : n29128;
  assign n29130 = pi16 ? n20208 : ~n1815;
  assign n29131 = pi15 ? n32 : n29130;
  assign n29132 = pi14 ? n18661 : n29131;
  assign n29133 = pi13 ? n18661 : n29132;
  assign n29134 = pi12 ? n29129 : n29133;
  assign n29135 = pi16 ? n20208 : ~n2137;
  assign n29136 = pi18 ? n6145 : n814;
  assign n29137 = pi17 ? n13946 : n29136;
  assign n29138 = pi16 ? n1471 : ~n29137;
  assign n29139 = pi15 ? n29135 : n29138;
  assign n29140 = pi19 ? n32 : n23644;
  assign n29141 = pi18 ? n940 : ~n29140;
  assign n29142 = pi17 ? n32 : n29141;
  assign n29143 = pi20 ? n5854 : n428;
  assign n29144 = pi19 ? n4670 : ~n29143;
  assign n29145 = pi20 ? n428 : n5854;
  assign n29146 = pi19 ? n29145 : n19598;
  assign n29147 = pi18 ? n29144 : ~n29146;
  assign n29148 = pi20 ? n357 : n310;
  assign n29149 = pi20 ? n2358 : n1611;
  assign n29150 = pi19 ? n29148 : ~n29149;
  assign n29151 = pi18 ? n29150 : ~n822;
  assign n29152 = pi17 ? n29147 : ~n29151;
  assign n29153 = pi16 ? n29142 : ~n29152;
  assign n29154 = pi15 ? n29153 : n18535;
  assign n29155 = pi14 ? n29139 : n29154;
  assign n29156 = pi14 ? n19334 : n32;
  assign n29157 = pi13 ? n29155 : n29156;
  assign n29158 = pi20 ? n9641 : n9194;
  assign n29159 = pi20 ? n9488 : ~n1611;
  assign n29160 = pi19 ? n29158 : n29159;
  assign n29161 = pi18 ? n1819 : n29160;
  assign n29162 = pi17 ? n32 : n29161;
  assign n29163 = pi16 ? n29162 : ~n2137;
  assign n29164 = pi18 ? n32 : n28071;
  assign n29165 = pi17 ? n32 : n29164;
  assign n29166 = pi20 ? n448 : ~n207;
  assign n29167 = pi19 ? n29166 : n267;
  assign n29168 = pi18 ? n29167 : n1757;
  assign n29169 = pi17 ? n29168 : n2136;
  assign n29170 = pi16 ? n29165 : ~n29169;
  assign n29171 = pi15 ? n29163 : n29170;
  assign n29172 = pi14 ? n32 : n29171;
  assign n29173 = pi20 ? n974 : n2180;
  assign n29174 = pi19 ? n29173 : n9491;
  assign n29175 = pi19 ? n9491 : n9194;
  assign n29176 = pi18 ? n29174 : n29175;
  assign n29177 = pi19 ? n28356 : n17652;
  assign n29178 = pi18 ? n29177 : n359;
  assign n29179 = pi17 ? n29176 : n29178;
  assign n29180 = pi16 ? n32 : n29179;
  assign n29181 = pi15 ? n29180 : n18294;
  assign n29182 = pi14 ? n29181 : n18590;
  assign n29183 = pi13 ? n29172 : n29182;
  assign n29184 = pi12 ? n29157 : n29183;
  assign n29185 = pi11 ? n29134 : n29184;
  assign n29186 = pi20 ? n1076 : ~n266;
  assign n29187 = pi19 ? n349 : ~n29186;
  assign n29188 = pi18 ? n29187 : n618;
  assign n29189 = pi17 ? n23052 : ~n29188;
  assign n29190 = pi16 ? n32 : n29189;
  assign n29191 = pi15 ? n29190 : n28916;
  assign n29192 = pi19 ? n5614 : n343;
  assign n29193 = pi18 ? n29192 : ~n3350;
  assign n29194 = pi17 ? n3282 : n29193;
  assign n29195 = pi16 ? n32 : n29194;
  assign n29196 = pi15 ? n29195 : n19544;
  assign n29197 = pi14 ? n29191 : n29196;
  assign n29198 = pi15 ? n18439 : n32;
  assign n29199 = pi14 ? n18594 : n29198;
  assign n29200 = pi13 ? n29197 : n29199;
  assign n29201 = pi18 ? n18402 : n32;
  assign n29202 = pi17 ? n32 : n29201;
  assign n29203 = pi16 ? n32 : n29202;
  assign n29204 = pi15 ? n29203 : n17885;
  assign n29205 = pi15 ? n17885 : n28632;
  assign n29206 = pi14 ? n29204 : n29205;
  assign n29207 = pi15 ? n32 : n18326;
  assign n29208 = pi14 ? n32 : n29207;
  assign n29209 = pi13 ? n29206 : n29208;
  assign n29210 = pi12 ? n29200 : n29209;
  assign n29211 = pi20 ? n1611 : ~n207;
  assign n29212 = pi19 ? n32 : n29211;
  assign n29213 = pi18 ? n29212 : n32;
  assign n29214 = pi17 ? n32 : n29213;
  assign n29215 = pi16 ? n32 : n29214;
  assign n29216 = pi20 ? n915 : n220;
  assign n29217 = pi19 ? n9345 : ~n29216;
  assign n29218 = pi18 ? n940 : n29217;
  assign n29219 = pi17 ? n32 : n29218;
  assign n29220 = pi18 ? n248 : n32;
  assign n29221 = pi19 ? n4126 : n6298;
  assign n29222 = pi18 ? n29221 : ~n32;
  assign n29223 = pi17 ? n29220 : n29222;
  assign n29224 = pi16 ? n29219 : ~n29223;
  assign n29225 = pi15 ? n29215 : n29224;
  assign n29226 = pi19 ? n247 : ~n18502;
  assign n29227 = pi18 ? n222 : ~n29226;
  assign n29228 = pi17 ? n32 : n29227;
  assign n29229 = pi19 ? n1508 : n267;
  assign n29230 = pi18 ? n29229 : n28164;
  assign n29231 = pi19 ? n1757 : n18722;
  assign n29232 = pi18 ? n29231 : ~n32;
  assign n29233 = pi17 ? n29230 : n29232;
  assign n29234 = pi16 ? n29228 : ~n29233;
  assign n29235 = pi18 ? n18210 : n32;
  assign n29236 = pi17 ? n32 : n29235;
  assign n29237 = pi16 ? n32 : n29236;
  assign n29238 = pi15 ? n29234 : n29237;
  assign n29239 = pi14 ? n29225 : n29238;
  assign n29240 = pi16 ? n1214 : ~n1581;
  assign n29241 = pi19 ? n208 : ~n5688;
  assign n29242 = pi18 ? n29241 : n32;
  assign n29243 = pi17 ? n32 : n29242;
  assign n29244 = pi16 ? n32 : n29243;
  assign n29245 = pi15 ? n29240 : n29244;
  assign n29246 = pi19 ? n18728 : n32;
  assign n29247 = pi18 ? n32 : n29246;
  assign n29248 = pi17 ? n32 : n29247;
  assign n29249 = pi19 ? n18396 : n7642;
  assign n29250 = pi19 ? n1757 : ~n9345;
  assign n29251 = pi18 ? n29249 : n29250;
  assign n29252 = pi19 ? n15405 : n343;
  assign n29253 = pi18 ? n29252 : ~n32;
  assign n29254 = pi17 ? n29251 : ~n29253;
  assign n29255 = pi16 ? n29248 : n29254;
  assign n29256 = pi15 ? n29255 : n32;
  assign n29257 = pi14 ? n29245 : n29256;
  assign n29258 = pi13 ? n29239 : n29257;
  assign n29259 = pi20 ? n174 : n274;
  assign n29260 = pi19 ? n32 : n29259;
  assign n29261 = pi20 ? n357 : ~n831;
  assign n29262 = pi20 ? n32 : ~n831;
  assign n29263 = pi19 ? n29261 : n29262;
  assign n29264 = pi18 ? n29260 : n29263;
  assign n29265 = pi17 ? n29264 : n19904;
  assign n29266 = pi16 ? n19234 : n29265;
  assign n29267 = pi15 ? n32 : n29266;
  assign n29268 = pi14 ? n32 : n29267;
  assign n29269 = pi20 ? n246 : n6621;
  assign n29270 = pi20 ? n175 : ~n207;
  assign n29271 = pi19 ? n29269 : n29270;
  assign n29272 = pi18 ? n936 : n29271;
  assign n29273 = pi17 ? n32 : n29272;
  assign n29274 = pi20 ? n287 : ~n18073;
  assign n29275 = pi20 ? n785 : ~n12884;
  assign n29276 = pi19 ? n29274 : ~n29275;
  assign n29277 = pi20 ? n6621 : ~n206;
  assign n29278 = pi20 ? n18415 : ~n13171;
  assign n29279 = pi19 ? n29277 : ~n29278;
  assign n29280 = pi18 ? n29276 : ~n29279;
  assign n29281 = pi19 ? n21011 : ~n32;
  assign n29282 = pi18 ? n29281 : ~n32;
  assign n29283 = pi17 ? n29280 : n29282;
  assign n29284 = pi16 ? n29273 : ~n29283;
  assign n29285 = pi20 ? n9863 : n9491;
  assign n29286 = pi20 ? n1076 : n428;
  assign n29287 = pi19 ? n29285 : n29286;
  assign n29288 = pi18 ? n858 : n29287;
  assign n29289 = pi17 ? n32 : n29288;
  assign n29290 = pi20 ? n274 : ~n17669;
  assign n29291 = pi20 ? n405 : n2385;
  assign n29292 = pi19 ? n29290 : ~n29291;
  assign n29293 = pi20 ? n310 : n12884;
  assign n29294 = pi20 ? n5854 : ~n12884;
  assign n29295 = pi19 ? n29293 : ~n29294;
  assign n29296 = pi18 ? n29292 : ~n29295;
  assign n29297 = pi20 ? n5854 : ~n207;
  assign n29298 = pi20 ? n32 : ~n9863;
  assign n29299 = pi19 ? n29297 : ~n29298;
  assign n29300 = pi18 ? n29299 : n32;
  assign n29301 = pi17 ? n29296 : n29300;
  assign n29302 = pi16 ? n29289 : n29301;
  assign n29303 = pi15 ? n29284 : n29302;
  assign n29304 = pi18 ? n209 : ~n20164;
  assign n29305 = pi17 ? n32 : n29304;
  assign n29306 = pi16 ? n29305 : ~n1471;
  assign n29307 = pi15 ? n28992 : n29306;
  assign n29308 = pi14 ? n29303 : n29307;
  assign n29309 = pi13 ? n29268 : n29308;
  assign n29310 = pi12 ? n29258 : n29309;
  assign n29311 = pi11 ? n29210 : n29310;
  assign n29312 = pi10 ? n29185 : n29311;
  assign n29313 = pi09 ? n32 : n29312;
  assign n29314 = pi14 ? n32 : n18657;
  assign n29315 = pi13 ? n32 : n29314;
  assign n29316 = pi19 ? n32 : n14845;
  assign n29317 = pi18 ? n29316 : ~n32;
  assign n29318 = pi17 ? n32 : n29317;
  assign n29319 = pi16 ? n29318 : ~n2137;
  assign n29320 = pi15 ? n32 : n29319;
  assign n29321 = pi14 ? n18657 : n29320;
  assign n29322 = pi13 ? n18657 : n29321;
  assign n29323 = pi12 ? n29315 : n29322;
  assign n29324 = pi20 ? n32 : n17287;
  assign n29325 = pi19 ? n32 : n29324;
  assign n29326 = pi18 ? n29325 : ~n32;
  assign n29327 = pi17 ? n32 : n29326;
  assign n29328 = pi16 ? n29327 : ~n29137;
  assign n29329 = pi15 ? n29319 : n29328;
  assign n29330 = pi14 ? n29329 : n29154;
  assign n29331 = pi13 ? n29330 : n29156;
  assign n29332 = pi20 ? n18129 : ~n1611;
  assign n29333 = pi19 ? n857 : n29332;
  assign n29334 = pi18 ? n32 : n29333;
  assign n29335 = pi17 ? n32 : n29334;
  assign n29336 = pi16 ? n29335 : ~n2137;
  assign n29337 = pi16 ? n32 : ~n29169;
  assign n29338 = pi15 ? n29336 : n29337;
  assign n29339 = pi14 ? n32 : n29338;
  assign n29340 = pi20 ? n428 : n2180;
  assign n29341 = pi19 ? n29340 : n9491;
  assign n29342 = pi18 ? n29341 : n29175;
  assign n29343 = pi18 ? n29177 : n18425;
  assign n29344 = pi17 ? n29342 : n29343;
  assign n29345 = pi16 ? n32 : n29344;
  assign n29346 = pi15 ? n29345 : n18688;
  assign n29347 = pi15 ? n18688 : n32;
  assign n29348 = pi14 ? n29346 : n29347;
  assign n29349 = pi13 ? n29339 : n29348;
  assign n29350 = pi12 ? n29331 : n29349;
  assign n29351 = pi11 ? n29323 : n29350;
  assign n29352 = pi18 ? n29192 : ~n237;
  assign n29353 = pi17 ? n3282 : n29352;
  assign n29354 = pi16 ? n32 : n29353;
  assign n29355 = pi18 ? n1575 : ~n237;
  assign n29356 = pi17 ? n32 : n29355;
  assign n29357 = pi16 ? n32 : n29356;
  assign n29358 = pi15 ? n29354 : n29357;
  assign n29359 = pi14 ? n29191 : n29358;
  assign n29360 = pi14 ? n18814 : n29198;
  assign n29361 = pi13 ? n29359 : n29360;
  assign n29362 = pi12 ? n29361 : n29209;
  assign n29363 = pi20 ? n32 : n18282;
  assign n29364 = pi19 ? n32 : n29363;
  assign n29365 = pi20 ? n5854 : ~n18073;
  assign n29366 = pi20 ? n18256 : n17652;
  assign n29367 = pi19 ? n29365 : ~n29366;
  assign n29368 = pi18 ? n29364 : n29367;
  assign n29369 = pi17 ? n32 : n29368;
  assign n29370 = pi20 ? n6822 : ~n18073;
  assign n29371 = pi19 ? n29370 : ~n29275;
  assign n29372 = pi20 ? n20944 : ~n6621;
  assign n29373 = pi20 ? n18415 : ~n18415;
  assign n29374 = pi19 ? n29372 : ~n29373;
  assign n29375 = pi18 ? n29371 : ~n29374;
  assign n29376 = pi20 ? n7939 : ~n207;
  assign n29377 = pi19 ? n19555 : ~n29376;
  assign n29378 = pi18 ? n29377 : ~n32;
  assign n29379 = pi17 ? n29375 : n29378;
  assign n29380 = pi16 ? n29369 : ~n29379;
  assign n29381 = pi15 ? n29380 : n29224;
  assign n29382 = pi14 ? n29381 : n29238;
  assign n29383 = pi13 ? n29382 : n29257;
  assign n29384 = pi18 ? n13949 : n32;
  assign n29385 = pi17 ? n16982 : n29384;
  assign n29386 = pi16 ? n32 : n29385;
  assign n29387 = pi15 ? n32 : n29386;
  assign n29388 = pi14 ? n32 : n29387;
  assign n29389 = pi20 ? n1331 : n9491;
  assign n29390 = pi19 ? n29389 : n29286;
  assign n29391 = pi18 ? n858 : n29390;
  assign n29392 = pi17 ? n32 : n29391;
  assign n29393 = pi19 ? n29290 : ~n206;
  assign n29394 = pi20 ? n371 : ~n6621;
  assign n29395 = pi19 ? n29394 : ~n18133;
  assign n29396 = pi18 ? n29393 : ~n29395;
  assign n29397 = pi20 ? n5854 : ~n339;
  assign n29398 = pi19 ? n29397 : ~n29298;
  assign n29399 = pi18 ? n29398 : n32;
  assign n29400 = pi17 ? n29396 : n29399;
  assign n29401 = pi16 ? n29392 : n29400;
  assign n29402 = pi15 ? n29284 : n29401;
  assign n29403 = pi16 ? n1214 : ~n1843;
  assign n29404 = pi16 ? n29305 : ~n1843;
  assign n29405 = pi15 ? n29403 : n29404;
  assign n29406 = pi14 ? n29402 : n29405;
  assign n29407 = pi13 ? n29388 : n29406;
  assign n29408 = pi12 ? n29383 : n29407;
  assign n29409 = pi11 ? n29362 : n29408;
  assign n29410 = pi10 ? n29351 : n29409;
  assign n29411 = pi09 ? n32 : n29410;
  assign n29412 = pi08 ? n29313 : n29411;
  assign n29413 = pi07 ? n29127 : n29412;
  assign n29414 = pi06 ? n28817 : n29413;
  assign n29415 = pi05 ? n28316 : n29414;
  assign n29416 = pi04 ? n32 : n29415;
  assign n29417 = pi20 ? n32 : n9488;
  assign n29418 = pi19 ? n32 : n29417;
  assign n29419 = pi20 ? n9488 : ~n354;
  assign n29420 = pi19 ? n19129 : n29419;
  assign n29421 = pi18 ? n29418 : n29420;
  assign n29422 = pi18 ? n18520 : ~n6867;
  assign n29423 = pi17 ? n29421 : ~n29422;
  assign n29424 = pi16 ? n28819 : n29423;
  assign n29425 = pi15 ? n32 : n29424;
  assign n29426 = pi17 ? n18518 : ~n29422;
  assign n29427 = pi16 ? n32 : n29426;
  assign n29428 = pi15 ? n18657 : n29427;
  assign n29429 = pi14 ? n29425 : n29428;
  assign n29430 = pi13 ? n32 : n29429;
  assign n29431 = pi15 ? n18657 : n18890;
  assign n29432 = pi14 ? n29431 : n18890;
  assign n29433 = pi18 ? n18893 : n814;
  assign n29434 = pi17 ? n18892 : n29433;
  assign n29435 = pi16 ? n1471 : ~n29434;
  assign n29436 = pi15 ? n20104 : n29435;
  assign n29437 = pi14 ? n19032 : n29436;
  assign n29438 = pi13 ? n29432 : n29437;
  assign n29439 = pi12 ? n29430 : n29438;
  assign n29440 = pi19 ? n1464 : n4670;
  assign n29441 = pi18 ? n940 : ~n29440;
  assign n29442 = pi17 ? n32 : n29441;
  assign n29443 = pi19 ? n18502 : ~n25120;
  assign n29444 = pi20 ? n246 : ~n206;
  assign n29445 = pi19 ? n16431 : n29444;
  assign n29446 = pi18 ? n29443 : ~n29445;
  assign n29447 = pi19 ? n28952 : n220;
  assign n29448 = pi18 ? n29447 : n18532;
  assign n29449 = pi17 ? n29446 : n29448;
  assign n29450 = pi16 ? n29442 : n29449;
  assign n29451 = pi15 ? n18676 : n29450;
  assign n29452 = pi21 ? n259 : n174;
  assign n29453 = pi20 ? n18834 : n2019;
  assign n29454 = pi19 ? n29452 : ~n29453;
  assign n29455 = pi18 ? n32 : n29454;
  assign n29456 = pi17 ? n32 : n29455;
  assign n29457 = pi21 ? n206 : n173;
  assign n29458 = pi20 ? n18282 : ~n29457;
  assign n29459 = pi19 ? n29458 : n358;
  assign n29460 = pi18 ? n29459 : n7221;
  assign n29461 = pi20 ? n274 : n6303;
  assign n29462 = pi19 ? n18741 : n29461;
  assign n29463 = pi18 ? n29462 : n32;
  assign n29464 = pi17 ? n29460 : n29463;
  assign n29465 = pi16 ? n29456 : n29464;
  assign n29466 = pi15 ? n29465 : n18661;
  assign n29467 = pi14 ? n29451 : n29466;
  assign n29468 = pi14 ? n18661 : n18663;
  assign n29469 = pi13 ? n29467 : n29468;
  assign n29470 = pi20 ? n17665 : n1076;
  assign n29471 = pi19 ? n29363 : n29470;
  assign n29472 = pi20 ? n1076 : n357;
  assign n29473 = pi20 ? n175 : ~n6050;
  assign n29474 = pi19 ? n29472 : n29473;
  assign n29475 = pi18 ? n29471 : n29474;
  assign n29476 = pi20 ? n266 : ~n17669;
  assign n29477 = pi20 ? n1324 : n17652;
  assign n29478 = pi19 ? n29476 : ~n29477;
  assign n29479 = pi18 ? n29478 : n1813;
  assign n29480 = pi17 ? n29475 : ~n29479;
  assign n29481 = pi16 ? n32 : n29480;
  assign n29482 = pi19 ? n29270 : n22525;
  assign n29483 = pi18 ? n858 : n29482;
  assign n29484 = pi19 ? n4670 : n18497;
  assign n29485 = pi18 ? n29484 : n1813;
  assign n29486 = pi17 ? n29483 : ~n29485;
  assign n29487 = pi16 ? n32 : n29486;
  assign n29488 = pi15 ? n29481 : n29487;
  assign n29489 = pi14 ? n19395 : n29488;
  assign n29490 = pi14 ? n18536 : n29050;
  assign n29491 = pi13 ? n29489 : n29490;
  assign n29492 = pi12 ? n29469 : n29491;
  assign n29493 = pi11 ? n29439 : n29492;
  assign n29494 = pi18 ? n936 : ~n237;
  assign n29495 = pi17 ? n32 : n29494;
  assign n29496 = pi16 ? n32 : n29495;
  assign n29497 = pi15 ? n18814 : n29496;
  assign n29498 = pi16 ? n32 : n239;
  assign n29499 = pi15 ? n29498 : n19172;
  assign n29500 = pi14 ? n29497 : n29499;
  assign n29501 = pi18 ? n858 : ~n237;
  assign n29502 = pi17 ? n32 : n29501;
  assign n29503 = pi16 ? n32 : n29502;
  assign n29504 = pi15 ? n18814 : n29503;
  assign n29505 = pi15 ? n32 : n18601;
  assign n29506 = pi14 ? n29504 : n29505;
  assign n29507 = pi13 ? n29500 : n29506;
  assign n29508 = pi15 ? n18439 : n18008;
  assign n29509 = pi14 ? n18439 : n29508;
  assign n29510 = pi18 ? n17118 : n32;
  assign n29511 = pi17 ? n32 : n29510;
  assign n29512 = pi16 ? n32 : n29511;
  assign n29513 = pi15 ? n32 : n29512;
  assign n29514 = pi20 ? n1817 : ~n501;
  assign n29515 = pi19 ? n32 : n29514;
  assign n29516 = pi18 ? n29515 : n32;
  assign n29517 = pi17 ? n32 : n29516;
  assign n29518 = pi16 ? n32 : n29517;
  assign n29519 = pi16 ? n1233 : ~n1471;
  assign n29520 = pi15 ? n29518 : n29519;
  assign n29521 = pi14 ? n29513 : n29520;
  assign n29522 = pi13 ? n29509 : n29521;
  assign n29523 = pi12 ? n29507 : n29522;
  assign n29524 = pi21 ? n140 : n174;
  assign n29525 = pi20 ? n32 : n29524;
  assign n29526 = pi19 ? n32 : n29525;
  assign n29527 = pi20 ? n17671 : n17652;
  assign n29528 = pi19 ? n24755 : ~n29527;
  assign n29529 = pi18 ? n29526 : ~n29528;
  assign n29530 = pi17 ? n32 : n29529;
  assign n29531 = pi20 ? n5854 : ~n18762;
  assign n29532 = pi19 ? n29531 : ~n5675;
  assign n29533 = pi20 ? n309 : ~n10644;
  assign n29534 = pi20 ? n1331 : n17669;
  assign n29535 = pi19 ? n29533 : n29534;
  assign n29536 = pi18 ? n29532 : ~n29535;
  assign n29537 = pi20 ? n1331 : n12884;
  assign n29538 = pi19 ? n29537 : n322;
  assign n29539 = pi18 ? n29538 : ~n32;
  assign n29540 = pi17 ? n29536 : ~n29539;
  assign n29541 = pi16 ? n29530 : n29540;
  assign n29542 = pi19 ? n32 : ~n594;
  assign n29543 = pi18 ? n29542 : n32;
  assign n29544 = pi17 ? n32 : n29543;
  assign n29545 = pi16 ? n32 : n29544;
  assign n29546 = pi15 ? n29541 : n29545;
  assign n29547 = pi19 ? n322 : ~n594;
  assign n29548 = pi18 ? n29547 : n32;
  assign n29549 = pi17 ? n32 : n29548;
  assign n29550 = pi16 ? n32 : n29549;
  assign n29551 = pi14 ? n29546 : n29550;
  assign n29552 = pi19 ? n322 : ~n507;
  assign n29553 = pi18 ? n29552 : n32;
  assign n29554 = pi17 ? n32 : n29553;
  assign n29555 = pi16 ? n32 : n29554;
  assign n29556 = pi19 ? n6398 : ~n236;
  assign n29557 = pi18 ? n29556 : n32;
  assign n29558 = pi17 ? n32 : n29557;
  assign n29559 = pi16 ? n32 : n29558;
  assign n29560 = pi15 ? n29555 : n29559;
  assign n29561 = pi14 ? n29560 : n17638;
  assign n29562 = pi13 ? n29551 : n29561;
  assign n29563 = pi18 ? n917 : n16847;
  assign n29564 = pi17 ? n32 : n29563;
  assign n29565 = pi16 ? n29564 : n32;
  assign n29566 = pi15 ? n17637 : n29565;
  assign n29567 = pi14 ? n29566 : n32;
  assign n29568 = pi19 ? n507 : n266;
  assign n29569 = pi18 ? n29568 : n32;
  assign n29570 = pi17 ? n32 : n29569;
  assign n29571 = pi16 ? n32 : n29570;
  assign n29572 = pi18 ? n16394 : n32;
  assign n29573 = pi17 ? n32 : n29572;
  assign n29574 = pi16 ? n32 : n29573;
  assign n29575 = pi15 ? n29571 : n29574;
  assign n29576 = pi18 ? n341 : ~n16449;
  assign n29577 = pi17 ? n32 : n29576;
  assign n29578 = pi16 ? n29577 : ~n1594;
  assign n29579 = pi18 ? n18710 : ~n15844;
  assign n29580 = pi17 ? n32 : n29579;
  assign n29581 = pi19 ? n322 : ~n5675;
  assign n29582 = pi18 ? n29581 : ~n32;
  assign n29583 = pi17 ? n32 : n29582;
  assign n29584 = pi16 ? n29580 : ~n29583;
  assign n29585 = pi15 ? n29578 : n29584;
  assign n29586 = pi14 ? n29575 : n29585;
  assign n29587 = pi13 ? n29567 : n29586;
  assign n29588 = pi12 ? n29562 : n29587;
  assign n29589 = pi11 ? n29523 : n29588;
  assign n29590 = pi10 ? n29493 : n29589;
  assign n29591 = pi09 ? n32 : n29590;
  assign n29592 = pi18 ? n618 : ~n18894;
  assign n29593 = pi17 ? n16982 : ~n29592;
  assign n29594 = pi16 ? n32 : n29593;
  assign n29595 = pi15 ? n32 : n29594;
  assign n29596 = pi15 ? n18904 : n29594;
  assign n29597 = pi14 ? n29595 : n29596;
  assign n29598 = pi13 ? n32 : n29597;
  assign n29599 = pi15 ? n18904 : n165;
  assign n29600 = pi14 ? n29599 : n165;
  assign n29601 = pi16 ? n1233 : ~n1808;
  assign n29602 = pi18 ? n18893 : n1813;
  assign n29603 = pi17 ? n18892 : n29602;
  assign n29604 = pi16 ? n1471 : ~n29603;
  assign n29605 = pi15 ? n29601 : n29604;
  assign n29606 = pi14 ? n20746 : n29605;
  assign n29607 = pi13 ? n29600 : n29606;
  assign n29608 = pi12 ? n29598 : n29607;
  assign n29609 = pi18 ? n29447 : n18521;
  assign n29610 = pi17 ? n29446 : n29609;
  assign n29611 = pi16 ? n29442 : n29610;
  assign n29612 = pi15 ? n18798 : n29611;
  assign n29613 = pi20 ? n6621 : n266;
  assign n29614 = pi20 ? n7939 : ~n4279;
  assign n29615 = pi19 ? n29613 : ~n29614;
  assign n29616 = pi18 ? n32 : n29615;
  assign n29617 = pi17 ? n32 : n29616;
  assign n29618 = pi20 ? n1817 : ~n6050;
  assign n29619 = pi19 ? n29618 : n32;
  assign n29620 = pi18 ? n29619 : n32;
  assign n29621 = pi17 ? n29620 : n17705;
  assign n29622 = pi16 ? n29617 : n29621;
  assign n29623 = pi15 ? n29622 : n18661;
  assign n29624 = pi14 ? n29612 : n29623;
  assign n29625 = pi14 ? n20583 : n18661;
  assign n29626 = pi13 ? n29624 : n29625;
  assign n29627 = pi19 ? n1818 : n29470;
  assign n29628 = pi18 ? n29627 : n29474;
  assign n29629 = pi17 ? n29628 : ~n29479;
  assign n29630 = pi16 ? n32 : n29629;
  assign n29631 = pi18 ? n32 : n29482;
  assign n29632 = pi17 ? n29631 : ~n29485;
  assign n29633 = pi16 ? n32 : n29632;
  assign n29634 = pi15 ? n29630 : n29633;
  assign n29635 = pi14 ? n18947 : n29634;
  assign n29636 = pi14 ? n18536 : n32;
  assign n29637 = pi13 ? n29635 : n29636;
  assign n29638 = pi12 ? n29626 : n29637;
  assign n29639 = pi11 ? n29608 : n29638;
  assign n29640 = pi18 ? n936 : ~n1942;
  assign n29641 = pi17 ? n32 : n29640;
  assign n29642 = pi16 ? n32 : n29641;
  assign n29643 = pi15 ? n19061 : n29642;
  assign n29644 = pi18 ? n209 : ~n1942;
  assign n29645 = pi17 ? n32 : n29644;
  assign n29646 = pi16 ? n32 : n29645;
  assign n29647 = pi15 ? n29646 : n19166;
  assign n29648 = pi14 ? n29643 : n29647;
  assign n29649 = pi18 ? n858 : ~n1942;
  assign n29650 = pi17 ? n32 : n29649;
  assign n29651 = pi16 ? n32 : n29650;
  assign n29652 = pi15 ? n19061 : n29651;
  assign n29653 = pi14 ? n29652 : n29505;
  assign n29654 = pi13 ? n29648 : n29653;
  assign n29655 = pi15 ? n18439 : n17894;
  assign n29656 = pi14 ? n18439 : n29655;
  assign n29657 = pi20 ? n32 : n6822;
  assign n29658 = pi19 ? n32 : n29657;
  assign n29659 = pi20 ? n6822 : ~n18281;
  assign n29660 = pi20 ? n10889 : n6822;
  assign n29661 = pi19 ? n29659 : ~n29660;
  assign n29662 = pi18 ? n29658 : n29661;
  assign n29663 = pi17 ? n32 : n29662;
  assign n29664 = pi20 ? n18832 : n18073;
  assign n29665 = pi20 ? n10889 : n20944;
  assign n29666 = pi19 ? n29664 : n29665;
  assign n29667 = pi20 ? n20396 : ~n18337;
  assign n29668 = pi20 ? n17669 : ~n17669;
  assign n29669 = pi19 ? n29667 : ~n29668;
  assign n29670 = pi18 ? n29666 : n29669;
  assign n29671 = pi20 ? n17669 : ~n12884;
  assign n29672 = pi19 ? n29671 : n13714;
  assign n29673 = pi18 ? n29672 : ~n32;
  assign n29674 = pi17 ? n29670 : ~n29673;
  assign n29675 = pi16 ? n29663 : n29674;
  assign n29676 = pi16 ? n1135 : ~n1471;
  assign n29677 = pi15 ? n29675 : n29676;
  assign n29678 = pi14 ? n29513 : n29677;
  assign n29679 = pi13 ? n29656 : n29678;
  assign n29680 = pi12 ? n29654 : n29679;
  assign n29681 = pi19 ? n32 : n6622;
  assign n29682 = pi20 ? n17669 : n310;
  assign n29683 = pi19 ? n29682 : ~n29527;
  assign n29684 = pi18 ? n29681 : ~n29683;
  assign n29685 = pi17 ? n32 : n29684;
  assign n29686 = pi20 ? n5854 : ~n18261;
  assign n29687 = pi20 ? n9491 : n371;
  assign n29688 = pi19 ? n29686 : ~n29687;
  assign n29689 = pi20 ? n206 : n5854;
  assign n29690 = pi19 ? n29689 : ~n29110;
  assign n29691 = pi18 ? n29688 : n29690;
  assign n29692 = pi20 ? n310 : ~n4279;
  assign n29693 = pi19 ? n29692 : n322;
  assign n29694 = pi18 ? n29693 : ~n32;
  assign n29695 = pi17 ? n29691 : ~n29694;
  assign n29696 = pi16 ? n29685 : n29695;
  assign n29697 = pi15 ? n29696 : n29545;
  assign n29698 = pi14 ? n29697 : n29550;
  assign n29699 = pi18 ? n20172 : n32;
  assign n29700 = pi17 ? n32 : n29699;
  assign n29701 = pi16 ? n32 : n29700;
  assign n29702 = pi15 ? n29555 : n29701;
  assign n29703 = pi14 ? n29702 : n17911;
  assign n29704 = pi13 ? n29698 : n29703;
  assign n29705 = pi20 ? n274 : n266;
  assign n29706 = pi19 ? n507 : n29705;
  assign n29707 = pi18 ? n29706 : n32;
  assign n29708 = pi17 ? n32 : n29707;
  assign n29709 = pi16 ? n32 : n29708;
  assign n29710 = pi15 ? n29709 : n29574;
  assign n29711 = pi14 ? n29710 : n29585;
  assign n29712 = pi13 ? n29567 : n29711;
  assign n29713 = pi12 ? n29704 : n29712;
  assign n29714 = pi11 ? n29680 : n29713;
  assign n29715 = pi10 ? n29639 : n29714;
  assign n29716 = pi09 ? n32 : n29715;
  assign n29717 = pi08 ? n29591 : n29716;
  assign n29718 = pi19 ? n18741 : n32;
  assign n29719 = pi18 ? n29718 : n162;
  assign n29720 = pi17 ? n20658 : n29719;
  assign n29721 = pi16 ? n32 : n29720;
  assign n29722 = pi15 ? n32 : n29721;
  assign n29723 = pi14 ? n29722 : n29721;
  assign n29724 = pi13 ? n32 : n29723;
  assign n29725 = pi15 ? n29721 : n165;
  assign n29726 = pi16 ? n17636 : n164;
  assign n29727 = pi15 ? n165 : n29726;
  assign n29728 = pi14 ? n29725 : n29727;
  assign n29729 = pi16 ? n1471 : ~n1808;
  assign n29730 = pi18 ? n19120 : ~n618;
  assign n29731 = pi17 ? n19118 : ~n29730;
  assign n29732 = pi16 ? n1471 : ~n29731;
  assign n29733 = pi15 ? n29729 : n29732;
  assign n29734 = pi14 ? n20746 : n29733;
  assign n29735 = pi13 ? n29728 : n29734;
  assign n29736 = pi12 ? n29724 : n29735;
  assign n29737 = pi18 ? n858 : n29454;
  assign n29738 = pi17 ? n32 : n29737;
  assign n29739 = pi20 ? n357 : n915;
  assign n29740 = pi19 ? n29458 : n29739;
  assign n29741 = pi20 ? n915 : n1368;
  assign n29742 = pi20 ? n29452 : n175;
  assign n29743 = pi19 ? n29741 : n29742;
  assign n29744 = pi18 ? n29740 : n29743;
  assign n29745 = pi19 ? n32 : n6303;
  assign n29746 = pi18 ? n29745 : n18532;
  assign n29747 = pi17 ? n29744 : n29746;
  assign n29748 = pi16 ? n29738 : n29747;
  assign n29749 = pi19 ? n267 : n18678;
  assign n29750 = pi18 ? n32 : n29749;
  assign n29751 = pi17 ? n32 : n29750;
  assign n29752 = pi17 ? n19904 : n32;
  assign n29753 = pi16 ? n29751 : n29752;
  assign n29754 = pi15 ? n29748 : n29753;
  assign n29755 = pi15 ? n32 : n18657;
  assign n29756 = pi14 ? n29754 : n29755;
  assign n29757 = pi14 ? n20960 : n32;
  assign n29758 = pi13 ? n29756 : n29757;
  assign n29759 = pi19 ? n32 : n175;
  assign n29760 = pi18 ? n32 : n29759;
  assign n29761 = pi20 ? n1817 : n246;
  assign n29762 = pi19 ? n18789 : n29761;
  assign n29763 = pi18 ? n29762 : ~n350;
  assign n29764 = pi17 ? n29760 : n29763;
  assign n29765 = pi16 ? n32 : n29764;
  assign n29766 = pi15 ? n29765 : n19531;
  assign n29767 = pi14 ? n19531 : n29766;
  assign n29768 = pi13 ? n29767 : n19163;
  assign n29769 = pi12 ? n29758 : n29768;
  assign n29770 = pi11 ? n29736 : n29769;
  assign n29771 = pi15 ? n19405 : n19166;
  assign n29772 = pi14 ? n18814 : n29771;
  assign n29773 = pi14 ? n19461 : n29505;
  assign n29774 = pi13 ? n29772 : n29773;
  assign n29775 = pi18 ? n2197 : n32;
  assign n29776 = pi17 ? n32 : n29775;
  assign n29777 = pi16 ? n32 : n29776;
  assign n29778 = pi15 ? n29777 : n32;
  assign n29779 = pi14 ? n19720 : n29778;
  assign n29780 = pi16 ? n1135 : ~n1214;
  assign n29781 = pi15 ? n32 : n29780;
  assign n29782 = pi16 ? n19200 : ~n1214;
  assign n29783 = pi20 ? n6822 : n3843;
  assign n29784 = pi19 ? n29783 : ~n5854;
  assign n29785 = pi18 ? n29086 : ~n29784;
  assign n29786 = pi17 ? n32 : n29785;
  assign n29787 = pi20 ? n18261 : n18073;
  assign n29788 = pi19 ? n29787 : n3523;
  assign n29789 = pi20 ? n357 : n405;
  assign n29790 = pi20 ? n32 : n18762;
  assign n29791 = pi19 ? n29789 : n29790;
  assign n29792 = pi18 ? n29788 : n29791;
  assign n29793 = pi20 ? n266 : n18762;
  assign n29794 = pi19 ? n29793 : n507;
  assign n29795 = pi18 ? n29794 : ~n32;
  assign n29796 = pi17 ? n29792 : n29795;
  assign n29797 = pi16 ? n29786 : ~n29796;
  assign n29798 = pi15 ? n29782 : n29797;
  assign n29799 = pi14 ? n29781 : n29798;
  assign n29800 = pi13 ? n29779 : n29799;
  assign n29801 = pi12 ? n29774 : n29800;
  assign n29802 = pi19 ? n32 : ~n322;
  assign n29803 = pi18 ? n29802 : n32;
  assign n29804 = pi17 ? n32 : n29803;
  assign n29805 = pi16 ? n32 : n29804;
  assign n29806 = pi15 ? n29805 : n18181;
  assign n29807 = pi19 ? n32 : ~n1574;
  assign n29808 = pi18 ? n29807 : n32;
  assign n29809 = pi17 ? n32 : n29808;
  assign n29810 = pi16 ? n32 : n29809;
  assign n29811 = pi15 ? n18181 : n29810;
  assign n29812 = pi14 ? n29806 : n29811;
  assign n29813 = pi15 ? n18181 : n32;
  assign n29814 = pi14 ? n29813 : n32;
  assign n29815 = pi13 ? n29812 : n29814;
  assign n29816 = pi15 ? n32 : n271;
  assign n29817 = pi14 ? n29816 : n32;
  assign n29818 = pi15 ? n28632 : n18040;
  assign n29819 = pi18 ? n209 : ~n16234;
  assign n29820 = pi17 ? n32 : n29819;
  assign n29821 = pi16 ? n29820 : ~n1594;
  assign n29822 = pi18 ? n940 : ~n16234;
  assign n29823 = pi17 ? n32 : n29822;
  assign n29824 = pi19 ? n322 : ~n1818;
  assign n29825 = pi18 ? n29824 : ~n32;
  assign n29826 = pi17 ? n32 : n29825;
  assign n29827 = pi16 ? n29823 : ~n29826;
  assign n29828 = pi15 ? n29821 : n29827;
  assign n29829 = pi14 ? n29818 : n29828;
  assign n29830 = pi13 ? n29817 : n29829;
  assign n29831 = pi12 ? n29815 : n29830;
  assign n29832 = pi11 ? n29801 : n29831;
  assign n29833 = pi10 ? n29770 : n29832;
  assign n29834 = pi09 ? n32 : n29833;
  assign n29835 = pi18 ? n29718 : n19232;
  assign n29836 = pi17 ? n20658 : n29835;
  assign n29837 = pi16 ? n32 : n29836;
  assign n29838 = pi15 ? n32 : n29837;
  assign n29839 = pi14 ? n29838 : n29837;
  assign n29840 = pi13 ? n32 : n29839;
  assign n29841 = pi15 ? n29837 : n19235;
  assign n29842 = pi16 ? n17636 : n19239;
  assign n29843 = pi15 ? n19235 : n29842;
  assign n29844 = pi14 ? n29841 : n29843;
  assign n29845 = pi16 ? n1471 : ~n3338;
  assign n29846 = pi15 ? n29845 : n29732;
  assign n29847 = pi14 ? n19326 : n29846;
  assign n29848 = pi13 ? n29844 : n29847;
  assign n29849 = pi12 ? n29840 : n29848;
  assign n29850 = pi18 ? n858 : n29615;
  assign n29851 = pi17 ? n32 : n29850;
  assign n29852 = pi19 ? n29618 : n267;
  assign n29853 = pi19 ? n23180 : n1757;
  assign n29854 = pi18 ? n29852 : n29853;
  assign n29855 = pi18 ? n28876 : n32;
  assign n29856 = pi17 ? n29854 : n29855;
  assign n29857 = pi16 ? n29851 : n29856;
  assign n29858 = pi15 ? n29857 : n29753;
  assign n29859 = pi14 ? n29858 : n29755;
  assign n29860 = pi13 ? n29859 : n29757;
  assign n29861 = pi17 ? n32 : n20448;
  assign n29862 = pi16 ? n32 : n29861;
  assign n29863 = pi15 ? n29862 : n19531;
  assign n29864 = pi14 ? n19531 : n29863;
  assign n29865 = pi14 ? n18531 : n32;
  assign n29866 = pi13 ? n29864 : n29865;
  assign n29867 = pi12 ? n29860 : n29866;
  assign n29868 = pi11 ? n29849 : n29867;
  assign n29869 = pi15 ? n19459 : n19264;
  assign n29870 = pi14 ? n19536 : n29869;
  assign n29871 = pi15 ? n19536 : n19264;
  assign n29872 = pi14 ? n29871 : n29505;
  assign n29873 = pi13 ? n29870 : n29872;
  assign n29874 = pi14 ? n19720 : n28507;
  assign n29875 = pi16 ? n1233 : ~n1214;
  assign n29876 = pi15 ? n32 : n29875;
  assign n29877 = pi20 ? n17652 : n310;
  assign n29878 = pi19 ? n29877 : ~n5854;
  assign n29879 = pi18 ? n29418 : ~n29878;
  assign n29880 = pi17 ? n32 : n29879;
  assign n29881 = pi20 ? n18261 : n9491;
  assign n29882 = pi20 ? n17669 : n246;
  assign n29883 = pi19 ? n29881 : n29882;
  assign n29884 = pi20 ? n21111 : ~n2385;
  assign n29885 = pi20 ? n309 : ~n5854;
  assign n29886 = pi19 ? n29884 : ~n29885;
  assign n29887 = pi18 ? n29883 : ~n29886;
  assign n29888 = pi20 ? n310 : ~n5854;
  assign n29889 = pi19 ? n29888 : n507;
  assign n29890 = pi18 ? n29889 : ~n32;
  assign n29891 = pi17 ? n29887 : n29890;
  assign n29892 = pi16 ? n29880 : ~n29891;
  assign n29893 = pi15 ? n29782 : n29892;
  assign n29894 = pi14 ? n29876 : n29893;
  assign n29895 = pi13 ? n29874 : n29894;
  assign n29896 = pi12 ? n29873 : n29895;
  assign n29897 = pi18 ? n15570 : ~n1676;
  assign n29898 = pi17 ? n32 : n29897;
  assign n29899 = pi16 ? n32 : n29898;
  assign n29900 = pi18 ? n702 : n32;
  assign n29901 = pi17 ? n32 : n29900;
  assign n29902 = pi16 ? n32 : n29901;
  assign n29903 = pi15 ? n29899 : n29902;
  assign n29904 = pi14 ? n29806 : n29903;
  assign n29905 = pi13 ? n29904 : n29814;
  assign n29906 = pi12 ? n29905 : n29830;
  assign n29907 = pi11 ? n29896 : n29906;
  assign n29908 = pi10 ? n29868 : n29907;
  assign n29909 = pi09 ? n32 : n29908;
  assign n29910 = pi08 ? n29834 : n29909;
  assign n29911 = pi07 ? n29717 : n29910;
  assign n29912 = pi20 ? n18129 : ~n6050;
  assign n29913 = pi19 ? n32 : n29912;
  assign n29914 = pi20 ? n207 : n314;
  assign n29915 = pi19 ? n19115 : n29914;
  assign n29916 = pi18 ? n29913 : ~n29915;
  assign n29917 = pi19 ? n18839 : ~n18763;
  assign n29918 = pi20 ? n17665 : n32;
  assign n29919 = pi19 ? n29918 : n32;
  assign n29920 = pi18 ? n29917 : ~n29919;
  assign n29921 = pi17 ? n29916 : ~n29920;
  assign n29922 = pi16 ? n32 : n29921;
  assign n29923 = pi15 ? n32 : n29922;
  assign n29924 = pi15 ? n19235 : n29922;
  assign n29925 = pi14 ? n29923 : n29924;
  assign n29926 = pi13 ? n32 : n29925;
  assign n29927 = pi19 ? n19115 : ~n11374;
  assign n29928 = pi18 ? n19130 : ~n29927;
  assign n29929 = pi17 ? n29928 : ~n29920;
  assign n29930 = pi16 ? n32 : n29929;
  assign n29931 = pi16 ? n13947 : n19234;
  assign n29932 = pi15 ? n29930 : n29931;
  assign n29933 = pi16 ? n17850 : n19234;
  assign n29934 = pi15 ? n19235 : n29933;
  assign n29935 = pi14 ? n29932 : n29934;
  assign n29936 = pi16 ? n20257 : n32;
  assign n29937 = pi17 ? n18482 : n32;
  assign n29938 = pi16 ? n17120 : n29937;
  assign n29939 = pi15 ? n29936 : n29938;
  assign n29940 = pi14 ? n19326 : n29939;
  assign n29941 = pi13 ? n29935 : n29940;
  assign n29942 = pi12 ? n29926 : n29941;
  assign n29943 = pi18 ? n248 : n18894;
  assign n29944 = pi17 ? n32 : n29943;
  assign n29945 = pi16 ? n32 : n29944;
  assign n29946 = pi15 ? n165 : n29945;
  assign n29947 = pi14 ? n166 : n29946;
  assign n29948 = pi13 ? n167 : n29947;
  assign n29949 = pi21 ? n259 : ~n140;
  assign n29950 = pi20 ? n29949 : n32;
  assign n29951 = pi19 ? n29950 : n32;
  assign n29952 = pi18 ? n32 : n29951;
  assign n29953 = pi17 ? n32 : n29952;
  assign n29954 = pi16 ? n32 : n29953;
  assign n29955 = pi15 ? n29954 : n19691;
  assign n29956 = pi14 ? n19691 : n29955;
  assign n29957 = pi13 ? n29956 : n32;
  assign n29958 = pi12 ? n29948 : n29957;
  assign n29959 = pi11 ? n29942 : n29958;
  assign n29960 = pi15 ? n19267 : n19264;
  assign n29961 = pi14 ? n19264 : n29960;
  assign n29962 = pi15 ? n19264 : n19172;
  assign n29963 = pi15 ? n19172 : n32;
  assign n29964 = pi14 ? n29962 : n29963;
  assign n29965 = pi13 ? n29961 : n29964;
  assign n29966 = pi15 ? n19172 : n18008;
  assign n29967 = pi15 ? n32 : n18019;
  assign n29968 = pi14 ? n29966 : n29967;
  assign n29969 = pi15 ? n32 : n28947;
  assign n29970 = pi18 ? n4868 : n32;
  assign n29971 = pi17 ? n32 : n29970;
  assign n29972 = pi16 ? n32 : n29971;
  assign n29973 = pi15 ? n28947 : n29972;
  assign n29974 = pi14 ? n29969 : n29973;
  assign n29975 = pi13 ? n29968 : n29974;
  assign n29976 = pi12 ? n29965 : n29975;
  assign n29977 = pi15 ? n17885 : n17903;
  assign n29978 = pi19 ? n32 : n6307;
  assign n29979 = pi18 ? n29978 : n32;
  assign n29980 = pi17 ? n32 : n29979;
  assign n29981 = pi16 ? n32 : n29980;
  assign n29982 = pi15 ? n29902 : n29981;
  assign n29983 = pi14 ? n29977 : n29982;
  assign n29984 = pi13 ? n29983 : n28398;
  assign n29985 = pi16 ? n32 : n919;
  assign n29986 = pi15 ? n32 : n29985;
  assign n29987 = pi14 ? n32 : n29986;
  assign n29988 = pi15 ? n17702 : n18326;
  assign n29989 = pi14 ? n29988 : n18326;
  assign n29990 = pi13 ? n29987 : n29989;
  assign n29991 = pi12 ? n29984 : n29990;
  assign n29992 = pi11 ? n29976 : n29991;
  assign n29993 = pi10 ? n29959 : n29992;
  assign n29994 = pi09 ? n32 : n29993;
  assign n29995 = pi20 ? n22458 : n32;
  assign n29996 = pi19 ? n29995 : n32;
  assign n29997 = pi18 ? n29917 : ~n29996;
  assign n29998 = pi17 ? n29916 : ~n29997;
  assign n29999 = pi16 ? n32 : n29998;
  assign n30000 = pi15 ? n32 : n29999;
  assign n30001 = pi15 ? n19235 : n29999;
  assign n30002 = pi14 ? n30000 : n30001;
  assign n30003 = pi13 ? n32 : n30002;
  assign n30004 = pi17 ? n29928 : ~n29997;
  assign n30005 = pi16 ? n32 : n30004;
  assign n30006 = pi16 ? n13947 : n90;
  assign n30007 = pi15 ? n30005 : n30006;
  assign n30008 = pi16 ? n17850 : n19383;
  assign n30009 = pi15 ? n19384 : n30008;
  assign n30010 = pi14 ? n30007 : n30009;
  assign n30011 = pi15 ? n19384 : n32;
  assign n30012 = pi14 ? n30011 : n29939;
  assign n30013 = pi13 ? n30010 : n30012;
  assign n30014 = pi12 ? n30003 : n30013;
  assign n30015 = pi13 ? n32 : n29947;
  assign n30016 = pi13 ? n19691 : n19394;
  assign n30017 = pi12 ? n30015 : n30016;
  assign n30018 = pi11 ? n30014 : n30017;
  assign n30019 = pi15 ? n19896 : n19398;
  assign n30020 = pi14 ? n19264 : n30019;
  assign n30021 = pi15 ? n19398 : n19172;
  assign n30022 = pi14 ? n30021 : n29963;
  assign n30023 = pi13 ? n30020 : n30022;
  assign n30024 = pi14 ? n19172 : n29967;
  assign n30025 = pi16 ? n1233 : ~n1581;
  assign n30026 = pi15 ? n32 : n30025;
  assign n30027 = pi15 ? n30025 : n29972;
  assign n30028 = pi14 ? n30026 : n30027;
  assign n30029 = pi13 ? n30024 : n30028;
  assign n30030 = pi12 ? n30023 : n30029;
  assign n30031 = pi16 ? n32 : n375;
  assign n30032 = pi15 ? n32 : n30031;
  assign n30033 = pi14 ? n32 : n30032;
  assign n30034 = pi13 ? n30033 : n18326;
  assign n30035 = pi12 ? n29984 : n30034;
  assign n30036 = pi11 ? n30030 : n30035;
  assign n30037 = pi10 ? n30018 : n30036;
  assign n30038 = pi09 ? n32 : n30037;
  assign n30039 = pi08 ? n29994 : n30038;
  assign n30040 = pi20 ? n9194 : ~n17652;
  assign n30041 = pi19 ? n28070 : ~n30040;
  assign n30042 = pi18 ? n32 : n30041;
  assign n30043 = pi17 ? n32 : n30042;
  assign n30044 = pi20 ? n9491 : n9488;
  assign n30045 = pi20 ? n6303 : n428;
  assign n30046 = pi19 ? n30044 : ~n30045;
  assign n30047 = pi18 ? n30046 : ~n29146;
  assign n30048 = pi20 ? n357 : n333;
  assign n30049 = pi19 ? n30048 : ~n28580;
  assign n30050 = pi18 ? n30049 : ~n29996;
  assign n30051 = pi17 ? n30047 : ~n30050;
  assign n30052 = pi16 ? n30043 : n30051;
  assign n30053 = pi15 ? n32 : n30052;
  assign n30054 = pi15 ? n91 : n30052;
  assign n30055 = pi14 ? n30053 : n30054;
  assign n30056 = pi13 ? n32 : n30055;
  assign n30057 = pi20 ? n3843 : n246;
  assign n30058 = pi19 ? n32 : n30057;
  assign n30059 = pi20 ? n206 : n501;
  assign n30060 = pi19 ? n30059 : ~n19116;
  assign n30061 = pi18 ? n30058 : ~n30060;
  assign n30062 = pi20 ? n1611 : n5854;
  assign n30063 = pi19 ? n30062 : ~n1611;
  assign n30064 = pi18 ? n30063 : ~n29996;
  assign n30065 = pi17 ? n30061 : ~n30064;
  assign n30066 = pi16 ? n32 : n30065;
  assign n30067 = pi15 ? n30066 : n30006;
  assign n30068 = pi16 ? n17850 : n90;
  assign n30069 = pi15 ? n91 : n30068;
  assign n30070 = pi14 ? n30067 : n30069;
  assign n30071 = pi15 ? n30008 : n19235;
  assign n30072 = pi14 ? n30071 : n32;
  assign n30073 = pi13 ? n30070 : n30072;
  assign n30074 = pi12 ? n30056 : n30073;
  assign n30075 = pi19 ? n311 : ~n322;
  assign n30076 = pi18 ? n30075 : ~n19811;
  assign n30077 = pi17 ? n4261 : ~n30076;
  assign n30078 = pi16 ? n32 : n30077;
  assign n30079 = pi15 ? n19235 : n30078;
  assign n30080 = pi14 ? n19235 : n30079;
  assign n30081 = pi13 ? n21122 : n30080;
  assign n30082 = pi13 ? n20646 : n19454;
  assign n30083 = pi12 ? n30081 : n30082;
  assign n30084 = pi11 ? n30074 : n30083;
  assign n30085 = pi19 ? n26777 : n32;
  assign n30086 = pi18 ? n32 : n30085;
  assign n30087 = pi17 ? n32 : n30086;
  assign n30088 = pi16 ? n32 : n30087;
  assign n30089 = pi14 ? n19399 : n30088;
  assign n30090 = pi22 ? n173 : n84;
  assign n30091 = pi21 ? n30090 : n32;
  assign n30092 = pi20 ? n30091 : n32;
  assign n30093 = pi19 ? n30092 : n32;
  assign n30094 = pi18 ? n32 : n30093;
  assign n30095 = pi17 ? n32 : n30094;
  assign n30096 = pi16 ? n32 : n30095;
  assign n30097 = pi17 ? n32 : n20024;
  assign n30098 = pi16 ? n32 : n30097;
  assign n30099 = pi15 ? n30096 : n30098;
  assign n30100 = pi14 ? n30099 : n19172;
  assign n30101 = pi13 ? n30089 : n30100;
  assign n30102 = pi18 ? n17848 : ~n237;
  assign n30103 = pi17 ? n32 : n30102;
  assign n30104 = pi16 ? n32 : n30103;
  assign n30105 = pi15 ? n19172 : n30104;
  assign n30106 = pi14 ? n30105 : n29967;
  assign n30107 = pi18 ? n16847 : n32;
  assign n30108 = pi17 ? n32 : n30107;
  assign n30109 = pi16 ? n32 : n30108;
  assign n30110 = pi15 ? n28947 : n30109;
  assign n30111 = pi14 ? n29969 : n30110;
  assign n30112 = pi13 ? n30106 : n30111;
  assign n30113 = pi12 ? n30101 : n30112;
  assign n30114 = pi18 ? n20166 : n32;
  assign n30115 = pi17 ? n32 : n30114;
  assign n30116 = pi16 ? n32 : n30115;
  assign n30117 = pi15 ? n29810 : n30116;
  assign n30118 = pi14 ? n18016 : n30117;
  assign n30119 = pi13 ? n30118 : n28398;
  assign n30120 = pi16 ? n32 : n278;
  assign n30121 = pi15 ? n30120 : n17936;
  assign n30122 = pi14 ? n32 : n30121;
  assign n30123 = pi15 ? n17825 : n17851;
  assign n30124 = pi14 ? n30123 : n18326;
  assign n30125 = pi13 ? n30122 : n30124;
  assign n30126 = pi12 ? n30119 : n30125;
  assign n30127 = pi11 ? n30113 : n30126;
  assign n30128 = pi10 ? n30084 : n30127;
  assign n30129 = pi09 ? n32 : n30128;
  assign n30130 = pi19 ? n12885 : n32;
  assign n30131 = pi18 ? n30049 : ~n30130;
  assign n30132 = pi17 ? n30047 : ~n30131;
  assign n30133 = pi16 ? n30043 : n30132;
  assign n30134 = pi15 ? n32 : n30133;
  assign n30135 = pi15 ? n91 : n30133;
  assign n30136 = pi14 ? n30134 : n30135;
  assign n30137 = pi13 ? n32 : n30136;
  assign n30138 = pi18 ? n30063 : ~n30130;
  assign n30139 = pi17 ? n30061 : ~n30138;
  assign n30140 = pi16 ? n32 : n30139;
  assign n30141 = pi16 ? n13947 : n18561;
  assign n30142 = pi15 ? n30140 : n30141;
  assign n30143 = pi16 ? n17850 : n18561;
  assign n30144 = pi15 ? n19503 : n30143;
  assign n30145 = pi14 ? n30142 : n30144;
  assign n30146 = pi16 ? n17850 : n19804;
  assign n30147 = pi15 ? n30146 : n19235;
  assign n30148 = pi14 ? n30147 : n32;
  assign n30149 = pi13 ? n30145 : n30148;
  assign n30150 = pi12 ? n30137 : n30149;
  assign n30151 = pi13 ? n32 : n30080;
  assign n30152 = pi19 ? n16370 : n32;
  assign n30153 = pi18 ? n32 : n30152;
  assign n30154 = pi17 ? n32 : n30153;
  assign n30155 = pi16 ? n32 : n30154;
  assign n30156 = pi15 ? n18657 : n18904;
  assign n30157 = pi14 ? n30156 : n18657;
  assign n30158 = pi13 ? n30155 : n30157;
  assign n30159 = pi12 ? n30151 : n30158;
  assign n30160 = pi11 ? n30150 : n30159;
  assign n30161 = pi14 ? n19698 : n19531;
  assign n30162 = pi14 ? n19173 : n19172;
  assign n30163 = pi13 ? n30161 : n30162;
  assign n30164 = pi15 ? n30025 : n30109;
  assign n30165 = pi14 ? n30026 : n30164;
  assign n30166 = pi13 ? n30024 : n30165;
  assign n30167 = pi12 ? n30163 : n30166;
  assign n30168 = pi15 ? n29545 : n30116;
  assign n30169 = pi14 ? n18016 : n30168;
  assign n30170 = pi13 ? n30169 : n28398;
  assign n30171 = pi15 ? n30120 : n28168;
  assign n30172 = pi14 ? n32 : n30171;
  assign n30173 = pi13 ? n30172 : n30124;
  assign n30174 = pi12 ? n30170 : n30173;
  assign n30175 = pi11 ? n30167 : n30174;
  assign n30176 = pi10 ? n30160 : n30175;
  assign n30177 = pi09 ? n32 : n30176;
  assign n30178 = pi08 ? n30129 : n30177;
  assign n30179 = pi07 ? n30039 : n30178;
  assign n30180 = pi06 ? n29911 : n30179;
  assign n30181 = pi18 ? n936 : n344;
  assign n30182 = pi17 ? n32 : n30181;
  assign n30183 = pi16 ? n30182 : ~n1934;
  assign n30184 = pi15 ? n19503 : n30183;
  assign n30185 = pi14 ? n19504 : n30184;
  assign n30186 = pi13 ? n32 : n30185;
  assign n30187 = pi16 ? n18325 : n18561;
  assign n30188 = pi15 ? n19503 : n30187;
  assign n30189 = pi14 ? n156 : n30188;
  assign n30190 = pi16 ? n17706 : n18561;
  assign n30191 = pi15 ? n30190 : n32;
  assign n30192 = pi14 ? n30191 : n32;
  assign n30193 = pi13 ? n30189 : n30192;
  assign n30194 = pi12 ? n30186 : n30193;
  assign n30195 = pi14 ? n91 : n19384;
  assign n30196 = pi13 ? n93 : n30195;
  assign n30197 = pi18 ? n32 : n19654;
  assign n30198 = pi17 ? n32 : n30197;
  assign n30199 = pi16 ? n32 : n30198;
  assign n30200 = pi15 ? n18657 : n30199;
  assign n30201 = pi14 ? n29755 : n30200;
  assign n30202 = pi13 ? n19384 : n30201;
  assign n30203 = pi12 ? n30196 : n30202;
  assign n30204 = pi11 ? n30194 : n30203;
  assign n30205 = pi18 ? n17848 : n6059;
  assign n30206 = pi17 ? n32 : n30205;
  assign n30207 = pi16 ? n32 : n30206;
  assign n30208 = pi15 ? n19531 : n30207;
  assign n30209 = pi15 ? n19531 : n32;
  assign n30210 = pi14 ? n30208 : n30209;
  assign n30211 = pi15 ? n32 : n19172;
  assign n30212 = pi15 ? n32 : n18142;
  assign n30213 = pi14 ? n30211 : n30212;
  assign n30214 = pi13 ? n30210 : n30213;
  assign n30215 = pi14 ? n29963 : n32;
  assign n30216 = pi15 ? n18979 : n17885;
  assign n30217 = pi14 ? n29969 : n30216;
  assign n30218 = pi13 ? n30215 : n30217;
  assign n30219 = pi12 ? n30214 : n30218;
  assign n30220 = pi19 ? n32 : n23944;
  assign n30221 = pi18 ? n30220 : n32;
  assign n30222 = pi17 ? n32 : n30221;
  assign n30223 = pi16 ? n32 : n30222;
  assign n30224 = pi15 ? n17885 : n30223;
  assign n30225 = pi18 ? n1249 : n32;
  assign n30226 = pi17 ? n32 : n30225;
  assign n30227 = pi16 ? n32 : n30226;
  assign n30228 = pi15 ? n19217 : n30227;
  assign n30229 = pi14 ? n30224 : n30228;
  assign n30230 = pi13 ? n30229 : n32;
  assign n30231 = pi17 ? n1219 : ~n1682;
  assign n30232 = pi16 ? n1471 : n30231;
  assign n30233 = pi18 ? n18402 : ~n32;
  assign n30234 = pi17 ? n1219 : ~n30233;
  assign n30235 = pi16 ? n1471 : n30234;
  assign n30236 = pi15 ? n30232 : n30235;
  assign n30237 = pi14 ? n32 : n30236;
  assign n30238 = pi14 ? n17822 : n17826;
  assign n30239 = pi13 ? n30237 : n30238;
  assign n30240 = pi12 ? n30230 : n30239;
  assign n30241 = pi11 ? n30219 : n30240;
  assign n30242 = pi10 ? n30204 : n30241;
  assign n30243 = pi09 ? n32 : n30242;
  assign n30244 = pi16 ? n30182 : ~n2306;
  assign n30245 = pi15 ? n156 : n30244;
  assign n30246 = pi14 ? n157 : n30245;
  assign n30247 = pi13 ? n32 : n30246;
  assign n30248 = pi16 ? n18325 : n115;
  assign n30249 = pi15 ? n116 : n30248;
  assign n30250 = pi14 ? n116 : n30249;
  assign n30251 = pi16 ? n17706 : n115;
  assign n30252 = pi15 ? n30251 : n156;
  assign n30253 = pi14 ? n30252 : n32;
  assign n30254 = pi13 ? n30250 : n30253;
  assign n30255 = pi12 ? n30247 : n30254;
  assign n30256 = pi13 ? n32 : n30195;
  assign n30257 = pi14 ? n19384 : n19806;
  assign n30258 = pi15 ? n20646 : n18657;
  assign n30259 = pi14 ? n30258 : n30200;
  assign n30260 = pi13 ? n30257 : n30259;
  assign n30261 = pi12 ? n30256 : n30260;
  assign n30262 = pi11 ? n30255 : n30261;
  assign n30263 = pi15 ? n19691 : n165;
  assign n30264 = pi14 ? n30208 : n30263;
  assign n30265 = pi14 ? n30211 : n19333;
  assign n30266 = pi13 ? n30264 : n30265;
  assign n30267 = pi12 ? n30266 : n30218;
  assign n30268 = pi11 ? n30267 : n30240;
  assign n30269 = pi10 ? n30262 : n30268;
  assign n30270 = pi09 ? n32 : n30269;
  assign n30271 = pi08 ? n30243 : n30270;
  assign n30272 = pi18 ? n863 : n344;
  assign n30273 = pi17 ? n32 : n30272;
  assign n30274 = pi16 ? n30273 : ~n2306;
  assign n30275 = pi15 ? n116 : n30274;
  assign n30276 = pi14 ? n117 : n30275;
  assign n30277 = pi13 ? n32 : n30276;
  assign n30278 = pi15 ? n116 : n19503;
  assign n30279 = pi14 ? n30278 : n32;
  assign n30280 = pi13 ? n116 : n30279;
  assign n30281 = pi12 ? n30277 : n30280;
  assign n30282 = pi14 ? n19925 : n19503;
  assign n30283 = pi18 ? n32 : n18402;
  assign n30284 = pi18 ? n6399 : n4689;
  assign n30285 = pi17 ? n30283 : n30284;
  assign n30286 = pi16 ? n32 : n30285;
  assign n30287 = pi15 ? n30286 : n19805;
  assign n30288 = pi14 ? n19805 : n30287;
  assign n30289 = pi13 ? n30282 : n30288;
  assign n30290 = pi15 ? n30207 : n19531;
  assign n30291 = pi14 ? n19235 : n30290;
  assign n30292 = pi13 ? n19805 : n30291;
  assign n30293 = pi12 ? n30289 : n30292;
  assign n30294 = pi11 ? n30281 : n30293;
  assign n30295 = pi19 ? n6057 : n462;
  assign n30296 = pi18 ? n30295 : n19688;
  assign n30297 = pi17 ? n32 : n30296;
  assign n30298 = pi16 ? n32 : n30297;
  assign n30299 = pi15 ? n19691 : n30298;
  assign n30300 = pi15 ? n19691 : n32;
  assign n30301 = pi14 ? n30299 : n30300;
  assign n30302 = pi14 ? n30211 : n19173;
  assign n30303 = pi13 ? n30301 : n30302;
  assign n30304 = pi16 ? n1214 : ~n1683;
  assign n30305 = pi15 ? n30304 : n32;
  assign n30306 = pi14 ? n30026 : n30305;
  assign n30307 = pi13 ? n29963 : n30306;
  assign n30308 = pi12 ? n30303 : n30307;
  assign n30309 = pi14 ? n32 : n29967;
  assign n30310 = pi13 ? n30309 : n32;
  assign n30311 = pi15 ? n32 : n18439;
  assign n30312 = pi18 ? n13080 : n32;
  assign n30313 = pi17 ? n30312 : n1682;
  assign n30314 = pi16 ? n20208 : ~n30313;
  assign n30315 = pi17 ? n1219 : ~n4381;
  assign n30316 = pi16 ? n1471 : n30315;
  assign n30317 = pi15 ? n30314 : n30316;
  assign n30318 = pi14 ? n30311 : n30317;
  assign n30319 = pi15 ? n17903 : n17825;
  assign n30320 = pi14 ? n30319 : n17825;
  assign n30321 = pi13 ? n30318 : n30320;
  assign n30322 = pi12 ? n30310 : n30321;
  assign n30323 = pi11 ? n30308 : n30322;
  assign n30324 = pi10 ? n30294 : n30323;
  assign n30325 = pi09 ? n32 : n30324;
  assign n30326 = pi19 ? n29363 : n28058;
  assign n30327 = pi18 ? n32 : n30326;
  assign n30328 = pi17 ? n32 : n30327;
  assign n30329 = pi19 ? n18778 : ~n17652;
  assign n30330 = pi20 ? n17652 : ~n18408;
  assign n30331 = pi20 ? n18282 : n18281;
  assign n30332 = pi19 ? n30330 : n30331;
  assign n30333 = pi18 ? n30329 : ~n30332;
  assign n30334 = pi20 ? n18415 : ~n18073;
  assign n30335 = pi19 ? n30334 : ~n18281;
  assign n30336 = pi20 ? n18281 : ~n32;
  assign n30337 = pi19 ? n30336 : ~n32;
  assign n30338 = pi18 ? n30335 : ~n30337;
  assign n30339 = pi17 ? n30333 : ~n30338;
  assign n30340 = pi16 ? n30328 : ~n30339;
  assign n30341 = pi16 ? n30273 : ~n2530;
  assign n30342 = pi15 ? n30340 : n30341;
  assign n30343 = pi14 ? n117 : n30342;
  assign n30344 = pi13 ? n32 : n30343;
  assign n30345 = pi15 ? n180 : n20315;
  assign n30346 = pi14 ? n30345 : n32;
  assign n30347 = pi13 ? n180 : n30346;
  assign n30348 = pi12 ? n30344 : n30347;
  assign n30349 = pi20 ? n175 : n1324;
  assign n30350 = pi19 ? n32 : n30349;
  assign n30351 = pi18 ? n32 : n30350;
  assign n30352 = pi19 ? n6398 : n275;
  assign n30353 = pi18 ? n30352 : n4689;
  assign n30354 = pi17 ? n30351 : n30353;
  assign n30355 = pi16 ? n32 : n30354;
  assign n30356 = pi15 ? n30355 : n19805;
  assign n30357 = pi14 ? n19805 : n30356;
  assign n30358 = pi13 ? n30282 : n30357;
  assign n30359 = pi15 ? n19805 : n19868;
  assign n30360 = pi14 ? n19805 : n30359;
  assign n30361 = pi14 ? n19621 : n30290;
  assign n30362 = pi13 ? n30360 : n30361;
  assign n30363 = pi12 ? n30358 : n30362;
  assign n30364 = pi11 ? n30348 : n30363;
  assign n30365 = pi18 ? n30295 : n19811;
  assign n30366 = pi17 ? n32 : n30365;
  assign n30367 = pi16 ? n32 : n30366;
  assign n30368 = pi15 ? n19814 : n30367;
  assign n30369 = pi15 ? n19814 : n32;
  assign n30370 = pi14 ? n30368 : n30369;
  assign n30371 = pi15 ? n41 : n19172;
  assign n30372 = pi14 ? n30371 : n19173;
  assign n30373 = pi13 ? n30370 : n30372;
  assign n30374 = pi14 ? n29969 : n30305;
  assign n30375 = pi13 ? n29963 : n30374;
  assign n30376 = pi12 ? n30373 : n30375;
  assign n30377 = pi15 ? n17903 : n17915;
  assign n30378 = pi14 ? n30377 : n17915;
  assign n30379 = pi13 ? n30318 : n30378;
  assign n30380 = pi12 ? n30310 : n30379;
  assign n30381 = pi11 ? n30376 : n30380;
  assign n30382 = pi10 ? n30364 : n30381;
  assign n30383 = pi09 ? n32 : n30382;
  assign n30384 = pi08 ? n30325 : n30383;
  assign n30385 = pi07 ? n30271 : n30384;
  assign n30386 = pi16 ? n1581 : ~n2530;
  assign n30387 = pi19 ? n5371 : ~n18678;
  assign n30388 = pi18 ? n863 : n30387;
  assign n30389 = pi17 ? n32 : n30388;
  assign n30390 = pi17 ? n19904 : n2410;
  assign n30391 = pi16 ? n30389 : ~n30390;
  assign n30392 = pi15 ? n30386 : n30391;
  assign n30393 = pi14 ? n32 : n30392;
  assign n30394 = pi13 ? n32 : n30393;
  assign n30395 = pi14 ? n180 : n32;
  assign n30396 = pi13 ? n180 : n30395;
  assign n30397 = pi12 ? n30394 : n30396;
  assign n30398 = pi14 ? n19504 : n117;
  assign n30399 = pi20 ? n2385 : n357;
  assign n30400 = pi20 ? n12884 : n17669;
  assign n30401 = pi19 ? n30399 : n30400;
  assign n30402 = pi18 ? n30401 : n20249;
  assign n30403 = pi17 ? n32 : n30402;
  assign n30404 = pi16 ? n32 : n30403;
  assign n30405 = pi20 ? n18129 : n357;
  assign n30406 = pi19 ? n30405 : n21413;
  assign n30407 = pi18 ? n30406 : n19865;
  assign n30408 = pi17 ? n32 : n30407;
  assign n30409 = pi16 ? n32 : n30408;
  assign n30410 = pi15 ? n30404 : n30409;
  assign n30411 = pi14 ? n19868 : n30410;
  assign n30412 = pi13 ? n30398 : n30411;
  assign n30413 = pi15 ? n30409 : n32;
  assign n30414 = pi14 ? n30413 : n19983;
  assign n30415 = pi20 ? n1817 : n12884;
  assign n30416 = pi19 ? n18741 : n30415;
  assign n30417 = pi18 ? n30416 : n19811;
  assign n30418 = pi17 ? n32 : n30417;
  assign n30419 = pi16 ? n32 : n30418;
  assign n30420 = pi15 ? n30419 : n19942;
  assign n30421 = pi14 ? n30011 : n30420;
  assign n30422 = pi13 ? n30414 : n30421;
  assign n30423 = pi12 ? n30412 : n30422;
  assign n30424 = pi11 ? n30397 : n30423;
  assign n30425 = pi18 ? n21255 : n19811;
  assign n30426 = pi17 ? n32 : n30425;
  assign n30427 = pi16 ? n32 : n30426;
  assign n30428 = pi19 ? n507 : n531;
  assign n30429 = pi18 ? n30428 : ~n1548;
  assign n30430 = pi17 ? n32 : n30429;
  assign n30431 = pi16 ? n32 : n30430;
  assign n30432 = pi15 ? n30427 : n30431;
  assign n30433 = pi20 ? n18282 : n13171;
  assign n30434 = pi19 ? n18741 : n30433;
  assign n30435 = pi19 ? n6683 : ~n32;
  assign n30436 = pi18 ? n30434 : ~n30435;
  assign n30437 = pi17 ? n32 : n30436;
  assign n30438 = pi16 ? n32 : n30437;
  assign n30439 = pi15 ? n30438 : n32;
  assign n30440 = pi14 ? n30432 : n30439;
  assign n30441 = pi14 ? n32 : n30211;
  assign n30442 = pi13 ? n30440 : n30441;
  assign n30443 = pi18 ? n4127 : ~n237;
  assign n30444 = pi17 ? n32 : n30443;
  assign n30445 = pi16 ? n32 : n30444;
  assign n30446 = pi15 ? n19172 : n30445;
  assign n30447 = pi17 ? n14395 : n32;
  assign n30448 = pi16 ? n32 : n30447;
  assign n30449 = pi15 ? n19172 : n30448;
  assign n30450 = pi14 ? n30446 : n30449;
  assign n30451 = pi14 ? n19100 : n18143;
  assign n30452 = pi13 ? n30450 : n30451;
  assign n30453 = pi12 ? n30442 : n30452;
  assign n30454 = pi15 ? n32 : n18814;
  assign n30455 = pi14 ? n32 : n30454;
  assign n30456 = pi21 ? n1392 : n32;
  assign n30457 = pi20 ? n32 : n30456;
  assign n30458 = pi19 ? n32 : n30457;
  assign n30459 = pi18 ? n30458 : n32;
  assign n30460 = pi17 ? n32 : n30459;
  assign n30461 = pi20 ? n1385 : n266;
  assign n30462 = pi19 ? n30461 : n32;
  assign n30463 = pi18 ? n30462 : n32;
  assign n30464 = pi17 ? n30463 : n32;
  assign n30465 = pi16 ? n30460 : n30464;
  assign n30466 = pi15 ? n32 : n30465;
  assign n30467 = pi14 ? n32 : n30466;
  assign n30468 = pi13 ? n30455 : n30467;
  assign n30469 = pi18 ? n6163 : n32;
  assign n30470 = pi17 ? n30469 : n2123;
  assign n30471 = pi16 ? n1471 : ~n30470;
  assign n30472 = pi17 ? n28445 : n2123;
  assign n30473 = pi16 ? n19652 : ~n30472;
  assign n30474 = pi15 ? n30471 : n30473;
  assign n30475 = pi18 ? n13668 : n32;
  assign n30476 = pi17 ? n30475 : n2123;
  assign n30477 = pi16 ? n1135 : ~n30476;
  assign n30478 = pi15 ? n30477 : n17903;
  assign n30479 = pi14 ? n30474 : n30478;
  assign n30480 = pi18 ? n6581 : ~n32;
  assign n30481 = pi17 ? n2531 : ~n30480;
  assign n30482 = pi16 ? n3165 : n30481;
  assign n30483 = pi15 ? n17903 : n30482;
  assign n30484 = pi14 ? n17903 : n30483;
  assign n30485 = pi13 ? n30479 : n30484;
  assign n30486 = pi12 ? n30468 : n30485;
  assign n30487 = pi11 ? n30453 : n30486;
  assign n30488 = pi10 ? n30424 : n30487;
  assign n30489 = pi09 ? n32 : n30488;
  assign n30490 = pi16 ? n1581 : ~n2300;
  assign n30491 = pi17 ? n19904 : n2299;
  assign n30492 = pi16 ? n30389 : ~n30491;
  assign n30493 = pi15 ? n30490 : n30492;
  assign n30494 = pi14 ? n32 : n30493;
  assign n30495 = pi13 ? n32 : n30494;
  assign n30496 = pi14 ? n13392 : n32;
  assign n30497 = pi13 ? n13392 : n30496;
  assign n30498 = pi12 ? n30495 : n30497;
  assign n30499 = pi18 ? n32 : n335;
  assign n30500 = pi20 ? n13171 : ~n6085;
  assign n30501 = pi20 ? n3695 : n2358;
  assign n30502 = pi19 ? n30500 : ~n30501;
  assign n30503 = pi18 ? n30502 : ~n20249;
  assign n30504 = pi17 ? n30499 : ~n30503;
  assign n30505 = pi16 ? n32 : n30504;
  assign n30506 = pi19 ? n30405 : n6049;
  assign n30507 = pi18 ? n30506 : n19865;
  assign n30508 = pi17 ? n32 : n30507;
  assign n30509 = pi16 ? n32 : n30508;
  assign n30510 = pi15 ? n30505 : n30509;
  assign n30511 = pi14 ? n19868 : n30510;
  assign n30512 = pi13 ? n117 : n30511;
  assign n30513 = pi15 ? n30509 : n116;
  assign n30514 = pi19 ? n25448 : n32;
  assign n30515 = pi18 ? n32 : n30514;
  assign n30516 = pi17 ? n32 : n30515;
  assign n30517 = pi16 ? n32 : n30516;
  assign n30518 = pi15 ? n30517 : n19868;
  assign n30519 = pi14 ? n30513 : n30518;
  assign n30520 = pi15 ? n19805 : n32;
  assign n30521 = pi20 ? n32 : n8644;
  assign n30522 = pi20 ? n9194 : n17669;
  assign n30523 = pi19 ? n30521 : n30522;
  assign n30524 = pi18 ? n30523 : n19933;
  assign n30525 = pi17 ? n32 : n30524;
  assign n30526 = pi16 ? n32 : n30525;
  assign n30527 = pi15 ? n30526 : n20157;
  assign n30528 = pi14 ? n30520 : n30527;
  assign n30529 = pi13 ? n30519 : n30528;
  assign n30530 = pi12 ? n30512 : n30529;
  assign n30531 = pi11 ? n30498 : n30530;
  assign n30532 = pi18 ? n21255 : n19933;
  assign n30533 = pi17 ? n32 : n30532;
  assign n30534 = pi16 ? n32 : n30533;
  assign n30535 = pi18 ? n30428 : ~n2318;
  assign n30536 = pi17 ? n32 : n30535;
  assign n30537 = pi16 ? n32 : n30536;
  assign n30538 = pi15 ? n30534 : n30537;
  assign n30539 = pi20 ? n17671 : n333;
  assign n30540 = pi19 ? n18741 : n30539;
  assign n30541 = pi18 ? n30540 : ~n316;
  assign n30542 = pi17 ? n32 : n30541;
  assign n30543 = pi16 ? n32 : n30542;
  assign n30544 = pi15 ? n30543 : n32;
  assign n30545 = pi14 ? n30538 : n30544;
  assign n30546 = pi13 ? n30545 : n30441;
  assign n30547 = pi14 ? n18979 : n18143;
  assign n30548 = pi13 ? n30450 : n30547;
  assign n30549 = pi12 ? n30546 : n30548;
  assign n30550 = pi16 ? n270 : n30464;
  assign n30551 = pi15 ? n32 : n30550;
  assign n30552 = pi14 ? n32 : n30551;
  assign n30553 = pi13 ? n30455 : n30552;
  assign n30554 = pi17 ? n30469 : n3351;
  assign n30555 = pi16 ? n1471 : ~n30554;
  assign n30556 = pi16 ? n1214 : ~n30472;
  assign n30557 = pi15 ? n30555 : n30556;
  assign n30558 = pi14 ? n30557 : n30478;
  assign n30559 = pi13 ? n30558 : n30484;
  assign n30560 = pi12 ? n30553 : n30559;
  assign n30561 = pi11 ? n30549 : n30560;
  assign n30562 = pi10 ? n30531 : n30561;
  assign n30563 = pi09 ? n32 : n30562;
  assign n30564 = pi08 ? n30489 : n30563;
  assign n30565 = pi16 ? n1594 : ~n2300;
  assign n30566 = pi19 ? n18678 : n9007;
  assign n30567 = pi18 ? n17848 : n30566;
  assign n30568 = pi17 ? n32 : n30567;
  assign n30569 = pi19 ? n23644 : ~n17649;
  assign n30570 = pi20 ? n357 : n4279;
  assign n30571 = pi20 ? n448 : n1331;
  assign n30572 = pi19 ? n30570 : n30571;
  assign n30573 = pi18 ? n30569 : ~n30572;
  assign n30574 = pi19 ? n32 : ~n207;
  assign n30575 = pi19 ? n12020 : ~n32;
  assign n30576 = pi18 ? n30574 : n30575;
  assign n30577 = pi17 ? n30573 : ~n30576;
  assign n30578 = pi16 ? n30568 : n30577;
  assign n30579 = pi15 ? n30565 : n30578;
  assign n30580 = pi14 ? n32 : n30579;
  assign n30581 = pi13 ? n32 : n30580;
  assign n30582 = pi15 ? n19969 : n72;
  assign n30583 = pi14 ? n30582 : n32;
  assign n30584 = pi13 ? n19969 : n30583;
  assign n30585 = pi12 ? n30581 : n30584;
  assign n30586 = pi14 ? n181 : n180;
  assign n30587 = pi20 ? n310 : ~n2180;
  assign n30588 = pi19 ? n30587 : ~n501;
  assign n30589 = pi18 ? n30588 : ~n20525;
  assign n30590 = pi17 ? n30283 : n30589;
  assign n30591 = pi16 ? n32 : n30590;
  assign n30592 = pi15 ? n20531 : n30591;
  assign n30593 = pi20 ? n310 : ~n785;
  assign n30594 = pi19 ? n30593 : ~n501;
  assign n30595 = pi18 ? n30594 : ~n20525;
  assign n30596 = pi17 ? n30283 : n30595;
  assign n30597 = pi16 ? n32 : n30596;
  assign n30598 = pi15 ? n30597 : n20531;
  assign n30599 = pi14 ? n30592 : n30598;
  assign n30600 = pi13 ? n30586 : n30599;
  assign n30601 = pi15 ? n19805 : n180;
  assign n30602 = pi14 ? n30601 : n19805;
  assign n30603 = pi15 ? n19805 : n17637;
  assign n30604 = pi18 ? n4519 : n6059;
  assign n30605 = pi17 ? n32 : n30604;
  assign n30606 = pi16 ? n32 : n30605;
  assign n30607 = pi19 ? n322 : n6307;
  assign n30608 = pi18 ? n30607 : ~n350;
  assign n30609 = pi17 ? n32 : n30608;
  assign n30610 = pi16 ? n32 : n30609;
  assign n30611 = pi15 ? n30606 : n30610;
  assign n30612 = pi14 ? n30603 : n30611;
  assign n30613 = pi13 ? n30602 : n30612;
  assign n30614 = pi12 ? n30600 : n30613;
  assign n30615 = pi11 ? n30585 : n30614;
  assign n30616 = pi19 ? n1165 : n23193;
  assign n30617 = pi18 ? n30616 : n19933;
  assign n30618 = pi17 ? n32 : n30617;
  assign n30619 = pi16 ? n32 : n30618;
  assign n30620 = pi15 ? n30619 : n30537;
  assign n30621 = pi14 ? n30620 : n28396;
  assign n30622 = pi15 ? n19264 : n32;
  assign n30623 = pi14 ? n32 : n30622;
  assign n30624 = pi13 ? n30621 : n30623;
  assign n30625 = pi18 ? n4380 : ~n237;
  assign n30626 = pi17 ? n32 : n30625;
  assign n30627 = pi16 ? n32 : n30626;
  assign n30628 = pi18 ? n2026 : ~n237;
  assign n30629 = pi17 ? n32 : n30628;
  assign n30630 = pi16 ? n32 : n30629;
  assign n30631 = pi15 ? n30627 : n30630;
  assign n30632 = pi19 ? n1464 : ~n236;
  assign n30633 = pi18 ? n32 : n30632;
  assign n30634 = pi17 ? n30633 : n19170;
  assign n30635 = pi16 ? n32 : n30634;
  assign n30636 = pi19 ? n221 : n267;
  assign n30637 = pi18 ? n32 : n30636;
  assign n30638 = pi17 ? n30637 : n32;
  assign n30639 = pi16 ? n32 : n30638;
  assign n30640 = pi15 ? n30635 : n30639;
  assign n30641 = pi14 ? n30631 : n30640;
  assign n30642 = pi14 ? n19100 : n30211;
  assign n30643 = pi13 ? n30641 : n30642;
  assign n30644 = pi12 ? n30624 : n30643;
  assign n30645 = pi15 ? n18535 : n18814;
  assign n30646 = pi14 ? n32 : n30645;
  assign n30647 = pi18 ? n5005 : n32;
  assign n30648 = pi17 ? n30647 : n32;
  assign n30649 = pi16 ? n270 : n30648;
  assign n30650 = pi15 ? n32 : n30649;
  assign n30651 = pi14 ? n32 : n30650;
  assign n30652 = pi13 ? n30646 : n30651;
  assign n30653 = pi17 ? n30469 : n2325;
  assign n30654 = pi16 ? n1471 : ~n30653;
  assign n30655 = pi18 ? n5731 : n32;
  assign n30656 = pi17 ? n30655 : n2325;
  assign n30657 = pi16 ? n1214 : ~n30656;
  assign n30658 = pi15 ? n30654 : n30657;
  assign n30659 = pi20 ? n32 : ~n1076;
  assign n30660 = pi19 ? n30659 : n32;
  assign n30661 = pi18 ? n30660 : n32;
  assign n30662 = pi17 ? n30661 : n2325;
  assign n30663 = pi16 ? n1214 : ~n30662;
  assign n30664 = pi15 ? n30663 : n19544;
  assign n30665 = pi14 ? n30658 : n30664;
  assign n30666 = pi15 ? n19544 : n19717;
  assign n30667 = pi17 ? n19886 : n18437;
  assign n30668 = pi16 ? n32 : n30667;
  assign n30669 = pi18 ? n6581 : n618;
  assign n30670 = pi17 ? n2531 : ~n30669;
  assign n30671 = pi16 ? n3165 : n30670;
  assign n30672 = pi15 ? n30668 : n30671;
  assign n30673 = pi14 ? n30666 : n30672;
  assign n30674 = pi13 ? n30665 : n30673;
  assign n30675 = pi12 ? n30652 : n30674;
  assign n30676 = pi11 ? n30644 : n30675;
  assign n30677 = pi10 ? n30615 : n30676;
  assign n30678 = pi09 ? n32 : n30677;
  assign n30679 = pi16 ? n1594 : ~n3625;
  assign n30680 = pi19 ? n23644 : ~n5748;
  assign n30681 = pi20 ? n207 : ~n206;
  assign n30682 = pi20 ? n501 : ~n1331;
  assign n30683 = pi19 ? n30681 : n30682;
  assign n30684 = pi18 ? n30680 : n30683;
  assign n30685 = pi18 ? n30574 : n423;
  assign n30686 = pi17 ? n30684 : ~n30685;
  assign n30687 = pi16 ? n30568 : n30686;
  assign n30688 = pi15 ? n30679 : n30687;
  assign n30689 = pi14 ? n32 : n30688;
  assign n30690 = pi13 ? n32 : n30689;
  assign n30691 = pi15 ? n20048 : n106;
  assign n30692 = pi14 ? n30691 : n106;
  assign n30693 = pi14 ? n107 : n32;
  assign n30694 = pi13 ? n30692 : n30693;
  assign n30695 = pi12 ? n30690 : n30694;
  assign n30696 = pi20 ? n32 : n17669;
  assign n30697 = pi19 ? n32 : n30696;
  assign n30698 = pi18 ? n32 : n30697;
  assign n30699 = pi20 ? n2180 : n1076;
  assign n30700 = pi19 ? n30587 : ~n30699;
  assign n30701 = pi20 ? n17671 : ~n32;
  assign n30702 = pi19 ? n30701 : ~n32;
  assign n30703 = pi18 ? n30700 : ~n30702;
  assign n30704 = pi17 ? n30698 : n30703;
  assign n30705 = pi16 ? n32 : n30704;
  assign n30706 = pi15 ? n20531 : n30705;
  assign n30707 = pi19 ? n30593 : ~n30699;
  assign n30708 = pi18 ? n30707 : ~n30702;
  assign n30709 = pi17 ? n30283 : n30708;
  assign n30710 = pi16 ? n32 : n30709;
  assign n30711 = pi15 ? n30710 : n20531;
  assign n30712 = pi14 ? n30706 : n30711;
  assign n30713 = pi13 ? n30586 : n30712;
  assign n30714 = pi15 ? n19805 : n20531;
  assign n30715 = pi14 ? n30601 : n30714;
  assign n30716 = pi15 ? n19868 : n17637;
  assign n30717 = pi14 ? n30716 : n30611;
  assign n30718 = pi13 ? n30715 : n30717;
  assign n30719 = pi12 ? n30713 : n30718;
  assign n30720 = pi11 ? n30695 : n30719;
  assign n30721 = pi18 ? n30616 : n4689;
  assign n30722 = pi17 ? n32 : n30721;
  assign n30723 = pi16 ? n32 : n30722;
  assign n30724 = pi18 ? n30428 : ~n344;
  assign n30725 = pi17 ? n32 : n30724;
  assign n30726 = pi16 ? n32 : n30725;
  assign n30727 = pi15 ? n30723 : n30726;
  assign n30728 = pi14 ? n30727 : n28396;
  assign n30729 = pi15 ? n19628 : n32;
  assign n30730 = pi14 ? n32 : n30729;
  assign n30731 = pi13 ? n30728 : n30730;
  assign n30732 = pi14 ? n18979 : n30211;
  assign n30733 = pi13 ? n30641 : n30732;
  assign n30734 = pi12 ? n30731 : n30733;
  assign n30735 = pi18 ? n5164 : n32;
  assign n30736 = pi17 ? n30735 : n32;
  assign n30737 = pi16 ? n270 : n30736;
  assign n30738 = pi15 ? n32 : n30737;
  assign n30739 = pi14 ? n32 : n30738;
  assign n30740 = pi13 ? n30646 : n30739;
  assign n30741 = pi18 ? n4983 : n32;
  assign n30742 = pi17 ? n30741 : n2325;
  assign n30743 = pi16 ? n1214 : ~n30742;
  assign n30744 = pi15 ? n30743 : n19717;
  assign n30745 = pi14 ? n30658 : n30744;
  assign n30746 = pi14 ? n19717 : n30672;
  assign n30747 = pi13 ? n30745 : n30746;
  assign n30748 = pi12 ? n30740 : n30747;
  assign n30749 = pi11 ? n30734 : n30748;
  assign n30750 = pi10 ? n30720 : n30749;
  assign n30751 = pi09 ? n32 : n30750;
  assign n30752 = pi08 ? n30678 : n30751;
  assign n30753 = pi07 ? n30564 : n30752;
  assign n30754 = pi06 ? n30385 : n30753;
  assign n30755 = pi05 ? n30180 : n30754;
  assign n30756 = pi20 ? n333 : ~n321;
  assign n30757 = pi19 ? n30756 : n1844;
  assign n30758 = pi18 ? n30757 : ~n23073;
  assign n30759 = pi17 ? n18533 : n30758;
  assign n30760 = pi16 ? n32 : n30759;
  assign n30761 = pi20 ? n333 : n32;
  assign n30762 = pi19 ? n30761 : n1844;
  assign n30763 = pi20 ? n831 : ~n32;
  assign n30764 = pi19 ? n30763 : ~n32;
  assign n30765 = pi18 ? n30762 : ~n30764;
  assign n30766 = pi17 ? n18533 : n30765;
  assign n30767 = pi16 ? n32 : n30766;
  assign n30768 = pi15 ? n30760 : n30767;
  assign n30769 = pi14 ? n32 : n30768;
  assign n30770 = pi13 ? n32 : n30769;
  assign n30771 = pi14 ? n20127 : n32;
  assign n30772 = pi13 ? n20048 : n30771;
  assign n30773 = pi12 ? n30770 : n30772;
  assign n30774 = pi14 ? n19862 : n32;
  assign n30775 = pi19 ? n11879 : ~n6307;
  assign n30776 = pi18 ? n30775 : n19848;
  assign n30777 = pi17 ? n32 : n30776;
  assign n30778 = pi16 ? n32 : n30777;
  assign n30779 = pi19 ? n9007 : ~n6307;
  assign n30780 = pi19 ? n27066 : n32;
  assign n30781 = pi18 ? n30779 : n30780;
  assign n30782 = pi17 ? n32 : n30781;
  assign n30783 = pi16 ? n32 : n30782;
  assign n30784 = pi15 ? n30778 : n30783;
  assign n30785 = pi14 ? n30784 : n13392;
  assign n30786 = pi13 ? n30774 : n30785;
  assign n30787 = pi15 ? n13392 : n20136;
  assign n30788 = pi15 ? n20136 : n32;
  assign n30789 = pi14 ? n30787 : n30788;
  assign n30790 = pi18 ? n32 : n20366;
  assign n30791 = pi17 ? n32 : n30790;
  assign n30792 = pi16 ? n32 : n30791;
  assign n30793 = pi15 ? n18657 : n30792;
  assign n30794 = pi18 ? n209 : n4689;
  assign n30795 = pi17 ? n32 : n30794;
  assign n30796 = pi16 ? n32 : n30795;
  assign n30797 = pi18 ? n7038 : ~n344;
  assign n30798 = pi17 ? n32 : n30797;
  assign n30799 = pi16 ? n32 : n30798;
  assign n30800 = pi15 ? n30796 : n30799;
  assign n30801 = pi14 ? n30793 : n30800;
  assign n30802 = pi13 ? n30789 : n30801;
  assign n30803 = pi12 ? n30786 : n30802;
  assign n30804 = pi11 ? n30773 : n30803;
  assign n30805 = pi18 ? n496 : ~n344;
  assign n30806 = pi17 ? n16103 : n30805;
  assign n30807 = pi16 ? n32 : n30806;
  assign n30808 = pi20 ? n342 : ~n14286;
  assign n30809 = pi19 ? n32 : n30808;
  assign n30810 = pi18 ? n30809 : ~n350;
  assign n30811 = pi17 ? n16103 : n30810;
  assign n30812 = pi16 ? n32 : n30811;
  assign n30813 = pi15 ? n30807 : n30812;
  assign n30814 = pi14 ? n30813 : n32;
  assign n30815 = pi13 ? n30814 : n32;
  assign n30816 = pi19 ? n507 : ~n4406;
  assign n30817 = pi18 ? n32 : n30816;
  assign n30818 = pi18 ? n268 : ~n237;
  assign n30819 = pi17 ? n30817 : n30818;
  assign n30820 = pi16 ? n32 : n30819;
  assign n30821 = pi19 ? n322 : ~n28179;
  assign n30822 = pi18 ? n32 : n30821;
  assign n30823 = pi19 ? n20006 : n4126;
  assign n30824 = pi18 ? n30823 : ~n237;
  assign n30825 = pi17 ? n30822 : n30824;
  assign n30826 = pi16 ? n32 : n30825;
  assign n30827 = pi15 ? n30820 : n30826;
  assign n30828 = pi19 ? n236 : ~n247;
  assign n30829 = pi18 ? n30828 : ~n28193;
  assign n30830 = pi19 ? n6307 : n13069;
  assign n30831 = pi18 ? n30830 : ~n350;
  assign n30832 = pi17 ? n30829 : ~n30831;
  assign n30833 = pi16 ? n19171 : ~n30832;
  assign n30834 = pi19 ? n321 : n18390;
  assign n30835 = pi18 ? n4127 : ~n30834;
  assign n30836 = pi17 ? n32 : n30835;
  assign n30837 = pi20 ? n266 : n518;
  assign n30838 = pi19 ? n30837 : n5748;
  assign n30839 = pi19 ? n236 : n349;
  assign n30840 = pi18 ? n30838 : ~n30839;
  assign n30841 = pi18 ? n684 : ~n6059;
  assign n30842 = pi17 ? n30840 : n30841;
  assign n30843 = pi16 ? n30836 : ~n30842;
  assign n30844 = pi15 ? n30833 : n30843;
  assign n30845 = pi14 ? n30827 : n30844;
  assign n30846 = pi18 ? n863 : n342;
  assign n30847 = pi17 ? n32 : n30846;
  assign n30848 = pi19 ? n18728 : n266;
  assign n30849 = pi20 ? n220 : ~n246;
  assign n30850 = pi19 ? n30849 : ~n17766;
  assign n30851 = pi18 ? n30848 : ~n30850;
  assign n30852 = pi19 ? n7642 : ~n9345;
  assign n30853 = pi18 ? n30852 : n32;
  assign n30854 = pi17 ? n30851 : n30853;
  assign n30855 = pi16 ? n30847 : n30854;
  assign n30856 = pi15 ? n19531 : n30855;
  assign n30857 = pi14 ? n29601 : n30856;
  assign n30858 = pi13 ? n30845 : n30857;
  assign n30859 = pi12 ? n30815 : n30858;
  assign n30860 = pi18 ? n268 : n18532;
  assign n30861 = pi17 ? n32 : n30860;
  assign n30862 = pi16 ? n32 : n30861;
  assign n30863 = pi15 ? n32 : n30862;
  assign n30864 = pi14 ? n32 : n30863;
  assign n30865 = pi19 ? n321 : n4342;
  assign n30866 = pi18 ? n940 : ~n30865;
  assign n30867 = pi17 ? n32 : n30866;
  assign n30868 = pi19 ? n4964 : ~n4342;
  assign n30869 = pi18 ? n30868 : ~n32;
  assign n30870 = pi17 ? n30869 : ~n5077;
  assign n30871 = pi16 ? n30867 : n30870;
  assign n30872 = pi15 ? n32 : n30871;
  assign n30873 = pi14 ? n30211 : n30872;
  assign n30874 = pi13 ? n30864 : n30873;
  assign n30875 = pi17 ? n28440 : n2325;
  assign n30876 = pi16 ? n1471 : ~n30875;
  assign n30877 = pi18 ? n6581 : n32;
  assign n30878 = pi17 ? n30877 : n2325;
  assign n30879 = pi16 ? n1471 : ~n30878;
  assign n30880 = pi15 ? n30876 : n30879;
  assign n30881 = pi17 ? n1542 : n19785;
  assign n30882 = pi16 ? n32 : n30881;
  assign n30883 = pi15 ? n30882 : n19172;
  assign n30884 = pi14 ? n30880 : n30883;
  assign n30885 = pi17 ? n16103 : n18437;
  assign n30886 = pi16 ? n32 : n30885;
  assign n30887 = pi15 ? n19717 : n30886;
  assign n30888 = pi18 ? n12890 : n618;
  assign n30889 = pi17 ? n15228 : ~n30888;
  assign n30890 = pi16 ? n32 : n30889;
  assign n30891 = pi18 ? n268 : n6059;
  assign n30892 = pi17 ? n32 : n30891;
  assign n30893 = pi17 ? n21275 : n2123;
  assign n30894 = pi16 ? n30892 : ~n30893;
  assign n30895 = pi15 ? n30890 : n30894;
  assign n30896 = pi14 ? n30887 : n30895;
  assign n30897 = pi13 ? n30884 : n30896;
  assign n30898 = pi12 ? n30874 : n30897;
  assign n30899 = pi11 ? n30859 : n30898;
  assign n30900 = pi10 ? n30804 : n30899;
  assign n30901 = pi09 ? n32 : n30900;
  assign n30902 = pi18 ? n14153 : ~n20680;
  assign n30903 = pi17 ? n32 : n30902;
  assign n30904 = pi16 ? n32 : n30903;
  assign n30905 = pi20 ? n339 : n141;
  assign n30906 = pi19 ? n30905 : ~n32;
  assign n30907 = pi18 ? n32 : ~n30906;
  assign n30908 = pi17 ? n32 : n30907;
  assign n30909 = pi16 ? n32 : n30908;
  assign n30910 = pi15 ? n30904 : n30909;
  assign n30911 = pi14 ? n32 : n30910;
  assign n30912 = pi13 ? n32 : n30911;
  assign n30913 = pi15 ? n146 : n13684;
  assign n30914 = pi14 ? n30913 : n13684;
  assign n30915 = pi15 ? n13684 : n32;
  assign n30916 = pi14 ? n30915 : n32;
  assign n30917 = pi13 ? n30914 : n30916;
  assign n30918 = pi12 ? n30912 : n30917;
  assign n30919 = pi14 ? n19862 : n19969;
  assign n30920 = pi13 ? n30919 : n30785;
  assign n30921 = pi15 ? n19972 : n32;
  assign n30922 = pi14 ? n13392 : n30921;
  assign n30923 = pi15 ? n18657 : n30517;
  assign n30924 = pi18 ? n209 : n20249;
  assign n30925 = pi17 ? n32 : n30924;
  assign n30926 = pi16 ? n32 : n30925;
  assign n30927 = pi18 ? n7038 : ~n2304;
  assign n30928 = pi17 ? n32 : n30927;
  assign n30929 = pi16 ? n32 : n30928;
  assign n30930 = pi15 ? n30926 : n30929;
  assign n30931 = pi14 ? n30923 : n30930;
  assign n30932 = pi13 ? n30922 : n30931;
  assign n30933 = pi12 ? n30920 : n30932;
  assign n30934 = pi11 ? n30918 : n30933;
  assign n30935 = pi18 ? n496 : ~n2304;
  assign n30936 = pi17 ? n16103 : n30935;
  assign n30937 = pi16 ? n32 : n30936;
  assign n30938 = pi15 ? n30937 : n30812;
  assign n30939 = pi14 ? n30938 : n32;
  assign n30940 = pi13 ? n30939 : n32;
  assign n30941 = pi16 ? n1135 : ~n1808;
  assign n30942 = pi14 ? n30941 : n30856;
  assign n30943 = pi13 ? n30845 : n30942;
  assign n30944 = pi12 ? n30940 : n30943;
  assign n30945 = pi18 ? n940 : n1942;
  assign n30946 = pi17 ? n30869 : ~n30945;
  assign n30947 = pi16 ? n30867 : n30946;
  assign n30948 = pi15 ? n32 : n30947;
  assign n30949 = pi14 ? n30211 : n30948;
  assign n30950 = pi13 ? n30864 : n30949;
  assign n30951 = pi17 ? n28440 : n2136;
  assign n30952 = pi16 ? n1471 : ~n30951;
  assign n30953 = pi17 ? n30877 : n1943;
  assign n30954 = pi16 ? n1471 : ~n30953;
  assign n30955 = pi15 ? n30952 : n30954;
  assign n30956 = pi15 ? n19787 : n19172;
  assign n30957 = pi14 ? n30955 : n30956;
  assign n30958 = pi17 ? n21275 : n3351;
  assign n30959 = pi16 ? n30892 : ~n30958;
  assign n30960 = pi15 ? n30890 : n30959;
  assign n30961 = pi14 ? n30887 : n30960;
  assign n30962 = pi13 ? n30957 : n30961;
  assign n30963 = pi12 ? n30950 : n30962;
  assign n30964 = pi11 ? n30944 : n30963;
  assign n30965 = pi10 ? n30934 : n30964;
  assign n30966 = pi09 ? n32 : n30965;
  assign n30967 = pi08 ? n30901 : n30966;
  assign n30968 = pi19 ? n11374 : n32;
  assign n30969 = pi20 ? n501 : n141;
  assign n30970 = pi19 ? n30969 : ~n32;
  assign n30971 = pi18 ? n30968 : ~n30970;
  assign n30972 = pi17 ? n32 : n30971;
  assign n30973 = pi16 ? n32 : n30972;
  assign n30974 = pi15 ? n30973 : n146;
  assign n30975 = pi14 ? n32 : n30974;
  assign n30976 = pi13 ? n32 : n30975;
  assign n30977 = pi15 ? n146 : n106;
  assign n30978 = pi14 ? n30977 : n20049;
  assign n30979 = pi13 ? n146 : n30978;
  assign n30980 = pi12 ? n30976 : n30979;
  assign n30981 = pi15 ? n19972 : n20048;
  assign n30982 = pi14 ? n32 : n30981;
  assign n30983 = pi20 ? n6621 : ~n6050;
  assign n30984 = pi20 ? n29457 : n310;
  assign n30985 = pi19 ? n30983 : ~n30984;
  assign n30986 = pi19 ? n12854 : n32;
  assign n30987 = pi18 ? n30985 : n30986;
  assign n30988 = pi17 ? n32 : n30987;
  assign n30989 = pi16 ? n32 : n30988;
  assign n30990 = pi19 ? n29473 : ~n30984;
  assign n30991 = pi18 ? n30990 : n30986;
  assign n30992 = pi17 ? n32 : n30991;
  assign n30993 = pi16 ? n32 : n30992;
  assign n30994 = pi15 ? n30989 : n30993;
  assign n30995 = pi14 ? n30994 : n30981;
  assign n30996 = pi13 ? n30982 : n30995;
  assign n30997 = pi18 ? n863 : n177;
  assign n30998 = pi17 ? n32 : n30997;
  assign n30999 = pi16 ? n32 : n30998;
  assign n31000 = pi15 ? n19972 : n30999;
  assign n31001 = pi14 ? n19972 : n31000;
  assign n31002 = pi20 ? n18762 : ~n32;
  assign n31003 = pi19 ? n31002 : ~n32;
  assign n31004 = pi18 ? n7623 : ~n31003;
  assign n31005 = pi17 ? n32 : n31004;
  assign n31006 = pi16 ? n32 : n31005;
  assign n31007 = pi15 ? n30999 : n31006;
  assign n31008 = pi18 ? n18710 : n20327;
  assign n31009 = pi17 ? n32 : n31008;
  assign n31010 = pi16 ? n32 : n31009;
  assign n31011 = pi19 ? n11546 : ~n32;
  assign n31012 = pi18 ? n880 : ~n31011;
  assign n31013 = pi17 ? n32 : n31012;
  assign n31014 = pi16 ? n32 : n31013;
  assign n31015 = pi15 ? n31010 : n31014;
  assign n31016 = pi14 ? n31007 : n31015;
  assign n31017 = pi13 ? n31001 : n31016;
  assign n31018 = pi12 ? n30996 : n31017;
  assign n31019 = pi11 ? n30980 : n31018;
  assign n31020 = pi18 ? n22885 : ~n31011;
  assign n31021 = pi17 ? n32 : n31020;
  assign n31022 = pi16 ? n32 : n31021;
  assign n31023 = pi18 ? n22885 : ~n350;
  assign n31024 = pi17 ? n16103 : n31023;
  assign n31025 = pi16 ? n32 : n31024;
  assign n31026 = pi15 ? n31022 : n31025;
  assign n31027 = pi14 ? n31026 : n32;
  assign n31028 = pi13 ? n31027 : n19236;
  assign n31029 = pi19 ? n236 : ~n4721;
  assign n31030 = pi18 ? n31029 : n1548;
  assign n31031 = pi17 ? n14983 : ~n31030;
  assign n31032 = pi16 ? n32 : n31031;
  assign n31033 = pi19 ? n322 : ~n1757;
  assign n31034 = pi18 ? n19811 : n31033;
  assign n31035 = pi19 ? n3692 : ~n507;
  assign n31036 = pi21 ? n7478 : ~n259;
  assign n31037 = pi20 ? n31036 : n32;
  assign n31038 = pi19 ? n31037 : n32;
  assign n31039 = pi18 ? n31035 : ~n31038;
  assign n31040 = pi17 ? n31034 : ~n31039;
  assign n31041 = pi16 ? n32 : n31040;
  assign n31042 = pi15 ? n31032 : n31041;
  assign n31043 = pi19 ? n5694 : ~n321;
  assign n31044 = pi18 ? n917 : ~n31043;
  assign n31045 = pi17 ? n32 : n31044;
  assign n31046 = pi19 ? n4342 : ~n21296;
  assign n31047 = pi18 ? n31046 : n248;
  assign n31048 = pi18 ? n209 : n1548;
  assign n31049 = pi17 ? n31047 : n31048;
  assign n31050 = pi16 ? n31045 : ~n31049;
  assign n31051 = pi18 ? n16847 : n1548;
  assign n31052 = pi17 ? n32 : n31051;
  assign n31053 = pi16 ? n1135 : ~n31052;
  assign n31054 = pi15 ? n31050 : n31053;
  assign n31055 = pi14 ? n31042 : n31054;
  assign n31056 = pi16 ? n19652 : ~n1808;
  assign n31057 = pi18 ? n32 : ~n19811;
  assign n31058 = pi17 ? n32 : n31057;
  assign n31059 = pi16 ? n1214 : ~n31058;
  assign n31060 = pi15 ? n31056 : n31059;
  assign n31061 = pi19 ? n30849 : ~n9007;
  assign n31062 = pi18 ? n30848 : ~n31061;
  assign n31063 = pi18 ? n30852 : n19232;
  assign n31064 = pi17 ? n31062 : n31063;
  assign n31065 = pi16 ? n30847 : n31064;
  assign n31066 = pi15 ? n19814 : n31065;
  assign n31067 = pi14 ? n31060 : n31066;
  assign n31068 = pi13 ? n31055 : n31067;
  assign n31069 = pi12 ? n31028 : n31068;
  assign n31070 = pi15 ? n32 : n19264;
  assign n31071 = pi19 ? n4964 : n531;
  assign n31072 = pi18 ? n31071 : ~n32;
  assign n31073 = pi18 ? n940 : n814;
  assign n31074 = pi17 ? n31072 : ~n31073;
  assign n31075 = pi16 ? n30867 : n31074;
  assign n31076 = pi15 ? n19267 : n31075;
  assign n31077 = pi14 ? n31070 : n31076;
  assign n31078 = pi13 ? n30864 : n31077;
  assign n31079 = pi18 ? n25595 : n32;
  assign n31080 = pi17 ? n31079 : n2136;
  assign n31081 = pi16 ? n20208 : ~n31080;
  assign n31082 = pi17 ? n30877 : n2136;
  assign n31083 = pi16 ? n1471 : ~n31082;
  assign n31084 = pi15 ? n31081 : n31083;
  assign n31085 = pi18 ? n880 : ~n814;
  assign n31086 = pi17 ? n32 : n31085;
  assign n31087 = pi16 ? n32 : n31086;
  assign n31088 = pi15 ? n31087 : n19172;
  assign n31089 = pi14 ? n31084 : n31088;
  assign n31090 = pi17 ? n16099 : n18812;
  assign n31091 = pi16 ? n32 : n31090;
  assign n31092 = pi15 ? n19172 : n31091;
  assign n31093 = pi19 ? n349 : ~n507;
  assign n31094 = pi18 ? n31093 : n237;
  assign n31095 = pi17 ? n16042 : ~n31094;
  assign n31096 = pi16 ? n32 : n31095;
  assign n31097 = pi19 ? n22698 : n175;
  assign n31098 = pi18 ? n268 : n31097;
  assign n31099 = pi17 ? n32 : n31098;
  assign n31100 = pi20 ? n32 : ~n17665;
  assign n31101 = pi19 ? n31100 : ~n23688;
  assign n31102 = pi19 ? n8611 : ~n32;
  assign n31103 = pi18 ? n31101 : ~n31102;
  assign n31104 = pi17 ? n31103 : n2325;
  assign n31105 = pi16 ? n31099 : ~n31104;
  assign n31106 = pi15 ? n31096 : n31105;
  assign n31107 = pi14 ? n31092 : n31106;
  assign n31108 = pi13 ? n31089 : n31107;
  assign n31109 = pi12 ? n31078 : n31108;
  assign n31110 = pi11 ? n31069 : n31109;
  assign n31111 = pi10 ? n31019 : n31110;
  assign n31112 = pi09 ? n32 : n31111;
  assign n31113 = pi19 ? n9890 : ~n32;
  assign n31114 = pi18 ? n30968 : ~n31113;
  assign n31115 = pi17 ? n32 : n31114;
  assign n31116 = pi16 ? n32 : n31115;
  assign n31117 = pi15 ? n31116 : n13952;
  assign n31118 = pi14 ? n32 : n31117;
  assign n31119 = pi13 ? n32 : n31118;
  assign n31120 = pi15 ? n13952 : n32;
  assign n31121 = pi14 ? n31120 : n32;
  assign n31122 = pi13 ? n13952 : n31121;
  assign n31123 = pi12 ? n31119 : n31122;
  assign n31124 = pi15 ? n20493 : n30999;
  assign n31125 = pi14 ? n21521 : n31124;
  assign n31126 = pi21 ? n309 : n100;
  assign n31127 = pi20 ? n31126 : ~n32;
  assign n31128 = pi19 ? n31127 : ~n32;
  assign n31129 = pi18 ? n7623 : ~n31128;
  assign n31130 = pi17 ? n32 : n31129;
  assign n31131 = pi16 ? n32 : n31130;
  assign n31132 = pi15 ? n30999 : n31131;
  assign n31133 = pi18 ? n880 : ~n20518;
  assign n31134 = pi17 ? n32 : n31133;
  assign n31135 = pi16 ? n32 : n31134;
  assign n31136 = pi15 ? n31010 : n31135;
  assign n31137 = pi14 ? n31132 : n31136;
  assign n31138 = pi13 ? n31125 : n31137;
  assign n31139 = pi12 ? n30996 : n31138;
  assign n31140 = pi11 ? n31123 : n31139;
  assign n31141 = pi18 ? n31035 : ~n29919;
  assign n31142 = pi17 ? n31034 : ~n31141;
  assign n31143 = pi16 ? n32 : n31142;
  assign n31144 = pi15 ? n31032 : n31143;
  assign n31145 = pi14 ? n31144 : n31054;
  assign n31146 = pi16 ? n1214 : ~n1808;
  assign n31147 = pi15 ? n31146 : n31059;
  assign n31148 = pi18 ? n30852 : n19318;
  assign n31149 = pi17 ? n31062 : n31148;
  assign n31150 = pi16 ? n30847 : n31149;
  assign n31151 = pi15 ? n19814 : n31150;
  assign n31152 = pi14 ? n31147 : n31151;
  assign n31153 = pi13 ? n31145 : n31152;
  assign n31154 = pi12 ? n31028 : n31153;
  assign n31155 = pi20 ? n16195 : ~n32;
  assign n31156 = pi19 ? n31155 : ~n32;
  assign n31157 = pi18 ? n32 : ~n31156;
  assign n31158 = pi17 ? n32 : n31157;
  assign n31159 = pi16 ? n32 : n31158;
  assign n31160 = pi15 ? n32 : n31159;
  assign n31161 = pi18 ? n940 : n1813;
  assign n31162 = pi17 ? n31072 : ~n31161;
  assign n31163 = pi16 ? n30867 : n31162;
  assign n31164 = pi15 ? n19267 : n31163;
  assign n31165 = pi14 ? n31160 : n31164;
  assign n31166 = pi13 ? n30864 : n31165;
  assign n31167 = pi12 ? n31166 : n31108;
  assign n31168 = pi11 ? n31154 : n31167;
  assign n31169 = pi10 ? n31140 : n31168;
  assign n31170 = pi09 ? n32 : n31169;
  assign n31171 = pi08 ? n31112 : n31170;
  assign n31172 = pi07 ? n30967 : n31171;
  assign n31173 = pi15 ? n13952 : n671;
  assign n31174 = pi14 ? n20416 : n31173;
  assign n31175 = pi13 ? n32 : n31174;
  assign n31176 = pi15 ? n671 : n13952;
  assign n31177 = pi14 ? n31176 : n13952;
  assign n31178 = pi13 ? n31177 : n31121;
  assign n31179 = pi12 ? n31175 : n31178;
  assign n31180 = pi15 ? n20048 : n13684;
  assign n31181 = pi14 ? n32 : n31180;
  assign n31182 = pi20 ? n3523 : ~n18282;
  assign n31183 = pi20 ? n18282 : n1817;
  assign n31184 = pi19 ? n31182 : ~n31183;
  assign n31185 = pi20 ? n820 : ~n141;
  assign n31186 = pi19 ? n31185 : n32;
  assign n31187 = pi18 ? n31184 : n31186;
  assign n31188 = pi17 ? n32 : n31187;
  assign n31189 = pi16 ? n32 : n31188;
  assign n31190 = pi20 ? n32 : ~n18253;
  assign n31191 = pi19 ? n31190 : ~n30699;
  assign n31192 = pi18 ? n31191 : n31186;
  assign n31193 = pi17 ? n32 : n31192;
  assign n31194 = pi16 ? n32 : n31193;
  assign n31195 = pi15 ? n31189 : n31194;
  assign n31196 = pi19 ? n28070 : ~n30699;
  assign n31197 = pi20 ? n18245 : ~n141;
  assign n31198 = pi19 ? n31197 : n32;
  assign n31199 = pi18 ? n31196 : n31198;
  assign n31200 = pi17 ? n32 : n31199;
  assign n31201 = pi16 ? n32 : n31200;
  assign n31202 = pi20 ? n2180 : n9491;
  assign n31203 = pi19 ? n6398 : ~n31202;
  assign n31204 = pi20 ? n18408 : ~n141;
  assign n31205 = pi19 ? n31204 : n32;
  assign n31206 = pi18 ? n31203 : n31205;
  assign n31207 = pi17 ? n32 : n31206;
  assign n31208 = pi16 ? n32 : n31207;
  assign n31209 = pi15 ? n31201 : n31208;
  assign n31210 = pi14 ? n31195 : n31209;
  assign n31211 = pi13 ? n31181 : n31210;
  assign n31212 = pi20 ? n67 : ~n141;
  assign n31213 = pi19 ? n31212 : n32;
  assign n31214 = pi18 ? n32 : n31213;
  assign n31215 = pi17 ? n32 : n31214;
  assign n31216 = pi16 ? n32 : n31215;
  assign n31217 = pi15 ? n13380 : n31216;
  assign n31218 = pi15 ? n20493 : n32;
  assign n31219 = pi14 ? n31217 : n31218;
  assign n31220 = pi15 ? n17903 : n20531;
  assign n31221 = pi21 ? n405 : n20130;
  assign n31222 = pi20 ? n31221 : n32;
  assign n31223 = pi19 ? n31222 : n32;
  assign n31224 = pi18 ? n268 : n31223;
  assign n31225 = pi17 ? n32 : n31224;
  assign n31226 = pi16 ? n32 : n31225;
  assign n31227 = pi18 ? n268 : n13086;
  assign n31228 = pi17 ? n32 : n31227;
  assign n31229 = pi16 ? n32 : n31228;
  assign n31230 = pi15 ? n31226 : n31229;
  assign n31231 = pi14 ? n31220 : n31230;
  assign n31232 = pi13 ? n31219 : n31231;
  assign n31233 = pi12 ? n31211 : n31232;
  assign n31234 = pi11 ? n31179 : n31233;
  assign n31235 = pi14 ? n20447 : n32;
  assign n31236 = pi13 ? n31235 : n32;
  assign n31237 = pi19 ? n6988 : n20555;
  assign n31238 = pi18 ? n31237 : ~n32;
  assign n31239 = pi17 ? n2736 : ~n31238;
  assign n31240 = pi16 ? n32 : n31239;
  assign n31241 = pi18 ? n20615 : n702;
  assign n31242 = pi17 ? n31241 : ~n4723;
  assign n31243 = pi16 ? n32 : n31242;
  assign n31244 = pi15 ? n31240 : n31243;
  assign n31245 = pi18 ? n16295 : n32;
  assign n31246 = pi17 ? n31245 : n1697;
  assign n31247 = pi16 ? n1471 : ~n31246;
  assign n31248 = pi17 ? n32 : n31048;
  assign n31249 = pi16 ? n1135 : ~n31248;
  assign n31250 = pi15 ? n31247 : n31249;
  assign n31251 = pi14 ? n31244 : n31250;
  assign n31252 = pi17 ? n32 : n4685;
  assign n31253 = pi16 ? n1135 : ~n31252;
  assign n31254 = pi18 ? n1054 : ~n32;
  assign n31255 = pi17 ? n32 : n31254;
  assign n31256 = pi16 ? n1471 : ~n31255;
  assign n31257 = pi15 ? n31253 : n31256;
  assign n31258 = pi17 ? n15850 : n28803;
  assign n31259 = pi16 ? n1214 : ~n31258;
  assign n31260 = pi18 ? n14982 : n496;
  assign n31261 = pi17 ? n31260 : n31072;
  assign n31262 = pi16 ? n1471 : ~n31261;
  assign n31263 = pi15 ? n31259 : n31262;
  assign n31264 = pi14 ? n31257 : n31263;
  assign n31265 = pi13 ? n31251 : n31264;
  assign n31266 = pi12 ? n31236 : n31265;
  assign n31267 = pi15 ? n18535 : n18798;
  assign n31268 = pi14 ? n32 : n31267;
  assign n31269 = pi13 ? n32 : n31268;
  assign n31270 = pi18 ? n16847 : ~n1813;
  assign n31271 = pi17 ? n32 : n31270;
  assign n31272 = pi16 ? n32 : n31271;
  assign n31273 = pi18 ? n268 : ~n1813;
  assign n31274 = pi17 ? n32 : n31273;
  assign n31275 = pi16 ? n32 : n31274;
  assign n31276 = pi15 ? n31272 : n31275;
  assign n31277 = pi17 ? n16848 : n19396;
  assign n31278 = pi16 ? n32 : n31277;
  assign n31279 = pi15 ? n31278 : n19264;
  assign n31280 = pi14 ? n31276 : n31279;
  assign n31281 = pi17 ? n32 : n30818;
  assign n31282 = pi16 ? n32 : n31281;
  assign n31283 = pi17 ? n15850 : n30818;
  assign n31284 = pi16 ? n32 : n31283;
  assign n31285 = pi15 ? n31282 : n31284;
  assign n31286 = pi19 ? n531 : n5371;
  assign n31287 = pi18 ? n31286 : n1942;
  assign n31288 = pi17 ? n3067 : ~n31287;
  assign n31289 = pi16 ? n32 : n31288;
  assign n31290 = pi19 ? n4342 : n9007;
  assign n31291 = pi18 ? n31290 : n323;
  assign n31292 = pi17 ? n31291 : ~n2325;
  assign n31293 = pi16 ? n32 : n31292;
  assign n31294 = pi15 ? n31289 : n31293;
  assign n31295 = pi14 ? n31285 : n31294;
  assign n31296 = pi13 ? n31280 : n31295;
  assign n31297 = pi12 ? n31269 : n31296;
  assign n31298 = pi11 ? n31266 : n31297;
  assign n31299 = pi10 ? n31234 : n31298;
  assign n31300 = pi09 ? n32 : n31299;
  assign n31301 = pi15 ? n32 : n671;
  assign n31302 = pi15 ? n20477 : n486;
  assign n31303 = pi14 ? n31301 : n31302;
  assign n31304 = pi13 ? n32 : n31303;
  assign n31305 = pi14 ? n22320 : n32;
  assign n31306 = pi13 ? n486 : n31305;
  assign n31307 = pi12 ? n31304 : n31306;
  assign n31308 = pi14 ? n20416 : n20301;
  assign n31309 = pi20 ? n17652 : n5854;
  assign n31310 = pi19 ? n31182 : ~n31309;
  assign n31311 = pi20 ? n17669 : ~n339;
  assign n31312 = pi19 ? n31311 : n32;
  assign n31313 = pi18 ? n31310 : n31312;
  assign n31314 = pi17 ? n32 : n31313;
  assign n31315 = pi16 ? n32 : n31314;
  assign n31316 = pi19 ? n31190 : ~n501;
  assign n31317 = pi18 ? n31316 : n31312;
  assign n31318 = pi17 ? n32 : n31317;
  assign n31319 = pi16 ? n32 : n31318;
  assign n31320 = pi15 ? n31315 : n31319;
  assign n31321 = pi19 ? n28070 : ~n501;
  assign n31322 = pi20 ? n12884 : ~n339;
  assign n31323 = pi19 ? n31322 : n32;
  assign n31324 = pi18 ? n31321 : n31323;
  assign n31325 = pi17 ? n32 : n31324;
  assign n31326 = pi16 ? n32 : n31325;
  assign n31327 = pi19 ? n6398 : ~n19426;
  assign n31328 = pi20 ? n17665 : ~n339;
  assign n31329 = pi19 ? n31328 : n32;
  assign n31330 = pi18 ? n31327 : n31329;
  assign n31331 = pi17 ? n32 : n31330;
  assign n31332 = pi16 ? n32 : n31331;
  assign n31333 = pi15 ? n31326 : n31332;
  assign n31334 = pi14 ? n31320 : n31333;
  assign n31335 = pi13 ? n31308 : n31334;
  assign n31336 = pi15 ? n13375 : n13952;
  assign n31337 = pi15 ? n20301 : n32;
  assign n31338 = pi14 ? n31336 : n31337;
  assign n31339 = pi15 ? n30999 : n20531;
  assign n31340 = pi19 ? n18116 : n32;
  assign n31341 = pi18 ? n268 : n31340;
  assign n31342 = pi17 ? n32 : n31341;
  assign n31343 = pi16 ? n32 : n31342;
  assign n31344 = pi18 ? n268 : n13080;
  assign n31345 = pi17 ? n32 : n31344;
  assign n31346 = pi16 ? n32 : n31345;
  assign n31347 = pi15 ? n31343 : n31346;
  assign n31348 = pi14 ? n31339 : n31347;
  assign n31349 = pi13 ? n31338 : n31348;
  assign n31350 = pi12 ? n31335 : n31349;
  assign n31351 = pi11 ? n31307 : n31350;
  assign n31352 = pi16 ? n1233 : ~n31248;
  assign n31353 = pi15 ? n31247 : n31352;
  assign n31354 = pi14 ? n31244 : n31353;
  assign n31355 = pi13 ? n31354 : n31264;
  assign n31356 = pi12 ? n31236 : n31355;
  assign n31357 = pi15 ? n18535 : n29729;
  assign n31358 = pi14 ? n32 : n31357;
  assign n31359 = pi13 ? n32 : n31358;
  assign n31360 = pi18 ? n16847 : ~n814;
  assign n31361 = pi17 ? n32 : n31360;
  assign n31362 = pi16 ? n32 : n31361;
  assign n31363 = pi18 ? n268 : ~n814;
  assign n31364 = pi17 ? n32 : n31363;
  assign n31365 = pi16 ? n32 : n31364;
  assign n31366 = pi15 ? n31362 : n31365;
  assign n31367 = pi17 ? n16848 : n19262;
  assign n31368 = pi16 ? n32 : n31367;
  assign n31369 = pi15 ? n31368 : n19264;
  assign n31370 = pi14 ? n31366 : n31369;
  assign n31371 = pi18 ? n31286 : n237;
  assign n31372 = pi17 ? n3067 : ~n31371;
  assign n31373 = pi16 ? n32 : n31372;
  assign n31374 = pi15 ? n31373 : n31293;
  assign n31375 = pi14 ? n31285 : n31374;
  assign n31376 = pi13 ? n31370 : n31375;
  assign n31377 = pi12 ? n31359 : n31376;
  assign n31378 = pi11 ? n31356 : n31377;
  assign n31379 = pi10 ? n31351 : n31378;
  assign n31380 = pi09 ? n32 : n31379;
  assign n31381 = pi08 ? n31300 : n31380;
  assign n31382 = pi14 ? n487 : n22320;
  assign n31383 = pi13 ? n32 : n31382;
  assign n31384 = pi12 ? n31383 : n32;
  assign n31385 = pi19 ? n4406 : ~n32;
  assign n31386 = pi18 ? n31385 : ~n2424;
  assign n31387 = pi17 ? n32 : n31386;
  assign n31388 = pi16 ? n32 : n31387;
  assign n31389 = pi15 ? n20477 : n31388;
  assign n31390 = pi14 ? n20478 : n31389;
  assign n31391 = pi18 ? n532 : ~n2424;
  assign n31392 = pi17 ? n32 : n31391;
  assign n31393 = pi16 ? n32 : n31392;
  assign n31394 = pi15 ? n31393 : n21755;
  assign n31395 = pi20 ? n246 : ~n243;
  assign n31396 = pi19 ? n31395 : n32;
  assign n31397 = pi18 ? n30574 : n31396;
  assign n31398 = pi17 ? n32 : n31397;
  assign n31399 = pi16 ? n32 : n31398;
  assign n31400 = pi18 ? n20172 : n20474;
  assign n31401 = pi17 ? n32 : n31400;
  assign n31402 = pi16 ? n32 : n31401;
  assign n31403 = pi15 ? n31399 : n31402;
  assign n31404 = pi14 ? n31394 : n31403;
  assign n31405 = pi13 ? n31390 : n31404;
  assign n31406 = pi15 ? n21254 : n13952;
  assign n31407 = pi14 ? n31406 : n31120;
  assign n31408 = pi20 ? n8644 : n32;
  assign n31409 = pi19 ? n31408 : n32;
  assign n31410 = pi18 ? n4127 : n31409;
  assign n31411 = pi17 ? n32 : n31410;
  assign n31412 = pi16 ? n32 : n31411;
  assign n31413 = pi18 ? n32 : n31409;
  assign n31414 = pi17 ? n32 : n31413;
  assign n31415 = pi16 ? n32 : n31414;
  assign n31416 = pi15 ? n31412 : n31415;
  assign n31417 = pi15 ? n20862 : n32;
  assign n31418 = pi14 ? n31416 : n31417;
  assign n31419 = pi13 ? n31407 : n31418;
  assign n31420 = pi12 ? n31405 : n31419;
  assign n31421 = pi11 ? n31384 : n31420;
  assign n31422 = pi14 ? n30520 : n20447;
  assign n31423 = pi14 ? n19503 : n32;
  assign n31424 = pi13 ? n31422 : n31423;
  assign n31425 = pi18 ? n6596 : ~n32;
  assign n31426 = pi17 ? n2733 : ~n31425;
  assign n31427 = pi16 ? n32 : n31426;
  assign n31428 = pi18 ? n13940 : n702;
  assign n31429 = pi17 ? n31428 : ~n1697;
  assign n31430 = pi16 ? n32 : n31429;
  assign n31431 = pi15 ? n31427 : n31430;
  assign n31432 = pi18 ? n25760 : n32;
  assign n31433 = pi18 ? n880 : ~n248;
  assign n31434 = pi17 ? n31432 : n31433;
  assign n31435 = pi16 ? n1471 : ~n31434;
  assign n31436 = pi18 ? n28178 : n1548;
  assign n31437 = pi17 ? n32 : n31436;
  assign n31438 = pi16 ? n1135 : ~n31437;
  assign n31439 = pi15 ? n31435 : n31438;
  assign n31440 = pi14 ? n31431 : n31439;
  assign n31441 = pi18 ? n4380 : n350;
  assign n31442 = pi17 ? n32 : n31441;
  assign n31443 = pi16 ? n1135 : ~n31442;
  assign n31444 = pi18 ? n1249 : ~n32;
  assign n31445 = pi17 ? n32 : n31444;
  assign n31446 = pi16 ? n1471 : ~n31445;
  assign n31447 = pi15 ? n31443 : n31446;
  assign n31448 = pi17 ? n16848 : n4381;
  assign n31449 = pi16 ? n1135 : ~n31448;
  assign n31450 = pi15 ? n31449 : n31262;
  assign n31451 = pi14 ? n31447 : n31450;
  assign n31452 = pi13 ? n31440 : n31451;
  assign n31453 = pi12 ? n31424 : n31452;
  assign n31454 = pi16 ? n32 : n30892;
  assign n31455 = pi15 ? n32 : n31454;
  assign n31456 = pi15 ? n19531 : n29729;
  assign n31457 = pi14 ? n31455 : n31456;
  assign n31458 = pi13 ? n32 : n31457;
  assign n31459 = pi18 ? n16847 : ~n350;
  assign n31460 = pi17 ? n32 : n31459;
  assign n31461 = pi16 ? n32 : n31460;
  assign n31462 = pi18 ? n268 : ~n350;
  assign n31463 = pi17 ? n32 : n31462;
  assign n31464 = pi16 ? n32 : n31463;
  assign n31465 = pi15 ? n31461 : n31464;
  assign n31466 = pi17 ? n16848 : n18487;
  assign n31467 = pi16 ? n32 : n31466;
  assign n31468 = pi15 ? n31467 : n19172;
  assign n31469 = pi14 ? n31465 : n31468;
  assign n31470 = pi17 ? n17346 : n31363;
  assign n31471 = pi16 ? n32 : n31470;
  assign n31472 = pi18 ? n32 : n4722;
  assign n31473 = pi19 ? n9007 : n267;
  assign n31474 = pi18 ? n31473 : ~n814;
  assign n31475 = pi17 ? n31472 : n31474;
  assign n31476 = pi16 ? n32 : n31475;
  assign n31477 = pi15 ? n31471 : n31476;
  assign n31478 = pi19 ? n208 : n5371;
  assign n31479 = pi18 ? n31478 : n814;
  assign n31480 = pi17 ? n2726 : ~n31479;
  assign n31481 = pi16 ? n32 : n31480;
  assign n31482 = pi20 ? n5854 : n220;
  assign n31483 = pi20 ? n274 : ~n2385;
  assign n31484 = pi19 ? n31482 : n31483;
  assign n31485 = pi18 ? n940 : n31484;
  assign n31486 = pi17 ? n32 : n31485;
  assign n31487 = pi20 ? n915 : n246;
  assign n31488 = pi20 ? n207 : n518;
  assign n31489 = pi19 ? n31487 : n31488;
  assign n31490 = pi20 ? n321 : n501;
  assign n31491 = pi19 ? n31490 : ~n32;
  assign n31492 = pi18 ? n31489 : ~n31491;
  assign n31493 = pi17 ? n31492 : n2325;
  assign n31494 = pi16 ? n31486 : ~n31493;
  assign n31495 = pi15 ? n31481 : n31494;
  assign n31496 = pi14 ? n31477 : n31495;
  assign n31497 = pi13 ? n31469 : n31496;
  assign n31498 = pi12 ? n31458 : n31497;
  assign n31499 = pi11 ? n31453 : n31498;
  assign n31500 = pi10 ? n31421 : n31499;
  assign n31501 = pi09 ? n32 : n31500;
  assign n31502 = pi15 ? n21254 : n20477;
  assign n31503 = pi14 ? n31502 : n31120;
  assign n31504 = pi20 ? n8644 : ~n141;
  assign n31505 = pi19 ? n31504 : n32;
  assign n31506 = pi18 ? n4127 : n31505;
  assign n31507 = pi17 ? n32 : n31506;
  assign n31508 = pi16 ? n32 : n31507;
  assign n31509 = pi18 ? n32 : n31505;
  assign n31510 = pi17 ? n32 : n31509;
  assign n31511 = pi16 ? n32 : n31510;
  assign n31512 = pi15 ? n31508 : n31511;
  assign n31513 = pi18 ? n4722 : n20769;
  assign n31514 = pi17 ? n32 : n31513;
  assign n31515 = pi16 ? n32 : n31514;
  assign n31516 = pi15 ? n31515 : n32;
  assign n31517 = pi14 ? n31512 : n31516;
  assign n31518 = pi13 ? n31503 : n31517;
  assign n31519 = pi12 ? n31405 : n31518;
  assign n31520 = pi11 ? n32 : n31519;
  assign n31521 = pi18 ? n880 : ~n19237;
  assign n31522 = pi17 ? n31428 : ~n31521;
  assign n31523 = pi16 ? n32 : n31522;
  assign n31524 = pi15 ? n31427 : n31523;
  assign n31525 = pi14 ? n31524 : n31439;
  assign n31526 = pi16 ? n1233 : ~n31442;
  assign n31527 = pi15 ? n31526 : n31446;
  assign n31528 = pi18 ? n4380 : ~n113;
  assign n31529 = pi17 ? n16848 : n31528;
  assign n31530 = pi16 ? n1233 : ~n31529;
  assign n31531 = pi18 ? n31071 : ~n113;
  assign n31532 = pi17 ? n31260 : n31531;
  assign n31533 = pi16 ? n1471 : ~n31532;
  assign n31534 = pi15 ? n31530 : n31533;
  assign n31535 = pi14 ? n31527 : n31534;
  assign n31536 = pi13 ? n31525 : n31535;
  assign n31537 = pi12 ? n31424 : n31536;
  assign n31538 = pi18 ? n268 : n441;
  assign n31539 = pi17 ? n17346 : n31538;
  assign n31540 = pi16 ? n32 : n31539;
  assign n31541 = pi18 ? n31473 : n441;
  assign n31542 = pi17 ? n31472 : n31541;
  assign n31543 = pi16 ? n32 : n31542;
  assign n31544 = pi15 ? n31540 : n31543;
  assign n31545 = pi18 ? n31478 : ~n441;
  assign n31546 = pi17 ? n2726 : ~n31545;
  assign n31547 = pi16 ? n32 : n31546;
  assign n31548 = pi20 ? n820 : n2385;
  assign n31549 = pi19 ? n31482 : ~n31548;
  assign n31550 = pi18 ? n940 : n31549;
  assign n31551 = pi17 ? n32 : n31550;
  assign n31552 = pi20 ? n439 : n246;
  assign n31553 = pi20 ? n287 : n14286;
  assign n31554 = pi19 ? n31552 : n31553;
  assign n31555 = pi18 ? n31554 : ~n31491;
  assign n31556 = pi17 ? n31555 : n2325;
  assign n31557 = pi16 ? n31551 : ~n31556;
  assign n31558 = pi15 ? n31547 : n31557;
  assign n31559 = pi14 ? n31544 : n31558;
  assign n31560 = pi13 ? n31469 : n31559;
  assign n31561 = pi12 ? n31458 : n31560;
  assign n31562 = pi11 ? n31537 : n31561;
  assign n31563 = pi10 ? n31520 : n31562;
  assign n31564 = pi09 ? n32 : n31563;
  assign n31565 = pi08 ? n31501 : n31564;
  assign n31566 = pi07 ? n31381 : n31565;
  assign n31567 = pi06 ? n31172 : n31566;
  assign n31568 = pi14 ? n32 : n20831;
  assign n31569 = pi13 ? n32 : n31568;
  assign n31570 = pi14 ? n20831 : n20838;
  assign n31571 = pi15 ? n20660 : n21232;
  assign n31572 = pi14 ? n20661 : n31571;
  assign n31573 = pi13 ? n31570 : n31572;
  assign n31574 = pi12 ? n31569 : n31573;
  assign n31575 = pi18 ? n237 : ~n605;
  assign n31576 = pi17 ? n32 : n31575;
  assign n31577 = pi16 ? n32 : n31576;
  assign n31578 = pi15 ? n13948 : n31577;
  assign n31579 = pi18 ? n20788 : ~n605;
  assign n31580 = pi17 ? n32 : n31579;
  assign n31581 = pi16 ? n32 : n31580;
  assign n31582 = pi17 ? n32 : n21897;
  assign n31583 = pi16 ? n32 : n31582;
  assign n31584 = pi15 ? n31581 : n31583;
  assign n31585 = pi14 ? n31578 : n31584;
  assign n31586 = pi18 ? n520 : ~n605;
  assign n31587 = pi17 ? n32 : n31586;
  assign n31588 = pi16 ? n32 : n31587;
  assign n31589 = pi15 ? n31588 : n13948;
  assign n31590 = pi14 ? n31589 : n13948;
  assign n31591 = pi13 ? n31585 : n31590;
  assign n31592 = pi20 ? n8644 : ~n339;
  assign n31593 = pi19 ? n31592 : n32;
  assign n31594 = pi18 ? n4127 : n31593;
  assign n31595 = pi17 ? n32 : n31594;
  assign n31596 = pi16 ? n32 : n31595;
  assign n31597 = pi15 ? n19972 : n31596;
  assign n31598 = pi14 ? n21558 : n31597;
  assign n31599 = pi18 ? n11489 : ~n532;
  assign n31600 = pi17 ? n32 : n31599;
  assign n31601 = pi16 ? n32 : n31600;
  assign n31602 = pi15 ? n12098 : n31601;
  assign n31603 = pi14 ? n31602 : n32;
  assign n31604 = pi13 ? n31598 : n31603;
  assign n31605 = pi12 ? n31591 : n31604;
  assign n31606 = pi11 ? n31574 : n31605;
  assign n31607 = pi18 ? n32 : ~n23312;
  assign n31608 = pi17 ? n32 : n31607;
  assign n31609 = pi16 ? n32 : n31608;
  assign n31610 = pi15 ? n146 : n31609;
  assign n31611 = pi20 ? n3523 : ~n141;
  assign n31612 = pi19 ? n31611 : n32;
  assign n31613 = pi18 ? n4380 : n31612;
  assign n31614 = pi17 ? n32 : n31613;
  assign n31615 = pi16 ? n32 : n31614;
  assign n31616 = pi15 ? n31615 : n146;
  assign n31617 = pi14 ? n31610 : n31616;
  assign n31618 = pi17 ? n23052 : n32;
  assign n31619 = pi16 ? n32 : n31618;
  assign n31620 = pi15 ? n32 : n31619;
  assign n31621 = pi14 ? n146 : n31620;
  assign n31622 = pi13 ? n31617 : n31621;
  assign n31623 = pi19 ? n322 : n531;
  assign n31624 = pi18 ? n31623 : ~n32;
  assign n31625 = pi17 ? n2726 : ~n31624;
  assign n31626 = pi16 ? n32 : n31625;
  assign n31627 = pi19 ? n6057 : n4342;
  assign n31628 = pi19 ? n18478 : n32;
  assign n31629 = pi18 ? n31627 : ~n31628;
  assign n31630 = pi18 ? n4127 : n31385;
  assign n31631 = pi17 ? n31629 : ~n31630;
  assign n31632 = pi16 ? n23442 : n31631;
  assign n31633 = pi15 ? n31626 : n31632;
  assign n31634 = pi18 ? n11028 : ~n248;
  assign n31635 = pi17 ? n30107 : n31634;
  assign n31636 = pi16 ? n1214 : ~n31635;
  assign n31637 = pi18 ? n4380 : n344;
  assign n31638 = pi17 ? n32 : n31637;
  assign n31639 = pi16 ? n1214 : ~n31638;
  assign n31640 = pi15 ? n31636 : n31639;
  assign n31641 = pi14 ? n31633 : n31640;
  assign n31642 = pi16 ? n1214 : ~n31448;
  assign n31643 = pi19 ? n266 : ~n207;
  assign n31644 = pi18 ? n32 : n31643;
  assign n31645 = pi17 ? n32 : n31644;
  assign n31646 = pi19 ? n16002 : ~n246;
  assign n31647 = pi20 ? n266 : ~n246;
  assign n31648 = pi19 ? n18728 : n31647;
  assign n31649 = pi18 ? n31646 : ~n31648;
  assign n31650 = pi19 ? n29444 : n7642;
  assign n31651 = pi18 ? n31650 : n32;
  assign n31652 = pi17 ? n31649 : ~n31651;
  assign n31653 = pi16 ? n31645 : ~n31652;
  assign n31654 = pi15 ? n31642 : n31653;
  assign n31655 = pi19 ? n1464 : n208;
  assign n31656 = pi18 ? n31655 : ~n32;
  assign n31657 = pi17 ? n2726 : n31656;
  assign n31658 = pi16 ? n1214 : ~n31657;
  assign n31659 = pi18 ? n14982 : n32;
  assign n31660 = pi17 ? n880 : ~n31659;
  assign n31661 = pi16 ? n1471 : ~n31660;
  assign n31662 = pi15 ? n31658 : n31661;
  assign n31663 = pi14 ? n31654 : n31662;
  assign n31664 = pi13 ? n31641 : n31663;
  assign n31665 = pi12 ? n31622 : n31664;
  assign n31666 = pi15 ? n32 : n29862;
  assign n31667 = pi14 ? n32 : n31666;
  assign n31668 = pi20 ? n246 : n1324;
  assign n31669 = pi19 ? n31668 : n428;
  assign n31670 = pi18 ? n32 : n31669;
  assign n31671 = pi17 ? n32 : n31670;
  assign n31672 = pi20 ? n428 : n246;
  assign n31673 = pi19 ? n31672 : n30983;
  assign n31674 = pi20 ? n207 : n310;
  assign n31675 = pi20 ? n17669 : n206;
  assign n31676 = pi19 ? n31674 : ~n31675;
  assign n31677 = pi18 ? n31673 : ~n31676;
  assign n31678 = pi20 ? n206 : n6621;
  assign n31679 = pi19 ? n31678 : ~n7642;
  assign n31680 = pi18 ? n31679 : ~n350;
  assign n31681 = pi17 ? n31677 : n31680;
  assign n31682 = pi16 ? n31671 : n31681;
  assign n31683 = pi17 ? n269 : n1807;
  assign n31684 = pi16 ? n1214 : ~n31683;
  assign n31685 = pi15 ? n31682 : n31684;
  assign n31686 = pi16 ? n19652 : ~n3338;
  assign n31687 = pi16 ? n1683 : ~n1808;
  assign n31688 = pi15 ? n31686 : n31687;
  assign n31689 = pi14 ? n31685 : n31688;
  assign n31690 = pi13 ? n31667 : n31689;
  assign n31691 = pi18 ? n5335 : n323;
  assign n31692 = pi17 ? n31691 : ~n1807;
  assign n31693 = pi16 ? n32 : n31692;
  assign n31694 = pi17 ? n3067 : ~n3337;
  assign n31695 = pi16 ? n32 : n31694;
  assign n31696 = pi15 ? n31693 : n31695;
  assign n31697 = pi15 ? n29954 : n30199;
  assign n31698 = pi14 ? n31696 : n31697;
  assign n31699 = pi17 ? n2959 : n19265;
  assign n31700 = pi16 ? n32 : n31699;
  assign n31701 = pi18 ? n508 : n814;
  assign n31702 = pi17 ? n2959 : ~n31701;
  assign n31703 = pi16 ? n32 : n31702;
  assign n31704 = pi15 ? n31700 : n31703;
  assign n31705 = pi17 ? n2750 : ~n2136;
  assign n31706 = pi16 ? n32 : n31705;
  assign n31707 = pi16 ? n1135 : ~n2326;
  assign n31708 = pi15 ? n31706 : n31707;
  assign n31709 = pi14 ? n31704 : n31708;
  assign n31710 = pi13 ? n31698 : n31709;
  assign n31711 = pi12 ? n31690 : n31710;
  assign n31712 = pi11 ? n31665 : n31711;
  assign n31713 = pi10 ? n31606 : n31712;
  assign n31714 = pi09 ? n32 : n31713;
  assign n31715 = pi14 ? n20837 : n20836;
  assign n31716 = pi13 ? n32 : n31715;
  assign n31717 = pi15 ? n32 : n21232;
  assign n31718 = pi14 ? n32 : n31717;
  assign n31719 = pi13 ? n20970 : n31718;
  assign n31720 = pi12 ? n31716 : n31719;
  assign n31721 = pi15 ? n21232 : n31577;
  assign n31722 = pi14 ? n31721 : n31584;
  assign n31723 = pi20 ? n3523 : n333;
  assign n31724 = pi19 ? n519 : ~n31723;
  assign n31725 = pi20 ? n18129 : n207;
  assign n31726 = pi19 ? n31725 : ~n32;
  assign n31727 = pi18 ? n31724 : ~n31726;
  assign n31728 = pi17 ? n32 : n31727;
  assign n31729 = pi16 ? n32 : n31728;
  assign n31730 = pi15 ? n31729 : n13948;
  assign n31731 = pi14 ? n31730 : n13948;
  assign n31732 = pi13 ? n31722 : n31731;
  assign n31733 = pi12 ? n31732 : n31604;
  assign n31734 = pi11 ? n31720 : n31733;
  assign n31735 = pi15 ? n32 : n20072;
  assign n31736 = pi18 ? n4380 : n9170;
  assign n31737 = pi17 ? n32 : n31736;
  assign n31738 = pi16 ? n32 : n31737;
  assign n31739 = pi15 ? n31738 : n32;
  assign n31740 = pi14 ? n31735 : n31739;
  assign n31741 = pi14 ? n32 : n31620;
  assign n31742 = pi13 ? n31740 : n31741;
  assign n31743 = pi12 ? n31742 : n31664;
  assign n31744 = pi15 ? n31146 : n31687;
  assign n31745 = pi14 ? n31685 : n31744;
  assign n31746 = pi13 ? n31667 : n31745;
  assign n31747 = pi21 ? n242 : ~n140;
  assign n31748 = pi20 ? n31747 : n32;
  assign n31749 = pi19 ? n31748 : n32;
  assign n31750 = pi18 ? n32 : n31749;
  assign n31751 = pi17 ? n32 : n31750;
  assign n31752 = pi16 ? n32 : n31751;
  assign n31753 = pi15 ? n31752 : n30199;
  assign n31754 = pi14 ? n31696 : n31753;
  assign n31755 = pi13 ? n31754 : n31709;
  assign n31756 = pi12 ? n31746 : n31755;
  assign n31757 = pi11 ? n31743 : n31756;
  assign n31758 = pi10 ? n31734 : n31757;
  assign n31759 = pi09 ? n32 : n31758;
  assign n31760 = pi08 ? n31714 : n31759;
  assign n31761 = pi13 ? n32 : n20836;
  assign n31762 = pi14 ? n32 : n20844;
  assign n31763 = pi13 ? n20836 : n31762;
  assign n31764 = pi12 ? n31761 : n31763;
  assign n31765 = pi18 ? n31385 : ~n2413;
  assign n31766 = pi17 ? n9311 : n31765;
  assign n31767 = pi16 ? n32 : n31766;
  assign n31768 = pi18 ? n23073 : ~n2413;
  assign n31769 = pi17 ? n32 : n31768;
  assign n31770 = pi16 ? n32 : n31769;
  assign n31771 = pi15 ? n31767 : n31770;
  assign n31772 = pi18 ? n605 : ~n2413;
  assign n31773 = pi17 ? n32 : n31772;
  assign n31774 = pi16 ? n32 : n31773;
  assign n31775 = pi18 ? n520 : ~n2413;
  assign n31776 = pi17 ? n32 : n31775;
  assign n31777 = pi16 ? n32 : n31776;
  assign n31778 = pi15 ? n31774 : n31777;
  assign n31779 = pi14 ? n31771 : n31778;
  assign n31780 = pi15 ? n20756 : n21232;
  assign n31781 = pi14 ? n31780 : n21232;
  assign n31782 = pi13 ? n31779 : n31781;
  assign n31783 = pi15 ? n21232 : n13948;
  assign n31784 = pi20 ? n8644 : ~n207;
  assign n31785 = pi19 ? n31784 : n32;
  assign n31786 = pi18 ? n268 : n31785;
  assign n31787 = pi17 ? n32 : n31786;
  assign n31788 = pi16 ? n32 : n31787;
  assign n31789 = pi18 ? n684 : n20848;
  assign n31790 = pi17 ? n32 : n31789;
  assign n31791 = pi16 ? n32 : n31790;
  assign n31792 = pi15 ? n31788 : n31791;
  assign n31793 = pi14 ? n31783 : n31792;
  assign n31794 = pi18 ? n11028 : ~n418;
  assign n31795 = pi17 ? n32 : n31794;
  assign n31796 = pi16 ? n32 : n31795;
  assign n31797 = pi15 ? n12098 : n31796;
  assign n31798 = pi14 ? n31797 : n28396;
  assign n31799 = pi13 ? n31793 : n31798;
  assign n31800 = pi12 ? n31782 : n31799;
  assign n31801 = pi11 ? n31764 : n31800;
  assign n31802 = pi18 ? n17848 : n9170;
  assign n31803 = pi17 ? n32 : n31802;
  assign n31804 = pi16 ? n32 : n31803;
  assign n31805 = pi15 ? n31804 : n32;
  assign n31806 = pi14 ? n31735 : n31805;
  assign n31807 = pi17 ? n3164 : n32;
  assign n31808 = pi16 ? n32 : n31807;
  assign n31809 = pi15 ? n32 : n31808;
  assign n31810 = pi14 ? n32 : n31809;
  assign n31811 = pi13 ? n31806 : n31810;
  assign n31812 = pi18 ? n15116 : n880;
  assign n31813 = pi19 ? n507 : n21065;
  assign n31814 = pi18 ? n31813 : ~n19750;
  assign n31815 = pi17 ? n31812 : ~n31814;
  assign n31816 = pi16 ? n32 : n31815;
  assign n31817 = pi19 ? n321 : ~n321;
  assign n31818 = pi18 ? n32 : n31817;
  assign n31819 = pi17 ? n32 : n31818;
  assign n31820 = pi19 ? n18390 : ~n23114;
  assign n31821 = pi18 ? n31820 : n4343;
  assign n31822 = pi17 ? n31821 : n31630;
  assign n31823 = pi16 ? n31819 : ~n31822;
  assign n31824 = pi15 ? n31816 : n31823;
  assign n31825 = pi18 ? n863 : ~n19750;
  assign n31826 = pi17 ? n32 : n31825;
  assign n31827 = pi16 ? n19652 : ~n31826;
  assign n31828 = pi16 ? n1135 : ~n2530;
  assign n31829 = pi15 ? n31827 : n31828;
  assign n31830 = pi14 ? n31824 : n31829;
  assign n31831 = pi15 ? n31642 : n29676;
  assign n31832 = pi19 ? n322 : n208;
  assign n31833 = pi18 ? n31832 : ~n32;
  assign n31834 = pi17 ? n2726 : n31833;
  assign n31835 = pi16 ? n1214 : ~n31834;
  assign n31836 = pi15 ? n31835 : n31661;
  assign n31837 = pi14 ? n31831 : n31836;
  assign n31838 = pi13 ? n31830 : n31837;
  assign n31839 = pi12 ? n31811 : n31838;
  assign n31840 = pi18 ? n18474 : n863;
  assign n31841 = pi20 ? n259 : n5854;
  assign n31842 = pi20 ? n7839 : ~n2358;
  assign n31843 = pi19 ? n31841 : n31842;
  assign n31844 = pi18 ? n31843 : ~n350;
  assign n31845 = pi17 ? n31840 : n31844;
  assign n31846 = pi16 ? n32 : n31845;
  assign n31847 = pi15 ? n32 : n31846;
  assign n31848 = pi14 ? n32 : n31847;
  assign n31849 = pi19 ? n4342 : n14963;
  assign n31850 = pi19 ? n4670 : ~n236;
  assign n31851 = pi18 ? n31849 : n31850;
  assign n31852 = pi17 ? n31851 : n2537;
  assign n31853 = pi16 ? n31819 : ~n31852;
  assign n31854 = pi16 ? n1135 : ~n2540;
  assign n31855 = pi15 ? n31853 : n31854;
  assign n31856 = pi16 ? n1214 : ~n2540;
  assign n31857 = pi16 ? n1683 : ~n2540;
  assign n31858 = pi15 ? n31856 : n31857;
  assign n31859 = pi14 ? n31855 : n31858;
  assign n31860 = pi13 ? n31848 : n31859;
  assign n31861 = pi17 ? n31691 : ~n2537;
  assign n31862 = pi16 ? n32 : n31861;
  assign n31863 = pi17 ? n3067 : ~n2537;
  assign n31864 = pi16 ? n32 : n31863;
  assign n31865 = pi15 ? n31862 : n31864;
  assign n31866 = pi18 ? n6145 : n19811;
  assign n31867 = pi17 ? n32 : n31866;
  assign n31868 = pi16 ? n32 : n31867;
  assign n31869 = pi15 ? n31868 : n30199;
  assign n31870 = pi14 ? n31865 : n31869;
  assign n31871 = pi18 ? n6145 : ~n350;
  assign n31872 = pi17 ? n2954 : n31871;
  assign n31873 = pi16 ? n32 : n31872;
  assign n31874 = pi18 ? n702 : n814;
  assign n31875 = pi17 ? n2954 : ~n31874;
  assign n31876 = pi16 ? n32 : n31875;
  assign n31877 = pi15 ? n31873 : n31876;
  assign n31878 = pi20 ? n785 : n342;
  assign n31879 = pi19 ? n1248 : n31878;
  assign n31880 = pi19 ? n31483 : ~n32;
  assign n31881 = pi18 ? n31879 : n31880;
  assign n31882 = pi17 ? n31881 : ~n2325;
  assign n31883 = pi16 ? n22436 : n31882;
  assign n31884 = pi15 ? n31883 : n20034;
  assign n31885 = pi14 ? n31877 : n31884;
  assign n31886 = pi13 ? n31870 : n31885;
  assign n31887 = pi12 ? n31860 : n31886;
  assign n31888 = pi11 ? n31839 : n31887;
  assign n31889 = pi10 ? n31801 : n31888;
  assign n31890 = pi09 ? n32 : n31889;
  assign n31891 = pi15 ? n21033 : n14613;
  assign n31892 = pi14 ? n21034 : n31891;
  assign n31893 = pi13 ? n32 : n31892;
  assign n31894 = pi14 ? n14613 : n21326;
  assign n31895 = pi13 ? n31894 : n31762;
  assign n31896 = pi12 ? n31893 : n31895;
  assign n31897 = pi18 ? n31385 : ~n797;
  assign n31898 = pi17 ? n9311 : n31897;
  assign n31899 = pi16 ? n32 : n31898;
  assign n31900 = pi18 ? n23073 : ~n605;
  assign n31901 = pi17 ? n32 : n31900;
  assign n31902 = pi16 ? n32 : n31901;
  assign n31903 = pi15 ? n31899 : n31902;
  assign n31904 = pi14 ? n31903 : n31778;
  assign n31905 = pi13 ? n31904 : n31781;
  assign n31906 = pi14 ? n21232 : n31792;
  assign n31907 = pi18 ? n11028 : ~n2424;
  assign n31908 = pi17 ? n32 : n31907;
  assign n31909 = pi16 ? n32 : n31908;
  assign n31910 = pi15 ? n12098 : n31909;
  assign n31911 = pi14 ? n31910 : n28396;
  assign n31912 = pi13 ? n31906 : n31911;
  assign n31913 = pi12 ? n31905 : n31912;
  assign n31914 = pi11 ? n31896 : n31913;
  assign n31915 = pi16 ? n1214 : ~n31826;
  assign n31916 = pi15 ? n31915 : n31828;
  assign n31917 = pi14 ? n31824 : n31916;
  assign n31918 = pi18 ? n4380 : ~n19966;
  assign n31919 = pi17 ? n16848 : n31918;
  assign n31920 = pi16 ? n1214 : ~n31919;
  assign n31921 = pi15 ? n31920 : n29676;
  assign n31922 = pi18 ? n31832 : ~n19966;
  assign n31923 = pi17 ? n2726 : n31922;
  assign n31924 = pi16 ? n1214 : ~n31923;
  assign n31925 = pi15 ? n31924 : n31661;
  assign n31926 = pi14 ? n31921 : n31925;
  assign n31927 = pi13 ? n31917 : n31926;
  assign n31928 = pi12 ? n31811 : n31927;
  assign n31929 = pi18 ? n8106 : n1548;
  assign n31930 = pi17 ? n32 : n31929;
  assign n31931 = pi16 ? n1683 : ~n31930;
  assign n31932 = pi15 ? n31856 : n31931;
  assign n31933 = pi14 ? n31855 : n31932;
  assign n31934 = pi13 ? n31848 : n31933;
  assign n31935 = pi15 ? n31868 : n29954;
  assign n31936 = pi14 ? n31865 : n31935;
  assign n31937 = pi20 ? n175 : n1385;
  assign n31938 = pi19 ? n31937 : n357;
  assign n31939 = pi18 ? n32 : n31938;
  assign n31940 = pi17 ? n32 : n31939;
  assign n31941 = pi20 ? n357 : ~n266;
  assign n31942 = pi19 ? n31941 : n31878;
  assign n31943 = pi18 ? n31942 : n31880;
  assign n31944 = pi17 ? n31943 : ~n2325;
  assign n31945 = pi16 ? n31940 : n31944;
  assign n31946 = pi15 ? n31945 : n20034;
  assign n31947 = pi14 ? n31877 : n31946;
  assign n31948 = pi13 ? n31936 : n31947;
  assign n31949 = pi12 ? n31934 : n31948;
  assign n31950 = pi11 ? n31928 : n31949;
  assign n31951 = pi10 ? n31914 : n31950;
  assign n31952 = pi09 ? n32 : n31951;
  assign n31953 = pi08 ? n31890 : n31952;
  assign n31954 = pi07 ? n31760 : n31953;
  assign n31955 = pi13 ? n32 : n14613;
  assign n31956 = pi20 ? n342 : n785;
  assign n31957 = pi19 ? n507 : n31956;
  assign n31958 = pi18 ? n32 : n31957;
  assign n31959 = pi19 ? n9345 : ~n32;
  assign n31960 = pi18 ? n31959 : ~n2291;
  assign n31961 = pi17 ? n31958 : n31960;
  assign n31962 = pi16 ? n32 : n31961;
  assign n31963 = pi15 ? n20660 : n31962;
  assign n31964 = pi14 ? n20844 : n31963;
  assign n31965 = pi13 ? n31894 : n31964;
  assign n31966 = pi12 ? n31955 : n31965;
  assign n31967 = pi18 ? n323 : ~n797;
  assign n31968 = pi17 ? n32 : n31967;
  assign n31969 = pi16 ? n32 : n31968;
  assign n31970 = pi15 ? n31969 : n20836;
  assign n31971 = pi20 ? n310 : ~n274;
  assign n31972 = pi19 ? n31971 : ~n32;
  assign n31973 = pi18 ? n268 : ~n31972;
  assign n31974 = pi17 ? n32 : n31973;
  assign n31975 = pi16 ? n32 : n31974;
  assign n31976 = pi15 ? n31975 : n20836;
  assign n31977 = pi14 ? n31970 : n31976;
  assign n31978 = pi15 ? n20836 : n13943;
  assign n31979 = pi14 ? n20836 : n31978;
  assign n31980 = pi13 ? n31977 : n31979;
  assign n31981 = pi15 ? n12095 : n21153;
  assign n31982 = pi14 ? n13948 : n31981;
  assign n31983 = pi18 ? n1249 : ~n532;
  assign n31984 = pi17 ? n32 : n31983;
  assign n31985 = pi16 ? n32 : n31984;
  assign n31986 = pi18 ? n4380 : ~n21257;
  assign n31987 = pi17 ? n32 : n31986;
  assign n31988 = pi16 ? n32 : n31987;
  assign n31989 = pi15 ? n31985 : n31988;
  assign n31990 = pi18 ? n4380 : n4671;
  assign n31991 = pi17 ? n32 : n31990;
  assign n31992 = pi16 ? n32 : n31991;
  assign n31993 = pi15 ? n31992 : n20692;
  assign n31994 = pi14 ? n31989 : n31993;
  assign n31995 = pi13 ? n31982 : n31994;
  assign n31996 = pi12 ? n31980 : n31995;
  assign n31997 = pi11 ? n31966 : n31996;
  assign n31998 = pi18 ? n17848 : ~n532;
  assign n31999 = pi17 ? n32 : n31998;
  assign n32000 = pi16 ? n32 : n31999;
  assign n32001 = pi15 ? n20997 : n32000;
  assign n32002 = pi15 ? n13375 : n32;
  assign n32003 = pi14 ? n32001 : n32002;
  assign n32004 = pi17 ? n32 : ~n1028;
  assign n32005 = pi16 ? n32 : n32004;
  assign n32006 = pi15 ? n32 : n32005;
  assign n32007 = pi14 ? n32 : n32006;
  assign n32008 = pi13 ? n32003 : n32007;
  assign n32009 = pi18 ? n15831 : n863;
  assign n32010 = pi17 ? n32009 : ~n2410;
  assign n32011 = pi16 ? n32 : n32010;
  assign n32012 = pi19 ? n5694 : ~n7089;
  assign n32013 = pi18 ? n32 : n32012;
  assign n32014 = pi17 ? n32 : n32013;
  assign n32015 = pi19 ? n220 : ~n594;
  assign n32016 = pi19 ? n18502 : ~n1757;
  assign n32017 = pi18 ? n32015 : n32016;
  assign n32018 = pi17 ? n32017 : ~n20914;
  assign n32019 = pi16 ? n32014 : n32018;
  assign n32020 = pi15 ? n32011 : n32019;
  assign n32021 = pi16 ? n1135 : ~n1934;
  assign n32022 = pi16 ? n19652 : ~n1934;
  assign n32023 = pi15 ? n32021 : n32022;
  assign n32024 = pi14 ? n32020 : n32023;
  assign n32025 = pi19 ? n9007 : ~n236;
  assign n32026 = pi18 ? n863 : n32025;
  assign n32027 = pi17 ? n32 : n32026;
  assign n32028 = pi19 ? n6339 : n1757;
  assign n32029 = pi18 ? n4380 : n32028;
  assign n32030 = pi18 ? n24063 : n32;
  assign n32031 = pi17 ? n32029 : n32030;
  assign n32032 = pi16 ? n32027 : n32031;
  assign n32033 = pi18 ? n20172 : n350;
  assign n32034 = pi17 ? n32 : n32033;
  assign n32035 = pi16 ? n19652 : ~n32034;
  assign n32036 = pi15 ? n32032 : n32035;
  assign n32037 = pi18 ? n21270 : ~n32;
  assign n32038 = pi17 ? n32 : n32037;
  assign n32039 = pi16 ? n1214 : ~n32038;
  assign n32040 = pi18 ? n863 : ~n350;
  assign n32041 = pi18 ? n21274 : ~n32;
  assign n32042 = pi17 ? n32040 : n32041;
  assign n32043 = pi16 ? n1214 : ~n32042;
  assign n32044 = pi15 ? n32039 : n32043;
  assign n32045 = pi14 ? n32036 : n32044;
  assign n32046 = pi13 ? n32024 : n32045;
  assign n32047 = pi12 ? n32008 : n32046;
  assign n32048 = pi18 ? n5657 : n936;
  assign n32049 = pi17 ? n32048 : ~n2537;
  assign n32050 = pi16 ? n32 : n32049;
  assign n32051 = pi15 ? n32 : n32050;
  assign n32052 = pi14 ? n32 : n32051;
  assign n32053 = pi19 ? n5694 : ~n22525;
  assign n32054 = pi18 ? n32 : n32053;
  assign n32055 = pi17 ? n32 : n32054;
  assign n32056 = pi19 ? n246 : ~n247;
  assign n32057 = pi19 ? n18478 : ~n247;
  assign n32058 = pi18 ? n32056 : n32057;
  assign n32059 = pi17 ? n32058 : ~n2537;
  assign n32060 = pi16 ? n32055 : n32059;
  assign n32061 = pi19 ? n246 : n32;
  assign n32062 = pi18 ? n18710 : ~n32061;
  assign n32063 = pi17 ? n32 : n32062;
  assign n32064 = pi17 ? n19170 : n2537;
  assign n32065 = pi16 ? n32063 : ~n32064;
  assign n32066 = pi15 ? n32060 : n32065;
  assign n32067 = pi18 ? n13945 : n1548;
  assign n32068 = pi17 ? n19170 : n32067;
  assign n32069 = pi16 ? n32063 : ~n32068;
  assign n32070 = pi20 ? n18261 : ~n246;
  assign n32071 = pi19 ? n32070 : ~n32;
  assign n32072 = pi18 ? n32 : n32071;
  assign n32073 = pi17 ? n32 : n32072;
  assign n32074 = pi18 ? n13945 : ~n19933;
  assign n32075 = pi17 ? n18812 : n32074;
  assign n32076 = pi16 ? n32073 : ~n32075;
  assign n32077 = pi15 ? n32069 : n32076;
  assign n32078 = pi14 ? n32066 : n32077;
  assign n32079 = pi13 ? n32052 : n32078;
  assign n32080 = pi20 ? n12882 : n32;
  assign n32081 = pi19 ? n6057 : n32080;
  assign n32082 = pi20 ? n266 : n3523;
  assign n32083 = pi20 ? n785 : n246;
  assign n32084 = pi19 ? n32082 : ~n32083;
  assign n32085 = pi18 ? n32081 : n32084;
  assign n32086 = pi19 ? n5004 : ~n5371;
  assign n32087 = pi18 ? n32086 : n2318;
  assign n32088 = pi17 ? n32085 : ~n32087;
  assign n32089 = pi16 ? n23483 : n32088;
  assign n32090 = pi20 ? n220 : ~n207;
  assign n32091 = pi19 ? n1464 : n32090;
  assign n32092 = pi19 ? n18489 : ~n32090;
  assign n32093 = pi18 ? n32091 : n32092;
  assign n32094 = pi18 ? n14153 : n2318;
  assign n32095 = pi17 ? n32093 : ~n32094;
  assign n32096 = pi16 ? n32 : n32095;
  assign n32097 = pi15 ? n32089 : n32096;
  assign n32098 = pi18 ? n24942 : n684;
  assign n32099 = pi17 ? n32098 : ~n20567;
  assign n32100 = pi16 ? n32 : n32099;
  assign n32101 = pi19 ? n13069 : n6997;
  assign n32102 = pi18 ? n32101 : n1548;
  assign n32103 = pi17 ? n32 : ~n32102;
  assign n32104 = pi16 ? n32 : n32103;
  assign n32105 = pi15 ? n32100 : n32104;
  assign n32106 = pi14 ? n32097 : n32105;
  assign n32107 = pi18 ? n5657 : n880;
  assign n32108 = pi19 ? n9007 : n28957;
  assign n32109 = pi18 ? n32108 : ~n18532;
  assign n32110 = pi17 ? n32107 : ~n32109;
  assign n32111 = pi16 ? n32 : n32110;
  assign n32112 = pi19 ? n221 : ~n1757;
  assign n32113 = pi18 ? n20384 : n32112;
  assign n32114 = pi19 ? n32 : n29444;
  assign n32115 = pi18 ? n32114 : n237;
  assign n32116 = pi17 ? n32113 : ~n32115;
  assign n32117 = pi16 ? n32 : n32116;
  assign n32118 = pi15 ? n32111 : n32117;
  assign n32119 = pi14 ? n32118 : n20034;
  assign n32120 = pi13 ? n32106 : n32119;
  assign n32121 = pi12 ? n32079 : n32120;
  assign n32122 = pi11 ? n32047 : n32121;
  assign n32123 = pi10 ? n31997 : n32122;
  assign n32124 = pi09 ? n32 : n32123;
  assign n32125 = pi15 ? n14613 : n21319;
  assign n32126 = pi14 ? n32125 : n21319;
  assign n32127 = pi13 ? n32 : n32126;
  assign n32128 = pi15 ? n21319 : n32;
  assign n32129 = pi14 ? n21319 : n32128;
  assign n32130 = pi13 ? n32129 : n31964;
  assign n32131 = pi12 ? n32127 : n32130;
  assign n32132 = pi18 ? n323 : ~n2291;
  assign n32133 = pi17 ? n32 : n32132;
  assign n32134 = pi16 ? n32 : n32133;
  assign n32135 = pi15 ? n32134 : n20836;
  assign n32136 = pi14 ? n32135 : n31976;
  assign n32137 = pi13 ? n32136 : n31979;
  assign n32138 = pi14 ? n13948 : n12095;
  assign n32139 = pi18 ? n4380 : ~n22705;
  assign n32140 = pi17 ? n32 : n32139;
  assign n32141 = pi16 ? n32 : n32140;
  assign n32142 = pi15 ? n31985 : n32141;
  assign n32143 = pi14 ? n32142 : n31993;
  assign n32144 = pi13 ? n32138 : n32143;
  assign n32145 = pi12 ? n32137 : n32144;
  assign n32146 = pi11 ? n32131 : n32145;
  assign n32147 = pi17 ? n32009 : ~n2531;
  assign n32148 = pi16 ? n32 : n32147;
  assign n32149 = pi18 ? n32 : n20788;
  assign n32150 = pi17 ? n32017 : ~n32149;
  assign n32151 = pi16 ? n32014 : n32150;
  assign n32152 = pi15 ? n32148 : n32151;
  assign n32153 = pi16 ? n1214 : ~n1934;
  assign n32154 = pi15 ? n32021 : n32153;
  assign n32155 = pi14 ? n32152 : n32154;
  assign n32156 = pi16 ? n1214 : ~n32034;
  assign n32157 = pi15 ? n32032 : n32156;
  assign n32158 = pi14 ? n32157 : n32044;
  assign n32159 = pi13 ? n32155 : n32158;
  assign n32160 = pi12 ? n32008 : n32159;
  assign n32161 = pi17 ? n32048 : ~n1933;
  assign n32162 = pi16 ? n32 : n32161;
  assign n32163 = pi15 ? n32 : n32162;
  assign n32164 = pi14 ? n32 : n32163;
  assign n32165 = pi18 ? n127 : n32053;
  assign n32166 = pi17 ? n32 : n32165;
  assign n32167 = pi17 ? n32058 : ~n1933;
  assign n32168 = pi16 ? n32166 : n32167;
  assign n32169 = pi18 ? n29316 : ~n32061;
  assign n32170 = pi17 ? n32 : n32169;
  assign n32171 = pi17 ? n19170 : n2319;
  assign n32172 = pi16 ? n32170 : ~n32171;
  assign n32173 = pi15 ? n32168 : n32172;
  assign n32174 = pi18 ? n13945 : n2318;
  assign n32175 = pi17 ? n19170 : n32174;
  assign n32176 = pi16 ? n32063 : ~n32175;
  assign n32177 = pi15 ? n32176 : n32076;
  assign n32178 = pi14 ? n32173 : n32177;
  assign n32179 = pi13 ? n32164 : n32178;
  assign n32180 = pi18 ? n32101 : n3336;
  assign n32181 = pi17 ? n32 : ~n32180;
  assign n32182 = pi16 ? n32 : n32181;
  assign n32183 = pi15 ? n32100 : n32182;
  assign n32184 = pi14 ? n32097 : n32183;
  assign n32185 = pi16 ? n1233 : ~n2137;
  assign n32186 = pi14 ? n32118 : n32185;
  assign n32187 = pi13 ? n32184 : n32186;
  assign n32188 = pi12 ? n32179 : n32187;
  assign n32189 = pi11 ? n32160 : n32188;
  assign n32190 = pi10 ? n32146 : n32189;
  assign n32191 = pi09 ? n32 : n32190;
  assign n32192 = pi08 ? n32124 : n32191;
  assign n32193 = pi13 ? n32 : n21319;
  assign n32194 = pi19 ? n6398 : ~n32;
  assign n32195 = pi18 ? n32194 : ~n797;
  assign n32196 = pi17 ? n32 : n32195;
  assign n32197 = pi16 ? n32 : n32196;
  assign n32198 = pi15 ? n32197 : n11423;
  assign n32199 = pi14 ? n20844 : n32198;
  assign n32200 = pi13 ? n32129 : n32199;
  assign n32201 = pi12 ? n32193 : n32200;
  assign n32202 = pi19 ? n32 : ~n17669;
  assign n32203 = pi20 ? n266 : ~n7487;
  assign n32204 = pi19 ? n32203 : ~n32;
  assign n32205 = pi18 ? n32202 : ~n32204;
  assign n32206 = pi17 ? n32 : n32205;
  assign n32207 = pi16 ? n32 : n32206;
  assign n32208 = pi18 ? n496 : ~n2291;
  assign n32209 = pi17 ? n32 : n32208;
  assign n32210 = pi16 ? n32 : n32209;
  assign n32211 = pi15 ? n32207 : n32210;
  assign n32212 = pi15 ? n21033 : n14405;
  assign n32213 = pi14 ? n32211 : n32212;
  assign n32214 = pi15 ? n14405 : n21033;
  assign n32215 = pi14 ? n32214 : n21033;
  assign n32216 = pi13 ? n32213 : n32215;
  assign n32217 = pi18 ? n880 : ~n797;
  assign n32218 = pi17 ? n32 : n32217;
  assign n32219 = pi16 ? n32 : n32218;
  assign n32220 = pi15 ? n32219 : n12095;
  assign n32221 = pi14 ? n20836 : n32220;
  assign n32222 = pi15 ? n20695 : n20692;
  assign n32223 = pi15 ? n32 : n13369;
  assign n32224 = pi14 ? n32222 : n32223;
  assign n32225 = pi13 ? n32221 : n32224;
  assign n32226 = pi12 ? n32216 : n32225;
  assign n32227 = pi11 ? n32201 : n32226;
  assign n32228 = pi18 ? n1592 : ~n532;
  assign n32229 = pi17 ? n32 : n32228;
  assign n32230 = pi16 ? n32 : n32229;
  assign n32231 = pi15 ? n32230 : n12788;
  assign n32232 = pi15 ? n20692 : n32;
  assign n32233 = pi14 ? n32231 : n32232;
  assign n32234 = pi18 ? n23571 : n32;
  assign n32235 = pi17 ? n32 : n32234;
  assign n32236 = pi16 ? n32 : n32235;
  assign n32237 = pi18 ? n29140 : ~n237;
  assign n32238 = pi17 ? n32 : n32237;
  assign n32239 = pi16 ? n32 : n32238;
  assign n32240 = pi15 ? n32236 : n32239;
  assign n32241 = pi14 ? n32 : n32240;
  assign n32242 = pi13 ? n32233 : n32241;
  assign n32243 = pi19 ? n236 : ~n4670;
  assign n32244 = pi18 ? n32243 : ~n532;
  assign n32245 = pi17 ? n32 : n32244;
  assign n32246 = pi16 ? n32 : n32245;
  assign n32247 = pi19 ? n6057 : n19129;
  assign n32248 = pi18 ? n463 : n32247;
  assign n32249 = pi17 ? n32 : n32248;
  assign n32250 = pi19 ? n175 : n24755;
  assign n32251 = pi20 ? n785 : n207;
  assign n32252 = pi20 ? n501 : n18415;
  assign n32253 = pi19 ? n32251 : n32252;
  assign n32254 = pi18 ? n32250 : ~n32253;
  assign n32255 = pi19 ? n12801 : ~n32;
  assign n32256 = pi18 ? n32255 : ~n344;
  assign n32257 = pi17 ? n32254 : n32256;
  assign n32258 = pi16 ? n32249 : n32257;
  assign n32259 = pi15 ? n32246 : n32258;
  assign n32260 = pi14 ? n32259 : n32023;
  assign n32261 = pi20 ? n17665 : n1331;
  assign n32262 = pi20 ? n1331 : n17665;
  assign n32263 = pi19 ? n32261 : n32262;
  assign n32264 = pi18 ? n1395 : ~n32263;
  assign n32265 = pi17 ? n32 : n32264;
  assign n32266 = pi20 ? n18762 : n32;
  assign n32267 = pi19 ? n17665 : n32266;
  assign n32268 = pi19 ? n6398 : n20937;
  assign n32269 = pi18 ? n32267 : n32268;
  assign n32270 = pi20 ? n17665 : ~n357;
  assign n32271 = pi20 ? n6050 : ~n1331;
  assign n32272 = pi19 ? n32270 : ~n32271;
  assign n32273 = pi18 ? n32272 : n237;
  assign n32274 = pi17 ? n32269 : n32273;
  assign n32275 = pi16 ? n32265 : ~n32274;
  assign n32276 = pi15 ? n32275 : n32035;
  assign n32277 = pi16 ? n19652 : ~n32038;
  assign n32278 = pi17 ? n30197 : n32041;
  assign n32279 = pi16 ? n19652 : ~n32278;
  assign n32280 = pi15 ? n32277 : n32279;
  assign n32281 = pi14 ? n32276 : n32280;
  assign n32282 = pi13 ? n32260 : n32281;
  assign n32283 = pi12 ? n32242 : n32282;
  assign n32284 = pi17 ? n32 : n29220;
  assign n32285 = pi16 ? n32 : n32284;
  assign n32286 = pi15 ? n32 : n32285;
  assign n32287 = pi19 ? n17766 : n4342;
  assign n32288 = pi18 ? n32287 : n19750;
  assign n32289 = pi17 ? n32 : n32288;
  assign n32290 = pi16 ? n32 : n32289;
  assign n32291 = pi18 ? n237 : ~n344;
  assign n32292 = pi17 ? n32 : n32291;
  assign n32293 = pi16 ? n32 : n32292;
  assign n32294 = pi15 ? n32290 : n32293;
  assign n32295 = pi14 ? n32286 : n32294;
  assign n32296 = pi17 ? n20570 : n32291;
  assign n32297 = pi16 ? n32 : n32296;
  assign n32298 = pi15 ? n32293 : n32297;
  assign n32299 = pi18 ? n29226 : ~n344;
  assign n32300 = pi17 ? n32 : n32299;
  assign n32301 = pi16 ? n32 : n32300;
  assign n32302 = pi20 ? n342 : ~n206;
  assign n32303 = pi19 ? n23644 : ~n32302;
  assign n32304 = pi18 ? n32303 : n4689;
  assign n32305 = pi17 ? n32 : n32304;
  assign n32306 = pi16 ? n32 : n32305;
  assign n32307 = pi15 ? n32301 : n32306;
  assign n32308 = pi14 ? n32298 : n32307;
  assign n32309 = pi13 ? n32295 : n32308;
  assign n32310 = pi19 ? n21349 : n18478;
  assign n32311 = pi18 ? n32310 : ~n344;
  assign n32312 = pi17 ? n32 : n32311;
  assign n32313 = pi16 ? n32 : n32312;
  assign n32314 = pi20 ? n32 : ~n13171;
  assign n32315 = pi19 ? n32 : n32314;
  assign n32316 = pi18 ? n16449 : n32315;
  assign n32317 = pi19 ? n19191 : ~n32;
  assign n32318 = pi18 ? n32317 : ~n344;
  assign n32319 = pi17 ? n32316 : n32318;
  assign n32320 = pi16 ? n32 : n32319;
  assign n32321 = pi15 ? n32313 : n32320;
  assign n32322 = pi17 ? n2726 : ~n20561;
  assign n32323 = pi16 ? n32 : n32322;
  assign n32324 = pi19 ? n4964 : n5356;
  assign n32325 = pi18 ? n32324 : n350;
  assign n32326 = pi17 ? n32 : ~n32325;
  assign n32327 = pi16 ? n32 : n32326;
  assign n32328 = pi15 ? n32323 : n32327;
  assign n32329 = pi14 ? n32321 : n32328;
  assign n32330 = pi18 ? n16295 : n880;
  assign n32331 = pi20 ? n266 : ~n342;
  assign n32332 = pi19 ? n9007 : n32331;
  assign n32333 = pi18 ? n32332 : ~n6059;
  assign n32334 = pi17 ? n32330 : ~n32333;
  assign n32335 = pi16 ? n32 : n32334;
  assign n32336 = pi20 ? n287 : ~n1817;
  assign n32337 = pi19 ? n9007 : ~n32336;
  assign n32338 = pi18 ? n32 : n32337;
  assign n32339 = pi17 ? n32 : n32338;
  assign n32340 = pi20 ? n342 : n339;
  assign n32341 = pi19 ? n19596 : ~n32340;
  assign n32342 = pi19 ? n18200 : ~n1757;
  assign n32343 = pi18 ? n32341 : n32342;
  assign n32344 = pi20 ? n1331 : n3523;
  assign n32345 = pi19 ? n9007 : n32344;
  assign n32346 = pi18 ? n32345 : n30435;
  assign n32347 = pi17 ? n32343 : ~n32346;
  assign n32348 = pi16 ? n32339 : n32347;
  assign n32349 = pi15 ? n32335 : n32348;
  assign n32350 = pi14 ? n32349 : n20034;
  assign n32351 = pi13 ? n32329 : n32350;
  assign n32352 = pi12 ? n32309 : n32351;
  assign n32353 = pi11 ? n32283 : n32352;
  assign n32354 = pi10 ? n32227 : n32353;
  assign n32355 = pi09 ? n32 : n32354;
  assign n32356 = pi14 ? n21390 : n21464;
  assign n32357 = pi13 ? n32 : n32356;
  assign n32358 = pi19 ? n11145 : n32;
  assign n32359 = pi18 ? n32 : n32358;
  assign n32360 = pi17 ? n32 : n32359;
  assign n32361 = pi16 ? n32 : n32360;
  assign n32362 = pi15 ? n32 : n32361;
  assign n32363 = pi18 ? n32194 : ~n323;
  assign n32364 = pi17 ? n32 : n32363;
  assign n32365 = pi16 ? n32 : n32364;
  assign n32366 = pi15 ? n32365 : n11423;
  assign n32367 = pi14 ? n32362 : n32366;
  assign n32368 = pi13 ? n21468 : n32367;
  assign n32369 = pi12 ? n32357 : n32368;
  assign n32370 = pi19 ? n32 : ~n2358;
  assign n32371 = pi20 ? n310 : ~n266;
  assign n32372 = pi19 ? n32371 : ~n32;
  assign n32373 = pi18 ? n32370 : ~n32372;
  assign n32374 = pi17 ? n32 : n32373;
  assign n32375 = pi16 ? n32 : n32374;
  assign n32376 = pi15 ? n32375 : n11856;
  assign n32377 = pi14 ? n32376 : n31891;
  assign n32378 = pi13 ? n32377 : n21033;
  assign n32379 = pi15 ? n32219 : n12091;
  assign n32380 = pi14 ? n21035 : n32379;
  assign n32381 = pi19 ? n8235 : ~n32;
  assign n32382 = pi18 ? n940 : ~n32381;
  assign n32383 = pi17 ? n32 : n32382;
  assign n32384 = pi16 ? n32 : n32383;
  assign n32385 = pi15 ? n32384 : n20692;
  assign n32386 = pi14 ? n32385 : n32223;
  assign n32387 = pi13 ? n32380 : n32386;
  assign n32388 = pi12 ? n32378 : n32387;
  assign n32389 = pi11 ? n32369 : n32388;
  assign n32390 = pi19 ? n9816 : ~n32;
  assign n32391 = pi18 ? n29140 : ~n32390;
  assign n32392 = pi17 ? n32 : n32391;
  assign n32393 = pi16 ? n32 : n32392;
  assign n32394 = pi15 ? n32236 : n32393;
  assign n32395 = pi14 ? n32 : n32394;
  assign n32396 = pi13 ? n32233 : n32395;
  assign n32397 = pi18 ? n32243 : ~n3786;
  assign n32398 = pi17 ? n32 : n32397;
  assign n32399 = pi16 ? n32 : n32398;
  assign n32400 = pi19 ? n32251 : n502;
  assign n32401 = pi18 ? n24756 : ~n32400;
  assign n32402 = pi18 ? n31385 : ~n344;
  assign n32403 = pi17 ? n32401 : n32402;
  assign n32404 = pi16 ? n32 : n32403;
  assign n32405 = pi15 ? n32399 : n32404;
  assign n32406 = pi14 ? n32405 : n32154;
  assign n32407 = pi18 ? n209 : ~n32263;
  assign n32408 = pi17 ? n32 : n32407;
  assign n32409 = pi19 ? n32270 : ~n9197;
  assign n32410 = pi18 ? n32409 : n30906;
  assign n32411 = pi17 ? n32269 : n32410;
  assign n32412 = pi16 ? n32408 : ~n32411;
  assign n32413 = pi19 ? n7993 : ~n32;
  assign n32414 = pi18 ? n20172 : n32413;
  assign n32415 = pi17 ? n32 : n32414;
  assign n32416 = pi16 ? n1214 : ~n32415;
  assign n32417 = pi15 ? n32412 : n32416;
  assign n32418 = pi18 ? n21270 : ~n143;
  assign n32419 = pi17 ? n32 : n32418;
  assign n32420 = pi16 ? n1214 : ~n32419;
  assign n32421 = pi18 ? n21274 : ~n143;
  assign n32422 = pi17 ? n30197 : n32421;
  assign n32423 = pi16 ? n1214 : ~n32422;
  assign n32424 = pi15 ? n32420 : n32423;
  assign n32425 = pi14 ? n32417 : n32424;
  assign n32426 = pi13 ? n32406 : n32425;
  assign n32427 = pi12 ? n32396 : n32426;
  assign n32428 = pi18 ? n237 : ~n2304;
  assign n32429 = pi17 ? n32 : n32428;
  assign n32430 = pi16 ? n32 : n32429;
  assign n32431 = pi15 ? n32290 : n32430;
  assign n32432 = pi14 ? n32286 : n32431;
  assign n32433 = pi13 ? n32432 : n32308;
  assign n32434 = pi18 ? n16449 : n2387;
  assign n32435 = pi17 ? n32434 : n32318;
  assign n32436 = pi16 ? n32 : n32435;
  assign n32437 = pi15 ? n32313 : n32436;
  assign n32438 = pi14 ? n32437 : n32328;
  assign n32439 = pi18 ? n936 : n32337;
  assign n32440 = pi17 ? n32 : n32439;
  assign n32441 = pi20 ? n342 : n314;
  assign n32442 = pi19 ? n19596 : ~n32441;
  assign n32443 = pi20 ? n6621 : n10644;
  assign n32444 = pi19 ? n32443 : ~n1757;
  assign n32445 = pi18 ? n32442 : n32444;
  assign n32446 = pi17 ? n32445 : ~n32346;
  assign n32447 = pi16 ? n32440 : n32446;
  assign n32448 = pi15 ? n32335 : n32447;
  assign n32449 = pi14 ? n32448 : n20034;
  assign n32450 = pi13 ? n32438 : n32449;
  assign n32451 = pi12 ? n32433 : n32450;
  assign n32452 = pi11 ? n32427 : n32451;
  assign n32453 = pi10 ? n32389 : n32452;
  assign n32454 = pi09 ? n32 : n32453;
  assign n32455 = pi08 ? n32355 : n32454;
  assign n32456 = pi07 ? n32192 : n32455;
  assign n32457 = pi06 ? n31954 : n32456;
  assign n32458 = pi05 ? n31567 : n32457;
  assign n32459 = pi04 ? n30755 : n32458;
  assign n32460 = pi03 ? n29416 : n32459;
  assign n32461 = pi13 ? n32 : n21464;
  assign n32462 = pi15 ? n11650 : n12079;
  assign n32463 = pi14 ? n14156 : n32462;
  assign n32464 = pi13 ? n21468 : n32463;
  assign n32465 = pi12 ? n32461 : n32464;
  assign n32466 = pi18 ? n684 : ~n323;
  assign n32467 = pi17 ? n32 : n32466;
  assign n32468 = pi16 ? n32 : n32467;
  assign n32469 = pi15 ? n21319 : n32468;
  assign n32470 = pi14 ? n32469 : n21319;
  assign n32471 = pi14 ? n21322 : n14397;
  assign n32472 = pi13 ? n32470 : n32471;
  assign n32473 = pi20 ? n206 : ~n749;
  assign n32474 = pi19 ? n32473 : n32;
  assign n32475 = pi18 ? n863 : n32474;
  assign n32476 = pi17 ? n32 : n32475;
  assign n32477 = pi16 ? n32 : n32476;
  assign n32478 = pi19 ? n28179 : n32;
  assign n32479 = pi18 ? n863 : n32478;
  assign n32480 = pi17 ? n32 : n32479;
  assign n32481 = pi16 ? n32 : n32480;
  assign n32482 = pi15 ? n32477 : n32481;
  assign n32483 = pi14 ? n32 : n32482;
  assign n32484 = pi15 ? n19972 : n19172;
  assign n32485 = pi18 ? n6989 : ~n2413;
  assign n32486 = pi17 ? n29510 : n32485;
  assign n32487 = pi16 ? n32 : n32486;
  assign n32488 = pi15 ? n32 : n32487;
  assign n32489 = pi14 ? n32484 : n32488;
  assign n32490 = pi13 ? n32483 : n32489;
  assign n32491 = pi12 ? n32472 : n32490;
  assign n32492 = pi11 ? n32465 : n32491;
  assign n32493 = pi18 ? n344 : ~n32381;
  assign n32494 = pi17 ? n29510 : n32493;
  assign n32495 = pi16 ? n32 : n32494;
  assign n32496 = pi19 ? n12435 : ~n23193;
  assign n32497 = pi18 ? n32496 : ~n2413;
  assign n32498 = pi17 ? n28638 : n32497;
  assign n32499 = pi16 ? n32 : n32498;
  assign n32500 = pi15 ? n32495 : n32499;
  assign n32501 = pi14 ? n32500 : n20831;
  assign n32502 = pi14 ? n32 : n19862;
  assign n32503 = pi13 ? n32501 : n32502;
  assign n32504 = pi19 ? n1464 : ~n6307;
  assign n32505 = pi18 ? n32504 : n6059;
  assign n32506 = pi17 ? n32 : n32505;
  assign n32507 = pi16 ? n32 : n32506;
  assign n32508 = pi15 ? n32507 : n21268;
  assign n32509 = pi20 ? n206 : n310;
  assign n32510 = pi19 ? n5675 : ~n32509;
  assign n32511 = pi18 ? n32510 : n31385;
  assign n32512 = pi17 ? n32 : n32511;
  assign n32513 = pi16 ? n1135 : ~n32512;
  assign n32514 = pi15 ? n19805 : n32513;
  assign n32515 = pi14 ? n32508 : n32514;
  assign n32516 = pi18 ? n341 : ~n276;
  assign n32517 = pi17 ? n32 : n32516;
  assign n32518 = pi20 ? n274 : ~n354;
  assign n32519 = pi19 ? n274 : n32518;
  assign n32520 = pi19 ? n17665 : n18566;
  assign n32521 = pi18 ? n32519 : n32520;
  assign n32522 = pi20 ? n4279 : n207;
  assign n32523 = pi19 ? n32522 : ~n32;
  assign n32524 = pi18 ? n32523 : ~n32;
  assign n32525 = pi17 ? n32521 : n32524;
  assign n32526 = pi16 ? n32517 : ~n32525;
  assign n32527 = pi15 ? n32 : n32526;
  assign n32528 = pi16 ? n1135 : ~n3428;
  assign n32529 = pi17 ? n20529 : n1215;
  assign n32530 = pi16 ? n1214 : ~n32529;
  assign n32531 = pi15 ? n32528 : n32530;
  assign n32532 = pi14 ? n32527 : n32531;
  assign n32533 = pi13 ? n32515 : n32532;
  assign n32534 = pi12 ? n32503 : n32533;
  assign n32535 = pi19 ? n6988 : n32;
  assign n32536 = pi18 ? n32535 : n177;
  assign n32537 = pi17 ? n32 : n32536;
  assign n32538 = pi16 ? n32 : n32537;
  assign n32539 = pi15 ? n32 : n32538;
  assign n32540 = pi18 ? n15849 : ~n344;
  assign n32541 = pi17 ? n32 : n32540;
  assign n32542 = pi16 ? n32 : n32541;
  assign n32543 = pi15 ? n32 : n32542;
  assign n32544 = pi14 ? n32539 : n32543;
  assign n32545 = pi18 ? n6989 : ~n344;
  assign n32546 = pi17 ? n32 : n32545;
  assign n32547 = pi16 ? n32 : n32546;
  assign n32548 = pi19 ? n531 : ~n322;
  assign n32549 = pi18 ? n32548 : ~n344;
  assign n32550 = pi17 ? n32 : n32549;
  assign n32551 = pi16 ? n32 : n32550;
  assign n32552 = pi15 ? n32547 : n32551;
  assign n32553 = pi18 ? n15844 : ~n344;
  assign n32554 = pi17 ? n32 : n32553;
  assign n32555 = pi16 ? n32 : n32554;
  assign n32556 = pi15 ? n32555 : n19868;
  assign n32557 = pi14 ? n32552 : n32556;
  assign n32558 = pi13 ? n32544 : n32557;
  assign n32559 = pi18 ? n323 : ~n2304;
  assign n32560 = pi17 ? n32 : n32559;
  assign n32561 = pi16 ? n32 : n32560;
  assign n32562 = pi20 ? n3523 : n321;
  assign n32563 = pi19 ? n32562 : ~n32;
  assign n32564 = pi18 ? n32563 : ~n2304;
  assign n32565 = pi17 ? n32 : n32564;
  assign n32566 = pi16 ? n32 : n32565;
  assign n32567 = pi15 ? n32561 : n32566;
  assign n32568 = pi17 ? n32 : ~n1933;
  assign n32569 = pi16 ? n32 : n32568;
  assign n32570 = pi19 ? n321 : ~n531;
  assign n32571 = pi18 ? n32570 : ~n350;
  assign n32572 = pi17 ? n32 : n32571;
  assign n32573 = pi16 ? n32 : n32572;
  assign n32574 = pi15 ? n32569 : n32573;
  assign n32575 = pi14 ? n32567 : n32574;
  assign n32576 = pi19 ? n507 : ~n9321;
  assign n32577 = pi19 ? n18678 : ~n267;
  assign n32578 = pi18 ? n32576 : n32577;
  assign n32579 = pi18 ? n1509 : n1353;
  assign n32580 = pi17 ? n32578 : ~n32579;
  assign n32581 = pi16 ? n24246 : n32580;
  assign n32582 = pi18 ? n940 : ~n268;
  assign n32583 = pi17 ? n32 : n32582;
  assign n32584 = pi19 ? n23644 : n32;
  assign n32585 = pi18 ? n32 : n32584;
  assign n32586 = pi17 ? n32585 : n1807;
  assign n32587 = pi16 ? n32583 : ~n32586;
  assign n32588 = pi15 ? n32581 : n32587;
  assign n32589 = pi17 ? n19529 : n1807;
  assign n32590 = pi16 ? n19652 : ~n32589;
  assign n32591 = pi15 ? n32590 : n31056;
  assign n32592 = pi14 ? n32588 : n32591;
  assign n32593 = pi13 ? n32575 : n32592;
  assign n32594 = pi12 ? n32558 : n32593;
  assign n32595 = pi11 ? n32534 : n32594;
  assign n32596 = pi10 ? n32492 : n32595;
  assign n32597 = pi09 ? n32 : n32596;
  assign n32598 = pi15 ? n21464 : n387;
  assign n32599 = pi14 ? n32598 : n387;
  assign n32600 = pi13 ? n32 : n32599;
  assign n32601 = pi14 ? n387 : n388;
  assign n32602 = pi15 ? n11646 : n12079;
  assign n32603 = pi14 ? n14156 : n32602;
  assign n32604 = pi13 ? n32601 : n32603;
  assign n32605 = pi12 ? n32600 : n32604;
  assign n32606 = pi15 ? n21389 : n32468;
  assign n32607 = pi14 ? n32606 : n21319;
  assign n32608 = pi13 ? n32607 : n32471;
  assign n32609 = pi20 ? n206 : ~n1475;
  assign n32610 = pi19 ? n32609 : n32;
  assign n32611 = pi18 ? n863 : n32610;
  assign n32612 = pi17 ? n32 : n32611;
  assign n32613 = pi16 ? n32 : n32612;
  assign n32614 = pi15 ? n32613 : n32477;
  assign n32615 = pi14 ? n32 : n32614;
  assign n32616 = pi18 ? n6989 : ~n605;
  assign n32617 = pi17 ? n29510 : n32616;
  assign n32618 = pi16 ? n32 : n32617;
  assign n32619 = pi15 ? n32 : n32618;
  assign n32620 = pi14 ? n32484 : n32619;
  assign n32621 = pi13 ? n32615 : n32620;
  assign n32622 = pi12 ? n32608 : n32621;
  assign n32623 = pi11 ? n32605 : n32622;
  assign n32624 = pi18 ? n344 : ~n532;
  assign n32625 = pi17 ? n29510 : n32624;
  assign n32626 = pi16 ? n32 : n32625;
  assign n32627 = pi18 ? n32496 : ~n605;
  assign n32628 = pi17 ? n28638 : n32627;
  assign n32629 = pi16 ? n32 : n32628;
  assign n32630 = pi15 ? n32626 : n32629;
  assign n32631 = pi14 ? n32630 : n32;
  assign n32632 = pi13 ? n32631 : n32502;
  assign n32633 = pi20 ? n339 : n2358;
  assign n32634 = pi19 ? n32 : ~n32633;
  assign n32635 = pi18 ? n356 : ~n32634;
  assign n32636 = pi17 ? n32 : n32635;
  assign n32637 = pi20 ? n266 : ~n6050;
  assign n32638 = pi19 ? n266 : n32637;
  assign n32639 = pi20 ? n9641 : n246;
  assign n32640 = pi19 ? n17665 : n32639;
  assign n32641 = pi18 ? n32638 : n32640;
  assign n32642 = pi20 ? n12884 : ~n207;
  assign n32643 = pi19 ? n32642 : n32;
  assign n32644 = pi18 ? n32643 : n32;
  assign n32645 = pi17 ? n32641 : ~n32644;
  assign n32646 = pi16 ? n32636 : ~n32645;
  assign n32647 = pi15 ? n32 : n32646;
  assign n32648 = pi14 ? n32647 : n32531;
  assign n32649 = pi13 ? n32515 : n32648;
  assign n32650 = pi12 ? n32632 : n32649;
  assign n32651 = pi15 ? n32555 : n19805;
  assign n32652 = pi14 ? n32552 : n32651;
  assign n32653 = pi13 ? n32544 : n32652;
  assign n32654 = pi17 ? n32 : ~n2305;
  assign n32655 = pi16 ? n32 : n32654;
  assign n32656 = pi15 ? n32655 : n32573;
  assign n32657 = pi14 ? n32567 : n32656;
  assign n32658 = pi16 ? n1214 : ~n32589;
  assign n32659 = pi15 ? n32658 : n31146;
  assign n32660 = pi14 ? n32588 : n32659;
  assign n32661 = pi13 ? n32657 : n32660;
  assign n32662 = pi12 ? n32653 : n32661;
  assign n32663 = pi11 ? n32650 : n32662;
  assign n32664 = pi10 ? n32623 : n32663;
  assign n32665 = pi09 ? n32 : n32664;
  assign n32666 = pi08 ? n32597 : n32665;
  assign n32667 = pi14 ? n21858 : n21543;
  assign n32668 = pi13 ? n32 : n32667;
  assign n32669 = pi14 ? n21543 : n23466;
  assign n32670 = pi15 ? n12079 : n12289;
  assign n32671 = pi14 ? n14156 : n32670;
  assign n32672 = pi13 ? n32669 : n32671;
  assign n32673 = pi12 ? n32668 : n32672;
  assign n32674 = pi20 ? n310 : ~n7388;
  assign n32675 = pi19 ? n32674 : ~n32;
  assign n32676 = pi18 ? n268 : ~n32675;
  assign n32677 = pi17 ? n32 : n32676;
  assign n32678 = pi16 ? n32 : n32677;
  assign n32679 = pi15 ? n12083 : n32678;
  assign n32680 = pi14 ? n32679 : n21389;
  assign n32681 = pi14 ? n21389 : n22784;
  assign n32682 = pi13 ? n32680 : n32681;
  assign n32683 = pi18 ? n32 : n32535;
  assign n32684 = pi17 ? n32 : n32683;
  assign n32685 = pi16 ? n32 : n32684;
  assign n32686 = pi15 ? n32 : n32685;
  assign n32687 = pi15 ? n21346 : n13948;
  assign n32688 = pi14 ? n32686 : n32687;
  assign n32689 = pi19 ? n12899 : ~n32;
  assign n32690 = pi18 ? n32 : ~n32689;
  assign n32691 = pi17 ? n32 : n32690;
  assign n32692 = pi16 ? n32 : n32691;
  assign n32693 = pi15 ? n32 : n32692;
  assign n32694 = pi20 ? n518 : ~n749;
  assign n32695 = pi19 ? n32694 : n32;
  assign n32696 = pi18 ? n32 : n32695;
  assign n32697 = pi17 ? n32 : n32696;
  assign n32698 = pi16 ? n32 : n32697;
  assign n32699 = pi18 ? n6596 : ~n797;
  assign n32700 = pi17 ? n32 : n32699;
  assign n32701 = pi16 ? n32 : n32700;
  assign n32702 = pi15 ? n32698 : n32701;
  assign n32703 = pi14 ? n32693 : n32702;
  assign n32704 = pi13 ? n32688 : n32703;
  assign n32705 = pi12 ? n32682 : n32704;
  assign n32706 = pi11 ? n32673 : n32705;
  assign n32707 = pi18 ? n532 : ~n532;
  assign n32708 = pi17 ? n32 : n32707;
  assign n32709 = pi16 ? n32 : n32708;
  assign n32710 = pi18 ? n344 : ~n605;
  assign n32711 = pi17 ? n32 : n32710;
  assign n32712 = pi16 ? n32 : n32711;
  assign n32713 = pi15 ? n32709 : n32712;
  assign n32714 = pi19 ? n2386 : ~n236;
  assign n32715 = pi18 ? n32714 : ~n30435;
  assign n32716 = pi17 ? n32 : n32715;
  assign n32717 = pi16 ? n32 : n32716;
  assign n32718 = pi19 ? n1165 : n23180;
  assign n32719 = pi18 ? n32718 : ~n237;
  assign n32720 = pi17 ? n32 : n32719;
  assign n32721 = pi16 ? n32 : n32720;
  assign n32722 = pi15 ? n32717 : n32721;
  assign n32723 = pi14 ? n32713 : n32722;
  assign n32724 = pi14 ? n32 : n19972;
  assign n32725 = pi13 ? n32723 : n32724;
  assign n32726 = pi15 ? n20608 : n20692;
  assign n32727 = pi19 ? n8044 : n32;
  assign n32728 = pi18 ? n32 : n32727;
  assign n32729 = pi17 ? n32 : n32728;
  assign n32730 = pi16 ? n32 : n32729;
  assign n32731 = pi15 ? n32730 : n19805;
  assign n32732 = pi14 ? n32726 : n32731;
  assign n32733 = pi20 ? n207 : n342;
  assign n32734 = pi19 ? n32 : ~n32733;
  assign n32735 = pi18 ? n222 : ~n32734;
  assign n32736 = pi17 ? n32 : n32735;
  assign n32737 = pi19 ? n220 : n9345;
  assign n32738 = pi19 ? n32 : ~n5371;
  assign n32739 = pi18 ? n32737 : ~n32738;
  assign n32740 = pi17 ? n32739 : ~n32;
  assign n32741 = pi16 ? n32736 : ~n32740;
  assign n32742 = pi15 ? n32 : n32741;
  assign n32743 = pi18 ? n323 : ~n13949;
  assign n32744 = pi17 ? n32 : n32743;
  assign n32745 = pi16 ? n1135 : ~n32744;
  assign n32746 = pi17 ? n21344 : n1215;
  assign n32747 = pi16 ? n1214 : ~n32746;
  assign n32748 = pi15 ? n32745 : n32747;
  assign n32749 = pi14 ? n32742 : n32748;
  assign n32750 = pi13 ? n32732 : n32749;
  assign n32751 = pi12 ? n32725 : n32750;
  assign n32752 = pi18 ? n14153 : n32;
  assign n32753 = pi17 ? n32 : n32752;
  assign n32754 = pi16 ? n32 : n32753;
  assign n32755 = pi15 ? n32 : n32754;
  assign n32756 = pi18 ? n15849 : ~n430;
  assign n32757 = pi17 ? n32 : n32756;
  assign n32758 = pi16 ? n32 : n32757;
  assign n32759 = pi15 ? n180 : n32758;
  assign n32760 = pi14 ? n32755 : n32759;
  assign n32761 = pi18 ? n6596 : ~n430;
  assign n32762 = pi17 ? n32 : n32761;
  assign n32763 = pi16 ? n32 : n32762;
  assign n32764 = pi19 ? n5694 : n4964;
  assign n32765 = pi18 ? n32764 : ~n430;
  assign n32766 = pi17 ? n32 : n32765;
  assign n32767 = pi16 ? n32 : n32766;
  assign n32768 = pi15 ? n32763 : n32767;
  assign n32769 = pi18 ? n15844 : ~n430;
  assign n32770 = pi17 ? n32 : n32769;
  assign n32771 = pi16 ? n32 : n32770;
  assign n32772 = pi18 ? n16449 : n19750;
  assign n32773 = pi17 ? n32 : n32772;
  assign n32774 = pi16 ? n32 : n32773;
  assign n32775 = pi15 ? n32771 : n32774;
  assign n32776 = pi14 ? n32768 : n32775;
  assign n32777 = pi13 ? n32760 : n32776;
  assign n32778 = pi18 ? n323 : ~n430;
  assign n32779 = pi17 ? n32 : n32778;
  assign n32780 = pi16 ? n32 : n32779;
  assign n32781 = pi18 ? n323 : ~n344;
  assign n32782 = pi17 ? n32 : n32781;
  assign n32783 = pi16 ? n32 : n32782;
  assign n32784 = pi15 ? n32780 : n32783;
  assign n32785 = pi18 ? n268 : n16389;
  assign n32786 = pi17 ? n32785 : ~n1933;
  assign n32787 = pi16 ? n32 : n32786;
  assign n32788 = pi19 ? n22864 : ~n531;
  assign n32789 = pi18 ? n32788 : ~n350;
  assign n32790 = pi17 ? n269 : n32789;
  assign n32791 = pi16 ? n32 : n32790;
  assign n32792 = pi15 ? n32787 : n32791;
  assign n32793 = pi14 ? n32784 : n32792;
  assign n32794 = pi20 ? n321 : n2385;
  assign n32795 = pi19 ? n29705 : ~n32794;
  assign n32796 = pi18 ? n32 : n32795;
  assign n32797 = pi17 ? n32 : n32796;
  assign n32798 = pi19 ? n28686 : n32;
  assign n32799 = pi19 ? n11879 : n6057;
  assign n32800 = pi18 ? n32798 : n32799;
  assign n32801 = pi18 ? n463 : n350;
  assign n32802 = pi17 ? n32800 : n32801;
  assign n32803 = pi16 ? n32797 : ~n32802;
  assign n32804 = pi16 ? n1471 : ~n32589;
  assign n32805 = pi15 ? n32803 : n32804;
  assign n32806 = pi16 ? n1233 : ~n3338;
  assign n32807 = pi18 ? n21775 : ~n32;
  assign n32808 = pi17 ? n464 : n32807;
  assign n32809 = pi16 ? n1233 : ~n32808;
  assign n32810 = pi15 ? n32806 : n32809;
  assign n32811 = pi14 ? n32805 : n32810;
  assign n32812 = pi13 ? n32793 : n32811;
  assign n32813 = pi12 ? n32777 : n32812;
  assign n32814 = pi11 ? n32751 : n32813;
  assign n32815 = pi10 ? n32706 : n32814;
  assign n32816 = pi09 ? n32 : n32815;
  assign n32817 = pi15 ? n387 : n21786;
  assign n32818 = pi14 ? n32817 : n21786;
  assign n32819 = pi13 ? n21682 : n32818;
  assign n32820 = pi14 ? n21786 : n21790;
  assign n32821 = pi15 ? n14156 : n14152;
  assign n32822 = pi15 ? n12076 : n12289;
  assign n32823 = pi14 ? n32821 : n32822;
  assign n32824 = pi13 ? n32820 : n32823;
  assign n32825 = pi12 ? n32819 : n32824;
  assign n32826 = pi18 ? n880 : ~n323;
  assign n32827 = pi17 ? n32 : n32826;
  assign n32828 = pi16 ? n32 : n32827;
  assign n32829 = pi18 ? n268 : ~n32372;
  assign n32830 = pi17 ? n32 : n32829;
  assign n32831 = pi16 ? n32 : n32830;
  assign n32832 = pi15 ? n32828 : n32831;
  assign n32833 = pi14 ? n32832 : n21389;
  assign n32834 = pi16 ? n32 : n2106;
  assign n32835 = pi15 ? n21389 : n32834;
  assign n32836 = pi15 ? n32834 : n21389;
  assign n32837 = pi14 ? n32835 : n32836;
  assign n32838 = pi13 ? n32833 : n32837;
  assign n32839 = pi15 ? n21464 : n32685;
  assign n32840 = pi14 ? n32839 : n32687;
  assign n32841 = pi13 ? n32840 : n32703;
  assign n32842 = pi12 ? n32838 : n32841;
  assign n32843 = pi11 ? n32825 : n32842;
  assign n32844 = pi18 ? n5667 : ~n30435;
  assign n32845 = pi17 ? n32 : n32844;
  assign n32846 = pi16 ? n32 : n32845;
  assign n32847 = pi20 ? n32 : n9491;
  assign n32848 = pi20 ? n266 : n18129;
  assign n32849 = pi19 ? n32847 : n32848;
  assign n32850 = pi18 ? n32849 : ~n237;
  assign n32851 = pi17 ? n32 : n32850;
  assign n32852 = pi16 ? n32 : n32851;
  assign n32853 = pi15 ? n32846 : n32852;
  assign n32854 = pi14 ? n32713 : n32853;
  assign n32855 = pi13 ? n32854 : n32724;
  assign n32856 = pi20 ? n246 : n481;
  assign n32857 = pi19 ? n32856 : n32;
  assign n32858 = pi18 ? n32 : n32857;
  assign n32859 = pi17 ? n32 : n32858;
  assign n32860 = pi16 ? n32 : n32859;
  assign n32861 = pi15 ? n32730 : n32860;
  assign n32862 = pi14 ? n32726 : n32861;
  assign n32863 = pi16 ? n1233 : ~n32744;
  assign n32864 = pi15 ? n32863 : n32747;
  assign n32865 = pi14 ? n32742 : n32864;
  assign n32866 = pi13 ? n32862 : n32865;
  assign n32867 = pi12 ? n32855 : n32866;
  assign n32868 = pi16 ? n1135 : ~n32808;
  assign n32869 = pi15 ? n30941 : n32868;
  assign n32870 = pi14 ? n32805 : n32869;
  assign n32871 = pi13 ? n32793 : n32870;
  assign n32872 = pi12 ? n32777 : n32871;
  assign n32873 = pi11 ? n32867 : n32872;
  assign n32874 = pi10 ? n32843 : n32873;
  assign n32875 = pi09 ? n32 : n32874;
  assign n32876 = pi08 ? n32816 : n32875;
  assign n32877 = pi07 ? n32666 : n32876;
  assign n32878 = pi13 ? n21788 : n21786;
  assign n32879 = pi18 ? n1965 : ~n520;
  assign n32880 = pi17 ? n32 : n32879;
  assign n32881 = pi16 ? n32 : n32880;
  assign n32882 = pi15 ? n19172 : n32881;
  assign n32883 = pi18 ? n880 : ~n2747;
  assign n32884 = pi17 ? n32 : n32883;
  assign n32885 = pi16 ? n32 : n32884;
  assign n32886 = pi15 ? n32885 : n12518;
  assign n32887 = pi14 ? n32882 : n32886;
  assign n32888 = pi13 ? n32820 : n32887;
  assign n32889 = pi12 ? n32878 : n32888;
  assign n32890 = pi15 ? n12289 : n21543;
  assign n32891 = pi14 ? n32890 : n21543;
  assign n32892 = pi14 ? n21543 : n25126;
  assign n32893 = pi13 ? n32891 : n32892;
  assign n32894 = pi20 ? n206 : ~n1839;
  assign n32895 = pi19 ? n32894 : n32;
  assign n32896 = pi18 ? n863 : n32895;
  assign n32897 = pi17 ? n32 : n32896;
  assign n32898 = pi16 ? n32 : n32897;
  assign n32899 = pi15 ? n32898 : n14156;
  assign n32900 = pi14 ? n32899 : n21558;
  assign n32901 = pi18 ? n605 : ~n797;
  assign n32902 = pi17 ? n32 : n32901;
  assign n32903 = pi16 ? n32 : n32902;
  assign n32904 = pi15 ? n20836 : n32903;
  assign n32905 = pi14 ? n32 : n32904;
  assign n32906 = pi13 ? n32900 : n32905;
  assign n32907 = pi12 ? n32893 : n32906;
  assign n32908 = pi11 ? n32889 : n32907;
  assign n32909 = pi19 ? n322 : ~n5694;
  assign n32910 = pi18 ? n32909 : n5164;
  assign n32911 = pi17 ? n32 : n32910;
  assign n32912 = pi16 ? n32 : n32911;
  assign n32913 = pi20 ? n17665 : n18762;
  assign n32914 = pi19 ? n21412 : n32913;
  assign n32915 = pi18 ? n32914 : n32474;
  assign n32916 = pi17 ? n32 : n32915;
  assign n32917 = pi16 ? n32 : n32916;
  assign n32918 = pi15 ? n32912 : n32917;
  assign n32919 = pi19 ? n11972 : ~n32;
  assign n32920 = pi18 ? n605 : ~n32919;
  assign n32921 = pi17 ? n32 : n32920;
  assign n32922 = pi16 ? n32 : n32921;
  assign n32923 = pi15 ? n13948 : n32922;
  assign n32924 = pi14 ? n32918 : n32923;
  assign n32925 = pi13 ? n32924 : n32;
  assign n32926 = pi15 ? n32 : n19972;
  assign n32927 = pi14 ? n13671 : n32926;
  assign n32928 = pi19 ? n4342 : ~n32;
  assign n32929 = pi18 ? n940 : ~n32928;
  assign n32930 = pi17 ? n32929 : n1219;
  assign n32931 = pi16 ? n1471 : ~n32930;
  assign n32932 = pi18 ? n940 : n14153;
  assign n32933 = pi17 ? n32932 : n2355;
  assign n32934 = pi16 ? n1214 : ~n32933;
  assign n32935 = pi15 ? n32931 : n32934;
  assign n32936 = pi17 ? n14392 : n1480;
  assign n32937 = pi16 ? n1135 : ~n32936;
  assign n32938 = pi17 ? n14392 : n1215;
  assign n32939 = pi16 ? n1135 : ~n32938;
  assign n32940 = pi15 ? n32937 : n32939;
  assign n32941 = pi14 ? n32935 : n32940;
  assign n32942 = pi13 ? n32927 : n32941;
  assign n32943 = pi12 ? n32925 : n32942;
  assign n32944 = pi18 ? n16389 : n4492;
  assign n32945 = pi17 ? n32 : n32944;
  assign n32946 = pi16 ? n32 : n32945;
  assign n32947 = pi15 ? n20048 : n32946;
  assign n32948 = pi18 ? n15844 : n177;
  assign n32949 = pi17 ? n32 : n32948;
  assign n32950 = pi16 ? n32 : n32949;
  assign n32951 = pi15 ? n32950 : n32780;
  assign n32952 = pi14 ? n32947 : n32951;
  assign n32953 = pi19 ? n1464 : ~n176;
  assign n32954 = pi18 ? n32953 : ~n430;
  assign n32955 = pi17 ? n32 : n32954;
  assign n32956 = pi16 ? n32 : n32955;
  assign n32957 = pi18 ? n20193 : ~n430;
  assign n32958 = pi17 ? n32 : n32957;
  assign n32959 = pi16 ? n32 : n32958;
  assign n32960 = pi15 ? n32956 : n32959;
  assign n32961 = pi18 ? n29802 : n13086;
  assign n32962 = pi17 ? n32 : n32961;
  assign n32963 = pi16 ? n32 : n32962;
  assign n32964 = pi18 ? n24932 : n13086;
  assign n32965 = pi17 ? n32 : n32964;
  assign n32966 = pi16 ? n32 : n32965;
  assign n32967 = pi15 ? n32963 : n32966;
  assign n32968 = pi14 ? n32960 : n32967;
  assign n32969 = pi13 ? n32952 : n32968;
  assign n32970 = pi19 ? n29397 : n32;
  assign n32971 = pi18 ? n32970 : n2298;
  assign n32972 = pi17 ? n32 : ~n32971;
  assign n32973 = pi16 ? n17486 : n32972;
  assign n32974 = pi18 ? n30435 : ~n430;
  assign n32975 = pi17 ? n18017 : n32974;
  assign n32976 = pi16 ? n32 : n32975;
  assign n32977 = pi15 ? n32973 : n32976;
  assign n32978 = pi18 ? n350 : ~n430;
  assign n32979 = pi17 ? n18017 : n32978;
  assign n32980 = pi16 ? n32 : n32979;
  assign n32981 = pi19 ? n14463 : n6139;
  assign n32982 = pi18 ? n1249 : n32981;
  assign n32983 = pi18 ? n20182 : ~n248;
  assign n32984 = pi17 ? n32982 : ~n32983;
  assign n32985 = pi16 ? n26461 : n32984;
  assign n32986 = pi15 ? n32980 : n32985;
  assign n32987 = pi14 ? n32977 : n32986;
  assign n32988 = pi18 ? n209 : ~n5009;
  assign n32989 = pi17 ? n32 : n32988;
  assign n32990 = pi16 ? n32989 : ~n2540;
  assign n32991 = pi17 ? n32 : n5758;
  assign n32992 = pi16 ? n32991 : ~n2540;
  assign n32993 = pi15 ? n32990 : n32992;
  assign n32994 = pi18 ? n16432 : n350;
  assign n32995 = pi17 ? n32 : n32994;
  assign n32996 = pi16 ? n1135 : ~n32995;
  assign n32997 = pi18 ? n15844 : n350;
  assign n32998 = pi17 ? n32 : n32997;
  assign n32999 = pi16 ? n1135 : ~n32998;
  assign n33000 = pi15 ? n32996 : n32999;
  assign n33001 = pi14 ? n32993 : n33000;
  assign n33002 = pi13 ? n32987 : n33001;
  assign n33003 = pi12 ? n32969 : n33002;
  assign n33004 = pi11 ? n32943 : n33003;
  assign n33005 = pi10 ? n32908 : n33004;
  assign n33006 = pi09 ? n32 : n33005;
  assign n33007 = pi14 ? n21929 : n21928;
  assign n33008 = pi13 ? n21788 : n33007;
  assign n33009 = pi14 ? n21928 : n22133;
  assign n33010 = pi18 ? n1965 : ~n2747;
  assign n33011 = pi17 ? n32 : n33010;
  assign n33012 = pi16 ? n32 : n33011;
  assign n33013 = pi15 ? n19172 : n33012;
  assign n33014 = pi14 ? n33013 : n32886;
  assign n33015 = pi13 ? n33009 : n33014;
  assign n33016 = pi12 ? n33008 : n33015;
  assign n33017 = pi19 ? n21282 : n32;
  assign n33018 = pi18 ? n863 : n33017;
  assign n33019 = pi17 ? n32 : n33018;
  assign n33020 = pi16 ? n32 : n33019;
  assign n33021 = pi15 ? n33020 : n14156;
  assign n33022 = pi14 ? n33021 : n21558;
  assign n33023 = pi13 ? n33022 : n32905;
  assign n33024 = pi12 ? n32893 : n33023;
  assign n33025 = pi11 ? n33016 : n33024;
  assign n33026 = pi19 ? n857 : n357;
  assign n33027 = pi20 ? n2385 : ~n749;
  assign n33028 = pi19 ? n33027 : n32;
  assign n33029 = pi18 ? n33026 : n33028;
  assign n33030 = pi17 ? n32 : n33029;
  assign n33031 = pi16 ? n32 : n33030;
  assign n33032 = pi15 ? n32912 : n33031;
  assign n33033 = pi15 ? n13948 : n31583;
  assign n33034 = pi14 ? n33032 : n33033;
  assign n33035 = pi13 ? n33034 : n32;
  assign n33036 = pi14 ? n21346 : n32926;
  assign n33037 = pi13 ? n33036 : n32941;
  assign n33038 = pi12 ? n33035 : n33037;
  assign n33039 = pi15 ? n20301 : n32946;
  assign n33040 = pi18 ? n323 : ~n2298;
  assign n33041 = pi17 ? n32 : n33040;
  assign n33042 = pi16 ? n32 : n33041;
  assign n33043 = pi15 ? n32950 : n33042;
  assign n33044 = pi14 ? n33039 : n33043;
  assign n33045 = pi18 ? n32953 : ~n2298;
  assign n33046 = pi17 ? n32 : n33045;
  assign n33047 = pi16 ? n32 : n33046;
  assign n33048 = pi18 ? n20193 : ~n2298;
  assign n33049 = pi17 ? n32 : n33048;
  assign n33050 = pi16 ? n32 : n33049;
  assign n33051 = pi15 ? n33047 : n33050;
  assign n33052 = pi14 ? n33051 : n32967;
  assign n33053 = pi13 ? n33044 : n33052;
  assign n33054 = pi19 ? n29002 : n275;
  assign n33055 = pi18 ? n858 : n33054;
  assign n33056 = pi17 ? n33055 : ~n32971;
  assign n33057 = pi16 ? n17486 : n33056;
  assign n33058 = pi18 ? n30435 : ~n2298;
  assign n33059 = pi17 ? n18017 : n33058;
  assign n33060 = pi16 ? n32 : n33059;
  assign n33061 = pi15 ? n33057 : n33060;
  assign n33062 = pi18 ? n350 : ~n2298;
  assign n33063 = pi17 ? n18017 : n33062;
  assign n33064 = pi16 ? n32 : n33063;
  assign n33065 = pi15 ? n33064 : n32985;
  assign n33066 = pi14 ? n33061 : n33065;
  assign n33067 = pi16 ? n32989 : ~n1934;
  assign n33068 = pi16 ? n32991 : ~n2320;
  assign n33069 = pi15 ? n33067 : n33068;
  assign n33070 = pi16 ? n1233 : ~n32995;
  assign n33071 = pi16 ? n1233 : ~n32998;
  assign n33072 = pi15 ? n33070 : n33071;
  assign n33073 = pi14 ? n33069 : n33072;
  assign n33074 = pi13 ? n33066 : n33073;
  assign n33075 = pi12 ? n33053 : n33074;
  assign n33076 = pi11 ? n33038 : n33075;
  assign n33077 = pi10 ? n33025 : n33076;
  assign n33078 = pi09 ? n32 : n33077;
  assign n33079 = pi08 ? n33006 : n33078;
  assign n33080 = pi13 ? n21930 : n476;
  assign n33081 = pi15 ? n19172 : n12283;
  assign n33082 = pi14 ? n33081 : n12515;
  assign n33083 = pi13 ? n476 : n33082;
  assign n33084 = pi12 ? n33080 : n33083;
  assign n33085 = pi15 ? n12518 : n21686;
  assign n33086 = pi14 ? n33085 : n21686;
  assign n33087 = pi13 ? n33086 : n21686;
  assign n33088 = pi15 ? n13920 : n14394;
  assign n33089 = pi14 ? n33088 : n32;
  assign n33090 = pi15 ? n22087 : n11202;
  assign n33091 = pi14 ? n14397 : n33090;
  assign n33092 = pi13 ? n33089 : n33091;
  assign n33093 = pi12 ? n33087 : n33092;
  assign n33094 = pi11 ? n33084 : n33093;
  assign n33095 = pi18 ? n32909 : n4343;
  assign n33096 = pi17 ? n32 : n33095;
  assign n33097 = pi16 ? n32 : n33096;
  assign n33098 = pi15 ? n33097 : n32;
  assign n33099 = pi18 ? n323 : ~n605;
  assign n33100 = pi17 ? n32 : n33099;
  assign n33101 = pi16 ? n32 : n33100;
  assign n33102 = pi15 ? n32 : n33101;
  assign n33103 = pi14 ? n33098 : n33102;
  assign n33104 = pi13 ? n33103 : n31762;
  assign n33105 = pi18 ? n32 : n23401;
  assign n33106 = pi17 ? n32 : n33105;
  assign n33107 = pi16 ? n32 : n33106;
  assign n33108 = pi15 ? n19972 : n33107;
  assign n33109 = pi15 ? n13948 : n20692;
  assign n33110 = pi14 ? n33108 : n33109;
  assign n33111 = pi16 ? n1135 : ~n4064;
  assign n33112 = pi15 ? n32931 : n33111;
  assign n33113 = pi17 ? n22823 : n1480;
  assign n33114 = pi16 ? n1214 : ~n33113;
  assign n33115 = pi19 ? n322 : ~n4982;
  assign n33116 = pi18 ? n33115 : ~n13668;
  assign n33117 = pi17 ? n22823 : n33116;
  assign n33118 = pi16 ? n1214 : ~n33117;
  assign n33119 = pi15 ? n33114 : n33118;
  assign n33120 = pi14 ? n33112 : n33119;
  assign n33121 = pi13 ? n33110 : n33120;
  assign n33122 = pi12 ? n33104 : n33121;
  assign n33123 = pi19 ? n32 : n28134;
  assign n33124 = pi18 ? n33123 : ~n31959;
  assign n33125 = pi17 ? n32 : n33124;
  assign n33126 = pi16 ? n32 : n33125;
  assign n33127 = pi15 ? n13671 : n33126;
  assign n33128 = pi18 ? n323 : ~n532;
  assign n33129 = pi17 ? n32 : n33128;
  assign n33130 = pi16 ? n32 : n33129;
  assign n33131 = pi15 ? n22097 : n33130;
  assign n33132 = pi14 ? n33127 : n33131;
  assign n33133 = pi18 ? n702 : ~n532;
  assign n33134 = pi17 ? n32 : n33133;
  assign n33135 = pi16 ? n32 : n33134;
  assign n33136 = pi18 ? n20193 : ~n532;
  assign n33137 = pi17 ? n32 : n33136;
  assign n33138 = pi16 ? n32 : n33137;
  assign n33139 = pi15 ? n33135 : n33138;
  assign n33140 = pi18 ? n29802 : n13080;
  assign n33141 = pi17 ? n32 : n33140;
  assign n33142 = pi16 ? n32 : n33141;
  assign n33143 = pi15 ? n33142 : n33135;
  assign n33144 = pi14 ? n33139 : n33143;
  assign n33145 = pi13 ? n33132 : n33144;
  assign n33146 = pi19 ? n4342 : n7089;
  assign n33147 = pi18 ? n18710 : n33146;
  assign n33148 = pi17 ? n32 : n33147;
  assign n33149 = pi19 ? n7089 : ~n220;
  assign n33150 = pi20 ? n260 : n321;
  assign n33151 = pi19 ? n9037 : ~n33150;
  assign n33152 = pi18 ? n33149 : n33151;
  assign n33153 = pi18 ? n6059 : n344;
  assign n33154 = pi17 ? n33152 : n33153;
  assign n33155 = pi16 ? n33148 : ~n33154;
  assign n33156 = pi18 ? n350 : ~n344;
  assign n33157 = pi17 ? n19170 : n33156;
  assign n33158 = pi16 ? n32 : n33157;
  assign n33159 = pi15 ? n33155 : n33158;
  assign n33160 = pi18 ? n463 : n940;
  assign n33161 = pi17 ? n32 : n33160;
  assign n33162 = pi19 ? n23895 : n5004;
  assign n33163 = pi18 ? n11884 : n33162;
  assign n33164 = pi18 ? n22107 : n31385;
  assign n33165 = pi17 ? n33163 : n33164;
  assign n33166 = pi16 ? n33161 : ~n33165;
  assign n33167 = pi15 ? n33158 : n33166;
  assign n33168 = pi14 ? n33159 : n33167;
  assign n33169 = pi18 ? n341 : ~n14153;
  assign n33170 = pi17 ? n32 : n33169;
  assign n33171 = pi16 ? n33170 : ~n1934;
  assign n33172 = pi18 ? n18710 : ~n5009;
  assign n33173 = pi17 ? n32 : n33172;
  assign n33174 = pi16 ? n33173 : ~n2540;
  assign n33175 = pi15 ? n33171 : n33174;
  assign n33176 = pi14 ? n33175 : n32999;
  assign n33177 = pi13 ? n33168 : n33176;
  assign n33178 = pi12 ? n33145 : n33177;
  assign n33179 = pi11 ? n33122 : n33178;
  assign n33180 = pi10 ? n33094 : n33179;
  assign n33181 = pi09 ? n32 : n33180;
  assign n33182 = pi13 ? n32 : n648;
  assign n33183 = pi13 ? n648 : n33082;
  assign n33184 = pi12 ? n33182 : n33183;
  assign n33185 = pi15 ? n14397 : n11202;
  assign n33186 = pi14 ? n14397 : n33185;
  assign n33187 = pi13 ? n33089 : n33186;
  assign n33188 = pi12 ? n33087 : n33187;
  assign n33189 = pi11 ? n33184 : n33188;
  assign n33190 = pi14 ? n20832 : n22976;
  assign n33191 = pi13 ? n33103 : n33190;
  assign n33192 = pi20 ? n321 : n52;
  assign n33193 = pi19 ? n33192 : n32;
  assign n33194 = pi18 ? n32 : n33193;
  assign n33195 = pi17 ? n32 : n33194;
  assign n33196 = pi16 ? n32 : n33195;
  assign n33197 = pi15 ? n21232 : n33196;
  assign n33198 = pi14 ? n33108 : n33197;
  assign n33199 = pi18 ? n532 : ~n20828;
  assign n33200 = pi17 ? n32929 : n33199;
  assign n33201 = pi16 ? n1471 : ~n33200;
  assign n33202 = pi18 ? n702 : ~n20828;
  assign n33203 = pi17 ? n32 : n33202;
  assign n33204 = pi16 ? n1233 : ~n33203;
  assign n33205 = pi15 ? n33201 : n33204;
  assign n33206 = pi17 ? n22823 : n33202;
  assign n33207 = pi16 ? n19652 : ~n33206;
  assign n33208 = pi18 ? n33115 : ~n21487;
  assign n33209 = pi17 ? n22823 : n33208;
  assign n33210 = pi16 ? n1214 : ~n33209;
  assign n33211 = pi15 ? n33207 : n33210;
  assign n33212 = pi14 ? n33205 : n33211;
  assign n33213 = pi13 ? n33198 : n33212;
  assign n33214 = pi12 ? n33191 : n33213;
  assign n33215 = pi20 ? n220 : n339;
  assign n33216 = pi19 ? n33215 : ~n32;
  assign n33217 = pi18 ? n33123 : ~n33216;
  assign n33218 = pi17 ? n32 : n33217;
  assign n33219 = pi16 ? n32 : n33218;
  assign n33220 = pi15 ? n13671 : n33219;
  assign n33221 = pi14 ? n33220 : n33131;
  assign n33222 = pi13 ? n33221 : n33144;
  assign n33223 = pi14 ? n33175 : n33071;
  assign n33224 = pi13 ? n33168 : n33223;
  assign n33225 = pi12 ? n33222 : n33224;
  assign n33226 = pi11 ? n33214 : n33225;
  assign n33227 = pi10 ? n33189 : n33226;
  assign n33228 = pi09 ? n32 : n33227;
  assign n33229 = pi08 ? n33181 : n33228;
  assign n33230 = pi07 ? n33079 : n33229;
  assign n33231 = pi06 ? n32877 : n33230;
  assign n33232 = pi20 ? n207 : ~n111;
  assign n33233 = pi19 ? n33232 : ~n32;
  assign n33234 = pi18 ? n32 : ~n33233;
  assign n33235 = pi17 ? n32 : n33234;
  assign n33236 = pi16 ? n32 : n33235;
  assign n33237 = pi15 ? n648 : n33236;
  assign n33238 = pi14 ? n648 : n33237;
  assign n33239 = pi19 ? n18502 : ~n32;
  assign n33240 = pi18 ? n32 : ~n33239;
  assign n33241 = pi17 ? n32 : n33240;
  assign n33242 = pi16 ? n32 : n33241;
  assign n33243 = pi15 ? n33242 : n12515;
  assign n33244 = pi18 ? n863 : n13335;
  assign n33245 = pi17 ? n32 : n33244;
  assign n33246 = pi16 ? n32 : n33245;
  assign n33247 = pi15 ? n12764 : n33246;
  assign n33248 = pi14 ? n33243 : n33247;
  assign n33249 = pi13 ? n33238 : n33248;
  assign n33250 = pi12 ? n33182 : n33249;
  assign n33251 = pi18 ? n863 : n8908;
  assign n33252 = pi17 ? n32 : n33251;
  assign n33253 = pi16 ? n32 : n33252;
  assign n33254 = pi15 ? n33253 : n21853;
  assign n33255 = pi14 ? n33254 : n21853;
  assign n33256 = pi15 ? n21853 : n21928;
  assign n33257 = pi14 ? n33256 : n22638;
  assign n33258 = pi13 ? n33255 : n33257;
  assign n33259 = pi15 ? n14397 : n21319;
  assign n33260 = pi14 ? n14394 : n33259;
  assign n33261 = pi18 ? n15844 : n21386;
  assign n33262 = pi17 ? n32 : n33261;
  assign n33263 = pi16 ? n32 : n33262;
  assign n33264 = pi18 ? n20359 : ~n2754;
  assign n33265 = pi17 ? n32 : n33264;
  assign n33266 = pi16 ? n32 : n33265;
  assign n33267 = pi15 ? n33263 : n33266;
  assign n33268 = pi14 ? n21319 : n33267;
  assign n33269 = pi13 ? n33260 : n33268;
  assign n33270 = pi12 ? n33258 : n33269;
  assign n33271 = pi11 ? n33250 : n33270;
  assign n33272 = pi20 ? n20396 : ~n428;
  assign n33273 = pi19 ? n32 : ~n33272;
  assign n33274 = pi18 ? n33273 : n21692;
  assign n33275 = pi17 ? n32 : n33274;
  assign n33276 = pi16 ? n32 : n33275;
  assign n33277 = pi15 ? n33276 : n32;
  assign n33278 = pi19 ? n32 : ~n221;
  assign n33279 = pi18 ? n33278 : n13080;
  assign n33280 = pi17 ? n32 : n33279;
  assign n33281 = pi16 ? n32 : n33280;
  assign n33282 = pi19 ? n32 : ~n4126;
  assign n33283 = pi18 ? n33282 : ~n6063;
  assign n33284 = pi17 ? n32 : n33283;
  assign n33285 = pi16 ? n32 : n33284;
  assign n33286 = pi15 ? n33281 : n33285;
  assign n33287 = pi14 ? n33277 : n33286;
  assign n33288 = pi18 ? n17118 : n13945;
  assign n33289 = pi17 ? n32 : n33288;
  assign n33290 = pi16 ? n32 : n33289;
  assign n33291 = pi15 ? n33290 : n13948;
  assign n33292 = pi18 ? n16847 : n13945;
  assign n33293 = pi17 ? n32 : n33292;
  assign n33294 = pi16 ? n32 : n33293;
  assign n33295 = pi14 ? n33291 : n33294;
  assign n33296 = pi13 ? n33287 : n33295;
  assign n33297 = pi18 ? n4722 : ~n2413;
  assign n33298 = pi17 ? n32 : n33297;
  assign n33299 = pi16 ? n32 : n33298;
  assign n33300 = pi18 ? n4127 : n21229;
  assign n33301 = pi17 ? n32 : n33300;
  assign n33302 = pi16 ? n32 : n33301;
  assign n33303 = pi15 ? n33299 : n33302;
  assign n33304 = pi19 ? n24349 : ~n32;
  assign n33305 = pi18 ? n4722 : ~n33304;
  assign n33306 = pi17 ? n32 : n33305;
  assign n33307 = pi16 ? n32 : n33306;
  assign n33308 = pi15 ? n33307 : n13948;
  assign n33309 = pi14 ? n33303 : n33308;
  assign n33310 = pi19 ? n531 : ~n321;
  assign n33311 = pi18 ? n14153 : n33310;
  assign n33312 = pi19 ? n321 : ~n32;
  assign n33313 = pi18 ? n33312 : ~n32;
  assign n33314 = pi17 ? n33311 : n33313;
  assign n33315 = pi16 ? n1471 : ~n33314;
  assign n33316 = pi16 ? n1135 : ~n4055;
  assign n33317 = pi15 ? n33315 : n33316;
  assign n33318 = pi18 ? n15406 : n237;
  assign n33319 = pi17 ? n23931 : n33318;
  assign n33320 = pi16 ? n1214 : ~n33319;
  assign n33321 = pi18 ? n20164 : n2413;
  assign n33322 = pi17 ? n14983 : n33321;
  assign n33323 = pi16 ? n1471 : ~n33322;
  assign n33324 = pi15 ? n33320 : n33323;
  assign n33325 = pi14 ? n33317 : n33324;
  assign n33326 = pi13 ? n33309 : n33325;
  assign n33327 = pi12 ? n33296 : n33326;
  assign n33328 = pi18 ? n16234 : ~n23073;
  assign n33329 = pi17 ? n32 : n33328;
  assign n33330 = pi16 ? n32 : n33329;
  assign n33331 = pi18 ? n15849 : n4343;
  assign n33332 = pi17 ? n32 : n33331;
  assign n33333 = pi16 ? n32 : n33332;
  assign n33334 = pi15 ? n33330 : n33333;
  assign n33335 = pi18 ? n18183 : ~n532;
  assign n33336 = pi17 ? n32 : n33335;
  assign n33337 = pi16 ? n32 : n33336;
  assign n33338 = pi19 ? n15923 : n32;
  assign n33339 = pi18 ? n15849 : n33338;
  assign n33340 = pi17 ? n32 : n33339;
  assign n33341 = pi16 ? n32 : n33340;
  assign n33342 = pi15 ? n33337 : n33341;
  assign n33343 = pi14 ? n33334 : n33342;
  assign n33344 = pi18 ? n496 : ~n3786;
  assign n33345 = pi17 ? n32 : n33344;
  assign n33346 = pi16 ? n32 : n33345;
  assign n33347 = pi18 ? n697 : ~n3786;
  assign n33348 = pi17 ? n32 : n33347;
  assign n33349 = pi16 ? n32 : n33348;
  assign n33350 = pi15 ? n33349 : n33135;
  assign n33351 = pi14 ? n33346 : n33350;
  assign n33352 = pi13 ? n33343 : n33351;
  assign n33353 = pi18 ? n209 : ~n14982;
  assign n33354 = pi17 ? n32 : n33353;
  assign n33355 = pi17 ? n20165 : n2531;
  assign n33356 = pi16 ? n33354 : ~n33355;
  assign n33357 = pi17 ? n20065 : n33128;
  assign n33358 = pi16 ? n32 : n33357;
  assign n33359 = pi15 ? n33356 : n33358;
  assign n33360 = pi17 ? n20065 : n32781;
  assign n33361 = pi16 ? n32 : n33360;
  assign n33362 = pi18 ? n209 : ~n13416;
  assign n33363 = pi17 ? n32 : n33362;
  assign n33364 = pi16 ? n33363 : ~n1934;
  assign n33365 = pi15 ? n33361 : n33364;
  assign n33366 = pi14 ? n33359 : n33365;
  assign n33367 = pi18 ? n222 : ~n17118;
  assign n33368 = pi17 ? n32 : n33367;
  assign n33369 = pi19 ? n32 : ~n22185;
  assign n33370 = pi18 ? n237 : ~n33369;
  assign n33371 = pi17 ? n33370 : ~n1933;
  assign n33372 = pi16 ? n33368 : n33371;
  assign n33373 = pi18 ? n22186 : ~n350;
  assign n33374 = pi17 ? n22184 : ~n33373;
  assign n33375 = pi16 ? n1214 : ~n33374;
  assign n33376 = pi15 ? n33372 : n33375;
  assign n33377 = pi18 ? n16801 : ~n6059;
  assign n33378 = pi17 ? n32 : n33377;
  assign n33379 = pi16 ? n1135 : ~n33378;
  assign n33380 = pi14 ? n33376 : n33379;
  assign n33381 = pi13 ? n33366 : n33380;
  assign n33382 = pi12 ? n33352 : n33381;
  assign n33383 = pi11 ? n33327 : n33382;
  assign n33384 = pi10 ? n33271 : n33383;
  assign n33385 = pi09 ? n32 : n33384;
  assign n33386 = pi14 ? n32 : n15127;
  assign n33387 = pi13 ? n33386 : n15123;
  assign n33388 = pi15 ? n15263 : n19172;
  assign n33389 = pi14 ? n15123 : n33388;
  assign n33390 = pi18 ? n209 : ~n2627;
  assign n33391 = pi17 ? n32 : n33390;
  assign n33392 = pi16 ? n32 : n33391;
  assign n33393 = pi15 ? n33242 : n33392;
  assign n33394 = pi18 ? n863 : ~n2627;
  assign n33395 = pi17 ? n32 : n33394;
  assign n33396 = pi16 ? n32 : n33395;
  assign n33397 = pi18 ? n863 : n22752;
  assign n33398 = pi17 ? n32 : n33397;
  assign n33399 = pi16 ? n32 : n33398;
  assign n33400 = pi15 ? n33396 : n33399;
  assign n33401 = pi14 ? n33393 : n33400;
  assign n33402 = pi13 ? n33389 : n33401;
  assign n33403 = pi12 ? n33387 : n33402;
  assign n33404 = pi15 ? n33246 : n21853;
  assign n33405 = pi14 ? n33404 : n21853;
  assign n33406 = pi15 ? n21928 : n21686;
  assign n33407 = pi14 ? n33256 : n33406;
  assign n33408 = pi13 ? n33405 : n33407;
  assign n33409 = pi15 ? n14394 : n22006;
  assign n33410 = pi14 ? n33409 : n33259;
  assign n33411 = pi18 ? n15844 : n21316;
  assign n33412 = pi17 ? n32 : n33411;
  assign n33413 = pi16 ? n32 : n33412;
  assign n33414 = pi18 ? n20359 : ~n323;
  assign n33415 = pi17 ? n32 : n33414;
  assign n33416 = pi16 ? n32 : n33415;
  assign n33417 = pi15 ? n33413 : n33416;
  assign n33418 = pi14 ? n21319 : n33417;
  assign n33419 = pi13 ? n33410 : n33418;
  assign n33420 = pi12 ? n33408 : n33419;
  assign n33421 = pi11 ? n33403 : n33420;
  assign n33422 = pi19 ? n32 : n428;
  assign n33423 = pi18 ? n33422 : n9012;
  assign n33424 = pi17 ? n32 : n33423;
  assign n33425 = pi16 ? n32 : n33424;
  assign n33426 = pi15 ? n33425 : n32;
  assign n33427 = pi14 ? n33426 : n33286;
  assign n33428 = pi13 ? n33427 : n33295;
  assign n33429 = pi18 ? n4722 : ~n797;
  assign n33430 = pi17 ? n32 : n33429;
  assign n33431 = pi16 ? n32 : n33430;
  assign n33432 = pi18 ? n4127 : n13940;
  assign n33433 = pi17 ? n32 : n33432;
  assign n33434 = pi16 ? n32 : n33433;
  assign n33435 = pi15 ? n33431 : n33434;
  assign n33436 = pi14 ? n33435 : n33308;
  assign n33437 = pi18 ? n20164 : n605;
  assign n33438 = pi17 ? n14983 : n33437;
  assign n33439 = pi16 ? n1471 : ~n33438;
  assign n33440 = pi15 ? n33320 : n33439;
  assign n33441 = pi14 ? n33317 : n33440;
  assign n33442 = pi13 ? n33436 : n33441;
  assign n33443 = pi12 ? n33428 : n33442;
  assign n33444 = pi15 ? n33337 : n33333;
  assign n33445 = pi14 ? n33334 : n33444;
  assign n33446 = pi18 ? n496 : ~n532;
  assign n33447 = pi17 ? n32 : n33446;
  assign n33448 = pi16 ? n32 : n33447;
  assign n33449 = pi18 ? n702 : ~n3786;
  assign n33450 = pi17 ? n32 : n33449;
  assign n33451 = pi16 ? n32 : n33450;
  assign n33452 = pi15 ? n33349 : n33451;
  assign n33453 = pi14 ? n33448 : n33452;
  assign n33454 = pi13 ? n33445 : n33453;
  assign n33455 = pi17 ? n20165 : n3787;
  assign n33456 = pi16 ? n33354 : ~n33455;
  assign n33457 = pi18 ? n323 : ~n3786;
  assign n33458 = pi17 ? n20065 : n33457;
  assign n33459 = pi16 ? n32 : n33458;
  assign n33460 = pi15 ? n33456 : n33459;
  assign n33461 = pi14 ? n33460 : n33365;
  assign n33462 = pi16 ? n1233 : ~n33378;
  assign n33463 = pi15 ? n33379 : n33462;
  assign n33464 = pi14 ? n33376 : n33463;
  assign n33465 = pi13 ? n33461 : n33464;
  assign n33466 = pi12 ? n33454 : n33465;
  assign n33467 = pi11 ? n33443 : n33466;
  assign n33468 = pi10 ? n33421 : n33467;
  assign n33469 = pi09 ? n32 : n33468;
  assign n33470 = pi08 ? n33385 : n33469;
  assign n33471 = pi14 ? n32 : n15390;
  assign n33472 = pi13 ? n33471 : n15123;
  assign n33473 = pi15 ? n15123 : n19172;
  assign n33474 = pi14 ? n15123 : n33473;
  assign n33475 = pi15 ? n33242 : n12764;
  assign n33476 = pi19 ? n19411 : ~n32;
  assign n33477 = pi18 ? n863 : ~n33476;
  assign n33478 = pi17 ? n32 : n33477;
  assign n33479 = pi16 ? n32 : n33478;
  assign n33480 = pi20 ? n785 : n7880;
  assign n33481 = pi19 ? n33480 : n32;
  assign n33482 = pi18 ? n32 : n33481;
  assign n33483 = pi17 ? n32 : n33482;
  assign n33484 = pi16 ? n32 : n33483;
  assign n33485 = pi15 ? n33479 : n33484;
  assign n33486 = pi14 ? n33475 : n33485;
  assign n33487 = pi13 ? n33474 : n33486;
  assign n33488 = pi12 ? n33472 : n33487;
  assign n33489 = pi20 ? n206 : n246;
  assign n33490 = pi19 ? n33489 : n32;
  assign n33491 = pi18 ? n32 : n33490;
  assign n33492 = pi17 ? n32 : n33491;
  assign n33493 = pi16 ? n32 : n33492;
  assign n33494 = pi20 ? n32 : n16650;
  assign n33495 = pi19 ? n33494 : n32;
  assign n33496 = pi18 ? n32 : n33495;
  assign n33497 = pi17 ? n32 : n33496;
  assign n33498 = pi16 ? n32 : n33497;
  assign n33499 = pi15 ? n33493 : n33498;
  assign n33500 = pi15 ? n33498 : n14973;
  assign n33501 = pi14 ? n33499 : n33500;
  assign n33502 = pi20 ? n428 : n25513;
  assign n33503 = pi19 ? n33502 : n32;
  assign n33504 = pi18 ? n32 : n33503;
  assign n33505 = pi17 ? n32 : n33504;
  assign n33506 = pi16 ? n32 : n33505;
  assign n33507 = pi15 ? n33506 : n14790;
  assign n33508 = pi19 ? n20006 : n32;
  assign n33509 = pi18 ? n936 : n33508;
  assign n33510 = pi17 ? n32 : n33509;
  assign n33511 = pi16 ? n32 : n33510;
  assign n33512 = pi15 ? n14790 : n33511;
  assign n33513 = pi14 ? n33507 : n33512;
  assign n33514 = pi13 ? n33501 : n33513;
  assign n33515 = pi18 ? n268 : n4983;
  assign n33516 = pi17 ? n32 : n33515;
  assign n33517 = pi16 ? n32 : n33516;
  assign n33518 = pi15 ? n33517 : n21319;
  assign n33519 = pi14 ? n33518 : n32;
  assign n33520 = pi20 ? n339 : ~n246;
  assign n33521 = pi19 ? n266 : ~n33520;
  assign n33522 = pi18 ? n32 : n33521;
  assign n33523 = pi17 ? n32 : n33522;
  assign n33524 = pi20 ? n5854 : ~n2385;
  assign n33525 = pi19 ? n33524 : ~n7939;
  assign n33526 = pi20 ? n207 : ~n1817;
  assign n33527 = pi19 ? n13714 : n33526;
  assign n33528 = pi18 ? n33525 : ~n33527;
  assign n33529 = pi19 ? n31490 : n32;
  assign n33530 = pi18 ? n33529 : n5351;
  assign n33531 = pi17 ? n33528 : n33530;
  assign n33532 = pi16 ? n33523 : n33531;
  assign n33533 = pi15 ? n14397 : n33532;
  assign n33534 = pi19 ? n22525 : ~n5371;
  assign n33535 = pi18 ? n14153 : n33534;
  assign n33536 = pi19 ? n321 : ~n221;
  assign n33537 = pi20 ? n266 : n1685;
  assign n33538 = pi19 ? n33537 : n32;
  assign n33539 = pi18 ? n33536 : n33538;
  assign n33540 = pi17 ? n33535 : n33539;
  assign n33541 = pi16 ? n32 : n33540;
  assign n33542 = pi19 ? n5675 : ~n5371;
  assign n33543 = pi18 ? n13945 : n33542;
  assign n33544 = pi20 ? n175 : n342;
  assign n33545 = pi19 ? n33544 : ~n267;
  assign n33546 = pi18 ? n33545 : ~n520;
  assign n33547 = pi17 ? n33543 : n33546;
  assign n33548 = pi16 ? n32 : n33547;
  assign n33549 = pi15 ? n33541 : n33548;
  assign n33550 = pi14 ? n33533 : n33549;
  assign n33551 = pi13 ? n33519 : n33550;
  assign n33552 = pi12 ? n33514 : n33551;
  assign n33553 = pi11 ? n33488 : n33552;
  assign n33554 = pi19 ? n15135 : n32;
  assign n33555 = pi18 ? n16041 : n33554;
  assign n33556 = pi17 ? n32 : n33555;
  assign n33557 = pi16 ? n32 : n33556;
  assign n33558 = pi19 ? n10120 : ~n32;
  assign n33559 = pi18 ? n697 : ~n33558;
  assign n33560 = pi17 ? n32 : n33559;
  assign n33561 = pi16 ? n32 : n33560;
  assign n33562 = pi15 ? n33557 : n33561;
  assign n33563 = pi14 ? n32128 : n33562;
  assign n33564 = pi18 ? n17118 : n5749;
  assign n33565 = pi17 ? n32 : n33564;
  assign n33566 = pi16 ? n32 : n33565;
  assign n33567 = pi18 ? n268 : n13945;
  assign n33568 = pi17 ? n32 : n33567;
  assign n33569 = pi16 ? n32 : n33568;
  assign n33570 = pi15 ? n33566 : n33569;
  assign n33571 = pi18 ? n268 : n13940;
  assign n33572 = pi17 ? n32 : n33571;
  assign n33573 = pi16 ? n32 : n33572;
  assign n33574 = pi15 ? n33294 : n33573;
  assign n33575 = pi14 ? n33570 : n33574;
  assign n33576 = pi13 ? n33563 : n33575;
  assign n33577 = pi15 ? n32219 : n13943;
  assign n33578 = pi20 ? n206 : n749;
  assign n33579 = pi19 ? n33578 : ~n32;
  assign n33580 = pi18 ? n880 : ~n33579;
  assign n33581 = pi17 ? n32 : n33580;
  assign n33582 = pi16 ? n32 : n33581;
  assign n33583 = pi15 ? n33582 : n13943;
  assign n33584 = pi14 ? n33577 : n33583;
  assign n33585 = pi16 ? n1233 : ~n4733;
  assign n33586 = pi15 ? n33315 : n33585;
  assign n33587 = pi18 ? n16394 : n5436;
  assign n33588 = pi17 ? n24698 : n33587;
  assign n33589 = pi16 ? n1135 : ~n33588;
  assign n33590 = pi15 ? n33589 : n33439;
  assign n33591 = pi14 ? n33586 : n33590;
  assign n33592 = pi13 ? n33584 : n33591;
  assign n33593 = pi12 ? n33576 : n33592;
  assign n33594 = pi19 ? n32 : n6997;
  assign n33595 = pi20 ? n246 : n243;
  assign n33596 = pi19 ? n33595 : ~n32;
  assign n33597 = pi18 ? n33594 : ~n33596;
  assign n33598 = pi17 ? n32 : n33597;
  assign n33599 = pi16 ? n32 : n33598;
  assign n33600 = pi18 ? n15849 : n13372;
  assign n33601 = pi17 ? n32 : n33600;
  assign n33602 = pi16 ? n32 : n33601;
  assign n33603 = pi15 ? n33599 : n33602;
  assign n33604 = pi18 ? n18183 : ~n418;
  assign n33605 = pi17 ? n32 : n33604;
  assign n33606 = pi16 ? n32 : n33605;
  assign n33607 = pi15 ? n33606 : n33602;
  assign n33608 = pi14 ? n33603 : n33607;
  assign n33609 = pi18 ? n496 : ~n418;
  assign n33610 = pi17 ? n32 : n33609;
  assign n33611 = pi16 ? n32 : n33610;
  assign n33612 = pi18 ? n496 : n21597;
  assign n33613 = pi17 ? n32 : n33612;
  assign n33614 = pi16 ? n32 : n33613;
  assign n33615 = pi15 ? n33611 : n33614;
  assign n33616 = pi18 ? n697 : ~n532;
  assign n33617 = pi17 ? n32 : n33616;
  assign n33618 = pi16 ? n32 : n33617;
  assign n33619 = pi15 ? n33618 : n33135;
  assign n33620 = pi14 ? n33615 : n33619;
  assign n33621 = pi13 ? n33608 : n33620;
  assign n33622 = pi18 ? n1395 : ~n14982;
  assign n33623 = pi17 ? n32 : n33622;
  assign n33624 = pi17 ? n25209 : n2531;
  assign n33625 = pi16 ? n33623 : ~n33624;
  assign n33626 = pi17 ? n18395 : n33128;
  assign n33627 = pi16 ? n32 : n33626;
  assign n33628 = pi15 ? n33625 : n33627;
  assign n33629 = pi17 ? n18395 : n32781;
  assign n33630 = pi16 ? n32 : n33629;
  assign n33631 = pi18 ? n341 : ~n14413;
  assign n33632 = pi17 ? n32 : n33631;
  assign n33633 = pi16 ? n33632 : ~n1934;
  assign n33634 = pi15 ? n33630 : n33633;
  assign n33635 = pi14 ? n33628 : n33634;
  assign n33636 = pi19 ? n22185 : ~n246;
  assign n33637 = pi19 ? n32 : ~n20555;
  assign n33638 = pi18 ? n33636 : ~n33637;
  assign n33639 = pi17 ? n33638 : ~n1933;
  assign n33640 = pi16 ? n33368 : n33639;
  assign n33641 = pi18 ? n1464 : n350;
  assign n33642 = pi17 ? n18560 : n33641;
  assign n33643 = pi16 ? n1135 : ~n33642;
  assign n33644 = pi15 ? n33640 : n33643;
  assign n33645 = pi18 ? n16801 : n237;
  assign n33646 = pi17 ? n32 : n33645;
  assign n33647 = pi16 ? n1135 : ~n33646;
  assign n33648 = pi18 ? n16389 : n1353;
  assign n33649 = pi17 ? n32 : n33648;
  assign n33650 = pi16 ? n1135 : ~n33649;
  assign n33651 = pi15 ? n33647 : n33650;
  assign n33652 = pi14 ? n33644 : n33651;
  assign n33653 = pi13 ? n33635 : n33652;
  assign n33654 = pi12 ? n33621 : n33653;
  assign n33655 = pi11 ? n33593 : n33654;
  assign n33656 = pi10 ? n33553 : n33655;
  assign n33657 = pi09 ? n32 : n33656;
  assign n33658 = pi14 ? n24193 : n22347;
  assign n33659 = pi13 ? n33471 : n33658;
  assign n33660 = pi15 ? n22347 : n19172;
  assign n33661 = pi14 ? n23179 : n33660;
  assign n33662 = pi20 ? n785 : n1385;
  assign n33663 = pi19 ? n33662 : n32;
  assign n33664 = pi18 ? n32 : n33663;
  assign n33665 = pi17 ? n32 : n33664;
  assign n33666 = pi16 ? n32 : n33665;
  assign n33667 = pi15 ? n33479 : n33666;
  assign n33668 = pi14 ? n33475 : n33667;
  assign n33669 = pi13 ? n33661 : n33668;
  assign n33670 = pi12 ? n33659 : n33669;
  assign n33671 = pi15 ? n33493 : n32;
  assign n33672 = pi15 ? n648 : n14973;
  assign n33673 = pi14 ? n33671 : n33672;
  assign n33674 = pi20 ? n3523 : ~n206;
  assign n33675 = pi19 ? n33674 : n32;
  assign n33676 = pi18 ? n936 : n33675;
  assign n33677 = pi17 ? n32 : n33676;
  assign n33678 = pi16 ? n32 : n33677;
  assign n33679 = pi15 ? n14790 : n33678;
  assign n33680 = pi14 ? n33507 : n33679;
  assign n33681 = pi13 ? n33673 : n33680;
  assign n33682 = pi14 ? n33518 : n659;
  assign n33683 = pi20 ? n266 : n6621;
  assign n33684 = pi19 ? n33683 : ~n33520;
  assign n33685 = pi18 ? n32 : n33684;
  assign n33686 = pi17 ? n32 : n33685;
  assign n33687 = pi19 ? n28862 : n18834;
  assign n33688 = pi20 ? n18834 : n321;
  assign n33689 = pi20 ? n10644 : ~n9641;
  assign n33690 = pi19 ? n33688 : n33689;
  assign n33691 = pi18 ? n33687 : n33690;
  assign n33692 = pi19 ? n501 : n32;
  assign n33693 = pi18 ? n33692 : n5351;
  assign n33694 = pi17 ? n33691 : ~n33693;
  assign n33695 = pi16 ? n33686 : ~n33694;
  assign n33696 = pi15 ? n14397 : n33695;
  assign n33697 = pi14 ? n33696 : n33549;
  assign n33698 = pi13 ? n33682 : n33697;
  assign n33699 = pi12 ? n33681 : n33698;
  assign n33700 = pi11 ? n33670 : n33699;
  assign n33701 = pi20 ? n206 : n1475;
  assign n33702 = pi19 ? n33701 : ~n32;
  assign n33703 = pi18 ? n880 : ~n33702;
  assign n33704 = pi17 ? n32 : n33703;
  assign n33705 = pi16 ? n32 : n33704;
  assign n33706 = pi15 ? n33705 : n13943;
  assign n33707 = pi14 ? n33577 : n33706;
  assign n33708 = pi16 ? n1135 : ~n4733;
  assign n33709 = pi15 ? n33315 : n33708;
  assign n33710 = pi18 ? n16394 : n23291;
  assign n33711 = pi17 ? n24698 : n33710;
  assign n33712 = pi16 ? n1135 : ~n33711;
  assign n33713 = pi15 ? n33712 : n33439;
  assign n33714 = pi14 ? n33709 : n33713;
  assign n33715 = pi13 ? n33707 : n33714;
  assign n33716 = pi12 ? n33576 : n33715;
  assign n33717 = pi18 ? n33594 : ~n5436;
  assign n33718 = pi17 ? n32 : n33717;
  assign n33719 = pi16 ? n32 : n33718;
  assign n33720 = pi15 ? n33719 : n33602;
  assign n33721 = pi14 ? n33720 : n33607;
  assign n33722 = pi13 ? n33721 : n33620;
  assign n33723 = pi16 ? n33354 : ~n33624;
  assign n33724 = pi15 ? n33723 : n33627;
  assign n33725 = pi14 ? n33724 : n33634;
  assign n33726 = pi16 ? n1233 : ~n33649;
  assign n33727 = pi15 ? n33647 : n33726;
  assign n33728 = pi14 ? n33644 : n33727;
  assign n33729 = pi13 ? n33725 : n33728;
  assign n33730 = pi12 ? n33722 : n33729;
  assign n33731 = pi11 ? n33716 : n33730;
  assign n33732 = pi10 ? n33700 : n33731;
  assign n33733 = pi09 ? n32 : n33732;
  assign n33734 = pi08 ? n33657 : n33733;
  assign n33735 = pi07 ? n33470 : n33734;
  assign n33736 = pi14 ? n32 : n22543;
  assign n33737 = pi21 ? n206 : n2076;
  assign n33738 = pi20 ? n32 : n33737;
  assign n33739 = pi19 ? n33738 : n32;
  assign n33740 = pi18 ? n32 : n33739;
  assign n33741 = pi17 ? n32 : n33740;
  assign n33742 = pi16 ? n32 : n33741;
  assign n33743 = pi15 ? n15389 : n33742;
  assign n33744 = pi14 ? n15389 : n33743;
  assign n33745 = pi13 ? n33736 : n33744;
  assign n33746 = pi14 ? n22252 : n15123;
  assign n33747 = pi13 ? n22426 : n33746;
  assign n33748 = pi12 ? n33745 : n33747;
  assign n33749 = pi15 ? n648 : n15123;
  assign n33750 = pi14 ? n33749 : n15123;
  assign n33751 = pi20 ? n18624 : ~n428;
  assign n33752 = pi19 ? n33751 : n32;
  assign n33753 = pi18 ? n863 : n33752;
  assign n33754 = pi17 ? n32 : n33753;
  assign n33755 = pi16 ? n32 : n33754;
  assign n33756 = pi20 ? n1685 : n206;
  assign n33757 = pi19 ? n33756 : ~n32;
  assign n33758 = pi18 ? n4380 : ~n33757;
  assign n33759 = pi17 ? n32 : n33758;
  assign n33760 = pi16 ? n32 : n33759;
  assign n33761 = pi15 ? n33755 : n33760;
  assign n33762 = pi14 ? n15123 : n33761;
  assign n33763 = pi13 ? n33750 : n33762;
  assign n33764 = pi14 ? n30211 : n21681;
  assign n33765 = pi18 ? n3496 : n22003;
  assign n33766 = pi17 ? n32 : n33765;
  assign n33767 = pi16 ? n32 : n33766;
  assign n33768 = pi15 ? n14394 : n33767;
  assign n33769 = pi19 ? n9037 : ~n5356;
  assign n33770 = pi18 ? n32 : n33769;
  assign n33771 = pi17 ? n32 : n33770;
  assign n33772 = pi18 ? n18668 : n18941;
  assign n33773 = pi20 ? n321 : ~n17712;
  assign n33774 = pi19 ? n33773 : ~n32;
  assign n33775 = pi18 ? n4671 : n33774;
  assign n33776 = pi17 ? n33772 : n33775;
  assign n33777 = pi16 ? n33771 : ~n33776;
  assign n33778 = pi15 ? n33777 : n21543;
  assign n33779 = pi14 ? n33768 : n33778;
  assign n33780 = pi13 ? n33764 : n33779;
  assign n33781 = pi12 ? n33763 : n33780;
  assign n33782 = pi11 ? n33748 : n33781;
  assign n33783 = pi19 ? n28623 : n32;
  assign n33784 = pi19 ? n4982 : ~n23813;
  assign n33785 = pi18 ? n33783 : n33784;
  assign n33786 = pi20 ? n342 : ~n310;
  assign n33787 = pi19 ? n33786 : n15405;
  assign n33788 = pi18 ? n33787 : n9578;
  assign n33789 = pi17 ? n33785 : n33788;
  assign n33790 = pi16 ? n32 : n33789;
  assign n33791 = pi15 ? n21686 : n33790;
  assign n33792 = pi19 ? n32 : n20555;
  assign n33793 = pi18 ? n33792 : n32;
  assign n33794 = pi17 ? n32 : n33793;
  assign n33795 = pi16 ? n32 : n33794;
  assign n33796 = pi20 ? n266 : ~n266;
  assign n33797 = pi19 ? n33796 : ~n32;
  assign n33798 = pi18 ? n496 : ~n33797;
  assign n33799 = pi17 ? n32 : n33798;
  assign n33800 = pi16 ? n32 : n33799;
  assign n33801 = pi15 ? n33795 : n33800;
  assign n33802 = pi14 ? n33791 : n33801;
  assign n33803 = pi15 ? n32 : n23404;
  assign n33804 = pi15 ? n13948 : n13943;
  assign n33805 = pi14 ? n33803 : n33804;
  assign n33806 = pi13 ? n33802 : n33805;
  assign n33807 = pi19 ? n32 : n6722;
  assign n33808 = pi18 ? n33807 : n17650;
  assign n33809 = pi17 ? n32 : n33808;
  assign n33810 = pi16 ? n32 : n33809;
  assign n33811 = pi15 ? n33810 : n13360;
  assign n33812 = pi18 ? n9012 : n863;
  assign n33813 = pi18 ? n5657 : n13940;
  assign n33814 = pi17 ? n33812 : n33813;
  assign n33815 = pi16 ? n32 : n33814;
  assign n33816 = pi15 ? n13360 : n33815;
  assign n33817 = pi14 ? n33811 : n33816;
  assign n33818 = pi19 ? n18396 : n18478;
  assign n33819 = pi18 ? n22497 : n33818;
  assign n33820 = pi18 ? n22502 : n32;
  assign n33821 = pi17 ? n33819 : ~n33820;
  assign n33822 = pi16 ? n28993 : ~n33821;
  assign n33823 = pi20 ? n246 : ~n274;
  assign n33824 = pi19 ? n33823 : ~n32;
  assign n33825 = pi18 ? n18710 : n33824;
  assign n33826 = pi17 ? n32 : n33825;
  assign n33827 = pi16 ? n1233 : ~n33826;
  assign n33828 = pi15 ? n33822 : n33827;
  assign n33829 = pi17 ? n25761 : n2408;
  assign n33830 = pi16 ? n1214 : ~n33829;
  assign n33831 = pi17 ? n15850 : n2119;
  assign n33832 = pi16 ? n1471 : ~n33831;
  assign n33833 = pi15 ? n33830 : n33832;
  assign n33834 = pi14 ? n33828 : n33833;
  assign n33835 = pi13 ? n33817 : n33834;
  assign n33836 = pi12 ? n33806 : n33835;
  assign n33837 = pi18 ? n1249 : n5005;
  assign n33838 = pi17 ? n32 : n33837;
  assign n33839 = pi16 ? n32 : n33838;
  assign n33840 = pi18 ? n880 : n13668;
  assign n33841 = pi17 ? n32 : n33840;
  assign n33842 = pi16 ? n32 : n33841;
  assign n33843 = pi15 ? n33839 : n33842;
  assign n33844 = pi14 ? n33843 : n13671;
  assign n33845 = pi19 ? n28639 : n32;
  assign n33846 = pi18 ? n880 : n33845;
  assign n33847 = pi17 ? n32 : n33846;
  assign n33848 = pi16 ? n32 : n33847;
  assign n33849 = pi15 ? n33848 : n12098;
  assign n33850 = pi20 ? n915 : n339;
  assign n33851 = pi19 ? n33850 : ~n32;
  assign n33852 = pi18 ? n880 : ~n33851;
  assign n33853 = pi17 ? n14395 : n33852;
  assign n33854 = pi16 ? n32 : n33853;
  assign n33855 = pi17 ? n21952 : n33609;
  assign n33856 = pi16 ? n32 : n33855;
  assign n33857 = pi15 ? n33854 : n33856;
  assign n33858 = pi14 ? n33849 : n33857;
  assign n33859 = pi13 ? n33844 : n33858;
  assign n33860 = pi19 ? n21740 : n236;
  assign n33861 = pi18 ? n222 : ~n33860;
  assign n33862 = pi17 ? n32 : n33861;
  assign n33863 = pi17 ? n16802 : n2531;
  assign n33864 = pi16 ? n33862 : ~n33863;
  assign n33865 = pi19 ? n5694 : ~n349;
  assign n33866 = pi18 ? n20020 : n33865;
  assign n33867 = pi19 ? n9007 : ~n32;
  assign n33868 = pi18 ? n33867 : ~n532;
  assign n33869 = pi17 ? n33866 : n33868;
  assign n33870 = pi16 ? n32 : n33869;
  assign n33871 = pi15 ? n33864 : n33870;
  assign n33872 = pi19 ? n247 : ~n1757;
  assign n33873 = pi18 ? n209 : ~n33872;
  assign n33874 = pi17 ? n32 : n33873;
  assign n33875 = pi19 ? n5707 : ~n207;
  assign n33876 = pi19 ? n22185 : ~n4342;
  assign n33877 = pi18 ? n33875 : ~n33876;
  assign n33878 = pi19 ? n5371 : ~n1464;
  assign n33879 = pi18 ? n33878 : ~n430;
  assign n33880 = pi17 ? n33877 : ~n33879;
  assign n33881 = pi16 ? n33874 : ~n33880;
  assign n33882 = pi15 ? n33135 : n33881;
  assign n33883 = pi14 ? n33871 : n33882;
  assign n33884 = pi18 ? n880 : n350;
  assign n33885 = pi17 ? n16450 : n33884;
  assign n33886 = pi16 ? n1135 : ~n33885;
  assign n33887 = pi18 ? n22526 : n350;
  assign n33888 = pi17 ? n32 : n33887;
  assign n33889 = pi16 ? n1135 : ~n33888;
  assign n33890 = pi15 ? n33886 : n33889;
  assign n33891 = pi14 ? n33890 : n30941;
  assign n33892 = pi13 ? n33883 : n33891;
  assign n33893 = pi12 ? n33859 : n33892;
  assign n33894 = pi11 ? n33836 : n33893;
  assign n33895 = pi10 ? n33782 : n33894;
  assign n33896 = pi09 ? n32 : n33895;
  assign n33897 = pi15 ? n22540 : n15389;
  assign n33898 = pi19 ? n23944 : n32;
  assign n33899 = pi18 ? n32 : n33898;
  assign n33900 = pi17 ? n32 : n33899;
  assign n33901 = pi16 ? n32 : n33900;
  assign n33902 = pi15 ? n22540 : n33901;
  assign n33903 = pi14 ? n33897 : n33902;
  assign n33904 = pi13 ? n33736 : n33903;
  assign n33905 = pi15 ? n15123 : n22347;
  assign n33906 = pi14 ? n22252 : n33905;
  assign n33907 = pi13 ? n22544 : n33906;
  assign n33908 = pi12 ? n33904 : n33907;
  assign n33909 = pi13 ? n15123 : n33762;
  assign n33910 = pi18 ? n3496 : n5351;
  assign n33911 = pi17 ? n32 : n33910;
  assign n33912 = pi16 ? n32 : n33911;
  assign n33913 = pi15 ? n14394 : n33912;
  assign n33914 = pi19 ? n13529 : ~n32;
  assign n33915 = pi18 ? n4671 : n33914;
  assign n33916 = pi17 ? n33772 : n33915;
  assign n33917 = pi16 ? n33771 : ~n33916;
  assign n33918 = pi15 ? n33917 : n21543;
  assign n33919 = pi14 ? n33913 : n33918;
  assign n33920 = pi13 ? n33764 : n33919;
  assign n33921 = pi12 ? n33909 : n33920;
  assign n33922 = pi11 ? n33908 : n33921;
  assign n33923 = pi20 ? n342 : n287;
  assign n33924 = pi19 ? n33923 : n32;
  assign n33925 = pi19 ? n4982 : ~n23806;
  assign n33926 = pi18 ? n33924 : n33925;
  assign n33927 = pi17 ? n33926 : n33788;
  assign n33928 = pi16 ? n32 : n33927;
  assign n33929 = pi15 ? n21543 : n33928;
  assign n33930 = pi14 ? n33929 : n33801;
  assign n33931 = pi15 ? n13948 : n14156;
  assign n33932 = pi14 ? n33803 : n33931;
  assign n33933 = pi13 ? n33930 : n33932;
  assign n33934 = pi18 ? n19082 : n17650;
  assign n33935 = pi17 ? n32 : n33934;
  assign n33936 = pi16 ? n32 : n33935;
  assign n33937 = pi18 ? n32 : n5009;
  assign n33938 = pi17 ? n32 : n33937;
  assign n33939 = pi16 ? n32 : n33938;
  assign n33940 = pi15 ? n33936 : n33939;
  assign n33941 = pi14 ? n33940 : n33816;
  assign n33942 = pi16 ? n1135 : ~n33826;
  assign n33943 = pi15 ? n33822 : n33942;
  assign n33944 = pi14 ? n33943 : n33833;
  assign n33945 = pi13 ? n33941 : n33944;
  assign n33946 = pi12 ? n33933 : n33945;
  assign n33947 = pi20 ? n749 : ~n243;
  assign n33948 = pi19 ? n33947 : n32;
  assign n33949 = pi18 ? n880 : n33948;
  assign n33950 = pi17 ? n32 : n33949;
  assign n33951 = pi16 ? n32 : n33950;
  assign n33952 = pi15 ? n33951 : n21153;
  assign n33953 = pi20 ? n915 : n243;
  assign n33954 = pi19 ? n33953 : ~n32;
  assign n33955 = pi18 ? n880 : ~n33954;
  assign n33956 = pi17 ? n14395 : n33955;
  assign n33957 = pi16 ? n32 : n33956;
  assign n33958 = pi15 ? n33957 : n33856;
  assign n33959 = pi14 ? n33952 : n33958;
  assign n33960 = pi13 ? n33844 : n33959;
  assign n33961 = pi12 ? n33960 : n33892;
  assign n33962 = pi11 ? n33946 : n33961;
  assign n33963 = pi10 ? n33922 : n33962;
  assign n33964 = pi09 ? n32 : n33963;
  assign n33965 = pi08 ? n33896 : n33964;
  assign n33966 = pi14 ? n32 : n22812;
  assign n33967 = pi19 ? n4126 : n32;
  assign n33968 = pi18 ? n32 : n33967;
  assign n33969 = pi17 ? n32 : n33968;
  assign n33970 = pi16 ? n32 : n33969;
  assign n33971 = pi15 ? n22817 : n33970;
  assign n33972 = pi14 ? n22540 : n33971;
  assign n33973 = pi13 ? n33966 : n33972;
  assign n33974 = pi13 ? n22544 : n22425;
  assign n33975 = pi12 ? n33973 : n33974;
  assign n33976 = pi14 ? n33905 : n22347;
  assign n33977 = pi19 ? n6355 : n32;
  assign n33978 = pi18 ? n32 : n33977;
  assign n33979 = pi17 ? n32 : n33978;
  assign n33980 = pi16 ? n32 : n33979;
  assign n33981 = pi15 ? n22347 : n33980;
  assign n33982 = pi17 ? n17346 : n22937;
  assign n33983 = pi16 ? n32 : n33982;
  assign n33984 = pi19 ? n22106 : ~n32;
  assign n33985 = pi18 ? n222 : ~n33984;
  assign n33986 = pi17 ? n32 : n33985;
  assign n33987 = pi16 ? n32 : n33986;
  assign n33988 = pi15 ? n33983 : n33987;
  assign n33989 = pi14 ? n33981 : n33988;
  assign n33990 = pi13 ? n33976 : n33989;
  assign n33991 = pi15 ? n32 : n14397;
  assign n33992 = pi15 ? n21853 : n21543;
  assign n33993 = pi14 ? n33991 : n33992;
  assign n33994 = pi18 ? n20172 : n15008;
  assign n33995 = pi19 ? n266 : n236;
  assign n33996 = pi20 ? n266 : n1817;
  assign n33997 = pi19 ? n33996 : n32;
  assign n33998 = pi18 ? n33995 : n33997;
  assign n33999 = pi17 ? n33994 : n33998;
  assign n34000 = pi16 ? n32 : n33999;
  assign n34001 = pi15 ? n34000 : n32;
  assign n34002 = pi14 ? n26580 : n34001;
  assign n34003 = pi13 ? n33993 : n34002;
  assign n34004 = pi12 ? n33990 : n34003;
  assign n34005 = pi11 ? n33975 : n34004;
  assign n34006 = pi19 ? n342 : n32;
  assign n34007 = pi19 ? n5694 : ~n1740;
  assign n34008 = pi18 ? n34006 : n34007;
  assign n34009 = pi19 ? n507 : n15405;
  assign n34010 = pi18 ? n34009 : n32;
  assign n34011 = pi17 ? n34008 : n34010;
  assign n34012 = pi16 ? n32 : n34011;
  assign n34013 = pi15 ? n32 : n34012;
  assign n34014 = pi18 ? n880 : ~n6019;
  assign n34015 = pi17 ? n32 : n34014;
  assign n34016 = pi16 ? n32 : n34015;
  assign n34017 = pi15 ? n19787 : n34016;
  assign n34018 = pi14 ? n34013 : n34017;
  assign n34019 = pi15 ? n32 : n21337;
  assign n34020 = pi15 ? n32 : n14156;
  assign n34021 = pi14 ? n34019 : n34020;
  assign n34022 = pi13 ? n34018 : n34021;
  assign n34023 = pi17 ? n22435 : n33937;
  assign n34024 = pi16 ? n32 : n34023;
  assign n34025 = pi15 ? n32 : n34024;
  assign n34026 = pi19 ? n16591 : n32;
  assign n34027 = pi18 ? n32 : n34026;
  assign n34028 = pi17 ? n15121 : n34027;
  assign n34029 = pi16 ? n32 : n34028;
  assign n34030 = pi19 ? n6018 : ~n220;
  assign n34031 = pi20 ? n220 : n206;
  assign n34032 = pi19 ? n34031 : ~n31488;
  assign n34033 = pi18 ? n34030 : ~n34032;
  assign n34034 = pi19 ? n32733 : n349;
  assign n34035 = pi18 ? n34034 : ~n13945;
  assign n34036 = pi17 ? n34033 : ~n34035;
  assign n34037 = pi16 ? n24246 : n34036;
  assign n34038 = pi15 ? n34029 : n34037;
  assign n34039 = pi14 ? n34025 : n34038;
  assign n34040 = pi19 ? n9592 : n32;
  assign n34041 = pi18 ? n20007 : ~n34040;
  assign n34042 = pi17 ? n32 : n34041;
  assign n34043 = pi16 ? n1135 : ~n34042;
  assign n34044 = pi16 ? n1233 : ~n2409;
  assign n34045 = pi15 ? n34043 : n34044;
  assign n34046 = pi17 ? n16395 : n2408;
  assign n34047 = pi16 ? n1214 : ~n34046;
  assign n34048 = pi17 ? n15850 : n2408;
  assign n34049 = pi16 ? n1471 : ~n34048;
  assign n34050 = pi15 ? n34047 : n34049;
  assign n34051 = pi14 ? n34045 : n34050;
  assign n34052 = pi13 ? n34039 : n34051;
  assign n34053 = pi12 ? n34022 : n34052;
  assign n34054 = pi18 ? n940 : ~n6019;
  assign n34055 = pi17 ? n32 : n34054;
  assign n34056 = pi16 ? n32 : n34055;
  assign n34057 = pi20 ? n260 : n207;
  assign n34058 = pi19 ? n34057 : ~n32;
  assign n34059 = pi18 ? n222 : ~n34058;
  assign n34060 = pi17 ? n32 : n34059;
  assign n34061 = pi16 ? n32 : n34060;
  assign n34062 = pi15 ? n34056 : n34061;
  assign n34063 = pi18 ? n32 : ~n6019;
  assign n34064 = pi17 ? n32 : n34063;
  assign n34065 = pi16 ? n32 : n34064;
  assign n34066 = pi15 ? n34065 : n23071;
  assign n34067 = pi14 ? n34062 : n34066;
  assign n34068 = pi18 ? n1965 : ~n22705;
  assign n34069 = pi17 ? n32 : n34068;
  assign n34070 = pi16 ? n32 : n34069;
  assign n34071 = pi15 ? n34070 : n12098;
  assign n34072 = pi17 ? n15121 : n22711;
  assign n34073 = pi16 ? n32 : n34072;
  assign n34074 = pi17 ? n22435 : n33604;
  assign n34075 = pi16 ? n32 : n34074;
  assign n34076 = pi15 ? n34073 : n34075;
  assign n34077 = pi14 ? n34071 : n34076;
  assign n34078 = pi13 ? n34067 : n34077;
  assign n34079 = pi18 ? n32 : n21425;
  assign n34080 = pi17 ? n32 : n34079;
  assign n34081 = pi17 ? n17284 : n2653;
  assign n34082 = pi16 ? n34080 : ~n34081;
  assign n34083 = pi20 ? n339 : n18762;
  assign n34084 = pi20 ? n1324 : ~n342;
  assign n34085 = pi19 ? n34083 : n34084;
  assign n34086 = pi18 ? n22696 : ~n34085;
  assign n34087 = pi19 ? n22701 : n32;
  assign n34088 = pi18 ? n34087 : n418;
  assign n34089 = pi17 ? n34086 : ~n34088;
  assign n34090 = pi16 ? n32 : n34089;
  assign n34091 = pi15 ? n34082 : n34090;
  assign n34092 = pi20 ? n206 : ~n342;
  assign n34093 = pi20 ? n915 : ~n339;
  assign n34094 = pi19 ? n34092 : n34093;
  assign n34095 = pi18 ? n29325 : n34094;
  assign n34096 = pi17 ? n32 : n34095;
  assign n34097 = pi20 ? n1331 : n2385;
  assign n34098 = pi19 ? n34097 : n342;
  assign n34099 = pi20 ? n342 : n18129;
  assign n34100 = pi20 ? n17665 : n9641;
  assign n34101 = pi19 ? n34099 : n34100;
  assign n34102 = pi18 ? n34098 : n34101;
  assign n34103 = pi19 ? n20940 : ~n22702;
  assign n34104 = pi18 ? n34103 : n6059;
  assign n34105 = pi17 ? n34102 : n34104;
  assign n34106 = pi16 ? n34096 : n34105;
  assign n34107 = pi15 ? n33135 : n34106;
  assign n34108 = pi14 ? n34091 : n34107;
  assign n34109 = pi18 ? n880 : ~n6059;
  assign n34110 = pi17 ? n15845 : n34109;
  assign n34111 = pi16 ? n1214 : ~n34110;
  assign n34112 = pi18 ? n4722 : n350;
  assign n34113 = pi17 ? n32 : n34112;
  assign n34114 = pi16 ? n19652 : ~n34113;
  assign n34115 = pi15 ? n34111 : n34114;
  assign n34116 = pi15 ? n32153 : n31146;
  assign n34117 = pi14 ? n34115 : n34116;
  assign n34118 = pi13 ? n34108 : n34117;
  assign n34119 = pi12 ? n34078 : n34118;
  assign n34120 = pi11 ? n34053 : n34119;
  assign n34121 = pi10 ? n34005 : n34120;
  assign n34122 = pi09 ? n32 : n34121;
  assign n34123 = pi14 ? n22540 : n25086;
  assign n34124 = pi13 ? n33966 : n34123;
  assign n34125 = pi14 ? n22540 : n22541;
  assign n34126 = pi13 ? n22813 : n34125;
  assign n34127 = pi12 ? n34124 : n34126;
  assign n34128 = pi11 ? n34127 : n34004;
  assign n34129 = pi20 ? n321 : ~n1839;
  assign n34130 = pi19 ? n34129 : n32;
  assign n34131 = pi18 ? n32 : n34130;
  assign n34132 = pi17 ? n22435 : n34131;
  assign n34133 = pi16 ? n32 : n34132;
  assign n34134 = pi15 ? n32 : n34133;
  assign n34135 = pi20 ? n518 : ~n7013;
  assign n34136 = pi19 ? n34135 : n32;
  assign n34137 = pi18 ? n32 : n34136;
  assign n34138 = pi17 ? n15121 : n34137;
  assign n34139 = pi16 ? n32 : n34138;
  assign n34140 = pi15 ? n34139 : n34037;
  assign n34141 = pi14 ? n34134 : n34140;
  assign n34142 = pi19 ? n6339 : n32;
  assign n34143 = pi18 ? n20007 : ~n34142;
  assign n34144 = pi17 ? n32 : n34143;
  assign n34145 = pi16 ? n1135 : ~n34144;
  assign n34146 = pi16 ? n1135 : ~n2409;
  assign n34147 = pi15 ? n34145 : n34146;
  assign n34148 = pi14 ? n34147 : n34050;
  assign n34149 = pi13 ? n34141 : n34148;
  assign n34150 = pi12 ? n34022 : n34149;
  assign n34151 = pi18 ? n222 : n5749;
  assign n34152 = pi17 ? n32 : n34151;
  assign n34153 = pi16 ? n32 : n34152;
  assign n34154 = pi15 ? n34056 : n34153;
  assign n34155 = pi14 ? n34154 : n34066;
  assign n34156 = pi13 ? n34155 : n34077;
  assign n34157 = pi18 ? n940 : n34094;
  assign n34158 = pi17 ? n32 : n34157;
  assign n34159 = pi20 ? n342 : n175;
  assign n34160 = pi19 ? n34159 : n32;
  assign n34161 = pi18 ? n34098 : n34160;
  assign n34162 = pi19 ? n32 : ~n22702;
  assign n34163 = pi18 ? n34162 : n6059;
  assign n34164 = pi17 ? n34161 : n34163;
  assign n34165 = pi16 ? n34158 : n34164;
  assign n34166 = pi15 ? n33135 : n34165;
  assign n34167 = pi14 ? n34091 : n34166;
  assign n34168 = pi16 ? n19652 : ~n34110;
  assign n34169 = pi15 ? n34168 : n34114;
  assign n34170 = pi15 ? n32022 : n31056;
  assign n34171 = pi14 ? n34169 : n34170;
  assign n34172 = pi13 ? n34167 : n34171;
  assign n34173 = pi12 ? n34156 : n34172;
  assign n34174 = pi11 ? n34150 : n34173;
  assign n34175 = pi10 ? n34128 : n34174;
  assign n34176 = pi09 ? n32 : n34175;
  assign n34177 = pi08 ? n34122 : n34176;
  assign n34178 = pi07 ? n33965 : n34177;
  assign n34179 = pi06 ? n33735 : n34178;
  assign n34180 = pi05 ? n33231 : n34179;
  assign n34181 = pi14 ? n32 : n22925;
  assign n34182 = pi13 ? n34181 : n1109;
  assign n34183 = pi13 ? n22813 : n22540;
  assign n34184 = pi12 ? n34182 : n34183;
  assign n34185 = pi15 ? n22817 : n24919;
  assign n34186 = pi14 ? n22817 : n34185;
  assign n34187 = pi15 ? n25846 : n13629;
  assign n34188 = pi20 ? n246 : ~n321;
  assign n34189 = pi19 ? n34188 : n32;
  assign n34190 = pi18 ? n32 : n34189;
  assign n34191 = pi17 ? n32 : n34190;
  assign n34192 = pi16 ? n32 : n34191;
  assign n34193 = pi18 ? n4380 : n6059;
  assign n34194 = pi17 ? n32 : n34193;
  assign n34195 = pi16 ? n32 : n34194;
  assign n34196 = pi15 ? n34192 : n34195;
  assign n34197 = pi14 ? n34187 : n34196;
  assign n34198 = pi13 ? n34186 : n34197;
  assign n34199 = pi18 ? n863 : n22653;
  assign n34200 = pi17 ? n32 : n34199;
  assign n34201 = pi16 ? n32 : n34200;
  assign n34202 = pi15 ? n34201 : n21853;
  assign n34203 = pi14 ? n34202 : n21853;
  assign n34204 = pi18 ? n22865 : ~n22857;
  assign n34205 = pi17 ? n32 : n34204;
  assign n34206 = pi16 ? n32 : n34205;
  assign n34207 = pi18 ? n32 : n24942;
  assign n34208 = pi19 ? n32 : n5371;
  assign n34209 = pi18 ? n34208 : ~n323;
  assign n34210 = pi17 ? n34207 : n34209;
  assign n34211 = pi16 ? n32 : n34210;
  assign n34212 = pi15 ? n34206 : n34211;
  assign n34213 = pi19 ? n8383 : ~n32;
  assign n34214 = pi18 ? n32 : ~n34213;
  assign n34215 = pi17 ? n32 : n34214;
  assign n34216 = pi16 ? n32 : n34215;
  assign n34217 = pi15 ? n648 : n34216;
  assign n34218 = pi14 ? n34212 : n34217;
  assign n34219 = pi13 ? n34203 : n34218;
  assign n34220 = pi12 ? n34198 : n34219;
  assign n34221 = pi11 ? n34184 : n34220;
  assign n34222 = pi18 ? n4722 : n32;
  assign n34223 = pi17 ? n32 : n34222;
  assign n34224 = pi16 ? n32 : n34223;
  assign n34225 = pi18 ? n4380 : n23401;
  assign n34226 = pi17 ? n32 : n34225;
  assign n34227 = pi16 ? n32 : n34226;
  assign n34228 = pi15 ? n34224 : n34227;
  assign n34229 = pi19 ? n4391 : ~n32;
  assign n34230 = pi18 ? n940 : ~n34229;
  assign n34231 = pi17 ? n32 : n34230;
  assign n34232 = pi16 ? n32 : n34231;
  assign n34233 = pi15 ? n34232 : n32;
  assign n34234 = pi14 ? n34228 : n34233;
  assign n34235 = pi14 ? n33991 : n21217;
  assign n34236 = pi13 ? n34234 : n34235;
  assign n34237 = pi18 ? n20164 : n18474;
  assign n34238 = pi19 ? n9037 : n32;
  assign n34239 = pi18 ? n34238 : n32;
  assign n34240 = pi17 ? n34237 : n34239;
  assign n34241 = pi16 ? n32 : n34240;
  assign n34242 = pi19 ? n349 : ~n321;
  assign n34243 = pi19 ? n4342 : n11027;
  assign n34244 = pi18 ? n34242 : ~n34243;
  assign n34245 = pi18 ? n7038 : ~n32;
  assign n34246 = pi17 ? n34244 : ~n34245;
  assign n34247 = pi16 ? n15846 : n34246;
  assign n34248 = pi15 ? n34241 : n34247;
  assign n34249 = pi14 ? n32 : n34248;
  assign n34250 = pi19 ? n22864 : ~n32;
  assign n34251 = pi18 ? n32 : n34250;
  assign n34252 = pi17 ? n32 : n34251;
  assign n34253 = pi16 ? n34252 : ~n3769;
  assign n34254 = pi19 ? n28144 : n32;
  assign n34255 = pi18 ? n32 : ~n34254;
  assign n34256 = pi17 ? n32 : n34255;
  assign n34257 = pi16 ? n34256 : ~n3769;
  assign n34258 = pi15 ? n34253 : n34257;
  assign n34259 = pi15 ? n32828 : n12095;
  assign n34260 = pi14 ? n34258 : n34259;
  assign n34261 = pi13 ? n34249 : n34260;
  assign n34262 = pi12 ? n34236 : n34261;
  assign n34263 = pi18 ? n209 : n19194;
  assign n34264 = pi17 ? n32 : n34263;
  assign n34265 = pi16 ? n32 : n34264;
  assign n34266 = pi18 ? n268 : ~n34229;
  assign n34267 = pi17 ? n32 : n34266;
  assign n34268 = pi16 ? n32 : n34267;
  assign n34269 = pi15 ? n34265 : n34268;
  assign n34270 = pi18 ? n268 : n19194;
  assign n34271 = pi17 ? n32 : n34270;
  assign n34272 = pi16 ? n32 : n34271;
  assign n34273 = pi18 ? n4380 : ~n34229;
  assign n34274 = pi17 ? n32 : n34273;
  assign n34275 = pi16 ? n32 : n34274;
  assign n34276 = pi15 ? n34272 : n34275;
  assign n34277 = pi14 ? n34269 : n34276;
  assign n34278 = pi18 ? n32 : n30574;
  assign n34279 = pi17 ? n34278 : n12093;
  assign n34280 = pi16 ? n32 : n34279;
  assign n34281 = pi15 ? n12304 : n34280;
  assign n34282 = pi18 ? n20172 : n30574;
  assign n34283 = pi19 ? n322 : n349;
  assign n34284 = pi18 ? n34283 : ~n605;
  assign n34285 = pi17 ? n34282 : n34284;
  assign n34286 = pi16 ? n32 : n34285;
  assign n34287 = pi18 ? n20172 : n6118;
  assign n34288 = pi19 ? n322 : n343;
  assign n34289 = pi18 ? n34288 : ~n423;
  assign n34290 = pi17 ? n34287 : n34289;
  assign n34291 = pi16 ? n32 : n34290;
  assign n34292 = pi15 ? n34286 : n34291;
  assign n34293 = pi14 ? n34281 : n34292;
  assign n34294 = pi13 ? n34277 : n34293;
  assign n34295 = pi20 ? n321 : ~n357;
  assign n34296 = pi19 ? n7089 : ~n34295;
  assign n34297 = pi19 ? n5707 : n322;
  assign n34298 = pi18 ? n34296 : ~n34297;
  assign n34299 = pi18 ? n5749 : n532;
  assign n34300 = pi17 ? n34298 : ~n34299;
  assign n34301 = pi16 ? n32 : n34300;
  assign n34302 = pi19 ? n1612 : n247;
  assign n34303 = pi18 ? n8106 : n34302;
  assign n34304 = pi20 ? n207 : ~n6621;
  assign n34305 = pi19 ? n34304 : ~n3507;
  assign n34306 = pi18 ? n34305 : n532;
  assign n34307 = pi17 ? n34303 : ~n34306;
  assign n34308 = pi16 ? n32 : n34307;
  assign n34309 = pi15 ? n34301 : n34308;
  assign n34310 = pi18 ? n10078 : ~n350;
  assign n34311 = pi17 ? n32 : n34310;
  assign n34312 = pi16 ? n32 : n34311;
  assign n34313 = pi20 ? n7939 : ~n266;
  assign n34314 = pi20 ? n2358 : n207;
  assign n34315 = pi19 ? n34313 : n34314;
  assign n34316 = pi18 ? n276 : ~n34315;
  assign n34317 = pi17 ? n32 : n34316;
  assign n34318 = pi19 ? n207 : ~n1817;
  assign n34319 = pi20 ? n1817 : ~n207;
  assign n34320 = pi19 ? n34319 : ~n12899;
  assign n34321 = pi18 ? n34318 : ~n34320;
  assign n34322 = pi19 ? n247 : n4491;
  assign n34323 = pi18 ? n34322 : n6867;
  assign n34324 = pi17 ? n34321 : ~n34323;
  assign n34325 = pi16 ? n34317 : ~n34324;
  assign n34326 = pi15 ? n34312 : n34325;
  assign n34327 = pi14 ? n34309 : n34326;
  assign n34328 = pi18 ? n4380 : ~n4689;
  assign n34329 = pi17 ? n32 : n34328;
  assign n34330 = pi16 ? n1471 : ~n34329;
  assign n34331 = pi18 ? n17118 : n430;
  assign n34332 = pi17 ? n32 : n34331;
  assign n34333 = pi16 ? n1135 : ~n34332;
  assign n34334 = pi15 ? n34330 : n34333;
  assign n34335 = pi18 ? n32 : ~n19750;
  assign n34336 = pi17 ? n32 : n34335;
  assign n34337 = pi16 ? n1135 : ~n34336;
  assign n34338 = pi15 ? n31828 : n34337;
  assign n34339 = pi14 ? n34334 : n34338;
  assign n34340 = pi13 ? n34327 : n34339;
  assign n34341 = pi12 ? n34294 : n34340;
  assign n34342 = pi11 ? n34262 : n34341;
  assign n34343 = pi10 ? n34221 : n34342;
  assign n34344 = pi09 ? n32 : n34343;
  assign n34345 = pi14 ? n32 : n24913;
  assign n34346 = pi14 ? n1110 : n24275;
  assign n34347 = pi13 ? n34345 : n34346;
  assign n34348 = pi15 ? n24274 : n22923;
  assign n34349 = pi14 ? n34348 : n32;
  assign n34350 = pi15 ? n22540 : n22728;
  assign n34351 = pi14 ? n34350 : n22728;
  assign n34352 = pi13 ? n34349 : n34351;
  assign n34353 = pi12 ? n34347 : n34352;
  assign n34354 = pi19 ? n1053 : n32;
  assign n34355 = pi18 ? n32 : n34354;
  assign n34356 = pi17 ? n32 : n34355;
  assign n34357 = pi16 ? n32 : n34356;
  assign n34358 = pi15 ? n34357 : n13629;
  assign n34359 = pi14 ? n34358 : n34196;
  assign n34360 = pi13 ? n34186 : n34359;
  assign n34361 = pi15 ? n34201 : n27035;
  assign n34362 = pi14 ? n34361 : n21853;
  assign n34363 = pi15 ? n32 : n19628;
  assign n34364 = pi14 ? n34212 : n34363;
  assign n34365 = pi13 ? n34362 : n34364;
  assign n34366 = pi12 ? n34360 : n34365;
  assign n34367 = pi11 ? n34353 : n34366;
  assign n34368 = pi17 ? n34278 : n12089;
  assign n34369 = pi16 ? n32 : n34368;
  assign n34370 = pi15 ? n12304 : n34369;
  assign n34371 = pi14 ? n34370 : n34292;
  assign n34372 = pi13 ? n34277 : n34371;
  assign n34373 = pi18 ? n17118 : n2304;
  assign n34374 = pi17 ? n32 : n34373;
  assign n34375 = pi16 ? n1135 : ~n34374;
  assign n34376 = pi15 ? n34330 : n34375;
  assign n34377 = pi16 ? n1135 : ~n2306;
  assign n34378 = pi18 ? n32 : ~n19865;
  assign n34379 = pi17 ? n32 : n34378;
  assign n34380 = pi16 ? n1135 : ~n34379;
  assign n34381 = pi15 ? n34377 : n34380;
  assign n34382 = pi14 ? n34376 : n34381;
  assign n34383 = pi13 ? n34327 : n34382;
  assign n34384 = pi12 ? n34372 : n34383;
  assign n34385 = pi11 ? n34262 : n34384;
  assign n34386 = pi10 ? n34367 : n34385;
  assign n34387 = pi09 ? n32 : n34386;
  assign n34388 = pi08 ? n34344 : n34387;
  assign n34389 = pi15 ? n15665 : n24274;
  assign n34390 = pi14 ? n32 : n34389;
  assign n34391 = pi14 ? n24274 : n22923;
  assign n34392 = pi13 ? n34390 : n34391;
  assign n34393 = pi15 ? n32 : n22728;
  assign n34394 = pi15 ? n23011 : n15119;
  assign n34395 = pi14 ? n34393 : n34394;
  assign n34396 = pi13 ? n23089 : n34395;
  assign n34397 = pi12 ? n34392 : n34396;
  assign n34398 = pi15 ? n23011 : n22728;
  assign n34399 = pi15 ? n22728 : n25001;
  assign n34400 = pi14 ? n34398 : n34399;
  assign n34401 = pi19 ? n343 : ~n1105;
  assign n34402 = pi18 ? n32 : n34401;
  assign n34403 = pi17 ? n32 : n34402;
  assign n34404 = pi16 ? n32 : n34403;
  assign n34405 = pi15 ? n34404 : n13629;
  assign n34406 = pi14 ? n34405 : n22252;
  assign n34407 = pi13 ? n34400 : n34406;
  assign n34408 = pi15 ? n21853 : n32;
  assign n34409 = pi14 ? n22437 : n34408;
  assign n34410 = pi18 ? n940 : ~n22857;
  assign n34411 = pi17 ? n32 : n34410;
  assign n34412 = pi16 ? n32 : n34411;
  assign n34413 = pi20 ? n342 : ~n5854;
  assign n34414 = pi19 ? n32 : n34413;
  assign n34415 = pi18 ? n32 : n34414;
  assign n34416 = pi20 ? n246 : n518;
  assign n34417 = pi19 ? n18665 : n34416;
  assign n34418 = pi18 ? n34417 : ~n323;
  assign n34419 = pi17 ? n34415 : n34418;
  assign n34420 = pi16 ? n32 : n34419;
  assign n34421 = pi15 ? n34412 : n34420;
  assign n34422 = pi14 ? n34421 : n34363;
  assign n34423 = pi13 ? n34409 : n34422;
  assign n34424 = pi12 ? n34407 : n34423;
  assign n34425 = pi11 ? n34397 : n34424;
  assign n34426 = pi18 ? n32 : n24647;
  assign n34427 = pi18 ? n684 : n32;
  assign n34428 = pi17 ? n34426 : n34427;
  assign n34429 = pi16 ? n32 : n34428;
  assign n34430 = pi18 ? n4380 : n34189;
  assign n34431 = pi17 ? n32 : n34430;
  assign n34432 = pi16 ? n32 : n34431;
  assign n34433 = pi15 ? n34429 : n34432;
  assign n34434 = pi18 ? n32 : n18941;
  assign n34435 = pi17 ? n32 : n34434;
  assign n34436 = pi16 ? n32 : n34435;
  assign n34437 = pi15 ? n34232 : n34436;
  assign n34438 = pi14 ? n34433 : n34437;
  assign n34439 = pi14 ? n32 : n32128;
  assign n34440 = pi13 ? n34438 : n34439;
  assign n34441 = pi17 ? n3497 : n30107;
  assign n34442 = pi16 ? n32 : n34441;
  assign n34443 = pi15 ? n32 : n34442;
  assign n34444 = pi20 ? n1324 : ~n175;
  assign n34445 = pi19 ? n267 : ~n34444;
  assign n34446 = pi19 ? n175 : ~n16431;
  assign n34447 = pi18 ? n34445 : n34446;
  assign n34448 = pi19 ? n321 : n1757;
  assign n34449 = pi18 ? n34448 : n32;
  assign n34450 = pi17 ? n34447 : n34449;
  assign n34451 = pi16 ? n17120 : n34450;
  assign n34452 = pi18 ? n34242 : ~n4993;
  assign n34453 = pi19 ? n349 : ~n20555;
  assign n34454 = pi18 ? n34453 : ~n33239;
  assign n34455 = pi17 ? n34452 : n34454;
  assign n34456 = pi16 ? n32 : n34455;
  assign n34457 = pi15 ? n34451 : n34456;
  assign n34458 = pi14 ? n34443 : n34457;
  assign n34459 = pi18 ? n32 : n22865;
  assign n34460 = pi17 ? n32 : n34459;
  assign n34461 = pi16 ? n34460 : ~n2756;
  assign n34462 = pi16 ? n3061 : ~n2756;
  assign n34463 = pi15 ? n34461 : n34462;
  assign n34464 = pi15 ? n12083 : n32828;
  assign n34465 = pi14 ? n34463 : n34464;
  assign n34466 = pi13 ? n34458 : n34465;
  assign n34467 = pi12 ? n34440 : n34466;
  assign n34468 = pi19 ? n8220 : ~n32;
  assign n34469 = pi18 ? n32 : ~n34468;
  assign n34470 = pi17 ? n32 : n34469;
  assign n34471 = pi16 ? n32 : n34470;
  assign n34472 = pi15 ? n12297 : n34471;
  assign n34473 = pi20 ? n266 : n439;
  assign n34474 = pi19 ? n34473 : n32;
  assign n34475 = pi18 ? n32 : n34474;
  assign n34476 = pi17 ? n32 : n34475;
  assign n34477 = pi16 ? n32 : n34476;
  assign n34478 = pi18 ? n32 : ~n6063;
  assign n34479 = pi17 ? n32 : n34478;
  assign n34480 = pi16 ? n32 : n34479;
  assign n34481 = pi15 ? n34477 : n34480;
  assign n34482 = pi14 ? n34472 : n34481;
  assign n34483 = pi17 ? n16317 : n12298;
  assign n34484 = pi16 ? n32 : n34483;
  assign n34485 = pi19 ? n267 : n1757;
  assign n34486 = pi19 ? n9037 : ~n1490;
  assign n34487 = pi18 ? n34485 : n34486;
  assign n34488 = pi19 ? n21296 : ~n4342;
  assign n34489 = pi18 ? n34488 : ~n2413;
  assign n34490 = pi17 ? n34487 : n34489;
  assign n34491 = pi16 ? n32 : n34490;
  assign n34492 = pi15 ? n34484 : n34491;
  assign n34493 = pi19 ? n9007 : ~n22525;
  assign n34494 = pi19 ? n321 : ~n1490;
  assign n34495 = pi18 ? n34493 : n34494;
  assign n34496 = pi19 ? n6396 : ~n32;
  assign n34497 = pi18 ? n34496 : ~n605;
  assign n34498 = pi17 ? n34495 : n34497;
  assign n34499 = pi16 ? n32 : n34498;
  assign n34500 = pi19 ? n322 : n11879;
  assign n34501 = pi18 ? n20164 : n34500;
  assign n34502 = pi20 ? n7839 : n321;
  assign n34503 = pi19 ? n34502 : ~n32;
  assign n34504 = pi18 ? n34503 : ~n605;
  assign n34505 = pi17 ? n34501 : n34504;
  assign n34506 = pi16 ? n32 : n34505;
  assign n34507 = pi15 ? n34499 : n34506;
  assign n34508 = pi14 ? n34492 : n34507;
  assign n34509 = pi13 ? n34482 : n34508;
  assign n34510 = pi19 ? n1508 : ~n349;
  assign n34511 = pi18 ? n34510 : n13982;
  assign n34512 = pi18 ? n32535 : n605;
  assign n34513 = pi17 ? n34511 : ~n34512;
  assign n34514 = pi16 ? n32 : n34513;
  assign n34515 = pi15 ? n34514 : n11860;
  assign n34516 = pi17 ? n15832 : n30107;
  assign n34517 = pi16 ? n32 : n34516;
  assign n34518 = pi15 ? n32 : n34517;
  assign n34519 = pi14 ? n34515 : n34518;
  assign n34520 = pi16 ? n20208 : ~n31638;
  assign n34521 = pi15 ? n34520 : n32021;
  assign n34522 = pi18 ? n32 : n31385;
  assign n34523 = pi17 ? n32 : n34522;
  assign n34524 = pi16 ? n1135 : ~n34523;
  assign n34525 = pi18 ? n4380 : ~n248;
  assign n34526 = pi17 ? n32 : n34525;
  assign n34527 = pi16 ? n1135 : ~n34526;
  assign n34528 = pi15 ? n34524 : n34527;
  assign n34529 = pi14 ? n34521 : n34528;
  assign n34530 = pi13 ? n34519 : n34529;
  assign n34531 = pi12 ? n34509 : n34530;
  assign n34532 = pi11 ? n34467 : n34531;
  assign n34533 = pi10 ? n34425 : n34532;
  assign n34534 = pi09 ? n32 : n34533;
  assign n34535 = pi15 ? n15518 : n22923;
  assign n34536 = pi14 ? n32 : n34535;
  assign n34537 = pi15 ? n22923 : n15518;
  assign n34538 = pi14 ? n34537 : n23828;
  assign n34539 = pi13 ? n34536 : n34538;
  assign n34540 = pi14 ? n23828 : n32;
  assign n34541 = pi15 ? n32 : n23340;
  assign n34542 = pi14 ? n34541 : n15119;
  assign n34543 = pi13 ? n34540 : n34542;
  assign n34544 = pi12 ? n34539 : n34543;
  assign n34545 = pi15 ? n22817 : n22540;
  assign n34546 = pi14 ? n34545 : n34399;
  assign n34547 = pi13 ? n34546 : n34406;
  assign n34548 = pi12 ? n34547 : n34423;
  assign n34549 = pi11 ? n34544 : n34548;
  assign n34550 = pi18 ? n16847 : n2093;
  assign n34551 = pi17 ? n3497 : n34550;
  assign n34552 = pi16 ? n32 : n34551;
  assign n34553 = pi15 ? n21786 : n34552;
  assign n34554 = pi18 ? n34448 : n2093;
  assign n34555 = pi17 ? n34447 : n34554;
  assign n34556 = pi16 ? n17120 : n34555;
  assign n34557 = pi15 ? n34556 : n34456;
  assign n34558 = pi14 ? n34553 : n34557;
  assign n34559 = pi16 ? n34460 : ~n2518;
  assign n34560 = pi16 ? n3061 : ~n2518;
  assign n34561 = pi15 ? n34559 : n34560;
  assign n34562 = pi15 ? n12289 : n32828;
  assign n34563 = pi14 ? n34561 : n34562;
  assign n34564 = pi13 ? n34558 : n34563;
  assign n34565 = pi12 ? n34440 : n34564;
  assign n34566 = pi17 ? n16317 : n12295;
  assign n34567 = pi16 ? n32 : n34566;
  assign n34568 = pi18 ? n34488 : ~n605;
  assign n34569 = pi17 ? n34487 : n34568;
  assign n34570 = pi16 ? n32 : n34569;
  assign n34571 = pi15 ? n34567 : n34570;
  assign n34572 = pi14 ? n34571 : n34507;
  assign n34573 = pi13 ? n34482 : n34572;
  assign n34574 = pi18 ? n32535 : n2413;
  assign n34575 = pi17 ? n34511 : ~n34574;
  assign n34576 = pi16 ? n32 : n34575;
  assign n34577 = pi18 ? n684 : ~n2413;
  assign n34578 = pi17 ? n32 : n34577;
  assign n34579 = pi16 ? n32 : n34578;
  assign n34580 = pi15 ? n34576 : n34579;
  assign n34581 = pi14 ? n34580 : n34518;
  assign n34582 = pi16 ? n1233 : ~n34523;
  assign n34583 = pi16 ? n1233 : ~n34526;
  assign n34584 = pi15 ? n34582 : n34583;
  assign n34585 = pi14 ? n34521 : n34584;
  assign n34586 = pi13 ? n34581 : n34585;
  assign n34587 = pi12 ? n34573 : n34586;
  assign n34588 = pi11 ? n34565 : n34587;
  assign n34589 = pi10 ? n34549 : n34588;
  assign n34590 = pi09 ? n32 : n34589;
  assign n34591 = pi08 ? n34534 : n34590;
  assign n34592 = pi07 ? n34388 : n34591;
  assign n34593 = pi14 ? n32 : n24397;
  assign n34594 = pi13 ? n34593 : n23160;
  assign n34595 = pi14 ? n22923 : n34537;
  assign n34596 = pi13 ? n23256 : n34595;
  assign n34597 = pi12 ? n34594 : n34596;
  assign n34598 = pi19 ? n23193 : ~n617;
  assign n34599 = pi18 ? n32 : n34598;
  assign n34600 = pi17 ? n32 : n34599;
  assign n34601 = pi16 ? n32 : n34600;
  assign n34602 = pi15 ? n22923 : n34601;
  assign n34603 = pi19 ? n4982 : ~n617;
  assign n34604 = pi18 ? n32 : n34603;
  assign n34605 = pi17 ? n32 : n34604;
  assign n34606 = pi16 ? n32 : n34605;
  assign n34607 = pi19 ? n18396 : ~n617;
  assign n34608 = pi18 ? n32 : n34607;
  assign n34609 = pi17 ? n32 : n34608;
  assign n34610 = pi16 ? n32 : n34609;
  assign n34611 = pi15 ? n34606 : n34610;
  assign n34612 = pi14 ? n34602 : n34611;
  assign n34613 = pi19 ? n343 : ~n617;
  assign n34614 = pi18 ? n32 : n34613;
  assign n34615 = pi17 ? n32 : n34614;
  assign n34616 = pi16 ? n32 : n34615;
  assign n34617 = pi15 ? n34616 : n22817;
  assign n34618 = pi14 ? n34617 : n22817;
  assign n34619 = pi13 ? n34612 : n34618;
  assign n34620 = pi14 ? n22817 : n32;
  assign n34621 = pi19 ? n23944 : ~n32;
  assign n34622 = pi18 ? n16847 : ~n34621;
  assign n34623 = pi17 ? n32 : n34622;
  assign n34624 = pi16 ? n32 : n34623;
  assign n34625 = pi15 ? n22437 : n34624;
  assign n34626 = pi14 ? n15127 : n34625;
  assign n34627 = pi13 ? n34620 : n34626;
  assign n34628 = pi12 ? n34619 : n34627;
  assign n34629 = pi11 ? n34597 : n34628;
  assign n34630 = pi18 ? n13182 : n595;
  assign n34631 = pi17 ? n2726 : ~n34630;
  assign n34632 = pi16 ? n32 : n34631;
  assign n34633 = pi19 ? n1757 : n531;
  assign n34634 = pi18 ? n34633 : ~n508;
  assign n34635 = pi17 ? n34459 : n34634;
  assign n34636 = pi16 ? n32 : n34635;
  assign n34637 = pi15 ? n34632 : n34636;
  assign n34638 = pi18 ? n1509 : ~n595;
  assign n34639 = pi17 ? n32 : n34638;
  assign n34640 = pi16 ? n32 : n34639;
  assign n34641 = pi18 ? n858 : n5502;
  assign n34642 = pi17 ? n32 : n34641;
  assign n34643 = pi16 ? n32 : n34642;
  assign n34644 = pi15 ? n34640 : n34643;
  assign n34645 = pi14 ? n34637 : n34644;
  assign n34646 = pi13 ? n34645 : n32;
  assign n34647 = pi20 ? n518 : n266;
  assign n34648 = pi19 ? n32 : n34647;
  assign n34649 = pi18 ? n32 : n34648;
  assign n34650 = pi17 ? n34649 : n17901;
  assign n34651 = pi16 ? n32 : n34650;
  assign n34652 = pi15 ? n32 : n34651;
  assign n34653 = pi19 ? n3692 : n9007;
  assign n34654 = pi18 ? n34653 : ~n8908;
  assign n34655 = pi17 ? n1215 : ~n34654;
  assign n34656 = pi16 ? n32 : n34655;
  assign n34657 = pi17 ? n1028 : ~n2517;
  assign n34658 = pi16 ? n32 : n34657;
  assign n34659 = pi15 ? n34656 : n34658;
  assign n34660 = pi14 ? n34652 : n34659;
  assign n34661 = pi17 ? n18482 : n2517;
  assign n34662 = pi16 ? n32 : ~n34661;
  assign n34663 = pi17 ? n1215 : ~n2517;
  assign n34664 = pi16 ? n32 : n34663;
  assign n34665 = pi15 ? n34662 : n34664;
  assign n34666 = pi18 ? n532 : ~n520;
  assign n34667 = pi17 ? n1978 : n34666;
  assign n34668 = pi16 ? n32 : n34667;
  assign n34669 = pi19 ? n531 : ~n1464;
  assign n34670 = pi18 ? n34669 : ~n323;
  assign n34671 = pi17 ? n1978 : n34670;
  assign n34672 = pi16 ? n32 : n34671;
  assign n34673 = pi15 ? n34668 : n34672;
  assign n34674 = pi14 ? n34665 : n34673;
  assign n34675 = pi13 ? n34660 : n34674;
  assign n34676 = pi12 ? n34646 : n34675;
  assign n34677 = pi18 ? n880 : ~n2291;
  assign n34678 = pi17 ? n32 : n34677;
  assign n34679 = pi16 ? n32 : n34678;
  assign n34680 = pi18 ? n863 : ~n23397;
  assign n34681 = pi17 ? n32 : n34680;
  assign n34682 = pi16 ? n32 : n34681;
  assign n34683 = pi15 ? n34679 : n34682;
  assign n34684 = pi19 ? n14877 : ~n32;
  assign n34685 = pi18 ? n863 : ~n34684;
  assign n34686 = pi17 ? n32 : n34685;
  assign n34687 = pi16 ? n32 : n34686;
  assign n34688 = pi15 ? n34687 : n12777;
  assign n34689 = pi14 ? n34683 : n34688;
  assign n34690 = pi19 ? n1464 : n4964;
  assign n34691 = pi18 ? n34690 : ~n32;
  assign n34692 = pi18 ? n248 : n605;
  assign n34693 = pi17 ? n34691 : ~n34692;
  assign n34694 = pi16 ? n32 : n34693;
  assign n34695 = pi15 ? n12777 : n34694;
  assign n34696 = pi19 ? n32090 : n32;
  assign n34697 = pi18 ? n34696 : n605;
  assign n34698 = pi17 ? n1978 : ~n34697;
  assign n34699 = pi16 ? n32 : n34698;
  assign n34700 = pi18 ? n6063 : ~n605;
  assign n34701 = pi17 ? n1978 : n34700;
  assign n34702 = pi16 ? n32 : n34701;
  assign n34703 = pi15 ? n34699 : n34702;
  assign n34704 = pi14 ? n34695 : n34703;
  assign n34705 = pi13 ? n34689 : n34704;
  assign n34706 = pi18 ? n237 : n33312;
  assign n34707 = pi17 ? n34706 : ~n2119;
  assign n34708 = pi16 ? n32 : n34707;
  assign n34709 = pi15 ? n34708 : n20831;
  assign n34710 = pi19 ? n267 : n32733;
  assign n34711 = pi18 ? n34710 : n702;
  assign n34712 = pi19 ? n5004 : ~n507;
  assign n34713 = pi18 ? n34712 : n248;
  assign n34714 = pi17 ? n34711 : n34713;
  assign n34715 = pi16 ? n32 : n34714;
  assign n34716 = pi15 ? n32 : n34715;
  assign n34717 = pi14 ? n34709 : n34716;
  assign n34718 = pi19 ? n1464 : n247;
  assign n34719 = pi18 ? n34718 : n8203;
  assign n34720 = pi19 ? n5748 : n18478;
  assign n34721 = pi18 ? n34720 : n177;
  assign n34722 = pi17 ? n34719 : n34721;
  assign n34723 = pi16 ? n3438 : n34722;
  assign n34724 = pi19 ? n6042 : ~n32;
  assign n34725 = pi18 ? n863 : n34724;
  assign n34726 = pi17 ? n32 : n34725;
  assign n34727 = pi16 ? n1214 : ~n34726;
  assign n34728 = pi15 ? n34723 : n34727;
  assign n34729 = pi18 ? n863 : n31959;
  assign n34730 = pi17 ? n32 : n34729;
  assign n34731 = pi16 ? n1214 : ~n34730;
  assign n34732 = pi18 ? n863 : ~n4671;
  assign n34733 = pi17 ? n32 : n34732;
  assign n34734 = pi16 ? n1214 : ~n34733;
  assign n34735 = pi15 ? n34731 : n34734;
  assign n34736 = pi14 ? n34728 : n34735;
  assign n34737 = pi13 ? n34717 : n34736;
  assign n34738 = pi12 ? n34705 : n34737;
  assign n34739 = pi11 ? n34676 : n34738;
  assign n34740 = pi10 ? n34629 : n34739;
  assign n34741 = pi09 ? n32 : n34740;
  assign n34742 = pi15 ? n23160 : n15655;
  assign n34743 = pi14 ? n34742 : n23250;
  assign n34744 = pi13 ? n23161 : n34743;
  assign n34745 = pi14 ? n34537 : n15518;
  assign n34746 = pi13 ? n23426 : n34745;
  assign n34747 = pi12 ? n34744 : n34746;
  assign n34748 = pi15 ? n24274 : n34601;
  assign n34749 = pi14 ? n34748 : n34611;
  assign n34750 = pi13 ? n34749 : n34618;
  assign n34751 = pi14 ? n34398 : n32;
  assign n34752 = pi13 ? n34751 : n34626;
  assign n34753 = pi12 ? n34750 : n34752;
  assign n34754 = pi11 ? n34747 : n34753;
  assign n34755 = pi18 ? n34653 : ~n13341;
  assign n34756 = pi17 ? n1215 : ~n34755;
  assign n34757 = pi16 ? n32 : n34756;
  assign n34758 = pi17 ? n1028 : ~n2748;
  assign n34759 = pi16 ? n32 : n34758;
  assign n34760 = pi15 ? n34757 : n34759;
  assign n34761 = pi14 ? n34652 : n34760;
  assign n34762 = pi17 ? n18482 : n2748;
  assign n34763 = pi16 ? n32 : ~n34762;
  assign n34764 = pi17 ? n1215 : ~n2748;
  assign n34765 = pi16 ? n32 : n34764;
  assign n34766 = pi15 ? n34763 : n34765;
  assign n34767 = pi18 ? n532 : ~n2747;
  assign n34768 = pi17 ? n1978 : n34767;
  assign n34769 = pi16 ? n32 : n34768;
  assign n34770 = pi18 ? n34669 : ~n520;
  assign n34771 = pi17 ? n1978 : n34770;
  assign n34772 = pi16 ? n32 : n34771;
  assign n34773 = pi15 ? n34769 : n34772;
  assign n34774 = pi14 ? n34766 : n34773;
  assign n34775 = pi13 ? n34761 : n34774;
  assign n34776 = pi12 ? n34646 : n34775;
  assign n34777 = pi15 ? n32219 : n34687;
  assign n34778 = pi18 ? n863 : ~n2291;
  assign n34779 = pi17 ? n32 : n34778;
  assign n34780 = pi16 ? n32 : n34779;
  assign n34781 = pi15 ? n34687 : n34780;
  assign n34782 = pi14 ? n34777 : n34781;
  assign n34783 = pi18 ? n248 : n32919;
  assign n34784 = pi17 ? n34691 : ~n34783;
  assign n34785 = pi16 ? n32 : n34784;
  assign n34786 = pi15 ? n34780 : n34785;
  assign n34787 = pi14 ? n34786 : n34703;
  assign n34788 = pi13 ? n34782 : n34787;
  assign n34789 = pi15 ? n34708 : n32;
  assign n34790 = pi14 ? n34789 : n34716;
  assign n34791 = pi13 ? n34790 : n34736;
  assign n34792 = pi12 ? n34788 : n34791;
  assign n34793 = pi11 ? n34776 : n34792;
  assign n34794 = pi10 ? n34754 : n34793;
  assign n34795 = pi09 ? n32 : n34794;
  assign n34796 = pi08 ? n34741 : n34795;
  assign n34797 = pi14 ? n23250 : n15836;
  assign n34798 = pi13 ? n23251 : n34797;
  assign n34799 = pi15 ? n15518 : n23484;
  assign n34800 = pi14 ? n23828 : n34799;
  assign n34801 = pi13 ? n23327 : n34800;
  assign n34802 = pi12 ? n34798 : n34801;
  assign n34803 = pi19 ? n462 : ~n2614;
  assign n34804 = pi18 ? n32 : n34803;
  assign n34805 = pi17 ? n32 : n34804;
  assign n34806 = pi16 ? n32 : n34805;
  assign n34807 = pi19 ? n221 : ~n2614;
  assign n34808 = pi18 ? n32 : n34807;
  assign n34809 = pi17 ? n32 : n34808;
  assign n34810 = pi16 ? n32 : n34809;
  assign n34811 = pi15 ? n34806 : n34810;
  assign n34812 = pi19 ? n4982 : ~n2614;
  assign n34813 = pi18 ? n32 : n34812;
  assign n34814 = pi17 ? n32 : n34813;
  assign n34815 = pi16 ? n32 : n34814;
  assign n34816 = pi19 ? n4670 : n15661;
  assign n34817 = pi18 ? n32 : n34816;
  assign n34818 = pi17 ? n32 : n34817;
  assign n34819 = pi16 ? n32 : n34818;
  assign n34820 = pi15 ? n34815 : n34819;
  assign n34821 = pi14 ? n34811 : n34820;
  assign n34822 = pi14 ? n34617 : n22540;
  assign n34823 = pi13 ? n34821 : n34822;
  assign n34824 = pi14 ? n23264 : n32;
  assign n34825 = pi19 ? n19151 : n4982;
  assign n34826 = pi18 ? n34825 : ~n595;
  assign n34827 = pi17 ? n17463 : n34826;
  assign n34828 = pi16 ? n32 : n34827;
  assign n34829 = pi15 ? n22437 : n34828;
  assign n34830 = pi14 ? n15127 : n34829;
  assign n34831 = pi13 ? n34824 : n34830;
  assign n34832 = pi12 ? n34823 : n34831;
  assign n34833 = pi11 ? n34802 : n34832;
  assign n34834 = pi19 ? n5356 : ~n343;
  assign n34835 = pi18 ? n34834 : n595;
  assign n34836 = pi17 ? n2726 : ~n34835;
  assign n34837 = pi16 ? n32 : n34836;
  assign n34838 = pi17 ? n2959 : n34634;
  assign n34839 = pi16 ? n32 : n34838;
  assign n34840 = pi15 ? n34837 : n34839;
  assign n34841 = pi21 ? n206 : ~n9326;
  assign n34842 = pi20 ? n32 : n34841;
  assign n34843 = pi19 ? n34842 : n32;
  assign n34844 = pi18 ? n32 : n34843;
  assign n34845 = pi17 ? n32 : n34844;
  assign n34846 = pi16 ? n32 : n34845;
  assign n34847 = pi15 ? n13040 : n34846;
  assign n34848 = pi14 ? n34840 : n34847;
  assign n34849 = pi19 ? n5675 : n32;
  assign n34850 = pi18 ? n32 : n34849;
  assign n34851 = pi17 ? n32 : n34850;
  assign n34852 = pi16 ? n32 : n34851;
  assign n34853 = pi15 ? n34852 : n21853;
  assign n34854 = pi14 ? n34853 : n32;
  assign n34855 = pi13 ? n34848 : n34854;
  assign n34856 = pi18 ? n4127 : n32;
  assign n34857 = pi17 ? n17346 : n34856;
  assign n34858 = pi16 ? n32 : n34857;
  assign n34859 = pi15 ? n32 : n34858;
  assign n34860 = pi19 ? n13667 : n23193;
  assign n34861 = pi18 ? n34860 : n520;
  assign n34862 = pi17 ? n1215 : ~n34861;
  assign n34863 = pi16 ? n32 : n34862;
  assign n34864 = pi17 ? n2355 : ~n2517;
  assign n34865 = pi16 ? n32 : n34864;
  assign n34866 = pi15 ? n34863 : n34865;
  assign n34867 = pi14 ? n34859 : n34866;
  assign n34868 = pi17 ? n1227 : ~n2517;
  assign n34869 = pi16 ? n32 : n34868;
  assign n34870 = pi15 ? n34869 : n34765;
  assign n34871 = pi19 ? n531 : ~n208;
  assign n34872 = pi18 ? n34871 : ~n24036;
  assign n34873 = pi17 ? n1978 : n34872;
  assign n34874 = pi16 ? n32 : n34873;
  assign n34875 = pi15 ? n34769 : n34874;
  assign n34876 = pi14 ? n34870 : n34875;
  assign n34877 = pi13 ? n34867 : n34876;
  assign n34878 = pi12 ? n34855 : n34877;
  assign n34879 = pi19 ? n14861 : ~n32;
  assign n34880 = pi18 ? n32 : ~n34879;
  assign n34881 = pi17 ? n32 : n34880;
  assign n34882 = pi16 ? n32 : n34881;
  assign n34883 = pi15 ? n32828 : n34882;
  assign n34884 = pi15 ? n34882 : n13052;
  assign n34885 = pi14 ? n34883 : n34884;
  assign n34886 = pi18 ? n16847 : ~n32;
  assign n34887 = pi18 ? n13372 : n2291;
  assign n34888 = pi17 ? n34886 : ~n34887;
  assign n34889 = pi16 ? n32 : n34888;
  assign n34890 = pi15 ? n34780 : n34889;
  assign n34891 = pi18 ? n6767 : ~n32;
  assign n34892 = pi17 ? n34891 : ~n34887;
  assign n34893 = pi16 ? n32 : n34892;
  assign n34894 = pi18 ? n22705 : ~n2291;
  assign n34895 = pi17 ? n1966 : n34894;
  assign n34896 = pi16 ? n32 : n34895;
  assign n34897 = pi15 ? n34893 : n34896;
  assign n34898 = pi14 ? n34890 : n34897;
  assign n34899 = pi13 ? n34885 : n34898;
  assign n34900 = pi18 ? n32 : n32919;
  assign n34901 = pi17 ? n34706 : ~n34900;
  assign n34902 = pi16 ? n16983 : n34901;
  assign n34903 = pi15 ? n34902 : n32;
  assign n34904 = pi19 ? n28853 : n22185;
  assign n34905 = pi19 ? n266 : ~n32;
  assign n34906 = pi18 ? n34904 : n34905;
  assign n34907 = pi20 ? n501 : ~n342;
  assign n34908 = pi19 ? n34907 : ~n594;
  assign n34909 = pi18 ? n34908 : n32;
  assign n34910 = pi17 ? n34906 : n34909;
  assign n34911 = pi16 ? n17038 : n34910;
  assign n34912 = pi15 ? n32 : n34911;
  assign n34913 = pi14 ? n34903 : n34912;
  assign n34914 = pi18 ? n32 : n28927;
  assign n34915 = pi17 ? n32 : n34914;
  assign n34916 = pi20 ? n274 : n17652;
  assign n34917 = pi20 ? n17652 : ~n17669;
  assign n34918 = pi19 ? n34916 : n34917;
  assign n34919 = pi19 ? n266 : n28041;
  assign n34920 = pi18 ? n34918 : n34919;
  assign n34921 = pi20 ? n4279 : ~n342;
  assign n34922 = pi19 ? n34921 : n13323;
  assign n34923 = pi18 ? n34922 : n4671;
  assign n34924 = pi17 ? n34920 : n34923;
  assign n34925 = pi16 ? n34915 : n34924;
  assign n34926 = pi18 ? n863 : n23073;
  assign n34927 = pi17 ? n32 : n34926;
  assign n34928 = pi16 ? n1135 : ~n34927;
  assign n34929 = pi15 ? n34925 : n34928;
  assign n34930 = pi16 ? n1135 : ~n34730;
  assign n34931 = pi15 ? n34930 : n28947;
  assign n34932 = pi14 ? n34929 : n34931;
  assign n34933 = pi13 ? n34913 : n34932;
  assign n34934 = pi12 ? n34899 : n34933;
  assign n34935 = pi11 ? n34878 : n34934;
  assign n34936 = pi10 ? n34833 : n34935;
  assign n34937 = pi09 ? n32 : n34936;
  assign n34938 = pi14 ? n32 : n15836;
  assign n34939 = pi15 ? n15836 : n23631;
  assign n34940 = pi14 ? n34939 : n16108;
  assign n34941 = pi13 ? n34938 : n34940;
  assign n34942 = pi15 ? n23250 : n15836;
  assign n34943 = pi14 ? n23743 : n34942;
  assign n34944 = pi14 ? n23485 : n23250;
  assign n34945 = pi13 ? n34943 : n34944;
  assign n34946 = pi12 ? n34941 : n34945;
  assign n34947 = pi19 ? n462 : ~n617;
  assign n34948 = pi18 ? n32 : n34947;
  assign n34949 = pi17 ? n32 : n34948;
  assign n34950 = pi16 ? n32 : n34949;
  assign n34951 = pi19 ? n221 : ~n617;
  assign n34952 = pi18 ? n32 : n34951;
  assign n34953 = pi17 ? n32 : n34952;
  assign n34954 = pi16 ? n32 : n34953;
  assign n34955 = pi15 ? n34950 : n34954;
  assign n34956 = pi19 ? n4670 : ~n2614;
  assign n34957 = pi18 ? n32 : n34956;
  assign n34958 = pi17 ? n32 : n34957;
  assign n34959 = pi16 ? n32 : n34958;
  assign n34960 = pi15 ? n34815 : n34959;
  assign n34961 = pi14 ? n34955 : n34960;
  assign n34962 = pi13 ? n34961 : n34822;
  assign n34963 = pi12 ? n34962 : n34831;
  assign n34964 = pi11 ? n34946 : n34963;
  assign n34965 = pi15 ? n13040 : n14389;
  assign n34966 = pi14 ? n34840 : n34965;
  assign n34967 = pi15 ? n34852 : n14790;
  assign n34968 = pi14 ? n34967 : n32;
  assign n34969 = pi13 ? n34966 : n34968;
  assign n34970 = pi18 ? n4127 : n645;
  assign n34971 = pi17 ? n17346 : n34970;
  assign n34972 = pi16 ? n32 : n34971;
  assign n34973 = pi15 ? n648 : n34972;
  assign n34974 = pi18 ? n34860 : n508;
  assign n34975 = pi17 ? n1215 : ~n34974;
  assign n34976 = pi16 ? n32 : n34975;
  assign n34977 = pi15 ? n34976 : n5843;
  assign n34978 = pi14 ? n34973 : n34977;
  assign n34979 = pi17 ? n1227 : ~n2512;
  assign n34980 = pi16 ? n32 : n34979;
  assign n34981 = pi17 ? n1215 : ~n2512;
  assign n34982 = pi16 ? n32 : n34981;
  assign n34983 = pi15 ? n34980 : n34982;
  assign n34984 = pi18 ? n34871 : ~n323;
  assign n34985 = pi17 ? n1978 : n34984;
  assign n34986 = pi16 ? n32 : n34985;
  assign n34987 = pi15 ? n34668 : n34986;
  assign n34988 = pi14 ? n34983 : n34987;
  assign n34989 = pi13 ? n34978 : n34988;
  assign n34990 = pi12 ? n34969 : n34989;
  assign n34991 = pi18 ? n32 : ~n28193;
  assign n34992 = pi17 ? n32 : n34991;
  assign n34993 = pi16 ? n32 : n34992;
  assign n34994 = pi15 ? n32828 : n34993;
  assign n34995 = pi15 ? n34993 : n23892;
  assign n34996 = pi14 ? n34994 : n34995;
  assign n34997 = pi18 ? n13372 : n797;
  assign n34998 = pi17 ? n34886 : ~n34997;
  assign n34999 = pi16 ? n32 : n34998;
  assign n35000 = pi15 ? n12777 : n34999;
  assign n35001 = pi18 ? n22705 : ~n797;
  assign n35002 = pi17 ? n1966 : n35001;
  assign n35003 = pi16 ? n32 : n35002;
  assign n35004 = pi15 ? n34893 : n35003;
  assign n35005 = pi14 ? n35000 : n35004;
  assign n35006 = pi13 ? n34996 : n35005;
  assign n35007 = pi16 ? n1233 : ~n34730;
  assign n35008 = pi15 ? n35007 : n30025;
  assign n35009 = pi14 ? n34929 : n35008;
  assign n35010 = pi13 ? n34913 : n35009;
  assign n35011 = pi12 ? n35006 : n35010;
  assign n35012 = pi11 ? n34990 : n35011;
  assign n35013 = pi10 ? n34964 : n35012;
  assign n35014 = pi09 ? n32 : n35013;
  assign n35015 = pi08 ? n34937 : n35014;
  assign n35016 = pi07 ? n34796 : n35015;
  assign n35017 = pi06 ? n34592 : n35016;
  assign n35018 = pi14 ? n23623 : n16108;
  assign n35019 = pi13 ? n35018 : n16108;
  assign n35020 = pi19 ? n2359 : ~n1941;
  assign n35021 = pi18 ? n32 : n35020;
  assign n35022 = pi17 ? n32 : n35021;
  assign n35023 = pi16 ? n32 : n35022;
  assign n35024 = pi15 ? n23250 : n35023;
  assign n35025 = pi14 ? n23484 : n35024;
  assign n35026 = pi13 ? n23423 : n35025;
  assign n35027 = pi12 ? n35019 : n35026;
  assign n35028 = pi18 ? n32 : n6405;
  assign n35029 = pi17 ? n32 : n35028;
  assign n35030 = pi16 ? n32 : n35029;
  assign n35031 = pi19 ? n221 : ~n236;
  assign n35032 = pi18 ? n32 : n35031;
  assign n35033 = pi17 ? n32 : n35032;
  assign n35034 = pi16 ? n32 : n35033;
  assign n35035 = pi15 ? n35030 : n35034;
  assign n35036 = pi18 ? n32 : n28667;
  assign n35037 = pi17 ? n32 : n35036;
  assign n35038 = pi16 ? n32 : n35037;
  assign n35039 = pi15 ? n23250 : n35038;
  assign n35040 = pi14 ? n35035 : n35039;
  assign n35041 = pi15 ? n25790 : n22817;
  assign n35042 = pi14 ? n35041 : n22540;
  assign n35043 = pi13 ? n35040 : n35042;
  assign n35044 = pi15 ? n15119 : n23340;
  assign n35045 = pi14 ? n35044 : n22540;
  assign n35046 = pi19 ? n21349 : n5004;
  assign n35047 = pi18 ? n35046 : n702;
  assign n35048 = pi17 ? n863 : ~n35047;
  assign n35049 = pi16 ? n32 : n35048;
  assign n35050 = pi18 ? n20020 : n702;
  assign n35051 = pi17 ? n1978 : ~n35050;
  assign n35052 = pi16 ? n32 : n35051;
  assign n35053 = pi15 ? n35049 : n35052;
  assign n35054 = pi14 ? n1110 : n35053;
  assign n35055 = pi13 ? n35045 : n35054;
  assign n35056 = pi12 ? n35043 : n35055;
  assign n35057 = pi11 ? n35027 : n35056;
  assign n35058 = pi20 ? n1385 : n1817;
  assign n35059 = pi19 ? n6158 : n35058;
  assign n35060 = pi18 ? n863 : ~n35059;
  assign n35061 = pi18 ? n23440 : n702;
  assign n35062 = pi17 ? n35060 : ~n35061;
  assign n35063 = pi16 ? n32 : n35062;
  assign n35064 = pi19 ? n17766 : ~n15405;
  assign n35065 = pi18 ? n35064 : ~n508;
  assign n35066 = pi17 ? n3164 : n35065;
  assign n35067 = pi16 ? n32 : n35066;
  assign n35068 = pi15 ? n35063 : n35067;
  assign n35069 = pi18 ? n12135 : n22857;
  assign n35070 = pi17 ? n32 : ~n35069;
  assign n35071 = pi16 ? n32 : n35070;
  assign n35072 = pi15 ? n35071 : n19531;
  assign n35073 = pi14 ? n35068 : n35072;
  assign n35074 = pi15 ? n22437 : n21928;
  assign n35075 = pi14 ? n35074 : n32;
  assign n35076 = pi13 ? n35073 : n35075;
  assign n35077 = pi19 ? n8818 : ~n322;
  assign n35078 = pi18 ? n35077 : n2627;
  assign n35079 = pi17 ? n3292 : ~n35078;
  assign n35080 = pi16 ? n32 : n35079;
  assign n35081 = pi15 ? n32 : n35080;
  assign n35082 = pi19 ? n32 : n22652;
  assign n35083 = pi18 ? n35082 : n32563;
  assign n35084 = pi18 ? n14153 : ~n22752;
  assign n35085 = pi17 ? n35083 : ~n35084;
  assign n35086 = pi16 ? n32 : n35085;
  assign n35087 = pi19 ? n32 : n24349;
  assign n35088 = pi18 ? n35087 : ~n32;
  assign n35089 = pi17 ? n35088 : ~n2628;
  assign n35090 = pi16 ? n32 : n35089;
  assign n35091 = pi15 ? n35086 : n35090;
  assign n35092 = pi14 ? n35081 : n35091;
  assign n35093 = pi18 ? n1758 : ~n32;
  assign n35094 = pi17 ? n35093 : ~n2628;
  assign n35095 = pi16 ? n32 : n35094;
  assign n35096 = pi17 ? n2519 : ~n2628;
  assign n35097 = pi16 ? n32 : n35096;
  assign n35098 = pi15 ? n35095 : n35097;
  assign n35099 = pi19 ? n15751 : n32;
  assign n35100 = pi18 ? n4983 : ~n35099;
  assign n35101 = pi17 ? n8859 : ~n35100;
  assign n35102 = pi16 ? n32 : n35101;
  assign n35103 = pi19 ? n531 : n4342;
  assign n35104 = pi18 ? n35103 : n520;
  assign n35105 = pi17 ? n3067 : ~n35104;
  assign n35106 = pi16 ? n32 : n35105;
  assign n35107 = pi15 ? n35102 : n35106;
  assign n35108 = pi14 ? n35098 : n35107;
  assign n35109 = pi13 ? n35092 : n35108;
  assign n35110 = pi12 ? n35076 : n35109;
  assign n35111 = pi19 ? n6800 : n32;
  assign n35112 = pi18 ? n32 : n35111;
  assign n35113 = pi17 ? n32 : n35112;
  assign n35114 = pi16 ? n32 : n35113;
  assign n35115 = pi15 ? n23892 : n35114;
  assign n35116 = pi20 ? n259 : ~n321;
  assign n35117 = pi19 ? n35116 : n32;
  assign n35118 = pi18 ? n32 : n35117;
  assign n35119 = pi17 ? n32 : n35118;
  assign n35120 = pi16 ? n32 : n35119;
  assign n35121 = pi18 ? n936 : ~n323;
  assign n35122 = pi17 ? n32 : n35121;
  assign n35123 = pi16 ? n32 : n35122;
  assign n35124 = pi15 ? n35120 : n35123;
  assign n35125 = pi14 ? n35115 : n35124;
  assign n35126 = pi18 ? n940 : ~n323;
  assign n35127 = pi17 ? n32 : n35126;
  assign n35128 = pi16 ? n32 : n35127;
  assign n35129 = pi19 ? n507 : n343;
  assign n35130 = pi18 ? n32 : n35129;
  assign n35131 = pi19 ? n5694 : ~n343;
  assign n35132 = pi18 ? n35131 : n323;
  assign n35133 = pi17 ? n35130 : ~n35132;
  assign n35134 = pi16 ? n32 : n35133;
  assign n35135 = pi15 ? n35128 : n35134;
  assign n35136 = pi18 ? n14153 : n323;
  assign n35137 = pi17 ? n2519 : ~n35136;
  assign n35138 = pi16 ? n32 : n35137;
  assign n35139 = pi19 ? n349 : ~n247;
  assign n35140 = pi18 ? n35139 : ~n32;
  assign n35141 = pi17 ? n35140 : ~n2519;
  assign n35142 = pi16 ? n32 : n35141;
  assign n35143 = pi15 ? n35138 : n35142;
  assign n35144 = pi14 ? n35135 : n35143;
  assign n35145 = pi13 ? n35125 : n35144;
  assign n35146 = pi18 ? n23539 : n32;
  assign n35147 = pi17 ? n23538 : ~n35146;
  assign n35148 = pi16 ? n1683 : ~n35147;
  assign n35149 = pi17 ? n17346 : n19803;
  assign n35150 = pi16 ? n32 : n35149;
  assign n35151 = pi15 ? n35148 : n35150;
  assign n35152 = pi17 ? n17346 : n238;
  assign n35153 = pi16 ? n32 : n35152;
  assign n35154 = pi20 ? n6621 : ~n32;
  assign n35155 = pi19 ? n1490 : n35154;
  assign n35156 = pi18 ? n35155 : n30839;
  assign n35157 = pi17 ? n35156 : ~n2325;
  assign n35158 = pi16 ? n26095 : n35157;
  assign n35159 = pi15 ? n35153 : n35158;
  assign n35160 = pi14 ? n35151 : n35159;
  assign n35161 = pi16 ? n1683 : ~n2326;
  assign n35162 = pi16 ? n1135 : ~n3625;
  assign n35163 = pi15 ? n35161 : n35162;
  assign n35164 = pi15 ? n30941 : n18979;
  assign n35165 = pi14 ? n35163 : n35164;
  assign n35166 = pi13 ? n35160 : n35165;
  assign n35167 = pi12 ? n35145 : n35166;
  assign n35168 = pi11 ? n35110 : n35167;
  assign n35169 = pi10 ? n35057 : n35168;
  assign n35170 = pi09 ? n32 : n35169;
  assign n35171 = pi15 ? n16108 : n23574;
  assign n35172 = pi14 ? n35171 : n23736;
  assign n35173 = pi13 ? n35018 : n35172;
  assign n35174 = pi15 ? n23569 : n32;
  assign n35175 = pi14 ? n35174 : n32;
  assign n35176 = pi15 ? n23484 : n23749;
  assign n35177 = pi15 ? n23631 : n35023;
  assign n35178 = pi14 ? n35176 : n35177;
  assign n35179 = pi13 ? n35175 : n35178;
  assign n35180 = pi12 ? n35173 : n35179;
  assign n35181 = pi14 ? n24614 : n22540;
  assign n35182 = pi14 ? n32 : n35053;
  assign n35183 = pi13 ? n35181 : n35182;
  assign n35184 = pi12 ? n35043 : n35183;
  assign n35185 = pi11 ? n35180 : n35184;
  assign n35186 = pi19 ? n1757 : ~n1105;
  assign n35187 = pi18 ? n32 : n35186;
  assign n35188 = pi17 ? n32 : n35187;
  assign n35189 = pi16 ? n32 : n35188;
  assign n35190 = pi15 ? n35071 : n35189;
  assign n35191 = pi14 ? n35068 : n35190;
  assign n35192 = pi13 ? n35191 : n35075;
  assign n35193 = pi18 ? n14153 : ~n13335;
  assign n35194 = pi17 ? n35083 : ~n35193;
  assign n35195 = pi16 ? n32 : n35194;
  assign n35196 = pi15 ? n35195 : n35090;
  assign n35197 = pi14 ? n35081 : n35196;
  assign n35198 = pi17 ? n35093 : ~n2512;
  assign n35199 = pi16 ? n32 : n35198;
  assign n35200 = pi15 ? n35199 : n35097;
  assign n35201 = pi20 ? n207 : ~n10889;
  assign n35202 = pi19 ? n35201 : n32;
  assign n35203 = pi18 ? n4983 : ~n35202;
  assign n35204 = pi17 ? n8859 : ~n35203;
  assign n35205 = pi16 ? n32 : n35204;
  assign n35206 = pi15 ? n35205 : n35106;
  assign n35207 = pi14 ? n35200 : n35206;
  assign n35208 = pi13 ? n35197 : n35207;
  assign n35209 = pi12 ? n35192 : n35208;
  assign n35210 = pi18 ? n936 : ~n2754;
  assign n35211 = pi17 ? n32 : n35210;
  assign n35212 = pi16 ? n32 : n35211;
  assign n35213 = pi15 ? n35120 : n35212;
  assign n35214 = pi14 ? n35115 : n35213;
  assign n35215 = pi13 ? n35214 : n35144;
  assign n35216 = pi12 ? n35215 : n35166;
  assign n35217 = pi11 ? n35209 : n35216;
  assign n35218 = pi10 ? n35185 : n35217;
  assign n35219 = pi09 ? n32 : n35218;
  assign n35220 = pi08 ? n35170 : n35219;
  assign n35221 = pi14 ? n23726 : n23569;
  assign n35222 = pi15 ? n23569 : n23574;
  assign n35223 = pi14 ? n35222 : n23574;
  assign n35224 = pi13 ? n35221 : n35223;
  assign n35225 = pi15 ? n23484 : n23631;
  assign n35226 = pi15 ? n23749 : n14570;
  assign n35227 = pi14 ? n35225 : n35226;
  assign n35228 = pi13 ? n23577 : n35227;
  assign n35229 = pi12 ? n35224 : n35228;
  assign n35230 = pi19 ? n221 : n7502;
  assign n35231 = pi18 ? n32 : n35230;
  assign n35232 = pi17 ? n32 : n35231;
  assign n35233 = pi16 ? n32 : n35232;
  assign n35234 = pi15 ? n35233 : n23631;
  assign n35235 = pi15 ? n23631 : n35030;
  assign n35236 = pi14 ? n35234 : n35235;
  assign n35237 = pi15 ? n25790 : n23340;
  assign n35238 = pi14 ? n35237 : n26258;
  assign n35239 = pi13 ? n35236 : n35238;
  assign n35240 = pi15 ? n15119 : n22540;
  assign n35241 = pi18 ? n32 : n18102;
  assign n35242 = pi19 ? n1757 : n1844;
  assign n35243 = pi18 ? n35242 : n32;
  assign n35244 = pi17 ? n35241 : n35243;
  assign n35245 = pi16 ? n32 : n35244;
  assign n35246 = pi15 ? n32 : n35245;
  assign n35247 = pi14 ? n35240 : n35246;
  assign n35248 = pi20 ? n1076 : n9491;
  assign n35249 = pi19 ? n32 : n35248;
  assign n35250 = pi20 ? n287 : ~n2180;
  assign n35251 = pi19 ? n35250 : ~n9491;
  assign n35252 = pi18 ? n35249 : ~n35251;
  assign n35253 = pi20 ? n266 : n1076;
  assign n35254 = pi19 ? n35253 : n17649;
  assign n35255 = pi18 ? n35254 : n702;
  assign n35256 = pi17 ? n35252 : ~n35255;
  assign n35257 = pi16 ? n32 : n35256;
  assign n35258 = pi17 ? n1978 : ~n2750;
  assign n35259 = pi16 ? n32 : n35258;
  assign n35260 = pi15 ? n35257 : n35259;
  assign n35261 = pi14 ? n32 : n35260;
  assign n35262 = pi13 ? n35247 : n35261;
  assign n35263 = pi12 ? n35239 : n35262;
  assign n35264 = pi11 ? n35229 : n35263;
  assign n35265 = pi19 ? n349 : n18390;
  assign n35266 = pi18 ? n863 : ~n35265;
  assign n35267 = pi18 ? n25244 : n702;
  assign n35268 = pi17 ? n35266 : ~n35267;
  assign n35269 = pi16 ? n32 : n35268;
  assign n35270 = pi19 ? n5694 : n322;
  assign n35271 = pi18 ? n35270 : ~n508;
  assign n35272 = pi17 ? n32 : n35271;
  assign n35273 = pi16 ? n32 : n35272;
  assign n35274 = pi15 ? n35269 : n35273;
  assign n35275 = pi19 ? n236 : ~n1464;
  assign n35276 = pi18 ? n35275 : ~n32584;
  assign n35277 = pi17 ? n32 : ~n35276;
  assign n35278 = pi16 ? n32 : n35277;
  assign n35279 = pi15 ? n35278 : n13948;
  assign n35280 = pi14 ? n35274 : n35279;
  assign n35281 = pi15 ? n24543 : n32;
  assign n35282 = pi14 ? n35281 : n32;
  assign n35283 = pi13 ? n35280 : n35282;
  assign n35284 = pi19 ? n33796 : ~n5688;
  assign n35285 = pi18 ? n35284 : n595;
  assign n35286 = pi17 ? n2954 : ~n35285;
  assign n35287 = pi16 ? n32 : n35286;
  assign n35288 = pi15 ? n20836 : n35287;
  assign n35289 = pi19 ? n17918 : n1325;
  assign n35290 = pi18 ? n35289 : n595;
  assign n35291 = pi17 ? n2519 : ~n35290;
  assign n35292 = pi16 ? n32 : n35291;
  assign n35293 = pi17 ? n2531 : ~n2618;
  assign n35294 = pi16 ? n32 : n35293;
  assign n35295 = pi15 ? n35292 : n35294;
  assign n35296 = pi14 ? n35288 : n35295;
  assign n35297 = pi20 ? n29457 : ~n357;
  assign n35298 = pi19 ? n35297 : ~n32;
  assign n35299 = pi18 ? n18102 : n35298;
  assign n35300 = pi17 ? n35299 : ~n2618;
  assign n35301 = pi16 ? n32 : n35300;
  assign n35302 = pi15 ? n35301 : n8327;
  assign n35303 = pi19 ? n1325 : n349;
  assign n35304 = pi18 ? n32 : n35303;
  assign n35305 = pi18 ? n4983 : ~n13335;
  assign n35306 = pi17 ? n35304 : ~n35305;
  assign n35307 = pi16 ? n32 : n35306;
  assign n35308 = pi15 ? n35307 : n35106;
  assign n35309 = pi14 ? n35302 : n35308;
  assign n35310 = pi13 ? n35296 : n35309;
  assign n35311 = pi12 ? n35283 : n35310;
  assign n35312 = pi15 ? n23892 : n23551;
  assign n35313 = pi18 ? n32 : n19194;
  assign n35314 = pi17 ? n32 : n35313;
  assign n35315 = pi16 ? n32 : n35314;
  assign n35316 = pi15 ? n35315 : n23889;
  assign n35317 = pi14 ? n35312 : n35316;
  assign n35318 = pi19 ? n24763 : ~n208;
  assign n35319 = pi18 ? n35318 : n2754;
  assign n35320 = pi17 ? n31472 : ~n35319;
  assign n35321 = pi16 ? n32 : n35320;
  assign n35322 = pi15 ? n12527 : n35321;
  assign n35323 = pi20 ? n339 : n6050;
  assign n35324 = pi19 ? n176 : ~n35323;
  assign n35325 = pi20 ? n220 : ~n9491;
  assign n35326 = pi19 ? n35325 : n32;
  assign n35327 = pi18 ? n35324 : ~n35326;
  assign n35328 = pi18 ? n5502 : n2754;
  assign n35329 = pi17 ? n35327 : ~n35328;
  assign n35330 = pi16 ? n32 : n35329;
  assign n35331 = pi18 ? n20912 : n323;
  assign n35332 = pi17 ? n1500 : ~n35331;
  assign n35333 = pi16 ? n32 : n35332;
  assign n35334 = pi15 ? n35330 : n35333;
  assign n35335 = pi14 ? n35322 : n35334;
  assign n35336 = pi13 ? n35317 : n35335;
  assign n35337 = pi19 ? n321 : ~n4342;
  assign n35338 = pi18 ? n35337 : ~n32;
  assign n35339 = pi17 ? n2733 : n35338;
  assign n35340 = pi16 ? n1683 : ~n35339;
  assign n35341 = pi17 ? n4128 : n248;
  assign n35342 = pi16 ? n32 : n35341;
  assign n35343 = pi15 ? n35340 : n35342;
  assign n35344 = pi20 ? n342 : n1817;
  assign n35345 = pi19 ? n32 : n35344;
  assign n35346 = pi19 ? n4342 : ~n5707;
  assign n35347 = pi18 ? n35345 : n35346;
  assign n35348 = pi19 ? n28134 : ~n4342;
  assign n35349 = pi18 ? n35348 : ~n237;
  assign n35350 = pi17 ? n35347 : n35349;
  assign n35351 = pi16 ? n32 : n35350;
  assign n35352 = pi19 ? n14022 : n8611;
  assign n35353 = pi19 ? n18665 : ~n349;
  assign n35354 = pi18 ? n35352 : ~n35353;
  assign n35355 = pi17 ? n35354 : ~n2325;
  assign n35356 = pi16 ? n32 : n35355;
  assign n35357 = pi15 ? n35351 : n35356;
  assign n35358 = pi14 ? n35343 : n35357;
  assign n35359 = pi16 ? n1233 : ~n3625;
  assign n35360 = pi15 ? n35161 : n35359;
  assign n35361 = pi20 ? n32 : n259;
  assign n35362 = pi19 ? n32 : n35361;
  assign n35363 = pi18 ? n35362 : ~n32;
  assign n35364 = pi17 ? n32 : n35363;
  assign n35365 = pi19 ? n32340 : ~n32;
  assign n35366 = pi18 ? n32 : n35365;
  assign n35367 = pi17 ? n32 : n35366;
  assign n35368 = pi16 ? n35364 : ~n35367;
  assign n35369 = pi18 ? n32 : ~n13949;
  assign n35370 = pi17 ? n23711 : n35369;
  assign n35371 = pi16 ? n1233 : ~n35370;
  assign n35372 = pi15 ? n35368 : n35371;
  assign n35373 = pi14 ? n35360 : n35372;
  assign n35374 = pi13 ? n35358 : n35373;
  assign n35375 = pi12 ? n35336 : n35374;
  assign n35376 = pi11 ? n35311 : n35375;
  assign n35377 = pi10 ? n35264 : n35376;
  assign n35378 = pi09 ? n32 : n35377;
  assign n35379 = pi14 ? n23726 : n23574;
  assign n35380 = pi15 ? n23574 : n23730;
  assign n35381 = pi14 ? n35380 : n23725;
  assign n35382 = pi13 ? n35379 : n35381;
  assign n35383 = pi15 ? n23484 : n24256;
  assign n35384 = pi15 ? n23933 : n14570;
  assign n35385 = pi14 ? n35383 : n35384;
  assign n35386 = pi13 ? n23795 : n35385;
  assign n35387 = pi12 ? n35382 : n35386;
  assign n35388 = pi15 ? n14389 : n16108;
  assign n35389 = pi15 ? n23741 : n35030;
  assign n35390 = pi14 ? n35388 : n35389;
  assign n35391 = pi18 ? n32 : n6132;
  assign n35392 = pi17 ? n32 : n35391;
  assign n35393 = pi16 ? n32 : n35392;
  assign n35394 = pi15 ? n35393 : n15386;
  assign n35395 = pi15 ? n23484 : n15386;
  assign n35396 = pi14 ? n35394 : n35395;
  assign n35397 = pi13 ? n35390 : n35396;
  assign n35398 = pi15 ? n24742 : n22540;
  assign n35399 = pi14 ? n35398 : n35246;
  assign n35400 = pi19 ? n32 : n31202;
  assign n35401 = pi18 ? n35400 : ~n35251;
  assign n35402 = pi17 ? n35401 : ~n35255;
  assign n35403 = pi16 ? n32 : n35402;
  assign n35404 = pi15 ? n35403 : n35259;
  assign n35405 = pi14 ? n32 : n35404;
  assign n35406 = pi13 ? n35399 : n35405;
  assign n35407 = pi12 ? n35397 : n35406;
  assign n35408 = pi11 ? n35387 : n35407;
  assign n35409 = pi21 ? n174 : n7107;
  assign n35410 = pi20 ? n32 : n35409;
  assign n35411 = pi19 ? n35410 : n32;
  assign n35412 = pi18 ? n32 : n35411;
  assign n35413 = pi17 ? n32 : n35412;
  assign n35414 = pi16 ? n32 : n35413;
  assign n35415 = pi15 ? n35414 : n35287;
  assign n35416 = pi14 ? n35415 : n35295;
  assign n35417 = pi13 ? n35416 : n35309;
  assign n35418 = pi12 ? n35283 : n35417;
  assign n35419 = pi18 ? n32 : n8908;
  assign n35420 = pi17 ? n32 : n35419;
  assign n35421 = pi16 ? n32 : n35420;
  assign n35422 = pi15 ? n13046 : n35421;
  assign n35423 = pi14 ? n35422 : n35316;
  assign n35424 = pi18 ? n5502 : n323;
  assign n35425 = pi17 ? n35327 : ~n35424;
  assign n35426 = pi16 ? n32 : n35425;
  assign n35427 = pi15 ? n35426 : n35333;
  assign n35428 = pi14 ? n35322 : n35427;
  assign n35429 = pi13 ? n35423 : n35428;
  assign n35430 = pi16 ? n1135 : ~n35370;
  assign n35431 = pi15 ? n35368 : n35430;
  assign n35432 = pi14 ? n35163 : n35431;
  assign n35433 = pi13 ? n35358 : n35432;
  assign n35434 = pi12 ? n35429 : n35433;
  assign n35435 = pi11 ? n35418 : n35434;
  assign n35436 = pi10 ? n35408 : n35435;
  assign n35437 = pi09 ? n32 : n35436;
  assign n35438 = pi08 ? n35378 : n35437;
  assign n35439 = pi07 ? n35220 : n35438;
  assign n35440 = pi14 ? n23924 : n23725;
  assign n35441 = pi13 ? n35440 : n23725;
  assign n35442 = pi15 ? n25657 : n23730;
  assign n35443 = pi14 ? n23574 : n35442;
  assign n35444 = pi13 ? n23795 : n35443;
  assign n35445 = pi12 ? n35441 : n35444;
  assign n35446 = pi19 ? n267 : ~n813;
  assign n35447 = pi18 ? n32 : n35446;
  assign n35448 = pi17 ? n32 : n35447;
  assign n35449 = pi16 ? n32 : n35448;
  assign n35450 = pi18 ? n32 : n5725;
  assign n35451 = pi17 ? n32 : n35450;
  assign n35452 = pi16 ? n32 : n35451;
  assign n35453 = pi15 ? n35449 : n35452;
  assign n35454 = pi14 ? n23574 : n35453;
  assign n35455 = pi19 ? n275 : ~n617;
  assign n35456 = pi18 ? n35455 : n24015;
  assign n35457 = pi17 ? n32 : n35456;
  assign n35458 = pi16 ? n32 : n35457;
  assign n35459 = pi15 ? n35458 : n23484;
  assign n35460 = pi14 ? n35459 : n23484;
  assign n35461 = pi13 ? n35454 : n35460;
  assign n35462 = pi20 ? n428 : n501;
  assign n35463 = pi19 ? n5371 : n35462;
  assign n35464 = pi18 ? n35463 : ~n1750;
  assign n35465 = pi17 ? n32 : n35464;
  assign n35466 = pi16 ? n32 : n35465;
  assign n35467 = pi17 ? n32 : n9073;
  assign n35468 = pi19 ? n23644 : n28134;
  assign n35469 = pi19 ? n13069 : n3523;
  assign n35470 = pi18 ? n35468 : ~n35469;
  assign n35471 = pi20 ? n1331 : ~n266;
  assign n35472 = pi19 ? n35471 : n9822;
  assign n35473 = pi18 ? n35472 : ~n1750;
  assign n35474 = pi17 ? n35470 : ~n35473;
  assign n35475 = pi16 ? n35467 : ~n35474;
  assign n35476 = pi15 ? n35466 : n35475;
  assign n35477 = pi14 ? n24327 : n35476;
  assign n35478 = pi13 ? n32 : n35477;
  assign n35479 = pi12 ? n35461 : n35478;
  assign n35480 = pi11 ? n35445 : n35479;
  assign n35481 = pi20 ? n342 : n9488;
  assign n35482 = pi20 ? n2180 : n1611;
  assign n35483 = pi19 ? n35481 : ~n35482;
  assign n35484 = pi20 ? n357 : n2180;
  assign n35485 = pi19 ? n35484 : n18832;
  assign n35486 = pi18 ? n35483 : ~n35485;
  assign n35487 = pi20 ? n17669 : n5854;
  assign n35488 = pi20 ? n8644 : n17665;
  assign n35489 = pi19 ? n35487 : ~n35488;
  assign n35490 = pi19 ? n267 : n617;
  assign n35491 = pi18 ? n35489 : n35490;
  assign n35492 = pi17 ? n35486 : ~n35491;
  assign n35493 = pi16 ? n32 : n35492;
  assign n35494 = pi19 ? n3692 : n3523;
  assign n35495 = pi18 ? n32 : n35494;
  assign n35496 = pi20 ? n2385 : n342;
  assign n35497 = pi19 ? n8611 : n35496;
  assign n35498 = pi18 ? n35497 : n23514;
  assign n35499 = pi17 ? n35495 : n35498;
  assign n35500 = pi16 ? n32 : n35499;
  assign n35501 = pi15 ? n35493 : n35500;
  assign n35502 = pi19 ? n3495 : n507;
  assign n35503 = pi19 ? n16189 : n32;
  assign n35504 = pi18 ? n35502 : n35503;
  assign n35505 = pi17 ? n32 : n35504;
  assign n35506 = pi16 ? n32 : n35505;
  assign n35507 = pi18 ? n6059 : n248;
  assign n35508 = pi17 ? n32 : n35507;
  assign n35509 = pi16 ? n32 : n35508;
  assign n35510 = pi15 ? n35506 : n35509;
  assign n35511 = pi14 ? n35501 : n35510;
  assign n35512 = pi13 ? n35511 : n21455;
  assign n35513 = pi20 ? n321 : ~n101;
  assign n35514 = pi19 ? n35513 : n32;
  assign n35515 = pi18 ? n32 : n35514;
  assign n35516 = pi17 ? n32 : n35515;
  assign n35517 = pi16 ? n32 : n35516;
  assign n35518 = pi19 ? n507 : ~n1464;
  assign n35519 = pi20 ? n12884 : n101;
  assign n35520 = pi19 ? n35519 : ~n32;
  assign n35521 = pi18 ? n35518 : n35520;
  assign n35522 = pi17 ? n16848 : ~n35521;
  assign n35523 = pi16 ? n32 : n35522;
  assign n35524 = pi15 ? n35517 : n35523;
  assign n35525 = pi19 ? n322 : n4391;
  assign n35526 = pi18 ? n35525 : n4098;
  assign n35527 = pi17 ? n2726 : ~n35526;
  assign n35528 = pi16 ? n32 : n35527;
  assign n35529 = pi18 ? n34283 : n4098;
  assign n35530 = pi17 ? n2726 : ~n35529;
  assign n35531 = pi16 ? n32 : n35530;
  assign n35532 = pi15 ? n35528 : n35531;
  assign n35533 = pi14 ? n35524 : n35532;
  assign n35534 = pi17 ? n2750 : ~n2618;
  assign n35535 = pi16 ? n32 : n35534;
  assign n35536 = pi20 ? n518 : ~n2385;
  assign n35537 = pi19 ? n35536 : n32;
  assign n35538 = pi18 ? n32 : n35537;
  assign n35539 = pi17 ? n32 : n35538;
  assign n35540 = pi16 ? n32 : n35539;
  assign n35541 = pi15 ? n35535 : n35540;
  assign n35542 = pi18 ? n6669 : n508;
  assign n35543 = pi17 ? n2959 : ~n35542;
  assign n35544 = pi16 ? n32 : n35543;
  assign n35545 = pi19 ? n11027 : ~n32;
  assign n35546 = pi18 ? n940 : ~n35545;
  assign n35547 = pi17 ? n32 : n35546;
  assign n35548 = pi16 ? n32 : n35547;
  assign n35549 = pi15 ? n35544 : n35548;
  assign n35550 = pi14 ? n35541 : n35549;
  assign n35551 = pi13 ? n35533 : n35550;
  assign n35552 = pi12 ? n35512 : n35551;
  assign n35553 = pi19 ? n35344 : n32;
  assign n35554 = pi18 ? n32 : n35553;
  assign n35555 = pi17 ? n32 : n35554;
  assign n35556 = pi16 ? n32 : n35555;
  assign n35557 = pi15 ? n33939 : n35556;
  assign n35558 = pi14 ? n35557 : n23874;
  assign n35559 = pi15 ? n23874 : n13046;
  assign n35560 = pi19 ? n32 : n207;
  assign n35561 = pi18 ? n35560 : ~n32;
  assign n35562 = pi17 ? n35561 : ~n1807;
  assign n35563 = pi16 ? n32 : n35562;
  assign n35564 = pi19 ? n4964 : ~n32;
  assign n35565 = pi18 ? n35564 : ~n222;
  assign n35566 = pi18 ? n23875 : n32;
  assign n35567 = pi17 ? n35565 : n35566;
  assign n35568 = pi16 ? n32 : n35567;
  assign n35569 = pi15 ? n35563 : n35568;
  assign n35570 = pi14 ? n35559 : n35569;
  assign n35571 = pi13 ? n35558 : n35570;
  assign n35572 = pi18 ? n32 : n4428;
  assign n35573 = pi17 ? n32 : n35572;
  assign n35574 = pi18 ? n23882 : n32;
  assign n35575 = pi17 ? n32 : ~n35574;
  assign n35576 = pi16 ? n35573 : ~n35575;
  assign n35577 = pi15 ? n35576 : n32;
  assign n35578 = pi20 ? n1324 : ~n321;
  assign n35579 = pi19 ? n35578 : n4342;
  assign n35580 = pi18 ? n32 : ~n35579;
  assign n35581 = pi19 ? n322 : n6988;
  assign n35582 = pi18 ? n35581 : ~n32;
  assign n35583 = pi17 ? n35580 : ~n35582;
  assign n35584 = pi16 ? n32 : n35583;
  assign n35585 = pi19 ? n321 : ~n4670;
  assign n35586 = pi18 ? n32 : n35585;
  assign n35587 = pi18 ? n5694 : ~n32;
  assign n35588 = pi17 ? n35586 : ~n35587;
  assign n35589 = pi16 ? n32 : n35588;
  assign n35590 = pi15 ? n35584 : n35589;
  assign n35591 = pi14 ? n35577 : n35590;
  assign n35592 = pi19 ? n20006 : n349;
  assign n35593 = pi18 ? n35592 : ~n23896;
  assign n35594 = pi18 ? n23899 : ~n32;
  assign n35595 = pi17 ? n35593 : ~n35594;
  assign n35596 = pi16 ? n32 : n35595;
  assign n35597 = pi18 ? n1190 : ~n32;
  assign n35598 = pi17 ? n32 : n35597;
  assign n35599 = pi16 ? n35598 : ~n1808;
  assign n35600 = pi15 ? n35596 : n35599;
  assign n35601 = pi20 ? n32 : n29452;
  assign n35602 = pi19 ? n32 : n35601;
  assign n35603 = pi18 ? n35602 : n237;
  assign n35604 = pi17 ? n32 : n35603;
  assign n35605 = pi18 ? n23906 : n350;
  assign n35606 = pi17 ? n23905 : n35605;
  assign n35607 = pi16 ? n35604 : ~n35606;
  assign n35608 = pi18 ? n1190 : n605;
  assign n35609 = pi17 ? n32 : n35608;
  assign n35610 = pi18 ? n16432 : ~n814;
  assign n35611 = pi17 ? n23912 : ~n35610;
  assign n35612 = pi16 ? n35609 : ~n35611;
  assign n35613 = pi15 ? n35607 : n35612;
  assign n35614 = pi14 ? n35600 : n35613;
  assign n35615 = pi13 ? n35591 : n35614;
  assign n35616 = pi12 ? n35571 : n35615;
  assign n35617 = pi11 ? n35552 : n35616;
  assign n35618 = pi10 ? n35480 : n35617;
  assign n35619 = pi09 ? n32 : n35618;
  assign n35620 = pi15 ? n23725 : n16319;
  assign n35621 = pi14 ? n35620 : n16319;
  assign n35622 = pi13 ? n35440 : n35621;
  assign n35623 = pi15 ? n15248 : n23730;
  assign n35624 = pi14 ? n35380 : n35623;
  assign n35625 = pi13 ? n16322 : n35624;
  assign n35626 = pi12 ? n35622 : n35625;
  assign n35627 = pi16 ? n4578 : ~n35474;
  assign n35628 = pi15 ? n35466 : n35627;
  assign n35629 = pi14 ? n24327 : n35628;
  assign n35630 = pi13 ? n32 : n35629;
  assign n35631 = pi12 ? n35461 : n35630;
  assign n35632 = pi11 ? n35626 : n35631;
  assign n35633 = pi19 ? n35484 : n18173;
  assign n35634 = pi18 ? n35483 : ~n35633;
  assign n35635 = pi20 ? n18415 : n5854;
  assign n35636 = pi20 ? n1076 : n17665;
  assign n35637 = pi19 ? n35635 : ~n35636;
  assign n35638 = pi18 ? n35637 : n35490;
  assign n35639 = pi17 ? n35634 : ~n35638;
  assign n35640 = pi16 ? n32 : n35639;
  assign n35641 = pi19 ? n531 : n35496;
  assign n35642 = pi18 ? n35641 : n23514;
  assign n35643 = pi17 ? n35495 : n35642;
  assign n35644 = pi16 ? n32 : n35643;
  assign n35645 = pi15 ? n35640 : n35644;
  assign n35646 = pi14 ? n35645 : n35510;
  assign n35647 = pi13 ? n35646 : n21455;
  assign n35648 = pi18 ? n32 : n6159;
  assign n35649 = pi17 ? n32 : n35648;
  assign n35650 = pi16 ? n32 : n35649;
  assign n35651 = pi20 ? n12884 : n428;
  assign n35652 = pi19 ? n35651 : ~n32;
  assign n35653 = pi18 ? n35518 : n35652;
  assign n35654 = pi17 ? n16848 : ~n35653;
  assign n35655 = pi16 ? n32 : n35654;
  assign n35656 = pi15 ? n35650 : n35655;
  assign n35657 = pi18 ? n35525 : n595;
  assign n35658 = pi17 ? n2726 : ~n35657;
  assign n35659 = pi16 ? n32 : n35658;
  assign n35660 = pi18 ? n34283 : n595;
  assign n35661 = pi17 ? n2726 : ~n35660;
  assign n35662 = pi16 ? n32 : n35661;
  assign n35663 = pi15 ? n35659 : n35662;
  assign n35664 = pi14 ? n35656 : n35663;
  assign n35665 = pi19 ? n32302 : n32;
  assign n35666 = pi18 ? n32 : n35665;
  assign n35667 = pi17 ? n32 : n35666;
  assign n35668 = pi16 ? n32 : n35667;
  assign n35669 = pi15 ? n35535 : n35668;
  assign n35670 = pi14 ? n35669 : n35549;
  assign n35671 = pi13 ? n35664 : n35670;
  assign n35672 = pi12 ? n35647 : n35671;
  assign n35673 = pi15 ? n35596 : n30941;
  assign n35674 = pi18 ? n35362 : n237;
  assign n35675 = pi17 ? n32 : n35674;
  assign n35676 = pi16 ? n35675 : ~n35606;
  assign n35677 = pi18 ? n833 : n605;
  assign n35678 = pi17 ? n32 : n35677;
  assign n35679 = pi16 ? n35678 : ~n35611;
  assign n35680 = pi15 ? n35676 : n35679;
  assign n35681 = pi14 ? n35673 : n35680;
  assign n35682 = pi13 ? n35591 : n35681;
  assign n35683 = pi12 ? n35571 : n35682;
  assign n35684 = pi11 ? n35672 : n35683;
  assign n35685 = pi10 ? n35632 : n35684;
  assign n35686 = pi09 ? n32 : n35685;
  assign n35687 = pi08 ? n35619 : n35686;
  assign n35688 = pi15 ? n32 : n16377;
  assign n35689 = pi14 ? n35688 : n16319;
  assign n35690 = pi13 ? n35689 : n23981;
  assign n35691 = pi15 ? n23981 : n32;
  assign n35692 = pi14 ? n35691 : n32;
  assign n35693 = pi15 ? n23725 : n14917;
  assign n35694 = pi15 ? n15080 : n16105;
  assign n35695 = pi14 ? n35693 : n35694;
  assign n35696 = pi13 ? n35692 : n35695;
  assign n35697 = pi12 ? n35690 : n35696;
  assign n35698 = pi19 ? n531 : ~n813;
  assign n35699 = pi18 ? n32 : n35698;
  assign n35700 = pi17 ? n32 : n35699;
  assign n35701 = pi16 ? n32 : n35700;
  assign n35702 = pi15 ? n24251 : n35701;
  assign n35703 = pi14 ? n32 : n35702;
  assign n35704 = pi19 ? n267 : n3523;
  assign n35705 = pi18 ? n32 : n35704;
  assign n35706 = pi20 ? n310 : n266;
  assign n35707 = pi20 ? n6050 : ~n246;
  assign n35708 = pi19 ? n35706 : ~n35707;
  assign n35709 = pi19 ? n4406 : ~n813;
  assign n35710 = pi18 ? n35708 : n35709;
  assign n35711 = pi17 ? n35705 : n35710;
  assign n35712 = pi16 ? n32 : n35711;
  assign n35713 = pi15 ? n35712 : n23933;
  assign n35714 = pi14 ? n35713 : n23933;
  assign n35715 = pi13 ? n35703 : n35714;
  assign n35716 = pi18 ? n22819 : ~n1750;
  assign n35717 = pi17 ? n32 : n35716;
  assign n35718 = pi16 ? n32 : n35717;
  assign n35719 = pi19 ? n1757 : ~n32;
  assign n35720 = pi18 ? n23440 : ~n35719;
  assign n35721 = pi17 ? n13946 : n35720;
  assign n35722 = pi16 ? n32 : n35721;
  assign n35723 = pi15 ? n35718 : n35722;
  assign n35724 = pi14 ? n32 : n35723;
  assign n35725 = pi13 ? n32 : n35724;
  assign n35726 = pi12 ? n35715 : n35725;
  assign n35727 = pi11 ? n35697 : n35726;
  assign n35728 = pi19 ? n5371 : ~n617;
  assign n35729 = pi18 ? n6145 : n35728;
  assign n35730 = pi17 ? n13946 : n35729;
  assign n35731 = pi16 ? n32 : n35730;
  assign n35732 = pi19 ? n34295 : n32;
  assign n35733 = pi18 ? n6145 : n35732;
  assign n35734 = pi17 ? n32 : n35733;
  assign n35735 = pi16 ? n32 : n35734;
  assign n35736 = pi15 ? n35731 : n35735;
  assign n35737 = pi14 ? n35736 : n30921;
  assign n35738 = pi19 ? n22864 : n32;
  assign n35739 = pi18 ? n32 : n35738;
  assign n35740 = pi17 ? n32 : n35739;
  assign n35741 = pi16 ? n32 : n35740;
  assign n35742 = pi15 ? n32 : n35741;
  assign n35743 = pi14 ? n32 : n35742;
  assign n35744 = pi13 ? n35737 : n35743;
  assign n35745 = pi18 ? n19232 : n6163;
  assign n35746 = pi17 ? n32 : n35745;
  assign n35747 = pi16 ? n32 : n35746;
  assign n35748 = pi18 ? n508 : n35719;
  assign n35749 = pi17 ? n16848 : ~n35748;
  assign n35750 = pi16 ? n32 : n35749;
  assign n35751 = pi15 ? n35747 : n35750;
  assign n35752 = pi19 ? n1464 : n5435;
  assign n35753 = pi18 ? n35752 : n702;
  assign n35754 = pi17 ? n2726 : ~n35753;
  assign n35755 = pi16 ? n32 : n35754;
  assign n35756 = pi18 ? n34283 : n702;
  assign n35757 = pi17 ? n2726 : ~n35756;
  assign n35758 = pi16 ? n32 : n35757;
  assign n35759 = pi15 ? n35755 : n35758;
  assign n35760 = pi14 ? n35751 : n35759;
  assign n35761 = pi17 ? n2750 : ~n2512;
  assign n35762 = pi16 ? n32 : n35761;
  assign n35763 = pi15 ? n35762 : n8901;
  assign n35764 = pi18 ? n940 : ~n25110;
  assign n35765 = pi17 ? n32 : n35764;
  assign n35766 = pi16 ? n32 : n35765;
  assign n35767 = pi15 ? n35544 : n35766;
  assign n35768 = pi14 ? n35763 : n35767;
  assign n35769 = pi13 ? n35760 : n35768;
  assign n35770 = pi12 ? n35744 : n35769;
  assign n35771 = pi15 ? n33939 : n34852;
  assign n35772 = pi20 ? n342 : ~n1319;
  assign n35773 = pi19 ? n35772 : n32;
  assign n35774 = pi18 ? n32 : n35773;
  assign n35775 = pi17 ? n32 : n35774;
  assign n35776 = pi16 ? n32 : n35775;
  assign n35777 = pi15 ? n35776 : n13636;
  assign n35778 = pi14 ? n35771 : n35777;
  assign n35779 = pi15 ? n35776 : n13043;
  assign n35780 = pi19 ? n32 : ~n9007;
  assign n35781 = pi18 ? n35780 : ~n268;
  assign n35782 = pi19 ? n1757 : n32083;
  assign n35783 = pi18 ? n35782 : ~n9578;
  assign n35784 = pi17 ? n35781 : ~n35783;
  assign n35785 = pi16 ? n32 : n35784;
  assign n35786 = pi18 ? n35564 : ~n32;
  assign n35787 = pi17 ? n35786 : ~n1580;
  assign n35788 = pi16 ? n32 : n35787;
  assign n35789 = pi15 ? n35785 : n35788;
  assign n35790 = pi14 ? n35779 : n35789;
  assign n35791 = pi13 ? n35778 : n35790;
  assign n35792 = pi18 ? n16603 : ~n6059;
  assign n35793 = pi17 ? n32 : n35792;
  assign n35794 = pi16 ? n2745 : ~n35793;
  assign n35795 = pi15 ? n35794 : n32;
  assign n35796 = pi19 ? n4964 : n4342;
  assign n35797 = pi18 ? n32 : ~n35796;
  assign n35798 = pi19 ? n322 : n4964;
  assign n35799 = pi18 ? n35798 : ~n32;
  assign n35800 = pi17 ? n35797 : ~n35799;
  assign n35801 = pi16 ? n32 : n35800;
  assign n35802 = pi19 ? n31490 : ~n4670;
  assign n35803 = pi18 ? n18085 : n35802;
  assign n35804 = pi19 ? n267 : n5694;
  assign n35805 = pi18 ? n35804 : ~n32;
  assign n35806 = pi17 ? n35803 : ~n35805;
  assign n35807 = pi16 ? n32 : n35806;
  assign n35808 = pi15 ? n35801 : n35807;
  assign n35809 = pi14 ? n35795 : n35808;
  assign n35810 = pi18 ? n7038 : n24056;
  assign n35811 = pi18 ? n24058 : ~n32;
  assign n35812 = pi17 ? n35810 : ~n35811;
  assign n35813 = pi16 ? n32 : n35812;
  assign n35814 = pi18 ? n222 : ~n23302;
  assign n35815 = pi17 ? n32 : n35814;
  assign n35816 = pi16 ? n35815 : ~n1808;
  assign n35817 = pi15 ? n35813 : n35816;
  assign n35818 = pi19 ? n35154 : ~n32;
  assign n35819 = pi18 ? n268 : n35818;
  assign n35820 = pi17 ? n32 : n35819;
  assign n35821 = pi18 ? n24066 : n32;
  assign n35822 = pi17 ? n24065 : ~n35821;
  assign n35823 = pi16 ? n35820 : ~n35822;
  assign n35824 = pi18 ? n222 : n605;
  assign n35825 = pi17 ? n32 : n35824;
  assign n35826 = pi18 ? n24072 : ~n237;
  assign n35827 = pi17 ? n24071 : ~n35826;
  assign n35828 = pi16 ? n35825 : ~n35827;
  assign n35829 = pi15 ? n35823 : n35828;
  assign n35830 = pi14 ? n35817 : n35829;
  assign n35831 = pi13 ? n35809 : n35830;
  assign n35832 = pi12 ? n35791 : n35831;
  assign n35833 = pi11 ? n35770 : n35832;
  assign n35834 = pi10 ? n35727 : n35833;
  assign n35835 = pi09 ? n32 : n35834;
  assign n35836 = pi15 ? n32 : n25070;
  assign n35837 = pi14 ? n35836 : n23981;
  assign n35838 = pi14 ? n35688 : n16377;
  assign n35839 = pi13 ? n35837 : n35838;
  assign n35840 = pi14 ? n16377 : n32;
  assign n35841 = pi15 ? n16319 : n14917;
  assign n35842 = pi14 ? n35841 : n35694;
  assign n35843 = pi13 ? n35840 : n35842;
  assign n35844 = pi12 ? n35839 : n35843;
  assign n35845 = pi11 ? n35844 : n35726;
  assign n35846 = pi19 ? n22864 : ~n1105;
  assign n35847 = pi18 ? n32 : n35846;
  assign n35848 = pi17 ? n32 : n35847;
  assign n35849 = pi16 ? n32 : n35848;
  assign n35850 = pi15 ? n32 : n35849;
  assign n35851 = pi14 ? n32 : n35850;
  assign n35852 = pi13 ? n35737 : n35851;
  assign n35853 = pi15 ? n13620 : n35750;
  assign n35854 = pi14 ? n35853 : n35759;
  assign n35855 = pi13 ? n35854 : n35768;
  assign n35856 = pi12 ? n35852 : n35855;
  assign n35857 = pi15 ? n13920 : n23874;
  assign n35858 = pi14 ? n35771 : n35857;
  assign n35859 = pi15 ? n13920 : n13043;
  assign n35860 = pi14 ? n35859 : n35789;
  assign n35861 = pi13 ? n35858 : n35860;
  assign n35862 = pi18 ? n268 : n289;
  assign n35863 = pi17 ? n32 : n35862;
  assign n35864 = pi18 ? n24066 : n20828;
  assign n35865 = pi17 ? n24065 : ~n35864;
  assign n35866 = pi16 ? n35863 : ~n35865;
  assign n35867 = pi20 ? n207 : ~n52;
  assign n35868 = pi19 ? n35867 : ~n32;
  assign n35869 = pi18 ? n24072 : ~n35868;
  assign n35870 = pi17 ? n24071 : ~n35869;
  assign n35871 = pi16 ? n35825 : ~n35870;
  assign n35872 = pi15 ? n35866 : n35871;
  assign n35873 = pi14 ? n35817 : n35872;
  assign n35874 = pi13 ? n35809 : n35873;
  assign n35875 = pi12 ? n35861 : n35874;
  assign n35876 = pi11 ? n35856 : n35875;
  assign n35877 = pi10 ? n35845 : n35876;
  assign n35878 = pi09 ? n32 : n35877;
  assign n35879 = pi08 ? n35835 : n35878;
  assign n35880 = pi07 ? n35687 : n35879;
  assign n35881 = pi06 ? n35439 : n35880;
  assign n35882 = pi05 ? n35017 : n35881;
  assign n35883 = pi04 ? n34180 : n35882;
  assign n35884 = pi14 ? n26994 : n16377;
  assign n35885 = pi13 ? n35884 : n16377;
  assign n35886 = pi19 ? n519 : ~n2848;
  assign n35887 = pi18 ? n32 : n35886;
  assign n35888 = pi17 ? n32 : n35887;
  assign n35889 = pi16 ? n32 : n35888;
  assign n35890 = pi15 ? n16105 : n35889;
  assign n35891 = pi15 ? n35889 : n24382;
  assign n35892 = pi14 ? n35890 : n35891;
  assign n35893 = pi13 ? n35840 : n35892;
  assign n35894 = pi12 ? n35885 : n35893;
  assign n35895 = pi18 ? n32 : n32025;
  assign n35896 = pi17 ? n32 : n35895;
  assign n35897 = pi16 ? n32 : n35896;
  assign n35898 = pi15 ? n35897 : n24659;
  assign n35899 = pi14 ? n25779 : n35898;
  assign n35900 = pi15 ? n35030 : n23484;
  assign n35901 = pi19 ? n267 : ~n1812;
  assign n35902 = pi18 ? n32 : n35901;
  assign n35903 = pi17 ? n32 : n35902;
  assign n35904 = pi16 ? n32 : n35903;
  assign n35905 = pi15 ? n14397 : n35904;
  assign n35906 = pi14 ? n35900 : n35905;
  assign n35907 = pi13 ? n35899 : n35906;
  assign n35908 = pi18 ? n4380 : n34142;
  assign n35909 = pi17 ? n32 : n35908;
  assign n35910 = pi16 ? n32 : n35909;
  assign n35911 = pi15 ? n32 : n35910;
  assign n35912 = pi20 ? n2358 : ~n321;
  assign n35913 = pi19 ? n35912 : n321;
  assign n35914 = pi18 ? n35913 : ~n1750;
  assign n35915 = pi17 ? n35241 : n35914;
  assign n35916 = pi16 ? n32 : n35915;
  assign n35917 = pi19 ? n4721 : ~n21282;
  assign n35918 = pi18 ? n35917 : ~n697;
  assign n35919 = pi17 ? n32 : n35918;
  assign n35920 = pi16 ? n32 : n35919;
  assign n35921 = pi15 ? n35916 : n35920;
  assign n35922 = pi14 ? n35911 : n35921;
  assign n35923 = pi13 ? n32 : n35922;
  assign n35924 = pi12 ? n35907 : n35923;
  assign n35925 = pi11 ? n35894 : n35924;
  assign n35926 = pi20 ? n32 : ~n18832;
  assign n35927 = pi19 ? n35926 : ~n28965;
  assign n35928 = pi18 ? n35927 : ~n1750;
  assign n35929 = pi17 ? n32 : n35928;
  assign n35930 = pi16 ? n32 : n35929;
  assign n35931 = pi18 ? n20172 : ~n702;
  assign n35932 = pi17 ? n32 : n35931;
  assign n35933 = pi16 ? n32 : n35932;
  assign n35934 = pi15 ? n35930 : n35933;
  assign n35935 = pi15 ? n20614 : n32;
  assign n35936 = pi14 ? n35934 : n35935;
  assign n35937 = pi18 ? n32 : n33508;
  assign n35938 = pi17 ? n32 : n35937;
  assign n35939 = pi16 ? n32 : n35938;
  assign n35940 = pi15 ? n35939 : n14131;
  assign n35941 = pi14 ? n32 : n35940;
  assign n35942 = pi13 ? n35936 : n35941;
  assign n35943 = pi15 ? n14131 : n34404;
  assign n35944 = pi19 ? n349 : ~n1105;
  assign n35945 = pi18 ? n32 : n35944;
  assign n35946 = pi17 ? n32 : n35945;
  assign n35947 = pi16 ? n32 : n35946;
  assign n35948 = pi19 ? n23895 : ~n6988;
  assign n35949 = pi18 ? n35948 : ~n13318;
  assign n35950 = pi17 ? n2954 : ~n35949;
  assign n35951 = pi16 ? n32 : n35950;
  assign n35952 = pi15 ? n35947 : n35951;
  assign n35953 = pi14 ? n35943 : n35952;
  assign n35954 = pi19 ? n23895 : n9037;
  assign n35955 = pi18 ? n35954 : ~n23514;
  assign n35956 = pi17 ? n2954 : ~n35955;
  assign n35957 = pi16 ? n32 : n35956;
  assign n35958 = pi18 ? n32 : n32315;
  assign n35959 = pi20 ? n274 : ~n2358;
  assign n35960 = pi20 ? n287 : n6050;
  assign n35961 = pi19 ? n35959 : ~n35960;
  assign n35962 = pi18 ? n35961 : ~n13335;
  assign n35963 = pi17 ? n35958 : ~n35962;
  assign n35964 = pi16 ? n32 : n35963;
  assign n35965 = pi15 ? n35957 : n35964;
  assign n35966 = pi19 ? n4126 : ~n429;
  assign n35967 = pi18 ? n35966 : n508;
  assign n35968 = pi17 ? n32 : ~n35967;
  assign n35969 = pi16 ? n32 : n35968;
  assign n35970 = pi19 ? n4670 : n429;
  assign n35971 = pi18 ? n35970 : ~n508;
  assign n35972 = pi17 ? n32 : n35971;
  assign n35973 = pi16 ? n32 : n35972;
  assign n35974 = pi15 ? n35969 : n35973;
  assign n35975 = pi14 ? n35965 : n35974;
  assign n35976 = pi13 ? n35953 : n35975;
  assign n35977 = pi12 ? n35942 : n35976;
  assign n35978 = pi15 ? n13040 : n13629;
  assign n35979 = pi14 ? n34965 : n35978;
  assign n35980 = pi19 ? n32 : n3524;
  assign n35981 = pi18 ? n32 : n35980;
  assign n35982 = pi17 ? n32 : n35981;
  assign n35983 = pi18 ? n32 : n6063;
  assign n35984 = pi17 ? n29510 : n35983;
  assign n35985 = pi16 ? n35982 : ~n35984;
  assign n35986 = pi15 ? n13913 : n35985;
  assign n35987 = pi18 ? n35270 : n32;
  assign n35988 = pi17 ? n32 : n35987;
  assign n35989 = pi16 ? n32 : n35988;
  assign n35990 = pi18 ? n268 : ~n6059;
  assign n35991 = pi17 ? n35990 : ~n2325;
  assign n35992 = pi16 ? n32 : n35991;
  assign n35993 = pi15 ? n35989 : n35992;
  assign n35994 = pi14 ? n35986 : n35993;
  assign n35995 = pi13 ? n35979 : n35994;
  assign n35996 = pi20 ? n246 : ~n342;
  assign n35997 = pi19 ? n9822 : ~n35996;
  assign n35998 = pi18 ? n32 : n35997;
  assign n35999 = pi19 ? n5371 : ~n18722;
  assign n36000 = pi18 ? n35999 : n237;
  assign n36001 = pi17 ? n35998 : ~n36000;
  assign n36002 = pi16 ? n32 : n36001;
  assign n36003 = pi15 ? n36002 : n32;
  assign n36004 = pi14 ? n36003 : n20969;
  assign n36005 = pi19 ? n531 : n343;
  assign n36006 = pi18 ? n32 : n36005;
  assign n36007 = pi17 ? n32 : n36006;
  assign n36008 = pi18 ? n32 : ~n6059;
  assign n36009 = pi17 ? n32 : n36008;
  assign n36010 = pi16 ? n36007 : ~n36009;
  assign n36011 = pi15 ? n32 : n36010;
  assign n36012 = pi19 ? n4670 : ~n5371;
  assign n36013 = pi18 ? n209 : ~n36012;
  assign n36014 = pi17 ? n32 : n36013;
  assign n36015 = pi18 ? n247 : ~n237;
  assign n36016 = pi17 ? n24225 : ~n36015;
  assign n36017 = pi16 ? n36014 : ~n36016;
  assign n36018 = pi19 ? n9007 : ~n813;
  assign n36019 = pi18 ? n209 : ~n36018;
  assign n36020 = pi17 ? n32 : n36019;
  assign n36021 = pi16 ? n36020 : ~n1808;
  assign n36022 = pi15 ? n36017 : n36021;
  assign n36023 = pi14 ? n36011 : n36022;
  assign n36024 = pi13 ? n36004 : n36023;
  assign n36025 = pi12 ? n35995 : n36024;
  assign n36026 = pi11 ? n35977 : n36025;
  assign n36027 = pi10 ? n35925 : n36026;
  assign n36028 = pi09 ? n32 : n36027;
  assign n36029 = pi13 ? n35884 : n24237;
  assign n36030 = pi14 ? n24237 : n32;
  assign n36031 = pi13 ? n36030 : n35892;
  assign n36032 = pi12 ? n36029 : n36031;
  assign n36033 = pi15 ? n14397 : n35449;
  assign n36034 = pi14 ? n35900 : n36033;
  assign n36035 = pi13 ? n35899 : n36034;
  assign n36036 = pi12 ? n36035 : n35923;
  assign n36037 = pi11 ? n36032 : n36036;
  assign n36038 = pi19 ? n35926 : ~n19249;
  assign n36039 = pi18 ? n36038 : ~n1750;
  assign n36040 = pi17 ? n32 : n36039;
  assign n36041 = pi16 ? n32 : n36040;
  assign n36042 = pi19 ? n32 : ~n53;
  assign n36043 = pi18 ? n20172 : ~n36042;
  assign n36044 = pi17 ? n32 : n36043;
  assign n36045 = pi16 ? n32 : n36044;
  assign n36046 = pi15 ? n36041 : n36045;
  assign n36047 = pi14 ? n36046 : n35935;
  assign n36048 = pi15 ? n22434 : n25346;
  assign n36049 = pi14 ? n32 : n36048;
  assign n36050 = pi13 ? n36047 : n36049;
  assign n36051 = pi15 ? n14138 : n34404;
  assign n36052 = pi15 ? n13620 : n35951;
  assign n36053 = pi14 ? n36051 : n36052;
  assign n36054 = pi18 ? n32 : n2387;
  assign n36055 = pi20 ? n287 : n220;
  assign n36056 = pi19 ? n2358 : n36055;
  assign n36057 = pi18 ? n36056 : n13335;
  assign n36058 = pi17 ? n36054 : n36057;
  assign n36059 = pi16 ? n32 : n36058;
  assign n36060 = pi15 ? n35957 : n36059;
  assign n36061 = pi14 ? n36060 : n35974;
  assign n36062 = pi13 ? n36053 : n36061;
  assign n36063 = pi12 ? n36050 : n36062;
  assign n36064 = pi16 ? n2958 : ~n35984;
  assign n36065 = pi15 ? n13913 : n36064;
  assign n36066 = pi14 ? n36065 : n35993;
  assign n36067 = pi13 ? n35979 : n36066;
  assign n36068 = pi19 ? n531 : ~n10632;
  assign n36069 = pi18 ? n32 : n36068;
  assign n36070 = pi17 ? n32 : n36069;
  assign n36071 = pi16 ? n36070 : ~n36009;
  assign n36072 = pi15 ? n32 : n36071;
  assign n36073 = pi20 ? n915 : n266;
  assign n36074 = pi19 ? n4670 : n36073;
  assign n36075 = pi18 ? n209 : ~n36074;
  assign n36076 = pi17 ? n32 : n36075;
  assign n36077 = pi16 ? n36076 : ~n36016;
  assign n36078 = pi19 ? n9007 : n358;
  assign n36079 = pi18 ? n209 : ~n36078;
  assign n36080 = pi17 ? n32 : n36079;
  assign n36081 = pi16 ? n36080 : ~n1808;
  assign n36082 = pi15 ? n36077 : n36081;
  assign n36083 = pi14 ? n36072 : n36082;
  assign n36084 = pi13 ? n36004 : n36083;
  assign n36085 = pi12 ? n36067 : n36084;
  assign n36086 = pi11 ? n36063 : n36085;
  assign n36087 = pi10 ? n36037 : n36086;
  assign n36088 = pi09 ? n32 : n36087;
  assign n36089 = pi08 ? n36028 : n36088;
  assign n36090 = pi14 ? n24368 : n24573;
  assign n36091 = pi13 ? n36090 : n24237;
  assign n36092 = pi19 ? n519 : ~n589;
  assign n36093 = pi18 ? n32 : n36092;
  assign n36094 = pi17 ? n32 : n36093;
  assign n36095 = pi16 ? n32 : n36094;
  assign n36096 = pi15 ? n16105 : n36095;
  assign n36097 = pi19 ? n507 : ~n589;
  assign n36098 = pi18 ? n32 : n36097;
  assign n36099 = pi17 ? n32 : n36098;
  assign n36100 = pi16 ? n32 : n36099;
  assign n36101 = pi15 ? n36100 : n24511;
  assign n36102 = pi14 ? n36096 : n36101;
  assign n36103 = pi13 ? n36030 : n36102;
  assign n36104 = pi12 ? n36091 : n36103;
  assign n36105 = pi15 ? n23484 : n14917;
  assign n36106 = pi14 ? n25779 : n36105;
  assign n36107 = pi18 ? n32 : n6600;
  assign n36108 = pi17 ? n32 : n36107;
  assign n36109 = pi16 ? n32 : n36108;
  assign n36110 = pi15 ? n36109 : n24247;
  assign n36111 = pi15 ? n16105 : n23484;
  assign n36112 = pi14 ? n36110 : n36111;
  assign n36113 = pi13 ? n36106 : n36112;
  assign n36114 = pi15 ? n32 : n33970;
  assign n36115 = pi19 ? n4964 : n321;
  assign n36116 = pi18 ? n36115 : ~n697;
  assign n36117 = pi17 ? n32 : n36116;
  assign n36118 = pi16 ? n32 : n36117;
  assign n36119 = pi19 ? n531 : ~n5694;
  assign n36120 = pi18 ? n36119 : ~n697;
  assign n36121 = pi17 ? n32 : n36120;
  assign n36122 = pi16 ? n32 : n36121;
  assign n36123 = pi15 ? n36118 : n36122;
  assign n36124 = pi14 ? n36114 : n36123;
  assign n36125 = pi13 ? n32 : n36124;
  assign n36126 = pi12 ? n36113 : n36125;
  assign n36127 = pi11 ? n36104 : n36126;
  assign n36128 = pi18 ? n30632 : ~n4428;
  assign n36129 = pi17 ? n32 : n36128;
  assign n36130 = pi16 ? n32 : n36129;
  assign n36131 = pi15 ? n36122 : n36130;
  assign n36132 = pi18 ? n20172 : n13070;
  assign n36133 = pi17 ? n32 : n36132;
  assign n36134 = pi16 ? n32 : n36133;
  assign n36135 = pi15 ? n36134 : n32;
  assign n36136 = pi14 ? n36131 : n36135;
  assign n36137 = pi18 ? n5158 : n6059;
  assign n36138 = pi17 ? n32 : n36137;
  assign n36139 = pi16 ? n32 : n36138;
  assign n36140 = pi15 ? n36139 : n32;
  assign n36141 = pi20 ? n2385 : ~n266;
  assign n36142 = pi19 ? n36141 : ~n617;
  assign n36143 = pi18 ? n32 : n36142;
  assign n36144 = pi17 ? n32 : n36143;
  assign n36145 = pi16 ? n32 : n36144;
  assign n36146 = pi19 ? n3507 : ~n617;
  assign n36147 = pi18 ? n32 : n36146;
  assign n36148 = pi17 ? n32 : n36147;
  assign n36149 = pi16 ? n32 : n36148;
  assign n36150 = pi15 ? n36145 : n36149;
  assign n36151 = pi14 ? n36140 : n36150;
  assign n36152 = pi13 ? n36136 : n36151;
  assign n36153 = pi18 ? n6114 : n25787;
  assign n36154 = pi17 ? n32 : n36153;
  assign n36155 = pi16 ? n32 : n36154;
  assign n36156 = pi15 ? n36149 : n36155;
  assign n36157 = pi18 ? n16847 : n6163;
  assign n36158 = pi17 ? n32 : n36157;
  assign n36159 = pi16 ? n32 : n36158;
  assign n36160 = pi15 ? n25790 : n36159;
  assign n36161 = pi14 ? n36156 : n36160;
  assign n36162 = pi19 ? n32 : ~n321;
  assign n36163 = pi18 ? n36162 : n6163;
  assign n36164 = pi17 ? n32 : n36163;
  assign n36165 = pi16 ? n32 : n36164;
  assign n36166 = pi18 ? n222 : n5357;
  assign n36167 = pi17 ? n32 : n36166;
  assign n36168 = pi16 ? n32 : n36167;
  assign n36169 = pi15 ? n36165 : n36168;
  assign n36170 = pi18 ? n14873 : n508;
  assign n36171 = pi17 ? n32 : ~n36170;
  assign n36172 = pi16 ? n32 : n36171;
  assign n36173 = pi15 ? n36172 : n12515;
  assign n36174 = pi14 ? n36169 : n36173;
  assign n36175 = pi13 ? n36161 : n36174;
  assign n36176 = pi12 ? n36152 : n36175;
  assign n36177 = pi15 ? n23189 : n13626;
  assign n36178 = pi14 ? n34965 : n36177;
  assign n36179 = pi18 ? n32 : n28053;
  assign n36180 = pi17 ? n32 : n36179;
  assign n36181 = pi20 ? n2180 : n9194;
  assign n36182 = pi20 ? n17652 : n9491;
  assign n36183 = pi19 ? n36181 : ~n36182;
  assign n36184 = pi20 ? n310 : ~n321;
  assign n36185 = pi19 ? n18502 : ~n36184;
  assign n36186 = pi18 ? n36183 : ~n36185;
  assign n36187 = pi19 ? n35496 : n4342;
  assign n36188 = pi18 ? n36187 : ~n32;
  assign n36189 = pi17 ? n36186 : n36188;
  assign n36190 = pi16 ? n36180 : ~n36189;
  assign n36191 = pi15 ? n14143 : n36190;
  assign n36192 = pi19 ? n349 : ~n9007;
  assign n36193 = pi18 ? n32 : n36192;
  assign n36194 = pi17 ? n36193 : ~n2325;
  assign n36195 = pi16 ? n32 : n36194;
  assign n36196 = pi15 ? n35989 : n36195;
  assign n36197 = pi14 ? n36191 : n36196;
  assign n36198 = pi13 ? n36178 : n36197;
  assign n36199 = pi20 ? n246 : ~n1076;
  assign n36200 = pi19 ? n9822 : ~n36199;
  assign n36201 = pi18 ? n32 : n36200;
  assign n36202 = pi20 ? n1385 : ~n266;
  assign n36203 = pi19 ? n36202 : n19601;
  assign n36204 = pi18 ? n36203 : n237;
  assign n36205 = pi17 ? n36201 : ~n36204;
  assign n36206 = pi16 ? n32 : n36205;
  assign n36207 = pi15 ? n36206 : n32;
  assign n36208 = pi14 ? n36207 : n32;
  assign n36209 = pi19 ? n531 : n32340;
  assign n36210 = pi18 ? n32 : n36209;
  assign n36211 = pi17 ? n32 : n36210;
  assign n36212 = pi17 ? n24345 : ~n32;
  assign n36213 = pi16 ? n36211 : ~n36212;
  assign n36214 = pi15 ? n32 : n36213;
  assign n36215 = pi20 ? n321 : n17669;
  assign n36216 = pi19 ? n4670 : ~n36215;
  assign n36217 = pi18 ? n341 : ~n36216;
  assign n36218 = pi17 ? n32 : n36217;
  assign n36219 = pi18 ? n24352 : n359;
  assign n36220 = pi17 ? n24351 : ~n36219;
  assign n36221 = pi16 ? n36218 : ~n36220;
  assign n36222 = pi18 ? n341 : ~n23571;
  assign n36223 = pi17 ? n32 : n36222;
  assign n36224 = pi16 ? n36223 : ~n1808;
  assign n36225 = pi15 ? n36221 : n36224;
  assign n36226 = pi14 ? n36214 : n36225;
  assign n36227 = pi13 ? n36208 : n36226;
  assign n36228 = pi12 ? n36198 : n36227;
  assign n36229 = pi11 ? n36176 : n36228;
  assign n36230 = pi10 ? n36127 : n36229;
  assign n36231 = pi09 ? n32 : n36230;
  assign n36232 = pi13 ? n36090 : n24367;
  assign n36233 = pi15 ? n24504 : n36095;
  assign n36234 = pi14 ? n36233 : n36101;
  assign n36235 = pi13 ? n24371 : n36234;
  assign n36236 = pi12 ? n36232 : n36235;
  assign n36237 = pi15 ? n16105 : n24382;
  assign n36238 = pi15 ? n24718 : n14917;
  assign n36239 = pi14 ? n36237 : n36238;
  assign n36240 = pi13 ? n36239 : n36112;
  assign n36241 = pi18 ? n32 : n6826;
  assign n36242 = pi17 ? n32 : n36241;
  assign n36243 = pi16 ? n32 : n36242;
  assign n36244 = pi15 ? n32 : n36243;
  assign n36245 = pi18 ? n36119 : ~n962;
  assign n36246 = pi17 ? n32 : n36245;
  assign n36247 = pi16 ? n32 : n36246;
  assign n36248 = pi15 ? n36118 : n36247;
  assign n36249 = pi14 ? n36244 : n36248;
  assign n36250 = pi13 ? n32 : n36249;
  assign n36251 = pi12 ? n36240 : n36250;
  assign n36252 = pi11 ? n36236 : n36251;
  assign n36253 = pi20 ? n18415 : ~n32;
  assign n36254 = pi19 ? n275 : ~n36253;
  assign n36255 = pi18 ? n36254 : n6059;
  assign n36256 = pi17 ? n32 : n36255;
  assign n36257 = pi16 ? n32 : n36256;
  assign n36258 = pi15 ? n36257 : n32;
  assign n36259 = pi14 ? n36258 : n36150;
  assign n36260 = pi13 ? n36136 : n36259;
  assign n36261 = pi12 ? n36260 : n36175;
  assign n36262 = pi15 ? n13040 : n22958;
  assign n36263 = pi14 ? n36262 : n36177;
  assign n36264 = pi16 ? n17486 : ~n36189;
  assign n36265 = pi15 ? n14143 : n36264;
  assign n36266 = pi14 ? n36265 : n36196;
  assign n36267 = pi13 ? n36263 : n36266;
  assign n36268 = pi16 ? n36007 : ~n36212;
  assign n36269 = pi15 ? n32 : n36268;
  assign n36270 = pi19 ? n4670 : ~n6997;
  assign n36271 = pi18 ? n341 : ~n36270;
  assign n36272 = pi17 ? n32 : n36271;
  assign n36273 = pi16 ? n36272 : ~n36220;
  assign n36274 = pi15 ? n36273 : n29601;
  assign n36275 = pi14 ? n36269 : n36274;
  assign n36276 = pi13 ? n36208 : n36275;
  assign n36277 = pi12 ? n36267 : n36276;
  assign n36278 = pi11 ? n36261 : n36277;
  assign n36279 = pi10 ? n36252 : n36278;
  assign n36280 = pi09 ? n32 : n36279;
  assign n36281 = pi08 ? n36231 : n36280;
  assign n36282 = pi07 ? n36089 : n36281;
  assign n36283 = pi14 ? n24563 : n25775;
  assign n36284 = pi13 ? n36283 : n24367;
  assign n36285 = pi15 ? n32 : n16105;
  assign n36286 = pi14 ? n24370 : n36285;
  assign n36287 = pi15 ? n24504 : n24640;
  assign n36288 = pi14 ? n36287 : n24640;
  assign n36289 = pi13 ? n36286 : n36288;
  assign n36290 = pi12 ? n36284 : n36289;
  assign n36291 = pi15 ? n26078 : n15244;
  assign n36292 = pi14 ? n36291 : n24719;
  assign n36293 = pi19 ? n1464 : ~n349;
  assign n36294 = pi18 ? n32 : n36293;
  assign n36295 = pi17 ? n32 : n36294;
  assign n36296 = pi16 ? n32 : n36295;
  assign n36297 = pi15 ? n24247 : n36296;
  assign n36298 = pi19 ? n750 : ~n236;
  assign n36299 = pi18 ? n32 : n36298;
  assign n36300 = pi17 ? n32 : n36299;
  assign n36301 = pi16 ? n32 : n36300;
  assign n36302 = pi15 ? n15244 : n36301;
  assign n36303 = pi14 ? n36297 : n36302;
  assign n36304 = pi13 ? n36292 : n36303;
  assign n36305 = pi14 ? n21217 : n32;
  assign n36306 = pi19 ? n32 : n26777;
  assign n36307 = pi18 ? n32 : n36306;
  assign n36308 = pi17 ? n32 : n36307;
  assign n36309 = pi16 ? n32 : n36308;
  assign n36310 = pi18 ? n323 : ~n962;
  assign n36311 = pi17 ? n32 : n36310;
  assign n36312 = pi16 ? n32 : n36311;
  assign n36313 = pi15 ? n36309 : n36312;
  assign n36314 = pi18 ? n532 : ~n962;
  assign n36315 = pi17 ? n32 : n36314;
  assign n36316 = pi16 ? n32 : n36315;
  assign n36317 = pi18 ? n532 : ~n8471;
  assign n36318 = pi17 ? n32 : n36317;
  assign n36319 = pi16 ? n32 : n36318;
  assign n36320 = pi15 ? n36316 : n36319;
  assign n36321 = pi14 ? n36313 : n36320;
  assign n36322 = pi13 ? n36305 : n36321;
  assign n36323 = pi12 ? n36304 : n36322;
  assign n36324 = pi11 ? n36290 : n36323;
  assign n36325 = pi18 ? n16449 : n13080;
  assign n36326 = pi17 ? n32 : n36325;
  assign n36327 = pi16 ? n32 : n36326;
  assign n36328 = pi15 ? n36316 : n36327;
  assign n36329 = pi19 ? n6342 : n32;
  assign n36330 = pi18 ? n32 : n36329;
  assign n36331 = pi17 ? n32 : n36330;
  assign n36332 = pi16 ? n32 : n36331;
  assign n36333 = pi15 ? n36332 : n32;
  assign n36334 = pi14 ? n36328 : n36333;
  assign n36335 = pi18 ? n24942 : n5005;
  assign n36336 = pi17 ? n32 : n36335;
  assign n36337 = pi16 ? n32 : n36336;
  assign n36338 = pi19 ? n3524 : ~n617;
  assign n36339 = pi18 ? n32 : n36338;
  assign n36340 = pi17 ? n32 : n36339;
  assign n36341 = pi16 ? n32 : n36340;
  assign n36342 = pi15 ? n36337 : n36341;
  assign n36343 = pi15 ? n36341 : n23832;
  assign n36344 = pi14 ? n36342 : n36343;
  assign n36345 = pi13 ? n36334 : n36344;
  assign n36346 = pi19 ? n531 : ~n2614;
  assign n36347 = pi18 ? n32 : n36346;
  assign n36348 = pi17 ? n32 : n36347;
  assign n36349 = pi16 ? n32 : n36348;
  assign n36350 = pi19 ? n1464 : ~n4391;
  assign n36351 = pi18 ? n36350 : n34613;
  assign n36352 = pi17 ? n32 : n36351;
  assign n36353 = pi16 ? n32 : n36352;
  assign n36354 = pi15 ? n36353 : n14138;
  assign n36355 = pi14 ? n36349 : n36354;
  assign n36356 = pi18 ? n36350 : n13901;
  assign n36357 = pi17 ? n32 : n36356;
  assign n36358 = pi16 ? n32 : n36357;
  assign n36359 = pi15 ? n36358 : n13629;
  assign n36360 = pi19 ? n1490 : ~n18041;
  assign n36361 = pi18 ? n36360 : ~n508;
  assign n36362 = pi17 ? n32 : n36361;
  assign n36363 = pi16 ? n32 : n36362;
  assign n36364 = pi19 ? n1464 : n519;
  assign n36365 = pi18 ? n36364 : ~n595;
  assign n36366 = pi17 ? n32 : n36365;
  assign n36367 = pi16 ? n32 : n36366;
  assign n36368 = pi15 ? n36363 : n36367;
  assign n36369 = pi14 ? n36359 : n36368;
  assign n36370 = pi13 ? n36355 : n36369;
  assign n36371 = pi12 ? n36345 : n36370;
  assign n36372 = pi14 ? n21853 : n24547;
  assign n36373 = pi19 ? n1464 : n322;
  assign n36374 = pi20 ? n220 : n16008;
  assign n36375 = pi19 ? n36374 : ~n32;
  assign n36376 = pi18 ? n36373 : ~n36375;
  assign n36377 = pi17 ? n32 : n36376;
  assign n36378 = pi16 ? n32 : n36377;
  assign n36379 = pi18 ? n940 : n9012;
  assign n36380 = pi17 ? n32 : n36379;
  assign n36381 = pi16 ? n32 : n36380;
  assign n36382 = pi15 ? n36378 : n36381;
  assign n36383 = pi19 ? n531 : n5688;
  assign n36384 = pi18 ? n36383 : ~n344;
  assign n36385 = pi17 ? n16848 : n36384;
  assign n36386 = pi16 ? n32 : n36385;
  assign n36387 = pi19 ? n5707 : ~n531;
  assign n36388 = pi18 ? n36387 : n532;
  assign n36389 = pi17 ? n8653 : ~n36388;
  assign n36390 = pi16 ? n32 : n36389;
  assign n36391 = pi15 ? n36386 : n36390;
  assign n36392 = pi14 ? n36382 : n36391;
  assign n36393 = pi13 ? n36372 : n36392;
  assign n36394 = pi18 ? n702 : ~n34250;
  assign n36395 = pi18 ? n22889 : n32;
  assign n36396 = pi17 ? n36394 : n36395;
  assign n36397 = pi16 ? n32 : n36396;
  assign n36398 = pi15 ? n36397 : n32;
  assign n36399 = pi18 ? n24025 : n4343;
  assign n36400 = pi17 ? n32 : n36399;
  assign n36401 = pi16 ? n32 : n36400;
  assign n36402 = pi19 ? n32 : ~n16002;
  assign n36403 = pi18 ? n32 : n36402;
  assign n36404 = pi19 ? n4721 : n208;
  assign n36405 = pi18 ? n36404 : n4343;
  assign n36406 = pi17 ? n36403 : n36405;
  assign n36407 = pi16 ? n32 : n36406;
  assign n36408 = pi15 ? n36401 : n36407;
  assign n36409 = pi14 ? n36398 : n36408;
  assign n36410 = pi18 ? n209 : n940;
  assign n36411 = pi17 ? n32 : n36410;
  assign n36412 = pi17 ? n1028 : ~n14611;
  assign n36413 = pi16 ? n36411 : ~n36412;
  assign n36414 = pi15 ? n212 : n36413;
  assign n36415 = pi19 ? n32 : n19116;
  assign n36416 = pi18 ? n341 : ~n36415;
  assign n36417 = pi17 ? n32 : n36416;
  assign n36418 = pi17 ? n18482 : n2653;
  assign n36419 = pi16 ? n36417 : ~n36418;
  assign n36420 = pi15 ? n36419 : n35359;
  assign n36421 = pi14 ? n36414 : n36420;
  assign n36422 = pi13 ? n36409 : n36421;
  assign n36423 = pi12 ? n36393 : n36422;
  assign n36424 = pi11 ? n36371 : n36423;
  assign n36425 = pi10 ? n36324 : n36424;
  assign n36426 = pi09 ? n32 : n36425;
  assign n36427 = pi15 ? n16606 : n24495;
  assign n36428 = pi14 ? n24495 : n36427;
  assign n36429 = pi13 ? n36283 : n36428;
  assign n36430 = pi14 ? n24498 : n36285;
  assign n36431 = pi13 ? n36430 : n36288;
  assign n36432 = pi12 ? n36429 : n36431;
  assign n36433 = pi18 ? n323 : ~n4244;
  assign n36434 = pi17 ? n32 : n36433;
  assign n36435 = pi16 ? n32 : n36434;
  assign n36436 = pi15 ? n23574 : n36435;
  assign n36437 = pi14 ? n36436 : n36320;
  assign n36438 = pi13 ? n36305 : n36437;
  assign n36439 = pi12 ? n36304 : n36438;
  assign n36440 = pi11 ? n36432 : n36439;
  assign n36441 = pi18 ? n532 : ~n4244;
  assign n36442 = pi17 ? n32 : n36441;
  assign n36443 = pi16 ? n32 : n36442;
  assign n36444 = pi15 ? n36443 : n36327;
  assign n36445 = pi14 ? n36444 : n36333;
  assign n36446 = pi14 ? n36342 : n23832;
  assign n36447 = pi13 ? n36445 : n36446;
  assign n36448 = pi15 ? n36353 : n25346;
  assign n36449 = pi14 ? n36349 : n36448;
  assign n36450 = pi18 ? n36364 : ~n4098;
  assign n36451 = pi17 ? n32 : n36450;
  assign n36452 = pi16 ? n32 : n36451;
  assign n36453 = pi15 ? n36363 : n36452;
  assign n36454 = pi14 ? n36359 : n36453;
  assign n36455 = pi13 ? n36449 : n36454;
  assign n36456 = pi12 ? n36447 : n36455;
  assign n36457 = pi15 ? n35650 : n24543;
  assign n36458 = pi14 ? n22437 : n36457;
  assign n36459 = pi18 ? n36373 : ~n6019;
  assign n36460 = pi17 ? n32 : n36459;
  assign n36461 = pi16 ? n32 : n36460;
  assign n36462 = pi15 ? n36461 : n36381;
  assign n36463 = pi14 ? n36462 : n36391;
  assign n36464 = pi13 ? n36458 : n36463;
  assign n36465 = pi16 ? n36411 : ~n1355;
  assign n36466 = pi15 ? n212 : n36465;
  assign n36467 = pi18 ? n366 : ~n36415;
  assign n36468 = pi17 ? n32 : n36467;
  assign n36469 = pi17 ? n19432 : n2119;
  assign n36470 = pi16 ? n36468 : ~n36469;
  assign n36471 = pi15 ? n36470 : n35359;
  assign n36472 = pi14 ? n36466 : n36471;
  assign n36473 = pi13 ? n36409 : n36472;
  assign n36474 = pi12 ? n36464 : n36473;
  assign n36475 = pi11 ? n36456 : n36474;
  assign n36476 = pi10 ? n36440 : n36475;
  assign n36477 = pi09 ? n32 : n36476;
  assign n36478 = pi08 ? n36426 : n36477;
  assign n36479 = pi14 ? n24627 : n16607;
  assign n36480 = pi13 ? n36479 : n16606;
  assign n36481 = pi15 ? n24247 : n24700;
  assign n36482 = pi14 ? n36481 : n24700;
  assign n36483 = pi13 ? n36430 : n36482;
  assign n36484 = pi12 ? n36480 : n36483;
  assign n36485 = pi15 ? n32 : n36100;
  assign n36486 = pi14 ? n36485 : n24504;
  assign n36487 = pi15 ? n15244 : n14917;
  assign n36488 = pi14 ? n24511 : n36487;
  assign n36489 = pi13 ? n36486 : n36488;
  assign n36490 = pi14 ? n32 : n36285;
  assign n36491 = pi18 ? n323 : ~n697;
  assign n36492 = pi17 ? n32 : n36491;
  assign n36493 = pi16 ? n32 : n36492;
  assign n36494 = pi15 ? n23933 : n36493;
  assign n36495 = pi18 ? n532 : ~n697;
  assign n36496 = pi17 ? n32 : n36495;
  assign n36497 = pi16 ? n32 : n36496;
  assign n36498 = pi18 ? n605 : ~n6235;
  assign n36499 = pi17 ? n32 : n36498;
  assign n36500 = pi16 ? n32 : n36499;
  assign n36501 = pi15 ? n36497 : n36500;
  assign n36502 = pi14 ? n36494 : n36501;
  assign n36503 = pi13 ? n36490 : n36502;
  assign n36504 = pi12 ? n36489 : n36503;
  assign n36505 = pi11 ? n36484 : n36504;
  assign n36506 = pi18 ? n605 : ~n697;
  assign n36507 = pi17 ? n32 : n36506;
  assign n36508 = pi16 ? n32 : n36507;
  assign n36509 = pi19 ? n594 : n18211;
  assign n36510 = pi20 ? n321 : n357;
  assign n36511 = pi19 ? n36510 : n32;
  assign n36512 = pi18 ? n36509 : n36511;
  assign n36513 = pi17 ? n32 : n36512;
  assign n36514 = pi16 ? n32 : n36513;
  assign n36515 = pi15 ? n36508 : n36514;
  assign n36516 = pi19 ? n594 : n23895;
  assign n36517 = pi18 ? n36516 : n248;
  assign n36518 = pi17 ? n32 : n36517;
  assign n36519 = pi16 ? n32 : n36518;
  assign n36520 = pi15 ? n36519 : n32;
  assign n36521 = pi14 ? n36515 : n36520;
  assign n36522 = pi19 ? n594 : n11879;
  assign n36523 = pi19 ? n33674 : ~n236;
  assign n36524 = pi18 ? n36522 : n36523;
  assign n36525 = pi17 ? n32 : n36524;
  assign n36526 = pi16 ? n32 : n36525;
  assign n36527 = pi15 ? n36526 : n14580;
  assign n36528 = pi14 ? n36527 : n14580;
  assign n36529 = pi13 ? n36521 : n36528;
  assign n36530 = pi19 ? n4721 : ~n2614;
  assign n36531 = pi18 ? n32 : n36530;
  assign n36532 = pi17 ? n32 : n36531;
  assign n36533 = pi16 ? n32 : n36532;
  assign n36534 = pi15 ? n36533 : n25346;
  assign n36535 = pi14 ? n36349 : n36534;
  assign n36536 = pi15 ? n13904 : n33939;
  assign n36537 = pi18 ? n6581 : ~n508;
  assign n36538 = pi17 ? n32 : n36537;
  assign n36539 = pi16 ? n32 : n36538;
  assign n36540 = pi18 ? n6145 : ~n595;
  assign n36541 = pi17 ? n32 : n36540;
  assign n36542 = pi16 ? n32 : n36541;
  assign n36543 = pi15 ? n36539 : n36542;
  assign n36544 = pi14 ? n36536 : n36543;
  assign n36545 = pi13 ? n36535 : n36544;
  assign n36546 = pi12 ? n36529 : n36545;
  assign n36547 = pi15 ? n35650 : n14593;
  assign n36548 = pi14 ? n22437 : n36547;
  assign n36549 = pi18 ? n322 : ~n605;
  assign n36550 = pi17 ? n32 : n36549;
  assign n36551 = pi16 ? n32 : n36550;
  assign n36552 = pi17 ? n32 : n32932;
  assign n36553 = pi16 ? n32 : n36552;
  assign n36554 = pi15 ? n36551 : n36553;
  assign n36555 = pi17 ? n16848 : n21271;
  assign n36556 = pi16 ? n32 : n36555;
  assign n36557 = pi19 ? n32 : ~n247;
  assign n36558 = pi18 ? n32 : n36557;
  assign n36559 = pi19 ? n4342 : ~n531;
  assign n36560 = pi18 ? n36559 : n532;
  assign n36561 = pi17 ? n36558 : ~n36560;
  assign n36562 = pi16 ? n32 : n36561;
  assign n36563 = pi15 ? n36556 : n36562;
  assign n36564 = pi14 ? n36554 : n36563;
  assign n36565 = pi13 ? n36548 : n36564;
  assign n36566 = pi19 ? n1508 : ~n342;
  assign n36567 = pi18 ? n2684 : ~n36566;
  assign n36568 = pi19 ? n32733 : n16431;
  assign n36569 = pi18 ? n36568 : n32;
  assign n36570 = pi17 ? n36567 : n36569;
  assign n36571 = pi16 ? n32 : n36570;
  assign n36572 = pi15 ? n36571 : n32;
  assign n36573 = pi18 ? n32 : n10078;
  assign n36574 = pi19 ? n29033 : n6057;
  assign n36575 = pi18 ? n36574 : n4343;
  assign n36576 = pi17 ? n36573 : n36575;
  assign n36577 = pi16 ? n32 : n36576;
  assign n36578 = pi19 ? n32 : ~n18497;
  assign n36579 = pi18 ? n32 : n36578;
  assign n36580 = pi19 ? n247 : ~n207;
  assign n36581 = pi18 ? n36580 : ~n4343;
  assign n36582 = pi17 ? n36579 : ~n36581;
  assign n36583 = pi16 ? n32 : n36582;
  assign n36584 = pi15 ? n36577 : n36583;
  assign n36585 = pi14 ? n36572 : n36584;
  assign n36586 = pi18 ? n341 : n940;
  assign n36587 = pi17 ? n32 : n36586;
  assign n36588 = pi20 ? n266 : n2358;
  assign n36589 = pi19 ? n36588 : ~n32;
  assign n36590 = pi18 ? n36589 : ~n32;
  assign n36591 = pi17 ? n36590 : ~n32;
  assign n36592 = pi16 ? n36587 : ~n36591;
  assign n36593 = pi15 ? n553 : n36592;
  assign n36594 = pi18 ? n209 : ~n16847;
  assign n36595 = pi17 ? n32 : n36594;
  assign n36596 = pi20 ? n266 : n17665;
  assign n36597 = pi19 ? n36596 : n32;
  assign n36598 = pi18 ? n36597 : n32;
  assign n36599 = pi17 ? n36598 : n2119;
  assign n36600 = pi16 ? n36595 : ~n36599;
  assign n36601 = pi16 ? n1233 : ~n2120;
  assign n36602 = pi15 ? n36600 : n36601;
  assign n36603 = pi14 ? n36593 : n36602;
  assign n36604 = pi13 ? n36585 : n36603;
  assign n36605 = pi12 ? n36565 : n36604;
  assign n36606 = pi11 ? n36546 : n36605;
  assign n36607 = pi10 ? n36505 : n36606;
  assign n36608 = pi09 ? n32 : n36607;
  assign n36609 = pi13 ? n36479 : n16786;
  assign n36610 = pi14 ? n16840 : n36285;
  assign n36611 = pi13 ? n36610 : n36482;
  assign n36612 = pi12 ? n36609 : n36611;
  assign n36613 = pi15 ? n32 : n24705;
  assign n36614 = pi14 ? n36613 : n27308;
  assign n36615 = pi13 ? n36614 : n36488;
  assign n36616 = pi15 ? n24247 : n36493;
  assign n36617 = pi14 ? n36616 : n36501;
  assign n36618 = pi13 ? n36490 : n36617;
  assign n36619 = pi12 ? n36615 : n36618;
  assign n36620 = pi11 ? n36612 : n36619;
  assign n36621 = pi19 ? n33674 : ~n1941;
  assign n36622 = pi18 ? n36522 : n36621;
  assign n36623 = pi17 ? n32 : n36622;
  assign n36624 = pi16 ? n32 : n36623;
  assign n36625 = pi15 ? n36624 : n35030;
  assign n36626 = pi14 ? n36625 : n35030;
  assign n36627 = pi13 ? n36521 : n36626;
  assign n36628 = pi19 ? n4721 : ~n617;
  assign n36629 = pi18 ? n32 : n36628;
  assign n36630 = pi17 ? n32 : n36629;
  assign n36631 = pi16 ? n32 : n36630;
  assign n36632 = pi15 ? n36631 : n25346;
  assign n36633 = pi14 ? n35452 : n36632;
  assign n36634 = pi13 ? n36633 : n36544;
  assign n36635 = pi12 ? n36627 : n36634;
  assign n36636 = pi15 ? n35517 : n14593;
  assign n36637 = pi14 ? n22437 : n36636;
  assign n36638 = pi13 ? n36637 : n36564;
  assign n36639 = pi18 ? n702 : ~n36566;
  assign n36640 = pi17 ? n36639 : n36569;
  assign n36641 = pi16 ? n32 : n36640;
  assign n36642 = pi15 ? n36641 : n32;
  assign n36643 = pi16 ? n17824 : n36582;
  assign n36644 = pi15 ? n36577 : n36643;
  assign n36645 = pi14 ? n36642 : n36644;
  assign n36646 = pi19 ? n5688 : ~n32;
  assign n36647 = pi18 ? n36646 : ~n32;
  assign n36648 = pi17 ? n36647 : ~n32;
  assign n36649 = pi16 ? n36587 : ~n36648;
  assign n36650 = pi15 ? n553 : n36649;
  assign n36651 = pi18 ? n32584 : n32;
  assign n36652 = pi17 ? n36651 : n2119;
  assign n36653 = pi16 ? n36595 : ~n36652;
  assign n36654 = pi15 ? n36653 : n36601;
  assign n36655 = pi14 ? n36650 : n36654;
  assign n36656 = pi13 ? n36645 : n36655;
  assign n36657 = pi12 ? n36638 : n36656;
  assign n36658 = pi11 ? n36635 : n36657;
  assign n36659 = pi10 ? n36620 : n36658;
  assign n36660 = pi09 ? n32 : n36659;
  assign n36661 = pi08 ? n36608 : n36660;
  assign n36662 = pi07 ? n36478 : n36661;
  assign n36663 = pi06 ? n36282 : n36662;
  assign n36664 = pi15 ? n16837 : n16786;
  assign n36665 = pi14 ? n24797 : n36664;
  assign n36666 = pi13 ? n36665 : n16786;
  assign n36667 = pi15 ? n16452 : n16520;
  assign n36668 = pi15 ? n16520 : n16786;
  assign n36669 = pi14 ? n36667 : n36668;
  assign n36670 = pi13 ? n24692 : n36669;
  assign n36671 = pi12 ? n36666 : n36670;
  assign n36672 = pi18 ? n16847 : n24810;
  assign n36673 = pi17 ? n32 : n36672;
  assign n36674 = pi16 ? n32 : n36673;
  assign n36675 = pi15 ? n24237 : n36674;
  assign n36676 = pi14 ? n26994 : n36675;
  assign n36677 = pi15 ? n36100 : n32;
  assign n36678 = pi19 ? n29514 : n32;
  assign n36679 = pi18 ? n5657 : n36678;
  assign n36680 = pi17 ? n32 : n36679;
  assign n36681 = pi16 ? n32 : n36680;
  assign n36682 = pi15 ? n32 : n36681;
  assign n36683 = pi14 ? n36677 : n36682;
  assign n36684 = pi13 ? n36676 : n36683;
  assign n36685 = pi14 ? n32 : n16105;
  assign n36686 = pi18 ? n702 : ~n1758;
  assign n36687 = pi17 ? n32 : n36686;
  assign n36688 = pi16 ? n32 : n36687;
  assign n36689 = pi15 ? n16105 : n36688;
  assign n36690 = pi20 ? n518 : ~n5854;
  assign n36691 = pi19 ? n32 : n36690;
  assign n36692 = pi18 ? n36691 : ~n702;
  assign n36693 = pi17 ? n32 : n36692;
  assign n36694 = pi16 ? n32 : n36693;
  assign n36695 = pi18 ? n32 : ~n697;
  assign n36696 = pi17 ? n32 : n36695;
  assign n36697 = pi16 ? n32 : n36696;
  assign n36698 = pi15 ? n36694 : n36697;
  assign n36699 = pi14 ? n36689 : n36698;
  assign n36700 = pi13 ? n36685 : n36699;
  assign n36701 = pi12 ? n36684 : n36700;
  assign n36702 = pi11 ? n36671 : n36701;
  assign n36703 = pi15 ? n13904 : n32;
  assign n36704 = pi15 ? n32 : n34852;
  assign n36705 = pi14 ? n36703 : n36704;
  assign n36706 = pi15 ? n24018 : n24659;
  assign n36707 = pi14 ? n36706 : n24659;
  assign n36708 = pi13 ? n36705 : n36707;
  assign n36709 = pi19 ? n507 : n24755;
  assign n36710 = pi19 ? n6800 : n236;
  assign n36711 = pi18 ? n36709 : ~n36710;
  assign n36712 = pi17 ? n32 : n36711;
  assign n36713 = pi16 ? n32 : n36712;
  assign n36714 = pi15 ? n24659 : n36713;
  assign n36715 = pi18 ? n16432 : n23440;
  assign n36716 = pi17 ? n32 : n36715;
  assign n36717 = pi16 ? n32 : n36716;
  assign n36718 = pi15 ? n23443 : n36717;
  assign n36719 = pi14 ? n36714 : n36718;
  assign n36720 = pi19 ? n507 : ~n1053;
  assign n36721 = pi19 ? n32331 : n32;
  assign n36722 = pi18 ? n36720 : n36721;
  assign n36723 = pi17 ? n32 : n36722;
  assign n36724 = pi16 ? n32 : n36723;
  assign n36725 = pi20 ? n246 : n5854;
  assign n36726 = pi19 ? n507 : n36725;
  assign n36727 = pi18 ? n36726 : n5335;
  assign n36728 = pi17 ? n32 : n36727;
  assign n36729 = pi16 ? n32 : n36728;
  assign n36730 = pi15 ? n36724 : n36729;
  assign n36731 = pi19 ? n32 : n32090;
  assign n36732 = pi19 ? n813 : n32;
  assign n36733 = pi18 ? n36731 : n36732;
  assign n36734 = pi17 ? n32 : n36733;
  assign n36735 = pi16 ? n32 : n36734;
  assign n36736 = pi14 ? n36730 : n36735;
  assign n36737 = pi13 ? n36719 : n36736;
  assign n36738 = pi12 ? n36708 : n36737;
  assign n36739 = pi15 ? n13913 : n21853;
  assign n36740 = pi15 ? n23094 : n14156;
  assign n36741 = pi14 ? n36739 : n36740;
  assign n36742 = pi18 ? n32 : n28193;
  assign n36743 = pi17 ? n1807 : ~n36742;
  assign n36744 = pi16 ? n32 : n36743;
  assign n36745 = pi15 ? n7359 : n36744;
  assign n36746 = pi18 ? n5335 : n32;
  assign n36747 = pi17 ? n32 : n36746;
  assign n36748 = pi16 ? n32 : n36747;
  assign n36749 = pi19 ? n4406 : ~n4964;
  assign n36750 = pi18 ? n32 : n36749;
  assign n36751 = pi18 ? n1758 : n20788;
  assign n36752 = pi17 ? n36750 : ~n36751;
  assign n36753 = pi16 ? n32 : n36752;
  assign n36754 = pi15 ? n36748 : n36753;
  assign n36755 = pi14 ? n36745 : n36754;
  assign n36756 = pi13 ? n36741 : n36755;
  assign n36757 = pi20 ? n1324 : ~n266;
  assign n36758 = pi19 ? n32 : n36757;
  assign n36759 = pi19 ? n349 : ~n4964;
  assign n36760 = pi18 ? n36758 : ~n36759;
  assign n36761 = pi19 ? n32 : n20925;
  assign n36762 = pi18 ? n36761 : ~n4343;
  assign n36763 = pi17 ? n36760 : ~n36762;
  assign n36764 = pi16 ? n32 : n36763;
  assign n36765 = pi20 ? n7839 : ~n9863;
  assign n36766 = pi19 ? n36765 : n33996;
  assign n36767 = pi18 ? n6767 : ~n36766;
  assign n36768 = pi20 ? n1076 : n246;
  assign n36769 = pi19 ? n36768 : ~n531;
  assign n36770 = pi20 ? n310 : ~n207;
  assign n36771 = pi19 ? n36770 : n32;
  assign n36772 = pi18 ? n36769 : ~n36771;
  assign n36773 = pi17 ? n36767 : ~n36772;
  assign n36774 = pi16 ? n32 : n36773;
  assign n36775 = pi15 ? n36764 : n36774;
  assign n36776 = pi18 ? n23548 : n20788;
  assign n36777 = pi17 ? n32 : ~n36776;
  assign n36778 = pi16 ? n32 : n36777;
  assign n36779 = pi18 ? n24775 : n32;
  assign n36780 = pi17 ? n32 : n36779;
  assign n36781 = pi16 ? n810 : n36780;
  assign n36782 = pi15 ? n36778 : n36781;
  assign n36783 = pi14 ? n36775 : n36782;
  assign n36784 = pi18 ? n209 : ~n532;
  assign n36785 = pi17 ? n32 : n36784;
  assign n36786 = pi18 ? n16847 : ~n237;
  assign n36787 = pi17 ? n32 : n36786;
  assign n36788 = pi16 ? n36785 : n36787;
  assign n36789 = pi18 ? n6645 : n32;
  assign n36790 = pi17 ? n36789 : n30107;
  assign n36791 = pi16 ? n810 : n36790;
  assign n36792 = pi15 ? n36788 : n36791;
  assign n36793 = pi19 ? n5694 : n1757;
  assign n36794 = pi18 ? n36793 : n32;
  assign n36795 = pi17 ? n36794 : n2119;
  assign n36796 = pi16 ? n1135 : ~n36795;
  assign n36797 = pi15 ? n36796 : n36601;
  assign n36798 = pi14 ? n36792 : n36797;
  assign n36799 = pi13 ? n36783 : n36798;
  assign n36800 = pi12 ? n36756 : n36799;
  assign n36801 = pi11 ? n36738 : n36800;
  assign n36802 = pi10 ? n36702 : n36801;
  assign n36803 = pi09 ? n32 : n36802;
  assign n36804 = pi13 ? n36665 : n16837;
  assign n36805 = pi13 ? n24800 : n36669;
  assign n36806 = pi12 ? n36804 : n36805;
  assign n36807 = pi15 ? n32 : n24572;
  assign n36808 = pi18 ? n16847 : n24971;
  assign n36809 = pi17 ? n32 : n36808;
  assign n36810 = pi16 ? n32 : n36809;
  assign n36811 = pi15 ? n24572 : n36810;
  assign n36812 = pi14 ? n36807 : n36811;
  assign n36813 = pi13 ? n36812 : n36683;
  assign n36814 = pi12 ? n36813 : n36700;
  assign n36815 = pi11 ? n36806 : n36814;
  assign n36816 = pi15 ? n24659 : n25466;
  assign n36817 = pi14 ? n36706 : n36816;
  assign n36818 = pi13 ? n36705 : n36817;
  assign n36819 = pi15 ? n25466 : n36713;
  assign n36820 = pi14 ? n36819 : n36718;
  assign n36821 = pi13 ? n36820 : n36736;
  assign n36822 = pi12 ? n36818 : n36821;
  assign n36823 = pi15 ? n22437 : n14156;
  assign n36824 = pi14 ? n36739 : n36823;
  assign n36825 = pi13 ? n36824 : n36755;
  assign n36826 = pi20 ? n9863 : ~n18256;
  assign n36827 = pi19 ? n36826 : n33996;
  assign n36828 = pi18 ? n6767 : ~n36827;
  assign n36829 = pi17 ? n36828 : ~n36772;
  assign n36830 = pi16 ? n32 : n36829;
  assign n36831 = pi15 ? n36764 : n36830;
  assign n36832 = pi14 ? n36831 : n36782;
  assign n36833 = pi17 ? n31079 : n30107;
  assign n36834 = pi16 ? n810 : n36833;
  assign n36835 = pi15 ? n36788 : n36834;
  assign n36836 = pi19 ? n5694 : n1844;
  assign n36837 = pi18 ? n36836 : n32;
  assign n36838 = pi17 ? n36837 : n2119;
  assign n36839 = pi16 ? n1135 : ~n36838;
  assign n36840 = pi15 ? n36839 : n36601;
  assign n36841 = pi14 ? n36835 : n36840;
  assign n36842 = pi13 ? n36832 : n36841;
  assign n36843 = pi12 ? n36825 : n36842;
  assign n36844 = pi11 ? n36822 : n36843;
  assign n36845 = pi10 ? n36815 : n36844;
  assign n36846 = pi09 ? n32 : n36845;
  assign n36847 = pi08 ? n36803 : n36846;
  assign n36848 = pi19 ? n32 : n68;
  assign n36849 = pi18 ? n32 : n36848;
  assign n36850 = pi17 ? n32 : n36849;
  assign n36851 = pi16 ? n32 : n36850;
  assign n36852 = pi15 ? n16899 : n36851;
  assign n36853 = pi14 ? n24962 : n36852;
  assign n36854 = pi13 ? n36853 : n36851;
  assign n36855 = pi15 ? n36851 : n16837;
  assign n36856 = pi14 ? n36855 : n25640;
  assign n36857 = pi14 ? n24874 : n25504;
  assign n36858 = pi13 ? n36856 : n36857;
  assign n36859 = pi12 ? n36854 : n36858;
  assign n36860 = pi18 ? n16847 : n20172;
  assign n36861 = pi17 ? n32 : n36860;
  assign n36862 = pi16 ? n32 : n36861;
  assign n36863 = pi15 ? n16452 : n36862;
  assign n36864 = pi14 ? n24691 : n36863;
  assign n36865 = pi15 ? n15362 : n32;
  assign n36866 = pi19 ? n32 : n32082;
  assign n36867 = pi18 ? n36866 : n32;
  assign n36868 = pi17 ? n32 : n36867;
  assign n36869 = pi16 ? n32 : n36868;
  assign n36870 = pi15 ? n32 : n36869;
  assign n36871 = pi14 ? n36865 : n36870;
  assign n36872 = pi13 ? n36864 : n36871;
  assign n36873 = pi14 ? n32 : n24578;
  assign n36874 = pi20 ? n9488 : ~n207;
  assign n36875 = pi19 ? n36874 : n1757;
  assign n36876 = pi18 ? n36875 : n702;
  assign n36877 = pi17 ? n32 : ~n36876;
  assign n36878 = pi16 ? n32 : n36877;
  assign n36879 = pi19 ? n32 : n18665;
  assign n36880 = pi19 ? n32 : n7014;
  assign n36881 = pi18 ? n36879 : ~n36880;
  assign n36882 = pi17 ? n32 : n36881;
  assign n36883 = pi16 ? n32 : n36882;
  assign n36884 = pi15 ? n36878 : n36883;
  assign n36885 = pi14 ? n36689 : n36884;
  assign n36886 = pi13 ? n36873 : n36885;
  assign n36887 = pi12 ? n36872 : n36886;
  assign n36888 = pi11 ? n36859 : n36887;
  assign n36889 = pi19 ? n4406 : n32;
  assign n36890 = pi18 ? n36879 : n36889;
  assign n36891 = pi17 ? n32 : n36890;
  assign n36892 = pi16 ? n32 : n36891;
  assign n36893 = pi15 ? n36892 : n32;
  assign n36894 = pi15 ? n32 : n35452;
  assign n36895 = pi14 ? n36893 : n36894;
  assign n36896 = pi15 ? n35452 : n24742;
  assign n36897 = pi14 ? n36896 : n24838;
  assign n36898 = pi13 ? n36895 : n36897;
  assign n36899 = pi18 ? n16834 : n20172;
  assign n36900 = pi17 ? n32 : n36899;
  assign n36901 = pi16 ? n32 : n36900;
  assign n36902 = pi15 ? n24838 : n36901;
  assign n36903 = pi20 ? n321 : ~n2358;
  assign n36904 = pi19 ? n32 : n36903;
  assign n36905 = pi19 ? n15405 : ~n32;
  assign n36906 = pi18 ? n36904 : ~n36905;
  assign n36907 = pi17 ? n32 : n36906;
  assign n36908 = pi16 ? n32 : n36907;
  assign n36909 = pi15 ? n23443 : n36908;
  assign n36910 = pi14 ? n36902 : n36909;
  assign n36911 = pi19 ? n507 : ~n1508;
  assign n36912 = pi20 ? n2358 : n342;
  assign n36913 = pi19 ? n36912 : ~n32;
  assign n36914 = pi18 ? n36911 : ~n36913;
  assign n36915 = pi17 ? n32 : n36914;
  assign n36916 = pi16 ? n32 : n36915;
  assign n36917 = pi19 ? n507 : ~n11879;
  assign n36918 = pi19 ? n8818 : n32;
  assign n36919 = pi18 ? n36917 : n36918;
  assign n36920 = pi17 ? n32 : n36919;
  assign n36921 = pi16 ? n32 : n36920;
  assign n36922 = pi15 ? n36916 : n36921;
  assign n36923 = pi18 ? n16449 : n34401;
  assign n36924 = pi17 ? n32 : n36923;
  assign n36925 = pi16 ? n32 : n36924;
  assign n36926 = pi14 ? n36922 : n36925;
  assign n36927 = pi13 ? n36910 : n36926;
  assign n36928 = pi12 ? n36898 : n36927;
  assign n36929 = pi15 ? n13904 : n23443;
  assign n36930 = pi15 ? n21853 : n14156;
  assign n36931 = pi14 ? n36929 : n36930;
  assign n36932 = pi18 ? n32 : n21270;
  assign n36933 = pi18 ? n1758 : ~n248;
  assign n36934 = pi17 ? n36932 : ~n36933;
  assign n36935 = pi16 ? n32 : n36934;
  assign n36936 = pi15 ? n36748 : n36935;
  assign n36937 = pi14 ? n36745 : n36936;
  assign n36938 = pi13 ? n36931 : n36937;
  assign n36939 = pi18 ? n18102 : ~n36759;
  assign n36940 = pi18 ? n24932 : ~n4343;
  assign n36941 = pi17 ? n36939 : ~n36940;
  assign n36942 = pi16 ? n32 : n36941;
  assign n36943 = pi19 ? n18678 : n32;
  assign n36944 = pi18 ? n18102 : ~n36943;
  assign n36945 = pi18 ? n14982 : n23543;
  assign n36946 = pi17 ? n36944 : ~n36945;
  assign n36947 = pi16 ? n32 : n36946;
  assign n36948 = pi15 ? n36942 : n36947;
  assign n36949 = pi18 ? n23548 : n532;
  assign n36950 = pi17 ? n32 : ~n36949;
  assign n36951 = pi16 ? n32 : n36950;
  assign n36952 = pi15 ? n36951 : n535;
  assign n36953 = pi14 ? n36948 : n36952;
  assign n36954 = pi20 ? n321 : ~n7839;
  assign n36955 = pi19 ? n16002 : ~n36954;
  assign n36956 = pi18 ? n36955 : n5436;
  assign n36957 = pi17 ? n32 : ~n36956;
  assign n36958 = pi16 ? n534 : n36957;
  assign n36959 = pi19 ? n322 : ~n21349;
  assign n36960 = pi18 ? n36959 : n32;
  assign n36961 = pi17 ? n36960 : n30107;
  assign n36962 = pi16 ? n534 : n36961;
  assign n36963 = pi15 ? n36958 : n36962;
  assign n36964 = pi19 ? n5694 : n266;
  assign n36965 = pi18 ? n36964 : n32;
  assign n36966 = pi17 ? n36965 : n2119;
  assign n36967 = pi16 ? n1135 : ~n36966;
  assign n36968 = pi15 ? n36967 : n36601;
  assign n36969 = pi14 ? n36963 : n36968;
  assign n36970 = pi13 ? n36953 : n36969;
  assign n36971 = pi12 ? n36938 : n36970;
  assign n36972 = pi11 ? n36928 : n36971;
  assign n36973 = pi10 ? n36888 : n36972;
  assign n36974 = pi09 ? n32 : n36973;
  assign n36975 = pi13 ? n26123 : n16973;
  assign n36976 = pi14 ? n25961 : n25640;
  assign n36977 = pi13 ? n36976 : n36857;
  assign n36978 = pi12 ? n36975 : n36977;
  assign n36979 = pi15 ? n24367 : n36862;
  assign n36980 = pi14 ? n36807 : n36979;
  assign n36981 = pi18 ? n5657 : n32;
  assign n36982 = pi17 ? n32 : n36981;
  assign n36983 = pi16 ? n32 : n36982;
  assign n36984 = pi15 ? n32 : n36983;
  assign n36985 = pi14 ? n36865 : n36984;
  assign n36986 = pi13 ? n36980 : n36985;
  assign n36987 = pi18 ? n36879 : ~n697;
  assign n36988 = pi17 ? n32 : n36987;
  assign n36989 = pi16 ? n32 : n36988;
  assign n36990 = pi15 ? n36878 : n36989;
  assign n36991 = pi14 ? n36689 : n36990;
  assign n36992 = pi13 ? n36873 : n36991;
  assign n36993 = pi12 ? n36986 : n36992;
  assign n36994 = pi11 ? n36978 : n36993;
  assign n36995 = pi14 ? n36896 : n25657;
  assign n36996 = pi13 ? n36895 : n36995;
  assign n36997 = pi14 ? n24743 : n36909;
  assign n36998 = pi18 ? n16449 : n34613;
  assign n36999 = pi17 ? n32 : n36998;
  assign n37000 = pi16 ? n32 : n36999;
  assign n37001 = pi14 ? n36922 : n37000;
  assign n37002 = pi13 ? n36997 : n37001;
  assign n37003 = pi12 ? n36996 : n37002;
  assign n37004 = pi20 ? n246 : ~n7939;
  assign n37005 = pi19 ? n32 : n37004;
  assign n37006 = pi18 ? n37005 : ~n36943;
  assign n37007 = pi17 ? n37006 : ~n36945;
  assign n37008 = pi16 ? n32 : n37007;
  assign n37009 = pi15 ? n36942 : n37008;
  assign n37010 = pi15 ? n36951 : n811;
  assign n37011 = pi14 ? n37009 : n37010;
  assign n37012 = pi16 ? n810 : n36957;
  assign n37013 = pi19 ? n322 : ~n24218;
  assign n37014 = pi18 ? n37013 : n32;
  assign n37015 = pi17 ? n37014 : n30107;
  assign n37016 = pi16 ? n810 : n37015;
  assign n37017 = pi15 ? n37012 : n37016;
  assign n37018 = pi19 ? n5694 : n17769;
  assign n37019 = pi18 ? n37018 : n32;
  assign n37020 = pi17 ? n37019 : n2119;
  assign n37021 = pi16 ? n1233 : ~n37020;
  assign n37022 = pi15 ? n37021 : n36601;
  assign n37023 = pi14 ? n37017 : n37022;
  assign n37024 = pi13 ? n37011 : n37023;
  assign n37025 = pi12 ? n36938 : n37024;
  assign n37026 = pi11 ? n37003 : n37025;
  assign n37027 = pi10 ? n36994 : n37026;
  assign n37028 = pi09 ? n32 : n37027;
  assign n37029 = pi08 ? n36974 : n37028;
  assign n37030 = pi07 ? n36847 : n37029;
  assign n37031 = pi13 ? n26165 : n16973;
  assign n37032 = pi14 ? n16973 : n16837;
  assign n37033 = pi15 ? n16973 : n16452;
  assign n37034 = pi14 ? n25037 : n37033;
  assign n37035 = pi13 ? n37032 : n37034;
  assign n37036 = pi12 ? n37031 : n37035;
  assign n37037 = pi15 ? n16452 : n16101;
  assign n37038 = pi19 ? n4126 : n3692;
  assign n37039 = pi18 ? n32 : n37038;
  assign n37040 = pi17 ? n32 : n37039;
  assign n37041 = pi16 ? n32 : n37040;
  assign n37042 = pi15 ? n16101 : n37041;
  assign n37043 = pi14 ? n37037 : n37042;
  assign n37044 = pi15 ? n36296 : n24247;
  assign n37045 = pi14 ? n37044 : n32;
  assign n37046 = pi13 ? n37043 : n37045;
  assign n37047 = pi14 ? n16319 : n32;
  assign n37048 = pi18 ? n16847 : n5725;
  assign n37049 = pi17 ? n32 : n37048;
  assign n37050 = pi16 ? n32 : n37049;
  assign n37051 = pi15 ? n16105 : n37050;
  assign n37052 = pi19 ? n30044 : ~n5855;
  assign n37053 = pi19 ? n1757 : n349;
  assign n37054 = pi18 ? n37052 : ~n37053;
  assign n37055 = pi17 ? n30283 : n37054;
  assign n37056 = pi16 ? n32 : n37055;
  assign n37057 = pi20 ? n1331 : ~n246;
  assign n37058 = pi19 ? n32 : n37057;
  assign n37059 = pi19 ? n349 : ~n288;
  assign n37060 = pi18 ? n37058 : n37059;
  assign n37061 = pi17 ? n32 : n37060;
  assign n37062 = pi16 ? n32 : n37061;
  assign n37063 = pi15 ? n37056 : n37062;
  assign n37064 = pi14 ? n37051 : n37063;
  assign n37065 = pi13 ? n37047 : n37064;
  assign n37066 = pi12 ? n37046 : n37065;
  assign n37067 = pi11 ? n37036 : n37066;
  assign n37068 = pi19 ? n5004 : ~n236;
  assign n37069 = pi18 ? n37058 : n37068;
  assign n37070 = pi17 ? n32 : n37069;
  assign n37071 = pi16 ? n32 : n37070;
  assign n37072 = pi15 ? n37071 : n35897;
  assign n37073 = pi19 ? n20006 : ~n236;
  assign n37074 = pi18 ? n32 : n37073;
  assign n37075 = pi17 ? n32 : n37074;
  assign n37076 = pi16 ? n32 : n37075;
  assign n37077 = pi15 ? n37076 : n24443;
  assign n37078 = pi14 ? n37072 : n37077;
  assign n37079 = pi19 ? n311 : ~n813;
  assign n37080 = pi18 ? n32 : n37079;
  assign n37081 = pi17 ? n32 : n37080;
  assign n37082 = pi16 ? n32 : n37081;
  assign n37083 = pi15 ? n24443 : n37082;
  assign n37084 = pi15 ? n24304 : n25598;
  assign n37085 = pi14 ? n37083 : n37084;
  assign n37086 = pi13 ? n37078 : n37085;
  assign n37087 = pi19 ? n4491 : ~n32;
  assign n37088 = pi18 ? n17118 : ~n37087;
  assign n37089 = pi17 ? n32 : n37088;
  assign n37090 = pi16 ? n32 : n37089;
  assign n37091 = pi15 ? n35030 : n37090;
  assign n37092 = pi14 ? n26656 : n37091;
  assign n37093 = pi19 ? n20006 : ~n32;
  assign n37094 = pi18 ? n7647 : ~n37093;
  assign n37095 = pi17 ? n32 : n37094;
  assign n37096 = pi16 ? n32 : n37095;
  assign n37097 = pi18 ? n702 : ~n702;
  assign n37098 = pi17 ? n32 : n37097;
  assign n37099 = pi16 ? n32 : n37098;
  assign n37100 = pi15 ? n37096 : n37099;
  assign n37101 = pi18 ? n9346 : ~n32928;
  assign n37102 = pi17 ? n32 : n37101;
  assign n37103 = pi16 ? n32 : n37102;
  assign n37104 = pi18 ? n7038 : n6384;
  assign n37105 = pi17 ? n32 : n37104;
  assign n37106 = pi16 ? n32 : n37105;
  assign n37107 = pi15 ? n37103 : n37106;
  assign n37108 = pi14 ? n37100 : n37107;
  assign n37109 = pi13 ? n37092 : n37108;
  assign n37110 = pi12 ? n37086 : n37109;
  assign n37111 = pi15 ? n14138 : n33970;
  assign n37112 = pi18 ? n29802 : n25116;
  assign n37113 = pi17 ? n32 : n37112;
  assign n37114 = pi16 ? n32 : n37113;
  assign n37115 = pi18 ? n29802 : n20020;
  assign n37116 = pi17 ? n32 : n37115;
  assign n37117 = pi16 ? n32 : n37116;
  assign n37118 = pi15 ? n37114 : n37117;
  assign n37119 = pi14 ? n37111 : n37118;
  assign n37120 = pi19 ? n32 : ~n1464;
  assign n37121 = pi18 ? n32 : n37120;
  assign n37122 = pi19 ? n5694 : n4342;
  assign n37123 = pi18 ? n37122 : n33312;
  assign n37124 = pi17 ? n37121 : ~n37123;
  assign n37125 = pi16 ? n32 : n37124;
  assign n37126 = pi18 ? n20164 : ~n5372;
  assign n37127 = pi17 ? n20165 : n37126;
  assign n37128 = pi16 ? n32 : n37127;
  assign n37129 = pi15 ? n37125 : n37128;
  assign n37130 = pi18 ? n32909 : ~n532;
  assign n37131 = pi17 ? n32 : n37130;
  assign n37132 = pi16 ? n32 : n37131;
  assign n37133 = pi18 ? n31290 : n237;
  assign n37134 = pi17 ? n32 : ~n37133;
  assign n37135 = pi16 ? n32 : n37134;
  assign n37136 = pi15 ? n37132 : n37135;
  assign n37137 = pi14 ? n37129 : n37136;
  assign n37138 = pi13 ? n37119 : n37137;
  assign n37139 = pi17 ? n15845 : n28415;
  assign n37140 = pi16 ? n32 : n37139;
  assign n37141 = pi18 ? n21274 : ~n5164;
  assign n37142 = pi17 ? n36742 : ~n37141;
  assign n37143 = pi16 ? n32 : n37142;
  assign n37144 = pi15 ? n37140 : n37143;
  assign n37145 = pi18 ? n9012 : ~n797;
  assign n37146 = pi17 ? n32 : n37145;
  assign n37147 = pi16 ? n32 : n37146;
  assign n37148 = pi16 ? n955 : n13947;
  assign n37149 = pi15 ? n37147 : n37148;
  assign n37150 = pi14 ? n37144 : n37149;
  assign n37151 = pi18 ? n20164 : ~n797;
  assign n37152 = pi17 ? n32 : n37151;
  assign n37153 = pi16 ? n955 : n37152;
  assign n37154 = pi18 ? n32053 : n4343;
  assign n37155 = pi17 ? n19071 : n37154;
  assign n37156 = pi16 ? n882 : n37155;
  assign n37157 = pi15 ? n37153 : n37156;
  assign n37158 = pi17 ? n20065 : n2519;
  assign n37159 = pi16 ? n1135 : ~n37158;
  assign n37160 = pi16 ? n1972 : ~n2120;
  assign n37161 = pi15 ? n37159 : n37160;
  assign n37162 = pi14 ? n37157 : n37161;
  assign n37163 = pi13 ? n37150 : n37162;
  assign n37164 = pi12 ? n37138 : n37163;
  assign n37165 = pi11 ? n37110 : n37164;
  assign n37166 = pi10 ? n37067 : n37165;
  assign n37167 = pi09 ? n32 : n37166;
  assign n37168 = pi14 ? n26163 : n17039;
  assign n37169 = pi13 ? n37168 : n17039;
  assign n37170 = pi14 ? n32 : n27450;
  assign n37171 = pi15 ? n25384 : n16899;
  assign n37172 = pi14 ? n37171 : n37033;
  assign n37173 = pi13 ? n37170 : n37172;
  assign n37174 = pi12 ? n37169 : n37173;
  assign n37175 = pi19 ? n1464 : ~n7230;
  assign n37176 = pi18 ? n32 : n37175;
  assign n37177 = pi17 ? n32 : n37176;
  assign n37178 = pi16 ? n32 : n37177;
  assign n37179 = pi19 ? n32 : ~n7230;
  assign n37180 = pi18 ? n32 : n37179;
  assign n37181 = pi17 ? n32 : n37180;
  assign n37182 = pi16 ? n32 : n37181;
  assign n37183 = pi15 ? n37178 : n37182;
  assign n37184 = pi14 ? n37183 : n16840;
  assign n37185 = pi13 ? n37043 : n37184;
  assign n37186 = pi12 ? n37185 : n37065;
  assign n37187 = pi11 ? n37174 : n37186;
  assign n37188 = pi18 ? n32 : n28433;
  assign n37189 = pi17 ? n32 : n37188;
  assign n37190 = pi16 ? n32 : n37189;
  assign n37191 = pi15 ? n37076 : n37190;
  assign n37192 = pi14 ? n37072 : n37191;
  assign n37193 = pi15 ? n37190 : n37082;
  assign n37194 = pi19 ? n322 : ~n1812;
  assign n37195 = pi18 ? n32 : n37194;
  assign n37196 = pi17 ? n32 : n37195;
  assign n37197 = pi16 ? n32 : n37196;
  assign n37198 = pi15 ? n24304 : n37197;
  assign n37199 = pi14 ? n37193 : n37198;
  assign n37200 = pi13 ? n37192 : n37199;
  assign n37201 = pi12 ? n37200 : n37109;
  assign n37202 = pi19 ? n31941 : ~n32;
  assign n37203 = pi18 ? n32 : n37202;
  assign n37204 = pi17 ? n37203 : ~n37141;
  assign n37205 = pi16 ? n32 : n37204;
  assign n37206 = pi15 ? n37140 : n37205;
  assign n37207 = pi16 ? n12460 : n13947;
  assign n37208 = pi15 ? n37147 : n37207;
  assign n37209 = pi14 ? n37206 : n37208;
  assign n37210 = pi16 ? n12460 : n37152;
  assign n37211 = pi16 ? n11454 : n37155;
  assign n37212 = pi15 ? n37210 : n37211;
  assign n37213 = pi18 ? n32 : n5856;
  assign n37214 = pi17 ? n37213 : n2519;
  assign n37215 = pi16 ? n1594 : ~n37214;
  assign n37216 = pi16 ? n1594 : ~n2120;
  assign n37217 = pi15 ? n37215 : n37216;
  assign n37218 = pi14 ? n37212 : n37217;
  assign n37219 = pi13 ? n37209 : n37218;
  assign n37220 = pi12 ? n37138 : n37219;
  assign n37221 = pi11 ? n37201 : n37220;
  assign n37222 = pi10 ? n37187 : n37221;
  assign n37223 = pi09 ? n32 : n37222;
  assign n37224 = pi08 ? n37167 : n37223;
  assign n37225 = pi15 ? n17188 : n17036;
  assign n37226 = pi14 ? n37225 : n17043;
  assign n37227 = pi13 ? n37226 : n17039;
  assign n37228 = pi14 ? n32 : n24962;
  assign n37229 = pi15 ? n25384 : n16392;
  assign n37230 = pi14 ? n37229 : n16974;
  assign n37231 = pi13 ? n37228 : n37230;
  assign n37232 = pi12 ? n37227 : n37231;
  assign n37233 = pi20 ? n32 : ~n7939;
  assign n37234 = pi19 ? n37233 : ~n343;
  assign n37235 = pi18 ? n936 : n37234;
  assign n37236 = pi17 ? n32 : n37235;
  assign n37237 = pi16 ? n32 : n37236;
  assign n37238 = pi15 ? n16606 : n37237;
  assign n37239 = pi18 ? n936 : n24697;
  assign n37240 = pi17 ? n32 : n37239;
  assign n37241 = pi16 ? n32 : n37240;
  assign n37242 = pi15 ? n37237 : n37241;
  assign n37243 = pi14 ? n37238 : n37242;
  assign n37244 = pi14 ? n16105 : n32;
  assign n37245 = pi13 ? n37243 : n37244;
  assign n37246 = pi19 ? n531 : ~n20266;
  assign n37247 = pi18 ? n32 : n37246;
  assign n37248 = pi17 ? n32 : n37247;
  assign n37249 = pi16 ? n32 : n37248;
  assign n37250 = pi15 ? n32 : n37249;
  assign n37251 = pi19 ? n349 : ~n2317;
  assign n37252 = pi18 ? n4380 : n37251;
  assign n37253 = pi17 ? n32 : n37252;
  assign n37254 = pi16 ? n32 : n37253;
  assign n37255 = pi19 ? n22525 : n19317;
  assign n37256 = pi18 ? n32 : n37255;
  assign n37257 = pi17 ? n32 : n37256;
  assign n37258 = pi16 ? n32 : n37257;
  assign n37259 = pi15 ? n37254 : n37258;
  assign n37260 = pi14 ? n37250 : n37259;
  assign n37261 = pi13 ? n32 : n37260;
  assign n37262 = pi12 ? n37245 : n37261;
  assign n37263 = pi11 ? n37232 : n37262;
  assign n37264 = pi19 ? n20006 : ~n349;
  assign n37265 = pi18 ? n32 : n37264;
  assign n37266 = pi17 ? n32 : n37265;
  assign n37267 = pi16 ? n32 : n37266;
  assign n37268 = pi15 ? n37267 : n37190;
  assign n37269 = pi14 ? n30921 : n37268;
  assign n37270 = pi15 ? n37190 : n24304;
  assign n37271 = pi19 ? n1464 : ~n1812;
  assign n37272 = pi18 ? n32 : n37271;
  assign n37273 = pi17 ? n32 : n37272;
  assign n37274 = pi16 ? n32 : n37273;
  assign n37275 = pi15 ? n24304 : n37274;
  assign n37276 = pi14 ? n37270 : n37275;
  assign n37277 = pi13 ? n37269 : n37276;
  assign n37278 = pi19 ? n1818 : ~n1812;
  assign n37279 = pi18 ? n32 : n37278;
  assign n37280 = pi17 ? n32 : n37279;
  assign n37281 = pi16 ? n32 : n37280;
  assign n37282 = pi15 ? n37281 : n24256;
  assign n37283 = pi19 ? n1165 : ~n813;
  assign n37284 = pi18 ? n32 : n37283;
  assign n37285 = pi17 ? n32 : n37284;
  assign n37286 = pi16 ? n32 : n37285;
  assign n37287 = pi15 ? n37286 : n36697;
  assign n37288 = pi14 ? n37282 : n37287;
  assign n37289 = pi19 ? n4126 : n236;
  assign n37290 = pi18 ? n880 : ~n37289;
  assign n37291 = pi17 ? n32 : n37290;
  assign n37292 = pi16 ? n32 : n37291;
  assign n37293 = pi19 ? n32 : ~n6171;
  assign n37294 = pi18 ? n37293 : ~n1750;
  assign n37295 = pi17 ? n32 : n37294;
  assign n37296 = pi16 ? n32 : n37295;
  assign n37297 = pi15 ? n37292 : n37296;
  assign n37298 = pi19 ? n4342 : n617;
  assign n37299 = pi18 ? n880 : ~n37298;
  assign n37300 = pi17 ? n32 : n37299;
  assign n37301 = pi16 ? n32 : n37300;
  assign n37302 = pi15 ? n37301 : n37106;
  assign n37303 = pi14 ? n37297 : n37302;
  assign n37304 = pi13 ? n37288 : n37303;
  assign n37305 = pi12 ? n37277 : n37304;
  assign n37306 = pi18 ? n4380 : n6384;
  assign n37307 = pi17 ? n32 : n37306;
  assign n37308 = pi16 ? n32 : n37307;
  assign n37309 = pi19 ? n857 : ~n617;
  assign n37310 = pi18 ? n32 : n37309;
  assign n37311 = pi17 ? n32 : n37310;
  assign n37312 = pi16 ? n32 : n37311;
  assign n37313 = pi15 ? n37308 : n37312;
  assign n37314 = pi18 ? n29802 : n20912;
  assign n37315 = pi17 ? n32 : n37314;
  assign n37316 = pi16 ? n32 : n37315;
  assign n37317 = pi18 ? n29802 : n14955;
  assign n37318 = pi17 ? n32 : n37317;
  assign n37319 = pi16 ? n32 : n37318;
  assign n37320 = pi15 ? n37316 : n37319;
  assign n37321 = pi14 ? n37313 : n37320;
  assign n37322 = pi19 ? n32 : ~n1740;
  assign n37323 = pi18 ? n32 : n37322;
  assign n37324 = pi20 ? n266 : n1324;
  assign n37325 = pi20 ? n1385 : ~n206;
  assign n37326 = pi19 ? n37324 : ~n37325;
  assign n37327 = pi18 ? n37326 : ~n33312;
  assign n37328 = pi17 ? n37323 : n37327;
  assign n37329 = pi16 ? n32 : n37328;
  assign n37330 = pi18 ? n20164 : ~n350;
  assign n37331 = pi17 ? n20165 : n37330;
  assign n37332 = pi16 ? n32 : n37331;
  assign n37333 = pi15 ? n37329 : n37332;
  assign n37334 = pi14 ? n37333 : n37136;
  assign n37335 = pi13 ? n37321 : n37334;
  assign n37336 = pi19 ? n2359 : n236;
  assign n37337 = pi18 ? n32 : n37336;
  assign n37338 = pi18 ? n21274 : ~n5009;
  assign n37339 = pi17 ? n37337 : ~n37338;
  assign n37340 = pi16 ? n32 : n37339;
  assign n37341 = pi15 ? n37140 : n37340;
  assign n37342 = pi16 ? n11684 : n14155;
  assign n37343 = pi15 ? n32 : n37342;
  assign n37344 = pi14 ? n37341 : n37343;
  assign n37345 = pi18 ? n20164 : n23548;
  assign n37346 = pi17 ? n32 : n37345;
  assign n37347 = pi16 ? n11684 : n37346;
  assign n37348 = pi19 ? n4721 : ~n4126;
  assign n37349 = pi18 ? n37348 : n4343;
  assign n37350 = pi17 ? n19071 : n37349;
  assign n37351 = pi16 ? n11684 : n37350;
  assign n37352 = pi15 ? n37347 : n37351;
  assign n37353 = pi18 ? n32 : n34142;
  assign n37354 = pi17 ? n37353 : n2519;
  assign n37355 = pi16 ? n1577 : ~n37354;
  assign n37356 = pi16 ? n1577 : ~n2120;
  assign n37357 = pi15 ? n37355 : n37356;
  assign n37358 = pi14 ? n37352 : n37357;
  assign n37359 = pi13 ? n37344 : n37358;
  assign n37360 = pi12 ? n37335 : n37359;
  assign n37361 = pi11 ? n37305 : n37360;
  assign n37362 = pi10 ? n37263 : n37361;
  assign n37363 = pi09 ? n32 : n37362;
  assign n37364 = pi14 ? n37225 : n17036;
  assign n37365 = pi15 ? n17039 : n17188;
  assign n37366 = pi14 ? n37365 : n17070;
  assign n37367 = pi13 ? n37364 : n37366;
  assign n37368 = pi14 ? n25291 : n32;
  assign n37369 = pi13 ? n37168 : n37368;
  assign n37370 = pi12 ? n37367 : n37369;
  assign n37371 = pi19 ? n531 : ~n288;
  assign n37372 = pi18 ? n32 : n37371;
  assign n37373 = pi17 ? n32 : n37372;
  assign n37374 = pi16 ? n32 : n37373;
  assign n37375 = pi15 ? n32 : n37374;
  assign n37376 = pi19 ? n349 : ~n589;
  assign n37377 = pi18 ? n4380 : n37376;
  assign n37378 = pi17 ? n32 : n37377;
  assign n37379 = pi16 ? n32 : n37378;
  assign n37380 = pi19 ? n22525 : n3495;
  assign n37381 = pi18 ? n32 : n37380;
  assign n37382 = pi17 ? n32 : n37381;
  assign n37383 = pi16 ? n32 : n37382;
  assign n37384 = pi15 ? n37379 : n37383;
  assign n37385 = pi14 ? n37375 : n37384;
  assign n37386 = pi13 ? n32 : n37385;
  assign n37387 = pi12 ? n37245 : n37386;
  assign n37388 = pi11 ? n37370 : n37387;
  assign n37389 = pi19 ? n20006 : ~n589;
  assign n37390 = pi18 ? n32 : n37389;
  assign n37391 = pi17 ? n32 : n37390;
  assign n37392 = pi16 ? n32 : n37391;
  assign n37393 = pi19 ? n208 : ~n2848;
  assign n37394 = pi18 ? n32 : n37393;
  assign n37395 = pi17 ? n32 : n37394;
  assign n37396 = pi16 ? n32 : n37395;
  assign n37397 = pi15 ? n37392 : n37396;
  assign n37398 = pi14 ? n30921 : n37397;
  assign n37399 = pi15 ? n37396 : n36296;
  assign n37400 = pi15 ? n36296 : n37274;
  assign n37401 = pi14 ? n37399 : n37400;
  assign n37402 = pi13 ? n37398 : n37401;
  assign n37403 = pi15 ? n37281 : n25331;
  assign n37404 = pi19 ? n1165 : ~n1812;
  assign n37405 = pi18 ? n32 : n37404;
  assign n37406 = pi17 ? n32 : n37405;
  assign n37407 = pi16 ? n32 : n37406;
  assign n37408 = pi18 ? n32 : ~n2730;
  assign n37409 = pi17 ? n32 : n37408;
  assign n37410 = pi16 ? n32 : n37409;
  assign n37411 = pi15 ? n37407 : n37410;
  assign n37412 = pi14 ? n37403 : n37411;
  assign n37413 = pi19 ? n4126 : n1941;
  assign n37414 = pi18 ? n880 : ~n37413;
  assign n37415 = pi17 ? n32 : n37414;
  assign n37416 = pi16 ? n32 : n37415;
  assign n37417 = pi15 ? n37416 : n37296;
  assign n37418 = pi19 ? n4342 : n236;
  assign n37419 = pi18 ? n880 : ~n37418;
  assign n37420 = pi17 ? n32 : n37419;
  assign n37421 = pi16 ? n32 : n37420;
  assign n37422 = pi15 ? n37421 : n37106;
  assign n37423 = pi14 ? n37417 : n37422;
  assign n37424 = pi13 ? n37412 : n37423;
  assign n37425 = pi12 ? n37402 : n37424;
  assign n37426 = pi19 ? n1785 : ~n617;
  assign n37427 = pi18 ? n32 : n37426;
  assign n37428 = pi17 ? n32 : n37427;
  assign n37429 = pi16 ? n32 : n37428;
  assign n37430 = pi15 ? n37308 : n37429;
  assign n37431 = pi18 ? n29802 : n14964;
  assign n37432 = pi17 ? n32 : n37431;
  assign n37433 = pi16 ? n32 : n37432;
  assign n37434 = pi15 ? n37316 : n37433;
  assign n37435 = pi14 ? n37430 : n37434;
  assign n37436 = pi13 ? n37435 : n37334;
  assign n37437 = pi16 ? n11886 : n14155;
  assign n37438 = pi15 ? n32 : n37437;
  assign n37439 = pi14 ? n37341 : n37438;
  assign n37440 = pi16 ? n11886 : n37346;
  assign n37441 = pi16 ? n12116 : n37350;
  assign n37442 = pi15 ? n37440 : n37441;
  assign n37443 = pi18 ? n32 : n34040;
  assign n37444 = pi17 ? n37443 : n2519;
  assign n37445 = pi16 ? n2137 : ~n37444;
  assign n37446 = pi16 ? n2137 : ~n2120;
  assign n37447 = pi15 ? n37445 : n37446;
  assign n37448 = pi14 ? n37442 : n37447;
  assign n37449 = pi13 ? n37439 : n37448;
  assign n37450 = pi12 ? n37436 : n37449;
  assign n37451 = pi11 ? n37425 : n37450;
  assign n37452 = pi10 ? n37388 : n37451;
  assign n37453 = pi09 ? n32 : n37452;
  assign n37454 = pi08 ? n37363 : n37453;
  assign n37455 = pi07 ? n37224 : n37454;
  assign n37456 = pi06 ? n37030 : n37455;
  assign n37457 = pi05 ? n36663 : n37456;
  assign n37458 = pi15 ? n17111 : n16984;
  assign n37459 = pi14 ? n37458 : n17188;
  assign n37460 = pi13 ? n37459 : n25290;
  assign n37461 = pi14 ? n26163 : n25378;
  assign n37462 = pi14 ? n16940 : n32;
  assign n37463 = pi13 ? n37461 : n37462;
  assign n37464 = pi12 ? n37460 : n37463;
  assign n37465 = pi19 ? n507 : n10879;
  assign n37466 = pi18 ? n32 : n37465;
  assign n37467 = pi17 ? n32 : n37466;
  assign n37468 = pi16 ? n32 : n37467;
  assign n37469 = pi15 ? n32 : n37468;
  assign n37470 = pi15 ? n16837 : n16452;
  assign n37471 = pi14 ? n37469 : n37470;
  assign n37472 = pi19 ? n23193 : ~n4406;
  assign n37473 = pi18 ? n32 : n37472;
  assign n37474 = pi17 ? n32 : n37473;
  assign n37475 = pi16 ? n32 : n37474;
  assign n37476 = pi15 ? n16452 : n37475;
  assign n37477 = pi14 ? n16452 : n37476;
  assign n37478 = pi13 ? n37471 : n37477;
  assign n37479 = pi14 ? n24633 : n32;
  assign n37480 = pi19 ? n6355 : ~n349;
  assign n37481 = pi18 ? n32 : n37480;
  assign n37482 = pi17 ? n32 : n37481;
  assign n37483 = pi16 ? n32 : n37482;
  assign n37484 = pi19 ? n343 : ~n589;
  assign n37485 = pi18 ? n32 : n37484;
  assign n37486 = pi17 ? n32 : n37485;
  assign n37487 = pi16 ? n32 : n37486;
  assign n37488 = pi15 ? n37483 : n37487;
  assign n37489 = pi19 ? n22864 : ~n349;
  assign n37490 = pi18 ? n32 : n37489;
  assign n37491 = pi17 ? n32 : n37490;
  assign n37492 = pi16 ? n32 : n37491;
  assign n37493 = pi15 ? n37492 : n36296;
  assign n37494 = pi14 ? n37488 : n37493;
  assign n37495 = pi13 ? n37479 : n37494;
  assign n37496 = pi12 ? n37478 : n37495;
  assign n37497 = pi11 ? n37464 : n37496;
  assign n37498 = pi19 ? n322 : ~n589;
  assign n37499 = pi18 ? n32 : n37498;
  assign n37500 = pi17 ? n32 : n37499;
  assign n37501 = pi16 ? n32 : n37500;
  assign n37502 = pi15 ? n23933 : n37501;
  assign n37503 = pi14 ? n37502 : n14917;
  assign n37504 = pi15 ? n15244 : n24582;
  assign n37505 = pi14 ? n37504 : n15244;
  assign n37506 = pi13 ? n37503 : n37505;
  assign n37507 = pi15 ? n23484 : n24742;
  assign n37508 = pi15 ? n36301 : n35452;
  assign n37509 = pi14 ? n37507 : n37508;
  assign n37510 = pi19 ? n1757 : n236;
  assign n37511 = pi18 ? n863 : ~n37510;
  assign n37512 = pi17 ? n32 : n37511;
  assign n37513 = pi16 ? n32 : n37512;
  assign n37514 = pi15 ? n35393 : n37513;
  assign n37515 = pi15 ? n35452 : n24659;
  assign n37516 = pi14 ? n37514 : n37515;
  assign n37517 = pi13 ? n37509 : n37516;
  assign n37518 = pi12 ? n37506 : n37517;
  assign n37519 = pi18 ? n8192 : n23440;
  assign n37520 = pi17 ? n32 : n37519;
  assign n37521 = pi16 ? n32 : n37520;
  assign n37522 = pi19 ? n32 : n18390;
  assign n37523 = pi18 ? n37522 : ~n23200;
  assign n37524 = pi17 ? n32 : n37523;
  assign n37525 = pi16 ? n32 : n37524;
  assign n37526 = pi15 ? n37521 : n37525;
  assign n37527 = pi14 ? n32 : n37526;
  assign n37528 = pi17 ? n32 : n14153;
  assign n37529 = pi16 ? n32 : n37528;
  assign n37530 = pi15 ? n37529 : n33939;
  assign n37531 = pi14 ? n37530 : n20883;
  assign n37532 = pi13 ? n37527 : n37531;
  assign n37533 = pi19 ? n18502 : ~n531;
  assign n37534 = pi18 ? n37533 : n32;
  assign n37535 = pi17 ? n2954 : n37534;
  assign n37536 = pi16 ? n32 : n37535;
  assign n37537 = pi19 ? n18502 : ~n343;
  assign n37538 = pi18 ? n37537 : n32;
  assign n37539 = pi17 ? n2954 : n37538;
  assign n37540 = pi16 ? n32 : n37539;
  assign n37541 = pi15 ? n37536 : n37540;
  assign n37542 = pi20 ? n207 : n266;
  assign n37543 = pi19 ? n37542 : n32;
  assign n37544 = pi18 ? n940 : n37543;
  assign n37545 = pi17 ? n32 : n37544;
  assign n37546 = pi16 ? n2320 : n37545;
  assign n37547 = pi15 ? n32 : n37546;
  assign n37548 = pi14 ? n37541 : n37547;
  assign n37549 = pi20 ? n274 : n321;
  assign n37550 = pi19 ? n37549 : ~n32;
  assign n37551 = pi18 ? n268 : ~n37550;
  assign n37552 = pi17 ? n32 : n37551;
  assign n37553 = pi16 ? n2320 : n37552;
  assign n37554 = pi16 ? n179 : n30108;
  assign n37555 = pi15 ? n37553 : n37554;
  assign n37556 = pi16 ? n2320 : ~n3769;
  assign n37557 = pi14 ? n37555 : n37556;
  assign n37558 = pi13 ? n37548 : n37557;
  assign n37559 = pi12 ? n37532 : n37558;
  assign n37560 = pi11 ? n37518 : n37559;
  assign n37561 = pi10 ? n37497 : n37560;
  assign n37562 = pi09 ? n32 : n37561;
  assign n37563 = pi15 ? n17188 : n16984;
  assign n37564 = pi14 ? n16984 : n37563;
  assign n37565 = pi15 ? n17111 : n32;
  assign n37566 = pi14 ? n16985 : n37565;
  assign n37567 = pi13 ? n37564 : n37566;
  assign n37568 = pi15 ? n32 : n17036;
  assign n37569 = pi15 ? n17039 : n16832;
  assign n37570 = pi14 ? n37568 : n37569;
  assign n37571 = pi14 ? n16832 : n17189;
  assign n37572 = pi13 ? n37570 : n37571;
  assign n37573 = pi12 ? n37567 : n37572;
  assign n37574 = pi15 ? n16520 : n32;
  assign n37575 = pi14 ? n37574 : n32;
  assign n37576 = pi13 ? n37575 : n37494;
  assign n37577 = pi12 ? n37478 : n37576;
  assign n37578 = pi11 ? n37573 : n37577;
  assign n37579 = pi14 ? n37502 : n37501;
  assign n37580 = pi15 ? n36100 : n24582;
  assign n37581 = pi14 ? n37580 : n15244;
  assign n37582 = pi13 ? n37579 : n37581;
  assign n37583 = pi19 ? n750 : ~n813;
  assign n37584 = pi18 ? n32 : n37583;
  assign n37585 = pi17 ? n32 : n37584;
  assign n37586 = pi16 ? n32 : n37585;
  assign n37587 = pi15 ? n37586 : n35452;
  assign n37588 = pi14 ? n37507 : n37587;
  assign n37589 = pi19 ? n349 : ~n1941;
  assign n37590 = pi18 ? n32 : n37589;
  assign n37591 = pi17 ? n32 : n37590;
  assign n37592 = pi16 ? n32 : n37591;
  assign n37593 = pi19 ? n1757 : n1941;
  assign n37594 = pi18 ? n863 : ~n37593;
  assign n37595 = pi17 ? n32 : n37594;
  assign n37596 = pi16 ? n32 : n37595;
  assign n37597 = pi15 ? n37592 : n37596;
  assign n37598 = pi14 ? n37597 : n37515;
  assign n37599 = pi13 ? n37588 : n37598;
  assign n37600 = pi12 ? n37582 : n37599;
  assign n37601 = pi16 ? n3625 : n37545;
  assign n37602 = pi15 ? n32 : n37601;
  assign n37603 = pi14 ? n37541 : n37602;
  assign n37604 = pi16 ? n3625 : n37552;
  assign n37605 = pi15 ? n37604 : n30109;
  assign n37606 = pi16 ? n3625 : ~n3769;
  assign n37607 = pi16 ? n2654 : ~n3769;
  assign n37608 = pi15 ? n37606 : n37607;
  assign n37609 = pi14 ? n37605 : n37608;
  assign n37610 = pi13 ? n37603 : n37609;
  assign n37611 = pi12 ? n37532 : n37610;
  assign n37612 = pi11 ? n37600 : n37611;
  assign n37613 = pi10 ? n37578 : n37612;
  assign n37614 = pi09 ? n32 : n37613;
  assign n37615 = pi08 ? n37562 : n37614;
  assign n37616 = pi15 ? n25556 : n26115;
  assign n37617 = pi14 ? n37616 : n37458;
  assign n37618 = pi14 ? n37458 : n17412;
  assign n37619 = pi13 ? n37617 : n37618;
  assign n37620 = pi15 ? n16832 : n16973;
  assign n37621 = pi14 ? n37620 : n32;
  assign n37622 = pi13 ? n25288 : n37621;
  assign n37623 = pi12 ? n37619 : n37622;
  assign n37624 = pi15 ? n36851 : n25576;
  assign n37625 = pi14 ? n37624 : n27678;
  assign n37626 = pi19 ? n32 : ~n8946;
  assign n37627 = pi18 ? n32 : n37626;
  assign n37628 = pi17 ? n32 : n37627;
  assign n37629 = pi16 ? n32 : n37628;
  assign n37630 = pi15 ? n37629 : n16452;
  assign n37631 = pi19 ? n32 : ~n11108;
  assign n37632 = pi18 ? n32 : n37631;
  assign n37633 = pi17 ? n32 : n37632;
  assign n37634 = pi16 ? n32 : n37633;
  assign n37635 = pi15 ? n16452 : n37634;
  assign n37636 = pi14 ? n37630 : n37635;
  assign n37637 = pi13 ? n37625 : n37636;
  assign n37638 = pi19 ? n208 : ~n2303;
  assign n37639 = pi18 ? n32 : n37638;
  assign n37640 = pi17 ? n32 : n37639;
  assign n37641 = pi16 ? n32 : n37640;
  assign n37642 = pi15 ? n32 : n37641;
  assign n37643 = pi17 ? n32 : n30633;
  assign n37644 = pi16 ? n32 : n37643;
  assign n37645 = pi14 ? n37642 : n37644;
  assign n37646 = pi13 ? n37479 : n37645;
  assign n37647 = pi12 ? n37637 : n37646;
  assign n37648 = pi11 ? n37623 : n37647;
  assign n37649 = pi15 ? n24813 : n37501;
  assign n37650 = pi14 ? n37649 : n37501;
  assign n37651 = pi19 ? n507 : n7693;
  assign n37652 = pi18 ? n32 : n37651;
  assign n37653 = pi17 ? n32 : n37652;
  assign n37654 = pi16 ? n32 : n37653;
  assign n37655 = pi15 ? n15244 : n37654;
  assign n37656 = pi14 ? n37504 : n37655;
  assign n37657 = pi13 ? n37650 : n37656;
  assign n37658 = pi19 ? n4721 : n440;
  assign n37659 = pi18 ? n32 : n37658;
  assign n37660 = pi17 ? n32 : n37659;
  assign n37661 = pi16 ? n32 : n37660;
  assign n37662 = pi15 ? n25598 : n37661;
  assign n37663 = pi14 ? n37507 : n37662;
  assign n37664 = pi19 ? n20555 : ~n236;
  assign n37665 = pi18 ? n32 : n37664;
  assign n37666 = pi17 ? n32 : n37665;
  assign n37667 = pi16 ? n32 : n37666;
  assign n37668 = pi15 ? n37667 : n35393;
  assign n37669 = pi14 ? n37668 : n37515;
  assign n37670 = pi13 ? n37663 : n37669;
  assign n37671 = pi12 ? n37657 : n37670;
  assign n37672 = pi18 ? n8192 : n20020;
  assign n37673 = pi17 ? n32 : n37672;
  assign n37674 = pi16 ? n32 : n37673;
  assign n37675 = pi19 ? n22185 : ~n32;
  assign n37676 = pi18 ? n37522 : ~n37675;
  assign n37677 = pi17 ? n32 : n37676;
  assign n37678 = pi16 ? n32 : n37677;
  assign n37679 = pi15 ? n37674 : n37678;
  assign n37680 = pi14 ? n21929 : n37679;
  assign n37681 = pi20 ? n342 : ~n1324;
  assign n37682 = pi19 ? n37681 : n32;
  assign n37683 = pi18 ? n14153 : n37682;
  assign n37684 = pi17 ? n32 : n37683;
  assign n37685 = pi16 ? n32 : n37684;
  assign n37686 = pi19 ? n35912 : n32;
  assign n37687 = pi18 ? n32 : n37686;
  assign n37688 = pi17 ? n32 : n37687;
  assign n37689 = pi16 ? n32 : n37688;
  assign n37690 = pi15 ? n37685 : n37689;
  assign n37691 = pi14 ? n37690 : n20883;
  assign n37692 = pi13 ? n37680 : n37691;
  assign n37693 = pi18 ? n14873 : n32;
  assign n37694 = pi17 ? n32 : n37693;
  assign n37695 = pi16 ? n32 : n37694;
  assign n37696 = pi19 ? n15533 : n32;
  assign n37697 = pi18 ? n940 : n37696;
  assign n37698 = pi17 ? n1028 : ~n37697;
  assign n37699 = pi16 ? n2293 : ~n37698;
  assign n37700 = pi15 ? n20660 : n37699;
  assign n37701 = pi14 ? n37695 : n37700;
  assign n37702 = pi18 ? n268 : ~n28193;
  assign n37703 = pi17 ? n1028 : ~n37702;
  assign n37704 = pi16 ? n2293 : ~n37703;
  assign n37705 = pi16 ? n21542 : n30108;
  assign n37706 = pi15 ? n37704 : n37705;
  assign n37707 = pi16 ? n2293 : ~n3769;
  assign n37708 = pi14 ? n37706 : n37707;
  assign n37709 = pi13 ? n37701 : n37708;
  assign n37710 = pi12 ? n37692 : n37709;
  assign n37711 = pi11 ? n37671 : n37710;
  assign n37712 = pi10 ? n37648 : n37711;
  assign n37713 = pi09 ? n32 : n37712;
  assign n37714 = pi14 ? n25867 : n17111;
  assign n37715 = pi15 ? n32 : n26115;
  assign n37716 = pi14 ? n37715 : n25625;
  assign n37717 = pi13 ? n37714 : n37716;
  assign n37718 = pi14 ? n16984 : n16985;
  assign n37719 = pi15 ? n25763 : n17066;
  assign n37720 = pi14 ? n37719 : n17412;
  assign n37721 = pi13 ? n37718 : n37720;
  assign n37722 = pi12 ? n37717 : n37721;
  assign n37723 = pi15 ? n32 : n25576;
  assign n37724 = pi14 ? n37723 : n27678;
  assign n37725 = pi13 ? n37724 : n37636;
  assign n37726 = pi15 ? n32 : n14207;
  assign n37727 = pi14 ? n37726 : n37644;
  assign n37728 = pi13 ? n37479 : n37727;
  assign n37729 = pi12 ? n37725 : n37728;
  assign n37730 = pi11 ? n37722 : n37729;
  assign n37731 = pi19 ? n32 : ~n8286;
  assign n37732 = pi18 ? n32 : n37731;
  assign n37733 = pi17 ? n32 : n37732;
  assign n37734 = pi16 ? n32 : n37733;
  assign n37735 = pi15 ? n37734 : n37501;
  assign n37736 = pi14 ? n37735 : n37501;
  assign n37737 = pi13 ? n37736 : n37504;
  assign n37738 = pi12 ? n37737 : n37670;
  assign n37739 = pi16 ? n2513 : ~n37698;
  assign n37740 = pi15 ? n20660 : n37739;
  assign n37741 = pi14 ? n37695 : n37740;
  assign n37742 = pi16 ? n2513 : ~n37703;
  assign n37743 = pi15 ? n37742 : n30109;
  assign n37744 = pi16 ? n2513 : ~n3769;
  assign n37745 = pi16 ? n4100 : ~n3769;
  assign n37746 = pi15 ? n37744 : n37745;
  assign n37747 = pi14 ? n37743 : n37746;
  assign n37748 = pi13 ? n37741 : n37747;
  assign n37749 = pi12 ? n37692 : n37748;
  assign n37750 = pi11 ? n37738 : n37749;
  assign n37751 = pi10 ? n37730 : n37750;
  assign n37752 = pi09 ? n32 : n37751;
  assign n37753 = pi08 ? n37713 : n37752;
  assign n37754 = pi07 ? n37615 : n37753;
  assign n37755 = pi14 ? n17435 : n25556;
  assign n37756 = pi13 ? n37755 : n25626;
  assign n37757 = pi14 ? n37719 : n17039;
  assign n37758 = pi13 ? n16984 : n37757;
  assign n37759 = pi12 ? n37756 : n37758;
  assign n37760 = pi15 ? n16392 : n14985;
  assign n37761 = pi20 ? n3695 : n32;
  assign n37762 = pi19 ? n32 : n37761;
  assign n37763 = pi18 ? n32 : n37762;
  assign n37764 = pi17 ? n32 : n37763;
  assign n37765 = pi16 ? n32 : n37764;
  assign n37766 = pi15 ? n15847 : n37765;
  assign n37767 = pi14 ? n37760 : n37766;
  assign n37768 = pi20 ? n246 : ~n141;
  assign n37769 = pi19 ? n32 : n37768;
  assign n37770 = pi18 ? n32 : n37769;
  assign n37771 = pi17 ? n32 : n37770;
  assign n37772 = pi16 ? n32 : n37771;
  assign n37773 = pi15 ? n23250 : n37772;
  assign n37774 = pi15 ? n16452 : n24874;
  assign n37775 = pi14 ? n37773 : n37774;
  assign n37776 = pi13 ? n37767 : n37775;
  assign n37777 = pi14 ? n32 : n24691;
  assign n37778 = pi17 ? n32 : n30817;
  assign n37779 = pi16 ? n32 : n37778;
  assign n37780 = pi15 ? n37779 : n26623;
  assign n37781 = pi15 ? n15230 : n16452;
  assign n37782 = pi14 ? n37780 : n37781;
  assign n37783 = pi13 ? n37777 : n37782;
  assign n37784 = pi12 ? n37776 : n37783;
  assign n37785 = pi11 ? n37759 : n37784;
  assign n37786 = pi15 ? n15230 : n15244;
  assign n37787 = pi15 ? n15244 : n24247;
  assign n37788 = pi14 ? n37786 : n37787;
  assign n37789 = pi15 ? n24247 : n24511;
  assign n37790 = pi14 ? n37789 : n26919;
  assign n37791 = pi13 ? n37788 : n37790;
  assign n37792 = pi19 ? n857 : ~n236;
  assign n37793 = pi18 ? n32 : n37792;
  assign n37794 = pi17 ? n32 : n37793;
  assign n37795 = pi16 ? n32 : n37794;
  assign n37796 = pi15 ? n25657 : n37795;
  assign n37797 = pi14 ? n16105 : n37796;
  assign n37798 = pi19 ? n267 : ~n236;
  assign n37799 = pi18 ? n32 : n37798;
  assign n37800 = pi17 ? n32 : n37799;
  assign n37801 = pi16 ? n32 : n37800;
  assign n37802 = pi15 ? n23484 : n37801;
  assign n37803 = pi15 ? n25598 : n24742;
  assign n37804 = pi14 ? n37802 : n37803;
  assign n37805 = pi13 ? n37797 : n37804;
  assign n37806 = pi12 ? n37791 : n37805;
  assign n37807 = pi18 ? n863 : ~n24548;
  assign n37808 = pi17 ? n32 : n37807;
  assign n37809 = pi16 ? n32 : n37808;
  assign n37810 = pi15 ? n21853 : n37809;
  assign n37811 = pi14 ? n32 : n37810;
  assign n37812 = pi18 ? n4127 : ~n508;
  assign n37813 = pi17 ? n32 : n37812;
  assign n37814 = pi16 ? n32 : n37813;
  assign n37815 = pi19 ? n32 : n37233;
  assign n37816 = pi18 ? n37815 : ~n508;
  assign n37817 = pi17 ? n32 : n37816;
  assign n37818 = pi16 ? n32 : n37817;
  assign n37819 = pi15 ? n37814 : n37818;
  assign n37820 = pi15 ? n13073 : n23551;
  assign n37821 = pi14 ? n37819 : n37820;
  assign n37822 = pi13 ? n37811 : n37821;
  assign n37823 = pi15 ? n21319 : n23551;
  assign n37824 = pi20 ? n749 : n1685;
  assign n37825 = pi19 ? n37824 : n32;
  assign n37826 = pi18 ? n863 : n37825;
  assign n37827 = pi17 ? n32 : n37826;
  assign n37828 = pi16 ? n32 : n37827;
  assign n37829 = pi18 ? n32 : n33538;
  assign n37830 = pi17 ? n2355 : ~n37829;
  assign n37831 = pi16 ? n2745 : ~n37830;
  assign n37832 = pi15 ? n37828 : n37831;
  assign n37833 = pi14 ? n37823 : n37832;
  assign n37834 = pi18 ? n19811 : n32;
  assign n37835 = pi20 ? n206 : n1817;
  assign n37836 = pi19 ? n37835 : n32;
  assign n37837 = pi18 ? n32 : n37836;
  assign n37838 = pi17 ? n37834 : n37837;
  assign n37839 = pi16 ? n15408 : n37838;
  assign n37840 = pi17 ? n1219 : ~n19529;
  assign n37841 = pi16 ? n2745 : ~n37840;
  assign n37842 = pi15 ? n37839 : n37841;
  assign n37843 = pi16 ? n2745 : ~n3769;
  assign n37844 = pi14 ? n37842 : n37843;
  assign n37845 = pi13 ? n37833 : n37844;
  assign n37846 = pi12 ? n37822 : n37845;
  assign n37847 = pi11 ? n37806 : n37846;
  assign n37848 = pi10 ? n37785 : n37847;
  assign n37849 = pi09 ? n32 : n37848;
  assign n37850 = pi15 ? n25749 : n17435;
  assign n37851 = pi14 ? n37850 : n25625;
  assign n37852 = pi14 ? n17578 : n25693;
  assign n37853 = pi13 ? n37851 : n37852;
  assign n37854 = pi14 ? n16984 : n27059;
  assign n37855 = pi15 ? n25814 : n17066;
  assign n37856 = pi14 ? n37855 : n17039;
  assign n37857 = pi13 ? n37854 : n37856;
  assign n37858 = pi12 ? n37853 : n37857;
  assign n37859 = pi15 ? n23250 : n16452;
  assign n37860 = pi14 ? n37859 : n37774;
  assign n37861 = pi13 ? n37767 : n37860;
  assign n37862 = pi15 ? n37779 : n23484;
  assign n37863 = pi14 ? n37862 : n37781;
  assign n37864 = pi13 ? n37777 : n37863;
  assign n37865 = pi12 ? n37861 : n37864;
  assign n37866 = pi11 ? n37858 : n37865;
  assign n37867 = pi15 ? n25598 : n25657;
  assign n37868 = pi14 ? n37802 : n37867;
  assign n37869 = pi13 ? n37797 : n37868;
  assign n37870 = pi12 ? n37791 : n37869;
  assign n37871 = pi20 ? n32 : ~n18834;
  assign n37872 = pi19 ? n32 : n37871;
  assign n37873 = pi18 ? n37872 : ~n508;
  assign n37874 = pi17 ? n32 : n37873;
  assign n37875 = pi16 ? n32 : n37874;
  assign n37876 = pi15 ? n37814 : n37875;
  assign n37877 = pi14 ? n37876 : n37820;
  assign n37878 = pi13 ? n37811 : n37877;
  assign n37879 = pi19 ? n28408 : n32;
  assign n37880 = pi18 ? n863 : n37879;
  assign n37881 = pi17 ? n32 : n37880;
  assign n37882 = pi16 ? n32 : n37881;
  assign n37883 = pi16 ? n2851 : ~n37830;
  assign n37884 = pi15 ? n37882 : n37883;
  assign n37885 = pi14 ? n37823 : n37884;
  assign n37886 = pi18 ? n6867 : n32;
  assign n37887 = pi17 ? n37886 : n37837;
  assign n37888 = pi16 ? n16396 : n37887;
  assign n37889 = pi16 ? n2851 : ~n37840;
  assign n37890 = pi15 ? n37888 : n37889;
  assign n37891 = pi16 ? n3061 : ~n3769;
  assign n37892 = pi16 ? n2837 : ~n3769;
  assign n37893 = pi15 ? n37891 : n37892;
  assign n37894 = pi14 ? n37890 : n37893;
  assign n37895 = pi13 ? n37885 : n37894;
  assign n37896 = pi12 ? n37878 : n37895;
  assign n37897 = pi11 ? n37870 : n37896;
  assign n37898 = pi10 ? n37866 : n37897;
  assign n37899 = pi09 ? n32 : n37898;
  assign n37900 = pi08 ? n37849 : n37899;
  assign n37901 = pi14 ? n17298 : n17435;
  assign n37902 = pi15 ? n25749 : n32;
  assign n37903 = pi14 ? n25753 : n37902;
  assign n37904 = pi13 ? n37901 : n37903;
  assign n37905 = pi14 ? n25557 : n25556;
  assign n37906 = pi15 ? n25814 : n17039;
  assign n37907 = pi14 ? n37906 : n25378;
  assign n37908 = pi13 ? n37905 : n37907;
  assign n37909 = pi12 ? n37904 : n37908;
  assign n37910 = pi15 ? n16452 : n14985;
  assign n37911 = pi15 ? n14985 : n16392;
  assign n37912 = pi14 ? n37910 : n37911;
  assign n37913 = pi14 ? n32 : n16392;
  assign n37914 = pi13 ? n37912 : n37913;
  assign n37915 = pi15 ? n16105 : n24874;
  assign n37916 = pi14 ? n32 : n37915;
  assign n37917 = pi13 ? n32 : n37916;
  assign n37918 = pi12 ? n37914 : n37917;
  assign n37919 = pi11 ? n37909 : n37918;
  assign n37920 = pi19 ? n507 : ~n2303;
  assign n37921 = pi18 ? n32 : n37920;
  assign n37922 = pi17 ? n32 : n37921;
  assign n37923 = pi16 ? n32 : n37922;
  assign n37924 = pi15 ? n37923 : n15230;
  assign n37925 = pi15 ? n15230 : n24700;
  assign n37926 = pi14 ? n37924 : n37925;
  assign n37927 = pi15 ? n24700 : n24511;
  assign n37928 = pi19 ? n32 : n10662;
  assign n37929 = pi18 ? n32 : n37928;
  assign n37930 = pi17 ? n32 : n37929;
  assign n37931 = pi16 ? n32 : n37930;
  assign n37932 = pi15 ? n24504 : n37931;
  assign n37933 = pi14 ? n37927 : n37932;
  assign n37934 = pi13 ? n37926 : n37933;
  assign n37935 = pi14 ? n26017 : n24161;
  assign n37936 = pi14 ? n23484 : n27028;
  assign n37937 = pi13 ? n37935 : n37936;
  assign n37938 = pi12 ? n37934 : n37937;
  assign n37939 = pi19 ? n32 : n24204;
  assign n37940 = pi18 ? n37939 : ~n34229;
  assign n37941 = pi17 ? n32 : n37940;
  assign n37942 = pi16 ? n32 : n37941;
  assign n37943 = pi15 ? n22817 : n37942;
  assign n37944 = pi14 ? n32 : n37943;
  assign n37945 = pi18 ? n28178 : ~n508;
  assign n37946 = pi17 ? n32 : n37945;
  assign n37947 = pi16 ? n32 : n37946;
  assign n37948 = pi15 ? n37947 : n13040;
  assign n37949 = pi14 ? n37948 : n33939;
  assign n37950 = pi13 ? n37944 : n37949;
  assign n37951 = pi15 ? n32 : n33939;
  assign n37952 = pi19 ? n1757 : n5688;
  assign n37953 = pi18 ? n32 : n37952;
  assign n37954 = pi19 ? n32 : n786;
  assign n37955 = pi18 ? n37954 : ~n36646;
  assign n37956 = pi17 ? n37953 : ~n37955;
  assign n37957 = pi16 ? n2958 : ~n37956;
  assign n37958 = pi17 ? n1718 : ~n14395;
  assign n37959 = pi16 ? n2958 : ~n37958;
  assign n37960 = pi15 ? n37957 : n37959;
  assign n37961 = pi14 ? n37951 : n37960;
  assign n37962 = pi16 ? n17366 : n34851;
  assign n37963 = pi20 ? n10644 : n207;
  assign n37964 = pi19 ? n37963 : ~n32;
  assign n37965 = pi18 ? n37964 : ~n32;
  assign n37966 = pi17 ? n37965 : ~n32;
  assign n37967 = pi16 ? n2958 : ~n37966;
  assign n37968 = pi15 ? n37962 : n37967;
  assign n37969 = pi16 ? n2958 : ~n2409;
  assign n37970 = pi16 ? n2958 : ~n3769;
  assign n37971 = pi15 ? n37969 : n37970;
  assign n37972 = pi14 ? n37968 : n37971;
  assign n37973 = pi13 ? n37961 : n37972;
  assign n37974 = pi12 ? n37950 : n37973;
  assign n37975 = pi11 ? n37938 : n37974;
  assign n37976 = pi10 ? n37919 : n37975;
  assign n37977 = pi09 ? n32 : n37976;
  assign n37978 = pi19 ? n32 : n22603;
  assign n37979 = pi18 ? n32 : n37978;
  assign n37980 = pi17 ? n32 : n37979;
  assign n37981 = pi16 ? n32 : n37980;
  assign n37982 = pi15 ? n37981 : n17298;
  assign n37983 = pi14 ? n37982 : n37902;
  assign n37984 = pi13 ? n37983 : n17336;
  assign n37985 = pi14 ? n17578 : n17435;
  assign n37986 = pi15 ? n16804 : n17039;
  assign n37987 = pi14 ? n37986 : n25378;
  assign n37988 = pi13 ? n37985 : n37987;
  assign n37989 = pi12 ? n37984 : n37988;
  assign n37990 = pi15 ? n16105 : n25384;
  assign n37991 = pi14 ? n32 : n37990;
  assign n37992 = pi13 ? n32 : n37991;
  assign n37993 = pi12 ? n37914 : n37992;
  assign n37994 = pi11 ? n37989 : n37993;
  assign n37995 = pi19 ? n507 : ~n429;
  assign n37996 = pi18 ? n32 : n37995;
  assign n37997 = pi17 ? n32 : n37996;
  assign n37998 = pi16 ? n32 : n37997;
  assign n37999 = pi15 ? n37998 : n15230;
  assign n38000 = pi14 ? n37999 : n37925;
  assign n38001 = pi19 ? n32 : n20354;
  assign n38002 = pi18 ? n32 : n38001;
  assign n38003 = pi17 ? n32 : n38002;
  assign n38004 = pi16 ? n32 : n38003;
  assign n38005 = pi15 ? n24504 : n38004;
  assign n38006 = pi14 ? n37927 : n38005;
  assign n38007 = pi13 ? n38000 : n38006;
  assign n38008 = pi21 ? n259 : n85;
  assign n38009 = pi20 ? n38008 : n32;
  assign n38010 = pi19 ? n32 : n38009;
  assign n38011 = pi18 ? n32 : n38010;
  assign n38012 = pi17 ? n32 : n38011;
  assign n38013 = pi16 ? n32 : n38012;
  assign n38014 = pi15 ? n38013 : n16105;
  assign n38015 = pi14 ? n38014 : n24161;
  assign n38016 = pi13 ? n38015 : n37936;
  assign n38017 = pi12 ? n38007 : n38016;
  assign n38018 = pi18 ? n1592 : ~n34229;
  assign n38019 = pi17 ? n32 : n38018;
  assign n38020 = pi16 ? n32 : n38019;
  assign n38021 = pi15 ? n22817 : n38020;
  assign n38022 = pi14 ? n32 : n38021;
  assign n38023 = pi13 ? n38022 : n37949;
  assign n38024 = pi18 ? n4127 : ~n36646;
  assign n38025 = pi17 ? n37953 : ~n38024;
  assign n38026 = pi16 ? n3588 : ~n38025;
  assign n38027 = pi16 ? n3588 : ~n37958;
  assign n38028 = pi15 ? n38026 : n38027;
  assign n38029 = pi14 ? n37951 : n38028;
  assign n38030 = pi20 ? n314 : ~n1685;
  assign n38031 = pi19 ? n38030 : ~n32;
  assign n38032 = pi18 ? n38031 : ~n32;
  assign n38033 = pi17 ? n38032 : ~n34850;
  assign n38034 = pi16 ? n3588 : ~n38033;
  assign n38035 = pi20 ? n207 : n339;
  assign n38036 = pi19 ? n38035 : ~n32;
  assign n38037 = pi18 ? n38036 : ~n32;
  assign n38038 = pi17 ? n38037 : ~n32;
  assign n38039 = pi16 ? n3165 : ~n38038;
  assign n38040 = pi15 ? n38034 : n38039;
  assign n38041 = pi16 ? n3047 : ~n2409;
  assign n38042 = pi16 ? n3047 : ~n3769;
  assign n38043 = pi15 ? n38041 : n38042;
  assign n38044 = pi14 ? n38040 : n38043;
  assign n38045 = pi13 ? n38029 : n38044;
  assign n38046 = pi12 ? n38023 : n38045;
  assign n38047 = pi11 ? n38017 : n38046;
  assign n38048 = pi10 ? n37994 : n38047;
  assign n38049 = pi09 ? n32 : n38048;
  assign n38050 = pi08 ? n37977 : n38049;
  assign n38051 = pi07 ? n37900 : n38050;
  assign n38052 = pi06 ? n37754 : n38051;
  assign n38053 = pi15 ? n25902 : n25904;
  assign n38054 = pi14 ? n38053 : n17336;
  assign n38055 = pi13 ? n38054 : n17336;
  assign n38056 = pi14 ? n17271 : n27675;
  assign n38057 = pi14 ? n17121 : n16393;
  assign n38058 = pi13 ? n38056 : n38057;
  assign n38059 = pi12 ? n38055 : n38058;
  assign n38060 = pi15 ? n32 : n25708;
  assign n38061 = pi20 ? n207 : ~n243;
  assign n38062 = pi19 ? n32 : n38061;
  assign n38063 = pi18 ? n32 : n38062;
  assign n38064 = pi17 ? n32 : n38063;
  assign n38065 = pi16 ? n32 : n38064;
  assign n38066 = pi15 ? n25708 : n38065;
  assign n38067 = pi14 ? n38060 : n38066;
  assign n38068 = pi19 ? n32 : n21167;
  assign n38069 = pi18 ? n32 : n38068;
  assign n38070 = pi17 ? n32 : n38069;
  assign n38071 = pi16 ? n32 : n38070;
  assign n38072 = pi15 ? n25563 : n38071;
  assign n38073 = pi14 ? n38072 : n26330;
  assign n38074 = pi13 ? n38067 : n38073;
  assign n38075 = pi15 ? n16837 : n25211;
  assign n38076 = pi14 ? n32 : n38075;
  assign n38077 = pi13 ? n32 : n38076;
  assign n38078 = pi12 ? n38074 : n38077;
  assign n38079 = pi11 ? n38059 : n38078;
  assign n38080 = pi15 ? n25211 : n16452;
  assign n38081 = pi14 ? n38080 : n16101;
  assign n38082 = pi15 ? n25044 : n16298;
  assign n38083 = pi19 ? n32 : n7853;
  assign n38084 = pi18 ? n32 : n38083;
  assign n38085 = pi17 ? n32 : n38084;
  assign n38086 = pi16 ? n32 : n38085;
  assign n38087 = pi15 ? n38086 : n16105;
  assign n38088 = pi14 ? n38082 : n38087;
  assign n38089 = pi13 ? n38081 : n38088;
  assign n38090 = pi15 ? n38004 : n37931;
  assign n38091 = pi15 ? n24247 : n24382;
  assign n38092 = pi14 ? n38090 : n38091;
  assign n38093 = pi15 ? n24247 : n23933;
  assign n38094 = pi14 ? n38093 : n22818;
  assign n38095 = pi13 ? n38092 : n38094;
  assign n38096 = pi12 ? n38089 : n38095;
  assign n38097 = pi20 ? n32 : ~n17712;
  assign n38098 = pi19 ? n38097 : n32;
  assign n38099 = pi18 ? n32 : n38098;
  assign n38100 = pi17 ? n32 : n38099;
  assign n38101 = pi16 ? n32 : n38100;
  assign n38102 = pi15 ? n14138 : n38101;
  assign n38103 = pi14 ? n22817 : n38102;
  assign n38104 = pi18 ? n268 : n23440;
  assign n38105 = pi17 ? n32 : n38104;
  assign n38106 = pi16 ? n32 : n38105;
  assign n38107 = pi15 ? n38106 : n22437;
  assign n38108 = pi15 ? n21853 : n14389;
  assign n38109 = pi14 ? n38107 : n38108;
  assign n38110 = pi13 ? n38103 : n38109;
  assign n38111 = pi18 ? n268 : n20020;
  assign n38112 = pi17 ? n32 : n38111;
  assign n38113 = pi16 ? n32 : n38112;
  assign n38114 = pi18 ? n268 : n5502;
  assign n38115 = pi17 ? n32 : n38114;
  assign n38116 = pi16 ? n32 : n38115;
  assign n38117 = pi15 ? n38113 : n38116;
  assign n38118 = pi18 ? n36119 : ~n9012;
  assign n38119 = pi17 ? n32 : n38118;
  assign n38120 = pi16 ? n3438 : ~n38119;
  assign n38121 = pi19 ? n5675 : n236;
  assign n38122 = pi18 ? n38121 : ~n32;
  assign n38123 = pi17 ? n38122 : ~n14395;
  assign n38124 = pi16 ? n3438 : ~n38123;
  assign n38125 = pi15 ? n38120 : n38124;
  assign n38126 = pi14 ? n38117 : n38125;
  assign n38127 = pi19 ? n4670 : n349;
  assign n38128 = pi18 ? n38127 : ~n32;
  assign n38129 = pi17 ? n38128 : ~n14387;
  assign n38130 = pi16 ? n3438 : ~n38129;
  assign n38131 = pi16 ? n3156 : n14388;
  assign n38132 = pi15 ? n38130 : n38131;
  assign n38133 = pi16 ? n3438 : ~n3769;
  assign n38134 = pi14 ? n38132 : n38133;
  assign n38135 = pi13 ? n38126 : n38134;
  assign n38136 = pi12 ? n38110 : n38135;
  assign n38137 = pi11 ? n38096 : n38136;
  assign n38138 = pi10 ? n38079 : n38137;
  assign n38139 = pi09 ? n32 : n38138;
  assign n38140 = pi14 ? n25904 : n32;
  assign n38141 = pi15 ? n25904 : n25902;
  assign n38142 = pi14 ? n38141 : n38053;
  assign n38143 = pi13 ? n38140 : n38142;
  assign n38144 = pi15 ? n17121 : n25997;
  assign n38145 = pi14 ? n26047 : n38144;
  assign n38146 = pi15 ? n17261 : n17298;
  assign n38147 = pi15 ? n17336 : n16392;
  assign n38148 = pi14 ? n38146 : n38147;
  assign n38149 = pi13 ? n38145 : n38148;
  assign n38150 = pi12 ? n38143 : n38149;
  assign n38151 = pi20 ? n67 : ~n243;
  assign n38152 = pi19 ? n32 : n38151;
  assign n38153 = pi18 ? n32 : n38152;
  assign n38154 = pi17 ? n32 : n38153;
  assign n38155 = pi16 ? n32 : n38154;
  assign n38156 = pi15 ? n38155 : n38071;
  assign n38157 = pi14 ? n38156 : n26330;
  assign n38158 = pi13 ? n38067 : n38157;
  assign n38159 = pi15 ? n16392 : n15403;
  assign n38160 = pi14 ? n32 : n38159;
  assign n38161 = pi13 ? n32 : n38160;
  assign n38162 = pi12 ? n38158 : n38161;
  assign n38163 = pi11 ? n38150 : n38162;
  assign n38164 = pi15 ? n15403 : n16452;
  assign n38165 = pi14 ? n38164 : n16101;
  assign n38166 = pi15 ? n16101 : n16298;
  assign n38167 = pi14 ? n38166 : n25215;
  assign n38168 = pi13 ? n38165 : n38167;
  assign n38169 = pi14 ? n37931 : n37789;
  assign n38170 = pi13 ? n38169 : n38094;
  assign n38171 = pi12 ? n38168 : n38170;
  assign n38172 = pi19 ? n4721 : n32;
  assign n38173 = pi18 ? n32 : n38172;
  assign n38174 = pi17 ? n32 : n38173;
  assign n38175 = pi16 ? n32 : n38174;
  assign n38176 = pi15 ? n14138 : n38175;
  assign n38177 = pi14 ? n22817 : n38176;
  assign n38178 = pi13 ? n38177 : n38109;
  assign n38179 = pi17 ? n3557 : ~n38118;
  assign n38180 = pi16 ? n32 : n38179;
  assign n38181 = pi20 ? n726 : ~n266;
  assign n38182 = pi19 ? n38181 : ~n236;
  assign n38183 = pi18 ? n38182 : n32;
  assign n38184 = pi17 ? n38183 : n14395;
  assign n38185 = pi16 ? n32 : n38184;
  assign n38186 = pi15 ? n38180 : n38185;
  assign n38187 = pi14 ? n38117 : n38186;
  assign n38188 = pi20 ? n726 : ~n32;
  assign n38189 = pi19 ? n38188 : ~n349;
  assign n38190 = pi18 ? n38189 : n32;
  assign n38191 = pi17 ? n38190 : n14387;
  assign n38192 = pi16 ? n32 : n38191;
  assign n38193 = pi18 ? n38 : n32;
  assign n38194 = pi17 ? n38193 : n14387;
  assign n38195 = pi16 ? n32 : n38194;
  assign n38196 = pi15 ? n38192 : n38195;
  assign n38197 = pi17 ? n1028 : ~n2519;
  assign n38198 = pi16 ? n32 : n38197;
  assign n38199 = pi14 ? n38196 : n38198;
  assign n38200 = pi13 ? n38187 : n38199;
  assign n38201 = pi12 ? n38178 : n38200;
  assign n38202 = pi11 ? n38171 : n38201;
  assign n38203 = pi10 ? n38163 : n38202;
  assign n38204 = pi09 ? n32 : n38203;
  assign n38205 = pi08 ? n38139 : n38204;
  assign n38206 = pi19 ? n32 : n14401;
  assign n38207 = pi18 ? n32 : n38206;
  assign n38208 = pi17 ? n32 : n38207;
  assign n38209 = pi16 ? n32 : n38208;
  assign n38210 = pi15 ? n25988 : n38209;
  assign n38211 = pi15 ? n38209 : n25902;
  assign n38212 = pi14 ? n38210 : n38211;
  assign n38213 = pi13 ? n38212 : n25904;
  assign n38214 = pi15 ? n32 : n25997;
  assign n38215 = pi14 ? n17271 : n38214;
  assign n38216 = pi15 ? n17261 : n32;
  assign n38217 = pi14 ? n38216 : n32;
  assign n38218 = pi13 ? n38215 : n38217;
  assign n38219 = pi12 ? n38213 : n38218;
  assign n38220 = pi15 ? n32 : n16237;
  assign n38221 = pi20 ? n3523 : ~n207;
  assign n38222 = pi19 ? n32 : n38221;
  assign n38223 = pi18 ? n32 : n38222;
  assign n38224 = pi17 ? n32 : n38223;
  assign n38225 = pi16 ? n32 : n38224;
  assign n38226 = pi15 ? n16237 : n38225;
  assign n38227 = pi14 ? n38220 : n38226;
  assign n38228 = pi15 ? n17121 : n15847;
  assign n38229 = pi14 ? n38228 : n16392;
  assign n38230 = pi13 ? n38227 : n38229;
  assign n38231 = pi14 ? n24563 : n24498;
  assign n38232 = pi14 ? n17188 : n38159;
  assign n38233 = pi13 ? n38231 : n38232;
  assign n38234 = pi12 ? n38230 : n38233;
  assign n38235 = pi11 ? n38219 : n38234;
  assign n38236 = pi15 ? n15403 : n27662;
  assign n38237 = pi14 ? n38236 : n27662;
  assign n38238 = pi15 ? n26880 : n16452;
  assign n38239 = pi15 ? n16298 : n16308;
  assign n38240 = pi14 ? n38238 : n38239;
  assign n38241 = pi13 ? n38237 : n38240;
  assign n38242 = pi15 ? n38086 : n16308;
  assign n38243 = pi14 ? n38242 : n24511;
  assign n38244 = pi14 ? n24247 : n22541;
  assign n38245 = pi13 ? n38243 : n38244;
  assign n38246 = pi12 ? n38241 : n38245;
  assign n38247 = pi19 ? n4867 : ~n236;
  assign n38248 = pi18 ? n32 : n38247;
  assign n38249 = pi17 ? n32 : n38248;
  assign n38250 = pi16 ? n32 : n38249;
  assign n38251 = pi15 ? n25346 : n38250;
  assign n38252 = pi14 ? n22543 : n38251;
  assign n38253 = pi15 ? n27466 : n25247;
  assign n38254 = pi19 ? n1325 : n32;
  assign n38255 = pi18 ? n32 : n38254;
  assign n38256 = pi17 ? n32 : n38255;
  assign n38257 = pi16 ? n32 : n38256;
  assign n38258 = pi15 ? n38257 : n33970;
  assign n38259 = pi14 ? n38253 : n38258;
  assign n38260 = pi13 ? n38252 : n38259;
  assign n38261 = pi15 ? n23443 : n22825;
  assign n38262 = pi17 ? n3704 : ~n38118;
  assign n38263 = pi16 ? n32 : n38262;
  assign n38264 = pi19 ? n5597 : n1844;
  assign n38265 = pi18 ? n38264 : n32;
  assign n38266 = pi17 ? n38265 : n14395;
  assign n38267 = pi16 ? n32 : n38266;
  assign n38268 = pi15 ? n38263 : n38267;
  assign n38269 = pi14 ? n38261 : n38268;
  assign n38270 = pi18 ? n12598 : n32;
  assign n38271 = pi17 ? n38270 : n20021;
  assign n38272 = pi16 ? n32 : n38271;
  assign n38273 = pi20 ? n1368 : n220;
  assign n38274 = pi19 ? n38273 : n32;
  assign n38275 = pi18 ? n32 : n38274;
  assign n38276 = pi17 ? n38265 : n38275;
  assign n38277 = pi16 ? n32 : n38276;
  assign n38278 = pi15 ? n38272 : n38277;
  assign n38279 = pi17 ? n4041 : ~n2519;
  assign n38280 = pi16 ? n32 : n38279;
  assign n38281 = pi17 ? n1500 : ~n2519;
  assign n38282 = pi16 ? n32 : n38281;
  assign n38283 = pi15 ? n38280 : n38282;
  assign n38284 = pi14 ? n38278 : n38283;
  assign n38285 = pi13 ? n38269 : n38284;
  assign n38286 = pi12 ? n38260 : n38285;
  assign n38287 = pi11 ? n38246 : n38286;
  assign n38288 = pi10 ? n38235 : n38287;
  assign n38289 = pi09 ? n32 : n38288;
  assign n38290 = pi15 ? n25988 : n25904;
  assign n38291 = pi14 ? n25984 : n38290;
  assign n38292 = pi14 ? n25988 : n25984;
  assign n38293 = pi13 ? n38291 : n38292;
  assign n38294 = pi15 ? n32 : n26479;
  assign n38295 = pi14 ? n26147 : n38294;
  assign n38296 = pi14 ? n27376 : n32;
  assign n38297 = pi13 ? n38295 : n38296;
  assign n38298 = pi12 ? n38293 : n38297;
  assign n38299 = pi15 ? n16832 : n15403;
  assign n38300 = pi14 ? n32 : n38299;
  assign n38301 = pi13 ? n38231 : n38300;
  assign n38302 = pi12 ? n38230 : n38301;
  assign n38303 = pi11 ? n38298 : n38302;
  assign n38304 = pi15 ? n15403 : n25384;
  assign n38305 = pi14 ? n38304 : n24874;
  assign n38306 = pi13 ? n38305 : n38240;
  assign n38307 = pi14 ? n38239 : n24511;
  assign n38308 = pi13 ? n38307 : n38244;
  assign n38309 = pi12 ? n38306 : n38308;
  assign n38310 = pi17 ? n3855 : ~n38118;
  assign n38311 = pi16 ? n32 : n38310;
  assign n38312 = pi20 ? n2140 : ~n8644;
  assign n38313 = pi19 ? n38312 : n19773;
  assign n38314 = pi18 ? n38313 : n32;
  assign n38315 = pi17 ? n38314 : n14395;
  assign n38316 = pi16 ? n32 : n38315;
  assign n38317 = pi15 ? n38311 : n38316;
  assign n38318 = pi14 ? n38261 : n38317;
  assign n38319 = pi18 ? n13137 : n32;
  assign n38320 = pi17 ? n38319 : n20021;
  assign n38321 = pi16 ? n32 : n38320;
  assign n38322 = pi18 ? n103 : n32;
  assign n38323 = pi20 ? n175 : n220;
  assign n38324 = pi19 ? n38323 : n32;
  assign n38325 = pi18 ? n32 : n38324;
  assign n38326 = pi17 ? n38322 : n38325;
  assign n38327 = pi16 ? n32 : n38326;
  assign n38328 = pi15 ? n38321 : n38327;
  assign n38329 = pi17 ? n4037 : ~n2519;
  assign n38330 = pi16 ? n32 : n38329;
  assign n38331 = pi17 ? n1605 : ~n2519;
  assign n38332 = pi16 ? n32 : n38331;
  assign n38333 = pi15 ? n38330 : n38332;
  assign n38334 = pi14 ? n38328 : n38333;
  assign n38335 = pi13 ? n38318 : n38334;
  assign n38336 = pi12 ? n38260 : n38335;
  assign n38337 = pi11 ? n38309 : n38336;
  assign n38338 = pi10 ? n38303 : n38337;
  assign n38339 = pi09 ? n32 : n38338;
  assign n38340 = pi08 ? n38289 : n38339;
  assign n38341 = pi07 ? n38205 : n38340;
  assign n38342 = pi15 ? n26096 : n25988;
  assign n38343 = pi14 ? n26096 : n38342;
  assign n38344 = pi13 ? n38343 : n26035;
  assign n38345 = pi14 ? n27376 : n17271;
  assign n38346 = pi13 ? n25904 : n38345;
  assign n38347 = pi12 ? n38344 : n38346;
  assign n38348 = pi15 ? n17121 : n17298;
  assign n38349 = pi14 ? n17121 : n38348;
  assign n38350 = pi15 ? n25997 : n32;
  assign n38351 = pi14 ? n38350 : n16392;
  assign n38352 = pi13 ? n38349 : n38351;
  assign n38353 = pi15 ? n16392 : n25763;
  assign n38354 = pi15 ? n17066 : n32;
  assign n38355 = pi14 ? n38353 : n38354;
  assign n38356 = pi14 ? n26163 : n15847;
  assign n38357 = pi13 ? n38355 : n38356;
  assign n38358 = pi12 ? n38352 : n38357;
  assign n38359 = pi11 ? n38347 : n38358;
  assign n38360 = pi15 ? n15847 : n24874;
  assign n38361 = pi14 ? n38360 : n24874;
  assign n38362 = pi15 ? n25384 : n16452;
  assign n38363 = pi14 ? n38362 : n16452;
  assign n38364 = pi13 ? n38361 : n38363;
  assign n38365 = pi15 ? n24237 : n24640;
  assign n38366 = pi15 ? n38086 : n24511;
  assign n38367 = pi14 ? n38365 : n38366;
  assign n38368 = pi19 ? n32 : ~n502;
  assign n38369 = pi18 ? n32 : n38368;
  assign n38370 = pi17 ? n32 : n38369;
  assign n38371 = pi16 ? n32 : n38370;
  assign n38372 = pi19 ? n32 : n2250;
  assign n38373 = pi18 ? n32 : n38372;
  assign n38374 = pi17 ? n32 : n38373;
  assign n38375 = pi16 ? n32 : n38374;
  assign n38376 = pi15 ? n38371 : n38375;
  assign n38377 = pi14 ? n24504 : n38376;
  assign n38378 = pi13 ? n38367 : n38377;
  assign n38379 = pi12 ? n38364 : n38378;
  assign n38380 = pi15 ? n23250 : n15655;
  assign n38381 = pi14 ? n38380 : n37507;
  assign n38382 = pi14 ? n24742 : n22817;
  assign n38383 = pi13 ? n38381 : n38382;
  assign n38384 = pi18 ? n2424 : ~n21888;
  assign n38385 = pi18 ? n23073 : ~n9012;
  assign n38386 = pi17 ? n38384 : ~n38385;
  assign n38387 = pi16 ? n32 : n38386;
  assign n38388 = pi20 ? n206 : ~n518;
  assign n38389 = pi19 ? n244 : n38388;
  assign n38390 = pi18 ? n38389 : n20020;
  assign n38391 = pi17 ? n38390 : n32;
  assign n38392 = pi16 ? n32 : n38391;
  assign n38393 = pi15 ? n38387 : n38392;
  assign n38394 = pi14 ? n32 : n38393;
  assign n38395 = pi19 ? n244 : n17194;
  assign n38396 = pi18 ? n38395 : n32;
  assign n38397 = pi17 ? n38396 : n32;
  assign n38398 = pi16 ? n32 : n38397;
  assign n38399 = pi21 ? n66 : n309;
  assign n38400 = pi20 ? n32 : n38399;
  assign n38401 = pi19 ? n38400 : n28976;
  assign n38402 = pi19 ? n18722 : n18728;
  assign n38403 = pi18 ? n38401 : ~n38402;
  assign n38404 = pi20 ? n174 : ~n10644;
  assign n38405 = pi20 ? n173 : n3897;
  assign n38406 = pi19 ? n38404 : n38405;
  assign n38407 = pi20 ? n11107 : ~n266;
  assign n38408 = pi19 ? n38407 : ~n32;
  assign n38409 = pi18 ? n38406 : n38408;
  assign n38410 = pi17 ? n38403 : ~n38409;
  assign n38411 = pi16 ? n32 : n38410;
  assign n38412 = pi15 ? n38398 : n38411;
  assign n38413 = pi17 ? n5541 : ~n2519;
  assign n38414 = pi16 ? n32 : n38413;
  assign n38415 = pi17 ? n2355 : ~n2519;
  assign n38416 = pi16 ? n32 : n38415;
  assign n38417 = pi15 ? n38414 : n38416;
  assign n38418 = pi14 ? n38412 : n38417;
  assign n38419 = pi13 ? n38394 : n38418;
  assign n38420 = pi12 ? n38383 : n38419;
  assign n38421 = pi11 ? n38379 : n38420;
  assign n38422 = pi10 ? n38359 : n38421;
  assign n38423 = pi09 ? n32 : n38422;
  assign n38424 = pi19 ? n32 : n654;
  assign n38425 = pi18 ? n32 : n38424;
  assign n38426 = pi17 ? n32 : n38425;
  assign n38427 = pi16 ? n32 : n38426;
  assign n38428 = pi15 ? n38427 : n25988;
  assign n38429 = pi14 ? n26096 : n38428;
  assign n38430 = pi13 ? n38429 : n26101;
  assign n38431 = pi15 ? n25904 : n25984;
  assign n38432 = pi14 ? n25904 : n38431;
  assign n38433 = pi15 ? n17216 : n25988;
  assign n38434 = pi15 ? n25988 : n17121;
  assign n38435 = pi14 ? n38433 : n38434;
  assign n38436 = pi13 ? n38432 : n38435;
  assign n38437 = pi12 ? n38430 : n38436;
  assign n38438 = pi14 ? n37568 : n16485;
  assign n38439 = pi13 ? n38355 : n38438;
  assign n38440 = pi12 ? n38352 : n38439;
  assign n38441 = pi11 ? n38437 : n38440;
  assign n38442 = pi15 ? n25384 : n26009;
  assign n38443 = pi20 ? n14953 : n32;
  assign n38444 = pi19 ? n32 : n38443;
  assign n38445 = pi18 ? n32 : n38444;
  assign n38446 = pi17 ? n32 : n38445;
  assign n38447 = pi16 ? n32 : n38446;
  assign n38448 = pi15 ? n38447 : n24874;
  assign n38449 = pi14 ? n38442 : n38448;
  assign n38450 = pi13 ? n25384 : n38449;
  assign n38451 = pi15 ? n26885 : n24511;
  assign n38452 = pi15 ? n24237 : n24511;
  assign n38453 = pi14 ? n38451 : n38452;
  assign n38454 = pi14 ? n26919 : n38376;
  assign n38455 = pi13 ? n38453 : n38454;
  assign n38456 = pi12 ? n38450 : n38455;
  assign n38457 = pi14 ? n23250 : n37507;
  assign n38458 = pi13 ? n38457 : n38382;
  assign n38459 = pi18 ? n2754 : ~n21888;
  assign n38460 = pi17 ? n38459 : ~n38385;
  assign n38461 = pi16 ? n32 : n38460;
  assign n38462 = pi19 ? n1840 : n38388;
  assign n38463 = pi18 ? n38462 : n20020;
  assign n38464 = pi17 ? n38463 : n32;
  assign n38465 = pi16 ? n32 : n38464;
  assign n38466 = pi15 ? n38461 : n38465;
  assign n38467 = pi14 ? n32 : n38466;
  assign n38468 = pi20 ? n274 : ~n10889;
  assign n38469 = pi19 ? n1840 : n38468;
  assign n38470 = pi18 ? n38469 : n32;
  assign n38471 = pi17 ? n38470 : n32;
  assign n38472 = pi16 ? n32 : n38471;
  assign n38473 = pi19 ? n6398 : n28686;
  assign n38474 = pi18 ? n38473 : ~n38402;
  assign n38475 = pi17 ? n38474 : ~n38409;
  assign n38476 = pi16 ? n32 : n38475;
  assign n38477 = pi15 ? n38472 : n38476;
  assign n38478 = pi17 ? n2461 : ~n2519;
  assign n38479 = pi16 ? n32 : n38478;
  assign n38480 = pi15 ? n5773 : n38479;
  assign n38481 = pi14 ? n38477 : n38480;
  assign n38482 = pi13 ? n38467 : n38481;
  assign n38483 = pi12 ? n38458 : n38482;
  assign n38484 = pi11 ? n38456 : n38483;
  assign n38485 = pi10 ? n38441 : n38484;
  assign n38486 = pi09 ? n32 : n38485;
  assign n38487 = pi08 ? n38423 : n38486;
  assign n38488 = pi15 ? n26183 : n26189;
  assign n38489 = pi15 ? n26183 : n26096;
  assign n38490 = pi14 ? n38488 : n38489;
  assign n38491 = pi15 ? n17348 : n32;
  assign n38492 = pi14 ? n26136 : n38491;
  assign n38493 = pi13 ? n38490 : n38492;
  assign n38494 = pi14 ? n25905 : n26031;
  assign n38495 = pi14 ? n26034 : n17271;
  assign n38496 = pi13 ? n38494 : n38495;
  assign n38497 = pi12 ? n38493 : n38496;
  assign n38498 = pi15 ? n17435 : n25904;
  assign n38499 = pi15 ? n17431 : n17061;
  assign n38500 = pi14 ? n38498 : n38499;
  assign n38501 = pi14 ? n27443 : n16392;
  assign n38502 = pi13 ? n38500 : n38501;
  assign n38503 = pi15 ? n16392 : n16984;
  assign n38504 = pi14 ? n38503 : n38354;
  assign n38505 = pi15 ? n17066 : n17039;
  assign n38506 = pi14 ? n38505 : n15847;
  assign n38507 = pi13 ? n38504 : n38506;
  assign n38508 = pi12 ? n38502 : n38507;
  assign n38509 = pi11 ? n38497 : n38508;
  assign n38510 = pi14 ? n16452 : n26806;
  assign n38511 = pi15 ? n16546 : n26009;
  assign n38512 = pi14 ? n38511 : n38448;
  assign n38513 = pi13 ? n38510 : n38512;
  assign n38514 = pi15 ? n16452 : n24247;
  assign n38515 = pi14 ? n24882 : n38514;
  assign n38516 = pi15 ? n24247 : n15834;
  assign n38517 = pi14 ? n16105 : n38516;
  assign n38518 = pi13 ? n38515 : n38517;
  assign n38519 = pi12 ? n38513 : n38518;
  assign n38520 = pi20 ? n321 : ~n6050;
  assign n38521 = pi19 ? n32 : n38520;
  assign n38522 = pi18 ? n595 : ~n38521;
  assign n38523 = pi18 ? n22159 : ~n9012;
  assign n38524 = pi17 ? n38522 : ~n38523;
  assign n38525 = pi16 ? n32 : n38524;
  assign n38526 = pi19 ? n247 : n6158;
  assign n38527 = pi18 ? n4098 : ~n38526;
  assign n38528 = pi18 ? n22159 : ~n32;
  assign n38529 = pi17 ? n38527 : ~n38528;
  assign n38530 = pi16 ? n32 : n38529;
  assign n38531 = pi15 ? n38525 : n38530;
  assign n38532 = pi14 ? n32 : n38531;
  assign n38533 = pi19 ? n1574 : ~n5741;
  assign n38534 = pi18 ? n38533 : n6059;
  assign n38535 = pi17 ? n38534 : n32;
  assign n38536 = pi16 ? n32 : n38535;
  assign n38537 = pi20 ? n17287 : n339;
  assign n38538 = pi19 ? n32 : n38537;
  assign n38539 = pi20 ? n6085 : n3523;
  assign n38540 = pi20 ? n3843 : n448;
  assign n38541 = pi19 ? n38539 : n38540;
  assign n38542 = pi18 ? n38538 : ~n38541;
  assign n38543 = pi20 ? n175 : n974;
  assign n38544 = pi19 ? n38543 : n32;
  assign n38545 = pi20 ? n3847 : n321;
  assign n38546 = pi19 ? n38545 : ~n32;
  assign n38547 = pi18 ? n38544 : n38546;
  assign n38548 = pi17 ? n38542 : ~n38547;
  assign n38549 = pi16 ? n32 : n38548;
  assign n38550 = pi15 ? n38536 : n38549;
  assign n38551 = pi17 ? n1480 : ~n2517;
  assign n38552 = pi16 ? n32 : n38551;
  assign n38553 = pi15 ? n5937 : n38552;
  assign n38554 = pi14 ? n38550 : n38553;
  assign n38555 = pi13 ? n38532 : n38554;
  assign n38556 = pi12 ? n38383 : n38555;
  assign n38557 = pi11 ? n38519 : n38556;
  assign n38558 = pi10 ? n38509 : n38557;
  assign n38559 = pi09 ? n32 : n38558;
  assign n38560 = pi15 ? n26183 : n32;
  assign n38561 = pi14 ? n26190 : n38560;
  assign n38562 = pi13 ? n38490 : n38561;
  assign n38563 = pi14 ? n25905 : n26097;
  assign n38564 = pi14 ? n26100 : n17271;
  assign n38565 = pi13 ? n38563 : n38564;
  assign n38566 = pi12 ? n38562 : n38565;
  assign n38567 = pi14 ? n26111 : n38071;
  assign n38568 = pi13 ? n38504 : n38567;
  assign n38569 = pi12 ? n38502 : n38568;
  assign n38570 = pi11 ? n38566 : n38569;
  assign n38571 = pi20 ? n518 : ~n220;
  assign n38572 = pi19 ? n32 : n38571;
  assign n38573 = pi18 ? n2730 : ~n38572;
  assign n38574 = pi20 ? n32 : ~n174;
  assign n38575 = pi19 ? n38574 : ~n32;
  assign n38576 = pi18 ? n38575 : ~n9012;
  assign n38577 = pi17 ? n38573 : ~n38576;
  assign n38578 = pi16 ? n32 : n38577;
  assign n38579 = pi19 ? n247 : n589;
  assign n38580 = pi18 ? n2730 : ~n38579;
  assign n38581 = pi18 ? n38575 : ~n32;
  assign n38582 = pi17 ? n38580 : ~n38581;
  assign n38583 = pi16 ? n32 : n38582;
  assign n38584 = pi15 ? n38578 : n38583;
  assign n38585 = pi14 ? n32 : n38584;
  assign n38586 = pi21 ? n1939 : ~n174;
  assign n38587 = pi20 ? n38586 : ~n260;
  assign n38588 = pi19 ? n32 : n38587;
  assign n38589 = pi18 ? n38588 : n19654;
  assign n38590 = pi17 ? n38589 : n21317;
  assign n38591 = pi16 ? n32 : n38590;
  assign n38592 = pi17 ? n2159 : ~n2519;
  assign n38593 = pi16 ? n32 : n38592;
  assign n38594 = pi15 ? n38591 : n38593;
  assign n38595 = pi17 ? n4659 : ~n2519;
  assign n38596 = pi16 ? n32 : n38595;
  assign n38597 = pi17 ? n2159 : ~n2517;
  assign n38598 = pi16 ? n32 : n38597;
  assign n38599 = pi15 ? n38596 : n38598;
  assign n38600 = pi14 ? n38594 : n38599;
  assign n38601 = pi13 ? n38585 : n38600;
  assign n38602 = pi12 ? n38383 : n38601;
  assign n38603 = pi11 ? n38519 : n38602;
  assign n38604 = pi10 ? n38570 : n38603;
  assign n38605 = pi09 ? n32 : n38604;
  assign n38606 = pi08 ? n38559 : n38605;
  assign n38607 = pi07 ? n38487 : n38606;
  assign n38608 = pi06 ? n38341 : n38607;
  assign n38609 = pi05 ? n38052 : n38608;
  assign n38610 = pi04 ? n37457 : n38609;
  assign n38611 = pi03 ? n35883 : n38610;
  assign n38612 = pi02 ? n32460 : n38611;
  assign n38613 = pi01 ? n32 : n38612;
  assign n38614 = pi15 ? n26269 : n26225;
  assign n38615 = pi14 ? n26269 : n38614;
  assign n38616 = pi15 ? n26225 : n32;
  assign n38617 = pi14 ? n26225 : n38616;
  assign n38618 = pi13 ? n38615 : n38617;
  assign n38619 = pi14 ? n26133 : n38491;
  assign n38620 = pi15 ? n17121 : n17435;
  assign n38621 = pi14 ? n38620 : n17121;
  assign n38622 = pi13 ? n38619 : n38621;
  assign n38623 = pi12 ? n38618 : n38622;
  assign n38624 = pi14 ? n16393 : n25984;
  assign n38625 = pi13 ? n38624 : n38296;
  assign n38626 = pi15 ? n17039 : n17336;
  assign n38627 = pi14 ? n38626 : n32;
  assign n38628 = pi15 ? n17061 : n17039;
  assign n38629 = pi14 ? n38628 : n16392;
  assign n38630 = pi13 ? n38627 : n38629;
  assign n38631 = pi12 ? n38625 : n38630;
  assign n38632 = pi11 ? n38623 : n38631;
  assign n38633 = pi14 ? n38353 : n16392;
  assign n38634 = pi15 ? n16546 : n16606;
  assign n38635 = pi15 ? n16515 : n16452;
  assign n38636 = pi14 ? n38634 : n38635;
  assign n38637 = pi13 ? n38633 : n38636;
  assign n38638 = pi15 ? n24700 : n24247;
  assign n38639 = pi14 ? n16452 : n38638;
  assign n38640 = pi14 ? n24247 : n38516;
  assign n38641 = pi13 ? n38639 : n38640;
  assign n38642 = pi12 ? n38637 : n38641;
  assign n38643 = pi15 ? n15834 : n15655;
  assign n38644 = pi14 ? n38643 : n37507;
  assign n38645 = pi15 ? n24742 : n24659;
  assign n38646 = pi14 ? n38645 : n23443;
  assign n38647 = pi13 ? n38644 : n38646;
  assign n38648 = pi18 ? n32 : ~n5335;
  assign n38649 = pi17 ? n1700 : ~n38648;
  assign n38650 = pi16 ? n32 : n38649;
  assign n38651 = pi18 ? n2835 : ~n936;
  assign n38652 = pi20 ? n1368 : n342;
  assign n38653 = pi19 ? n38652 : ~n19191;
  assign n38654 = pi20 ? n342 : ~n10644;
  assign n38655 = pi19 ? n38654 : ~n32;
  assign n38656 = pi18 ? n38653 : n38655;
  assign n38657 = pi17 ? n38651 : ~n38656;
  assign n38658 = pi16 ? n32 : n38657;
  assign n38659 = pi15 ? n38650 : n38658;
  assign n38660 = pi14 ? n23443 : n38659;
  assign n38661 = pi20 ? n1319 : n260;
  assign n38662 = pi19 ? n32 : n38661;
  assign n38663 = pi19 ? n6342 : ~n24349;
  assign n38664 = pi18 ? n38662 : n38663;
  assign n38665 = pi19 ? n17194 : n1757;
  assign n38666 = pi18 ? n38665 : n25116;
  assign n38667 = pi17 ? n38664 : n38666;
  assign n38668 = pi16 ? n32 : n38667;
  assign n38669 = pi15 ? n38668 : n6434;
  assign n38670 = pi17 ? n4804 : ~n2517;
  assign n38671 = pi16 ? n32 : n38670;
  assign n38672 = pi17 ? n1706 : ~n2517;
  assign n38673 = pi16 ? n32 : n38672;
  assign n38674 = pi15 ? n38671 : n38673;
  assign n38675 = pi14 ? n38669 : n38674;
  assign n38676 = pi13 ? n38660 : n38675;
  assign n38677 = pi12 ? n38647 : n38676;
  assign n38678 = pi11 ? n38642 : n38677;
  assign n38679 = pi10 ? n38632 : n38678;
  assign n38680 = pi09 ? n32 : n38679;
  assign n38681 = pi13 ? n38615 : n26269;
  assign n38682 = pi19 ? n32 : n22778;
  assign n38683 = pi18 ? n32 : n38682;
  assign n38684 = pi17 ? n32 : n38683;
  assign n38685 = pi16 ? n32 : n38684;
  assign n38686 = pi21 ? n309 : ~n140;
  assign n38687 = pi20 ? n32 : n38686;
  assign n38688 = pi19 ? n32 : n38687;
  assign n38689 = pi18 ? n32 : n38688;
  assign n38690 = pi17 ? n32 : n38689;
  assign n38691 = pi16 ? n32 : n38690;
  assign n38692 = pi15 ? n38685 : n38691;
  assign n38693 = pi14 ? n38692 : n17121;
  assign n38694 = pi13 ? n38619 : n38693;
  assign n38695 = pi12 ? n38681 : n38694;
  assign n38696 = pi14 ? n25133 : n32;
  assign n38697 = pi13 ? n38696 : n38629;
  assign n38698 = pi12 ? n38625 : n38697;
  assign n38699 = pi11 ? n38695 : n38698;
  assign n38700 = pi15 ? n24742 : n25247;
  assign n38701 = pi14 ? n38700 : n23443;
  assign n38702 = pi13 ? n38644 : n38701;
  assign n38703 = pi17 ? n1232 : ~n38648;
  assign n38704 = pi16 ? n32 : n38703;
  assign n38705 = pi20 ? n357 : n17671;
  assign n38706 = pi19 ? n38705 : n507;
  assign n38707 = pi18 ? n366 : ~n38706;
  assign n38708 = pi19 ? n38652 : ~n18478;
  assign n38709 = pi18 ? n38708 : n38655;
  assign n38710 = pi17 ? n38707 : ~n38709;
  assign n38711 = pi16 ? n32 : n38710;
  assign n38712 = pi15 ? n38704 : n38711;
  assign n38713 = pi14 ? n23443 : n38712;
  assign n38714 = pi19 ? n13074 : ~n24349;
  assign n38715 = pi18 ? n728 : n38714;
  assign n38716 = pi17 ? n38715 : n38666;
  assign n38717 = pi16 ? n32 : n38716;
  assign n38718 = pi17 ? n1134 : ~n2512;
  assign n38719 = pi16 ? n32 : n38718;
  assign n38720 = pi15 ? n38717 : n38719;
  assign n38721 = pi17 ? n930 : ~n2517;
  assign n38722 = pi16 ? n32 : n38721;
  assign n38723 = pi17 ? n1134 : ~n2517;
  assign n38724 = pi16 ? n32 : n38723;
  assign n38725 = pi15 ? n38722 : n38724;
  assign n38726 = pi14 ? n38720 : n38725;
  assign n38727 = pi13 ? n38713 : n38726;
  assign n38728 = pi12 ? n38702 : n38727;
  assign n38729 = pi11 ? n38642 : n38728;
  assign n38730 = pi10 ? n38699 : n38729;
  assign n38731 = pi09 ? n32 : n38730;
  assign n38732 = pi08 ? n38680 : n38731;
  assign n38733 = pi15 ? n17531 : n26354;
  assign n38734 = pi15 ? n26354 : n26269;
  assign n38735 = pi14 ? n38733 : n38734;
  assign n38736 = pi13 ? n38735 : n26269;
  assign n38737 = pi15 ? n17348 : n16984;
  assign n38738 = pi14 ? n26133 : n38737;
  assign n38739 = pi15 ? n16984 : n17435;
  assign n38740 = pi14 ? n38739 : n17435;
  assign n38741 = pi13 ? n38738 : n38740;
  assign n38742 = pi12 ? n38736 : n38741;
  assign n38743 = pi14 ? n17121 : n16850;
  assign n38744 = pi15 ? n16850 : n32;
  assign n38745 = pi14 ? n38744 : n26163;
  assign n38746 = pi13 ? n38743 : n38745;
  assign n38747 = pi19 ? n32 : n20940;
  assign n38748 = pi18 ? n32 : n38747;
  assign n38749 = pi17 ? n32 : n38748;
  assign n38750 = pi16 ? n32 : n38749;
  assign n38751 = pi20 ? n428 : n7487;
  assign n38752 = pi19 ? n32 : n38751;
  assign n38753 = pi18 ? n32 : n38752;
  assign n38754 = pi17 ? n32 : n38753;
  assign n38755 = pi16 ? n32 : n38754;
  assign n38756 = pi15 ? n38750 : n38755;
  assign n38757 = pi15 ? n38750 : n17061;
  assign n38758 = pi14 ? n38756 : n38757;
  assign n38759 = pi14 ? n38628 : n24799;
  assign n38760 = pi13 ? n38758 : n38759;
  assign n38761 = pi12 ? n38746 : n38760;
  assign n38762 = pi11 ? n38742 : n38761;
  assign n38763 = pi14 ? n24799 : n26330;
  assign n38764 = pi13 ? n38763 : n38636;
  assign n38765 = pi14 ? n16452 : n37786;
  assign n38766 = pi13 ? n38765 : n24247;
  assign n38767 = pi12 ? n38764 : n38766;
  assign n38768 = pi20 ? n632 : n32;
  assign n38769 = pi19 ? n32 : n38768;
  assign n38770 = pi18 ? n32 : n38769;
  assign n38771 = pi17 ? n32 : n38770;
  assign n38772 = pi16 ? n32 : n38771;
  assign n38773 = pi15 ? n24247 : n38772;
  assign n38774 = pi14 ? n38773 : n26656;
  assign n38775 = pi15 ? n23340 : n25247;
  assign n38776 = pi14 ? n38775 : n27431;
  assign n38777 = pi13 ? n38774 : n38776;
  assign n38778 = pi20 ? n32 : n8943;
  assign n38779 = pi19 ? n32 : n38778;
  assign n38780 = pi18 ? n38779 : ~n32;
  assign n38781 = pi17 ? n38780 : ~n38648;
  assign n38782 = pi16 ? n32 : n38781;
  assign n38783 = pi21 ? n100 : ~n174;
  assign n38784 = pi20 ? n32 : n38783;
  assign n38785 = pi19 ? n32 : n38784;
  assign n38786 = pi18 ? n38785 : ~n32;
  assign n38787 = pi19 ? n4670 : n267;
  assign n38788 = pi18 ? n38787 : n7090;
  assign n38789 = pi17 ? n38786 : ~n38788;
  assign n38790 = pi16 ? n32 : n38789;
  assign n38791 = pi15 ? n38782 : n38790;
  assign n38792 = pi14 ? n23443 : n38791;
  assign n38793 = pi19 ? n32 : n28686;
  assign n38794 = pi18 ? n38785 : ~n38793;
  assign n38795 = pi20 ? n246 : n206;
  assign n38796 = pi19 ? n28686 : n38795;
  assign n38797 = pi18 ? n38796 : ~n5502;
  assign n38798 = pi17 ? n38794 : ~n38797;
  assign n38799 = pi16 ? n32 : n38798;
  assign n38800 = pi17 ? n1842 : ~n2512;
  assign n38801 = pi16 ? n32 : n38800;
  assign n38802 = pi15 ? n38799 : n38801;
  assign n38803 = pi17 ? n1842 : ~n2519;
  assign n38804 = pi16 ? n32 : n38803;
  assign n38805 = pi17 ? n1842 : ~n2517;
  assign n38806 = pi16 ? n32 : n38805;
  assign n38807 = pi15 ? n38804 : n38806;
  assign n38808 = pi14 ? n38802 : n38807;
  assign n38809 = pi13 ? n38792 : n38808;
  assign n38810 = pi12 ? n38777 : n38809;
  assign n38811 = pi11 ? n38767 : n38810;
  assign n38812 = pi10 ? n38762 : n38811;
  assign n38813 = pi09 ? n32 : n38812;
  assign n38814 = pi15 ? n17531 : n32;
  assign n38815 = pi14 ? n38733 : n38814;
  assign n38816 = pi14 ? n26354 : n38734;
  assign n38817 = pi13 ? n38815 : n38816;
  assign n38818 = pi12 ? n38817 : n38741;
  assign n38819 = pi11 ? n38818 : n38761;
  assign n38820 = pi14 ? n38093 : n26656;
  assign n38821 = pi13 ? n38820 : n38776;
  assign n38822 = pi17 ? n2143 : ~n38648;
  assign n38823 = pi16 ? n32 : n38822;
  assign n38824 = pi17 ? n2143 : ~n38788;
  assign n38825 = pi16 ? n32 : n38824;
  assign n38826 = pi15 ? n38823 : n38825;
  assign n38827 = pi14 ? n23443 : n38826;
  assign n38828 = pi18 ? n936 : ~n38793;
  assign n38829 = pi17 ? n38828 : ~n38797;
  assign n38830 = pi16 ? n32 : n38829;
  assign n38831 = pi15 ? n38830 : n7289;
  assign n38832 = pi17 ? n1576 : ~n2519;
  assign n38833 = pi16 ? n32 : n38832;
  assign n38834 = pi17 ? n1833 : ~n2517;
  assign n38835 = pi16 ? n32 : n38834;
  assign n38836 = pi15 ? n38833 : n38835;
  assign n38837 = pi14 ? n38831 : n38836;
  assign n38838 = pi13 ? n38827 : n38837;
  assign n38839 = pi12 ? n38821 : n38838;
  assign n38840 = pi11 ? n38767 : n38839;
  assign n38841 = pi10 ? n38819 : n38840;
  assign n38842 = pi09 ? n32 : n38841;
  assign n38843 = pi08 ? n38813 : n38842;
  assign n38844 = pi07 ? n38732 : n38843;
  assign n38845 = pi18 ? n32 : n17719;
  assign n38846 = pi17 ? n32 : n38845;
  assign n38847 = pi16 ? n32 : n38846;
  assign n38848 = pi15 ? n38847 : n26269;
  assign n38849 = pi14 ? n17514 : n38848;
  assign n38850 = pi13 ? n26462 : n38849;
  assign n38851 = pi20 ? n32 : n17665;
  assign n38852 = pi19 ? n32 : n38851;
  assign n38853 = pi18 ? n32 : n38852;
  assign n38854 = pi17 ? n32 : n38853;
  assign n38855 = pi16 ? n32 : n38854;
  assign n38856 = pi15 ? n26269 : n38855;
  assign n38857 = pi14 ? n38856 : n38855;
  assign n38858 = pi13 ? n38857 : n32;
  assign n38859 = pi12 ? n38850 : n38858;
  assign n38860 = pi14 ? n32 : n26163;
  assign n38861 = pi13 ? n25491 : n38860;
  assign n38862 = pi15 ? n38750 : n26322;
  assign n38863 = pi14 ? n17039 : n38862;
  assign n38864 = pi14 ? n17061 : n32;
  assign n38865 = pi13 ? n38863 : n38864;
  assign n38866 = pi12 ? n38861 : n38865;
  assign n38867 = pi11 ? n38859 : n38866;
  assign n38868 = pi15 ? n15847 : n16606;
  assign n38869 = pi14 ? n38868 : n38635;
  assign n38870 = pi13 ? n38763 : n38869;
  assign n38871 = pi15 ? n24700 : n16105;
  assign n38872 = pi14 ? n16452 : n38871;
  assign n38873 = pi14 ? n25779 : n24247;
  assign n38874 = pi13 ? n38872 : n38873;
  assign n38875 = pi12 ? n38870 : n38874;
  assign n38876 = pi15 ? n24247 : n32;
  assign n38877 = pi15 ? n22817 : n25247;
  assign n38878 = pi14 ? n38876 : n38877;
  assign n38879 = pi15 ? n22817 : n15119;
  assign n38880 = pi14 ? n38879 : n23443;
  assign n38881 = pi13 ? n38878 : n38880;
  assign n38882 = pi17 ? n2123 : ~n2512;
  assign n38883 = pi16 ? n32 : n38882;
  assign n38884 = pi15 ? n14147 : n38883;
  assign n38885 = pi18 ? n268 : n22307;
  assign n38886 = pi17 ? n2123 : ~n38885;
  assign n38887 = pi16 ? n32 : n38886;
  assign n38888 = pi18 ? n32 : n24548;
  assign n38889 = pi17 ? n3351 : ~n38888;
  assign n38890 = pi16 ? n32 : n38889;
  assign n38891 = pi15 ? n38887 : n38890;
  assign n38892 = pi14 ? n38884 : n38891;
  assign n38893 = pi21 ? n242 : n259;
  assign n38894 = pi20 ? n38893 : ~n32;
  assign n38895 = pi19 ? n38894 : ~n32;
  assign n38896 = pi18 ? n32 : n38895;
  assign n38897 = pi18 ? n32 : n33312;
  assign n38898 = pi17 ? n38896 : ~n38897;
  assign n38899 = pi16 ? n32 : n38898;
  assign n38900 = pi17 ? n2325 : ~n2519;
  assign n38901 = pi16 ? n32 : n38900;
  assign n38902 = pi15 ? n38899 : n38901;
  assign n38903 = pi17 ? n1943 : ~n2519;
  assign n38904 = pi16 ? n32 : n38903;
  assign n38905 = pi14 ? n38902 : n38904;
  assign n38906 = pi13 ? n38892 : n38905;
  assign n38907 = pi12 ? n38881 : n38906;
  assign n38908 = pi11 ? n38875 : n38907;
  assign n38909 = pi10 ? n38867 : n38908;
  assign n38910 = pi09 ? n32 : n38909;
  assign n38911 = pi18 ? n32 : n17699;
  assign n38912 = pi17 ? n32 : n38911;
  assign n38913 = pi16 ? n32 : n38912;
  assign n38914 = pi15 ? n26462 : n38913;
  assign n38915 = pi14 ? n26462 : n38914;
  assign n38916 = pi15 ? n26272 : n26269;
  assign n38917 = pi14 ? n26428 : n38916;
  assign n38918 = pi13 ? n38915 : n38917;
  assign n38919 = pi20 ? n32 : n22458;
  assign n38920 = pi19 ? n32 : n38919;
  assign n38921 = pi18 ? n32 : n38920;
  assign n38922 = pi17 ? n32 : n38921;
  assign n38923 = pi16 ? n32 : n38922;
  assign n38924 = pi15 ? n26269 : n38923;
  assign n38925 = pi21 ? n1009 : ~n242;
  assign n38926 = pi20 ? n32 : n38925;
  assign n38927 = pi19 ? n32 : n38926;
  assign n38928 = pi18 ? n32 : n38927;
  assign n38929 = pi17 ? n32 : n38928;
  assign n38930 = pi16 ? n32 : n38929;
  assign n38931 = pi14 ? n38924 : n38930;
  assign n38932 = pi21 ? n124 : n85;
  assign n38933 = pi20 ? n32 : n38932;
  assign n38934 = pi19 ? n32 : n38933;
  assign n38935 = pi18 ? n32 : n38934;
  assign n38936 = pi17 ? n32 : n38935;
  assign n38937 = pi16 ? n32 : n38936;
  assign n38938 = pi15 ? n38937 : n17111;
  assign n38939 = pi14 ? n38937 : n38938;
  assign n38940 = pi13 ? n38931 : n38939;
  assign n38941 = pi12 ? n38918 : n38940;
  assign n38942 = pi14 ? n17412 : n26163;
  assign n38943 = pi13 ? n16984 : n38942;
  assign n38944 = pi12 ? n38943 : n38865;
  assign n38945 = pi11 ? n38941 : n38944;
  assign n38946 = pi17 ? n1814 : ~n2512;
  assign n38947 = pi16 ? n32 : n38946;
  assign n38948 = pi15 ? n14147 : n38947;
  assign n38949 = pi17 ? n1814 : ~n38885;
  assign n38950 = pi16 ? n32 : n38949;
  assign n38951 = pi17 ? n1807 : ~n38888;
  assign n38952 = pi16 ? n32 : n38951;
  assign n38953 = pi15 ? n38950 : n38952;
  assign n38954 = pi14 ? n38948 : n38953;
  assign n38955 = pi17 ? n2537 : ~n38897;
  assign n38956 = pi16 ? n32 : n38955;
  assign n38957 = pi17 ? n2537 : ~n2519;
  assign n38958 = pi16 ? n32 : n38957;
  assign n38959 = pi15 ? n38956 : n38958;
  assign n38960 = pi14 ? n38959 : n38958;
  assign n38961 = pi13 ? n38954 : n38960;
  assign n38962 = pi12 ? n38881 : n38961;
  assign n38963 = pi11 ? n38875 : n38962;
  assign n38964 = pi10 ? n38945 : n38963;
  assign n38965 = pi09 ? n32 : n38964;
  assign n38966 = pi08 ? n38910 : n38965;
  assign n38967 = pi15 ? n32 : n26951;
  assign n38968 = pi14 ? n32 : n38967;
  assign n38969 = pi13 ? n32 : n38968;
  assign n38970 = pi12 ? n32 : n38969;
  assign n38971 = pi11 ? n32 : n38970;
  assign n38972 = pi10 ? n32 : n38971;
  assign n38973 = pi15 ? n38913 : n26462;
  assign n38974 = pi14 ? n38913 : n38973;
  assign n38975 = pi14 ? n17465 : n38491;
  assign n38976 = pi13 ? n38974 : n38975;
  assign n38977 = pi14 ? n17531 : n38814;
  assign n38978 = pi13 ? n26350 : n38977;
  assign n38979 = pi12 ? n38976 : n38978;
  assign n38980 = pi15 ? n16984 : n17198;
  assign n38981 = pi14 ? n16984 : n38980;
  assign n38982 = pi14 ? n17178 : n26163;
  assign n38983 = pi13 ? n38981 : n38982;
  assign n38984 = pi15 ? n17039 : n17061;
  assign n38985 = pi14 ? n17039 : n38984;
  assign n38986 = pi14 ? n17061 : n24799;
  assign n38987 = pi13 ? n38985 : n38986;
  assign n38988 = pi12 ? n38983 : n38987;
  assign n38989 = pi11 ? n38979 : n38988;
  assign n38990 = pi13 ? n37913 : n38869;
  assign n38991 = pi12 ? n38990 : n38874;
  assign n38992 = pi15 ? n23484 : n32;
  assign n38993 = pi14 ? n38992 : n24914;
  assign n38994 = pi13 ? n38993 : n38880;
  assign n38995 = pi17 ? n35983 : ~n2512;
  assign n38996 = pi16 ? n32 : n38995;
  assign n38997 = pi15 ? n14147 : n38996;
  assign n38998 = pi20 ? n428 : n18173;
  assign n38999 = pi19 ? n38998 : ~n1508;
  assign n39000 = pi18 ? n32 : n38999;
  assign n39001 = pi20 ? n266 : n274;
  assign n39002 = pi19 ? n39001 : n23644;
  assign n39003 = pi18 ? n39002 : n22307;
  assign n39004 = pi17 ? n39000 : ~n39003;
  assign n39005 = pi16 ? n32 : n39004;
  assign n39006 = pi20 ? n101 : n339;
  assign n39007 = pi19 ? n39006 : ~n32;
  assign n39008 = pi18 ? n32 : n39007;
  assign n39009 = pi17 ? n39008 : ~n38888;
  assign n39010 = pi16 ? n32 : n39009;
  assign n39011 = pi15 ? n39005 : n39010;
  assign n39012 = pi14 ? n38997 : n39011;
  assign n39013 = pi17 ? n2299 : ~n38897;
  assign n39014 = pi16 ? n32 : n39013;
  assign n39015 = pi17 ? n2299 : ~n2519;
  assign n39016 = pi16 ? n32 : n39015;
  assign n39017 = pi15 ? n39014 : n39016;
  assign n39018 = pi17 ? n2299 : ~n2408;
  assign n39019 = pi16 ? n32 : n39018;
  assign n39020 = pi15 ? n39016 : n39019;
  assign n39021 = pi14 ? n39017 : n39020;
  assign n39022 = pi13 ? n39012 : n39021;
  assign n39023 = pi12 ? n38994 : n39022;
  assign n39024 = pi11 ? n38991 : n39023;
  assign n39025 = pi10 ? n38989 : n39024;
  assign n39026 = pi09 ? n38972 : n39025;
  assign n39027 = pi21 ? n259 : n51;
  assign n39028 = pi20 ? n32 : n39027;
  assign n39029 = pi19 ? n32 : n39028;
  assign n39030 = pi18 ? n32 : n39029;
  assign n39031 = pi17 ? n32 : n39030;
  assign n39032 = pi16 ? n32 : n39031;
  assign n39033 = pi15 ? n39032 : n32;
  assign n39034 = pi14 ? n17618 : n39033;
  assign n39035 = pi13 ? n38974 : n39034;
  assign n39036 = pi12 ? n39035 : n32;
  assign n39037 = pi15 ? n17188 : n17198;
  assign n39038 = pi14 ? n17188 : n39037;
  assign n39039 = pi13 ? n39038 : n38982;
  assign n39040 = pi12 ? n39039 : n38987;
  assign n39041 = pi11 ? n39036 : n39040;
  assign n39042 = pi15 ? n15847 : n16452;
  assign n39043 = pi14 ? n39042 : n38635;
  assign n39044 = pi13 ? n37913 : n39043;
  assign n39045 = pi15 ? n16452 : n16298;
  assign n39046 = pi14 ? n39045 : n38871;
  assign n39047 = pi13 ? n39046 : n38873;
  assign n39048 = pi12 ? n39044 : n39047;
  assign n39049 = pi17 ? n2425 : ~n2512;
  assign n39050 = pi16 ? n32 : n39049;
  assign n39051 = pi15 ? n14147 : n39050;
  assign n39052 = pi19 ? n786 : ~n38571;
  assign n39053 = pi18 ? n32 : n39052;
  assign n39054 = pi20 ? n266 : n7839;
  assign n39055 = pi19 ? n266 : n39054;
  assign n39056 = pi18 ? n39055 : n22307;
  assign n39057 = pi17 ? n39053 : ~n39056;
  assign n39058 = pi16 ? n32 : n39057;
  assign n39059 = pi17 ? n2425 : ~n38888;
  assign n39060 = pi16 ? n32 : n39059;
  assign n39061 = pi15 ? n39058 : n39060;
  assign n39062 = pi14 ? n39051 : n39061;
  assign n39063 = pi17 ? n2425 : ~n38897;
  assign n39064 = pi16 ? n32 : n39063;
  assign n39065 = pi17 ? n2119 : ~n2519;
  assign n39066 = pi16 ? n32 : n39065;
  assign n39067 = pi15 ? n39064 : n39066;
  assign n39068 = pi17 ? n2408 : ~n2408;
  assign n39069 = pi16 ? n32 : n39068;
  assign n39070 = pi15 ? n39066 : n39069;
  assign n39071 = pi14 ? n39067 : n39070;
  assign n39072 = pi13 ? n39062 : n39071;
  assign n39073 = pi12 ? n38994 : n39072;
  assign n39074 = pi11 ? n39048 : n39073;
  assign n39075 = pi10 ? n39041 : n39074;
  assign n39076 = pi09 ? n38972 : n39075;
  assign n39077 = pi08 ? n39026 : n39076;
  assign n39078 = pi07 ? n38966 : n39077;
  assign n39079 = pi06 ? n38844 : n39078;
  assign n39080 = pi15 ? n17487 : n32;
  assign n39081 = pi14 ? n17487 : n39080;
  assign n39082 = pi13 ? n39081 : n32;
  assign n39083 = pi15 ? n17278 : n17111;
  assign n39084 = pi14 ? n17278 : n39083;
  assign n39085 = pi13 ? n17278 : n39084;
  assign n39086 = pi12 ? n39082 : n39085;
  assign n39087 = pi15 ? n17188 : n17286;
  assign n39088 = pi14 ? n17188 : n39087;
  assign n39089 = pi14 ? n16850 : n26163;
  assign n39090 = pi13 ? n39088 : n39089;
  assign n39091 = pi15 ? n26322 : n17061;
  assign n39092 = pi14 ? n17039 : n39091;
  assign n39093 = pi13 ? n39092 : n38986;
  assign n39094 = pi12 ? n39090 : n39093;
  assign n39095 = pi11 ? n39086 : n39094;
  assign n39096 = pi14 ? n38060 : n15847;
  assign n39097 = pi14 ? n32 : n38635;
  assign n39098 = pi13 ? n39096 : n39097;
  assign n39099 = pi15 ? n15230 : n16101;
  assign n39100 = pi14 ? n39099 : n38871;
  assign n39101 = pi14 ? n24247 : n38876;
  assign n39102 = pi13 ? n39100 : n39101;
  assign n39103 = pi12 ? n39098 : n39102;
  assign n39104 = pi15 ? n23484 : n22817;
  assign n39105 = pi14 ? n39104 : n22817;
  assign n39106 = pi15 ? n22817 : n14580;
  assign n39107 = pi15 ? n23443 : n35939;
  assign n39108 = pi14 ? n39106 : n39107;
  assign n39109 = pi13 ? n39105 : n39108;
  assign n39110 = pi19 ? n32 : n34188;
  assign n39111 = pi18 ? n39110 : n24548;
  assign n39112 = pi17 ? n2292 : ~n39111;
  assign n39113 = pi16 ? n32 : n39112;
  assign n39114 = pi15 ? n14147 : n39113;
  assign n39115 = pi17 ? n35572 : ~n2512;
  assign n39116 = pi16 ? n32 : n39115;
  assign n39117 = pi15 ? n14147 : n39116;
  assign n39118 = pi14 ? n39114 : n39117;
  assign n39119 = pi17 ? n35572 : ~n2519;
  assign n39120 = pi16 ? n32 : n39119;
  assign n39121 = pi17 ? n2748 : ~n2119;
  assign n39122 = pi16 ? n32 : n39121;
  assign n39123 = pi15 ? n39120 : n39122;
  assign n39124 = pi17 ? n2517 : ~n2119;
  assign n39125 = pi16 ? n32 : n39124;
  assign n39126 = pi14 ? n39123 : n39125;
  assign n39127 = pi13 ? n39118 : n39126;
  assign n39128 = pi12 ? n39109 : n39127;
  assign n39129 = pi11 ? n39103 : n39128;
  assign n39130 = pi10 ? n39095 : n39129;
  assign n39131 = pi09 ? n32 : n39130;
  assign n39132 = pi14 ? n17487 : n32;
  assign n39133 = pi13 ? n39132 : n32;
  assign n39134 = pi14 ? n17278 : n17279;
  assign n39135 = pi13 ? n17278 : n39134;
  assign n39136 = pi12 ? n39133 : n39135;
  assign n39137 = pi11 ? n39136 : n39094;
  assign n39138 = pi17 ? n2512 : ~n39111;
  assign n39139 = pi16 ? n32 : n39138;
  assign n39140 = pi15 ? n14147 : n39139;
  assign n39141 = pi15 ? n14147 : n8493;
  assign n39142 = pi14 ? n39140 : n39141;
  assign n39143 = pi17 ? n4099 : ~n2408;
  assign n39144 = pi16 ? n32 : n39143;
  assign n39145 = pi17 ? n4099 : ~n2119;
  assign n39146 = pi16 ? n32 : n39145;
  assign n39147 = pi15 ? n39144 : n39146;
  assign n39148 = pi14 ? n39147 : n39146;
  assign n39149 = pi13 ? n39142 : n39148;
  assign n39150 = pi12 ? n39109 : n39149;
  assign n39151 = pi11 ? n39103 : n39150;
  assign n39152 = pi10 ? n39137 : n39151;
  assign n39153 = pi09 ? n32 : n39152;
  assign n39154 = pi08 ? n39131 : n39153;
  assign n39155 = pi15 ? n17278 : n17367;
  assign n39156 = pi14 ? n17278 : n39155;
  assign n39157 = pi13 ? n17465 : n39156;
  assign n39158 = pi12 ? n32 : n39157;
  assign n39159 = pi14 ? n16850 : n17039;
  assign n39160 = pi13 ? n39088 : n39159;
  assign n39161 = pi14 ? n16804 : n16837;
  assign n39162 = pi13 ? n39092 : n39161;
  assign n39163 = pi12 ? n39160 : n39162;
  assign n39164 = pi11 ? n39158 : n39163;
  assign n39165 = pi15 ? n15230 : n16298;
  assign n39166 = pi14 ? n39165 : n38871;
  assign n39167 = pi13 ? n39166 : n39101;
  assign n39168 = pi12 ? n39098 : n39167;
  assign n39169 = pi15 ? n26623 : n22540;
  assign n39170 = pi14 ? n39169 : n22817;
  assign n39171 = pi15 ? n22817 : n22825;
  assign n39172 = pi15 ? n23443 : n14147;
  assign n39173 = pi14 ? n39171 : n39172;
  assign n39174 = pi13 ? n39170 : n39173;
  assign n39175 = pi21 ? n7659 : n313;
  assign n39176 = pi20 ? n39175 : ~n915;
  assign n39177 = pi19 ? n32 : n39176;
  assign n39178 = pi18 ? n32 : n39177;
  assign n39179 = pi20 ? n310 : n246;
  assign n39180 = pi19 ? n28957 : ~n39179;
  assign n39181 = pi20 ? n1076 : n342;
  assign n39182 = pi19 ? n39181 : ~n32;
  assign n39183 = pi18 ? n39180 : n39182;
  assign n39184 = pi17 ? n39178 : ~n39183;
  assign n39185 = pi16 ? n32 : n39184;
  assign n39186 = pi15 ? n14147 : n39185;
  assign n39187 = pi15 ? n14147 : n8703;
  assign n39188 = pi14 ? n39186 : n39187;
  assign n39189 = pi17 ? n2616 : ~n2517;
  assign n39190 = pi16 ? n32 : n39189;
  assign n39191 = pi17 ? n2736 : ~n2119;
  assign n39192 = pi16 ? n32 : n39191;
  assign n39193 = pi15 ? n39190 : n39192;
  assign n39194 = pi17 ? n2724 : ~n2119;
  assign n39195 = pi16 ? n32 : n39194;
  assign n39196 = pi15 ? n39192 : n39195;
  assign n39197 = pi14 ? n39193 : n39196;
  assign n39198 = pi13 ? n39188 : n39197;
  assign n39199 = pi12 ? n39174 : n39198;
  assign n39200 = pi11 ? n39168 : n39199;
  assign n39201 = pi10 ? n39164 : n39200;
  assign n39202 = pi09 ? n32 : n39201;
  assign n39203 = pi14 ? n39169 : n22931;
  assign n39204 = pi13 ? n39203 : n39173;
  assign n39205 = pi18 ? n32 : n11923;
  assign n39206 = pi20 ? n321 : n206;
  assign n39207 = pi19 ? n39206 : n39179;
  assign n39208 = pi18 ? n39207 : ~n39182;
  assign n39209 = pi17 ? n39205 : n39208;
  assign n39210 = pi16 ? n32 : n39209;
  assign n39211 = pi15 ? n14147 : n39210;
  assign n39212 = pi17 ? n3067 : ~n2517;
  assign n39213 = pi16 ? n32 : n39212;
  assign n39214 = pi15 ? n14147 : n39213;
  assign n39215 = pi14 ? n39211 : n39214;
  assign n39216 = pi17 ? n2836 : ~n2119;
  assign n39217 = pi16 ? n32 : n39216;
  assign n39218 = pi15 ? n39213 : n39217;
  assign n39219 = pi14 ? n39218 : n39217;
  assign n39220 = pi13 ? n39215 : n39219;
  assign n39221 = pi12 ? n39204 : n39220;
  assign n39222 = pi11 ? n39168 : n39221;
  assign n39223 = pi10 ? n39164 : n39222;
  assign n39224 = pi09 ? n32 : n39223;
  assign n39225 = pi08 ? n39202 : n39224;
  assign n39226 = pi07 ? n39154 : n39225;
  assign n39227 = pi13 ? n32 : n39084;
  assign n39228 = pi12 ? n32 : n39227;
  assign n39229 = pi15 ? n17188 : n16850;
  assign n39230 = pi14 ? n17188 : n39229;
  assign n39231 = pi13 ? n39230 : n39159;
  assign n39232 = pi14 ? n17039 : n17061;
  assign n39233 = pi14 ? n26250 : n16837;
  assign n39234 = pi13 ? n39232 : n39233;
  assign n39235 = pi12 ? n39231 : n39234;
  assign n39236 = pi11 ? n39228 : n39235;
  assign n39237 = pi14 ? n16393 : n16452;
  assign n39238 = pi14 ? n16452 : n39045;
  assign n39239 = pi13 ? n39237 : n39238;
  assign n39240 = pi19 ? n322 : n3692;
  assign n39241 = pi18 ? n32 : n39240;
  assign n39242 = pi17 ? n32 : n39241;
  assign n39243 = pi16 ? n32 : n39242;
  assign n39244 = pi19 ? n322 : n9724;
  assign n39245 = pi18 ? n32 : n39244;
  assign n39246 = pi17 ? n32 : n39245;
  assign n39247 = pi16 ? n32 : n39246;
  assign n39248 = pi15 ? n39243 : n39247;
  assign n39249 = pi15 ? n24582 : n15244;
  assign n39250 = pi14 ? n39248 : n39249;
  assign n39251 = pi15 ? n15244 : n25657;
  assign n39252 = pi15 ? n23933 : n25657;
  assign n39253 = pi14 ? n39251 : n39252;
  assign n39254 = pi13 ? n39250 : n39253;
  assign n39255 = pi12 ? n39239 : n39254;
  assign n39256 = pi15 ? n24742 : n23447;
  assign n39257 = pi14 ? n39256 : n24914;
  assign n39258 = pi15 ? n14389 : n14147;
  assign n39259 = pi14 ? n38261 : n39258;
  assign n39260 = pi13 ? n39257 : n39259;
  assign n39261 = pi15 ? n14147 : n14152;
  assign n39262 = pi19 ? n6339 : n18678;
  assign n39263 = pi19 ? n34416 : ~n32;
  assign n39264 = pi18 ? n39262 : ~n39263;
  assign n39265 = pi17 ? n32 : n39264;
  assign n39266 = pi16 ? n32 : n39265;
  assign n39267 = pi17 ? n2963 : ~n2408;
  assign n39268 = pi16 ? n32 : n39267;
  assign n39269 = pi15 ? n39266 : n39268;
  assign n39270 = pi14 ? n39261 : n39269;
  assign n39271 = pi17 ? n2963 : ~n2292;
  assign n39272 = pi16 ? n32 : n39271;
  assign n39273 = pi17 ? n2726 : ~n2292;
  assign n39274 = pi16 ? n32 : n39273;
  assign n39275 = pi15 ? n39272 : n39274;
  assign n39276 = pi17 ? n2726 : ~n2531;
  assign n39277 = pi16 ? n32 : n39276;
  assign n39278 = pi17 ? n2963 : ~n2119;
  assign n39279 = pi16 ? n32 : n39278;
  assign n39280 = pi15 ? n39277 : n39279;
  assign n39281 = pi14 ? n39275 : n39280;
  assign n39282 = pi13 ? n39270 : n39281;
  assign n39283 = pi12 ? n39260 : n39282;
  assign n39284 = pi11 ? n39255 : n39283;
  assign n39285 = pi10 ? n39236 : n39284;
  assign n39286 = pi09 ? n32 : n39285;
  assign n39287 = pi13 ? n32 : n39134;
  assign n39288 = pi12 ? n32 : n39287;
  assign n39289 = pi11 ? n39288 : n39235;
  assign n39290 = pi14 ? n16452 : n16299;
  assign n39291 = pi13 ? n39237 : n39290;
  assign n39292 = pi12 ? n39291 : n39254;
  assign n39293 = pi17 ? n2959 : ~n2408;
  assign n39294 = pi16 ? n32 : n39293;
  assign n39295 = pi15 ? n39266 : n39294;
  assign n39296 = pi14 ? n39261 : n39295;
  assign n39297 = pi15 ? n9435 : n39294;
  assign n39298 = pi17 ? n3046 : ~n2531;
  assign n39299 = pi16 ? n32 : n39298;
  assign n39300 = pi17 ? n2959 : ~n2119;
  assign n39301 = pi16 ? n32 : n39300;
  assign n39302 = pi15 ? n39299 : n39301;
  assign n39303 = pi14 ? n39297 : n39302;
  assign n39304 = pi13 ? n39296 : n39303;
  assign n39305 = pi12 ? n39260 : n39304;
  assign n39306 = pi11 ? n39292 : n39305;
  assign n39307 = pi10 ? n39289 : n39306;
  assign n39308 = pi09 ? n32 : n39307;
  assign n39309 = pi08 ? n39286 : n39308;
  assign n39310 = pi14 ? n16852 : n17039;
  assign n39311 = pi13 ? n39230 : n39310;
  assign n39312 = pi13 ? n39232 : n16837;
  assign n39313 = pi12 ? n39311 : n39312;
  assign n39314 = pi11 ? n39288 : n39313;
  assign n39315 = pi14 ? n39247 : n39249;
  assign n39316 = pi19 ? n519 : ~n813;
  assign n39317 = pi18 ? n32 : n39316;
  assign n39318 = pi17 ? n32 : n39317;
  assign n39319 = pi16 ? n32 : n39318;
  assign n39320 = pi15 ? n39319 : n24742;
  assign n39321 = pi14 ? n25657 : n39320;
  assign n39322 = pi13 ? n39315 : n39321;
  assign n39323 = pi12 ? n39291 : n39322;
  assign n39324 = pi15 ? n24742 : n15263;
  assign n39325 = pi15 ? n14967 : n22437;
  assign n39326 = pi14 ? n39324 : n39325;
  assign n39327 = pi15 ? n14593 : n14143;
  assign n39328 = pi14 ? n27435 : n39327;
  assign n39329 = pi13 ? n39326 : n39328;
  assign n39330 = pi20 ? n10644 : ~n32;
  assign n39331 = pi19 ? n9007 : ~n39330;
  assign n39332 = pi18 ? n39331 : n23543;
  assign n39333 = pi17 ? n32 : ~n39332;
  assign n39334 = pi16 ? n32 : n39333;
  assign n39335 = pi17 ? n30283 : ~n2519;
  assign n39336 = pi16 ? n32 : n39335;
  assign n39337 = pi15 ? n39334 : n39336;
  assign n39338 = pi14 ? n39261 : n39337;
  assign n39339 = pi17 ? n3728 : ~n2119;
  assign n39340 = pi16 ? n32 : n39339;
  assign n39341 = pi17 ? n2954 : ~n2531;
  assign n39342 = pi16 ? n32 : n39341;
  assign n39343 = pi17 ? n3728 : ~n2653;
  assign n39344 = pi16 ? n32 : n39343;
  assign n39345 = pi15 ? n39342 : n39344;
  assign n39346 = pi14 ? n39340 : n39345;
  assign n39347 = pi13 ? n39338 : n39346;
  assign n39348 = pi12 ? n39329 : n39347;
  assign n39349 = pi11 ? n39323 : n39348;
  assign n39350 = pi10 ? n39314 : n39349;
  assign n39351 = pi09 ? n32 : n39350;
  assign n39352 = pi18 ? n32 : n6108;
  assign n39353 = pi17 ? n32 : n39352;
  assign n39354 = pi16 ? n32 : n39353;
  assign n39355 = pi15 ? n39354 : n24742;
  assign n39356 = pi14 ? n25657 : n39355;
  assign n39357 = pi13 ? n39315 : n39356;
  assign n39358 = pi12 ? n39291 : n39357;
  assign n39359 = pi15 ? n22437 : n14593;
  assign n39360 = pi15 ? n14593 : n24543;
  assign n39361 = pi14 ? n39359 : n39360;
  assign n39362 = pi13 ? n39326 : n39361;
  assign n39363 = pi17 ? n3569 : ~n39332;
  assign n39364 = pi16 ? n32 : n39363;
  assign n39365 = pi17 ? n3569 : ~n2519;
  assign n39366 = pi16 ? n32 : n39365;
  assign n39367 = pi15 ? n39364 : n39366;
  assign n39368 = pi14 ? n39261 : n39367;
  assign n39369 = pi17 ? n32 : ~n2119;
  assign n39370 = pi16 ? n32 : n39369;
  assign n39371 = pi17 ? n32 : ~n2531;
  assign n39372 = pi16 ? n32 : n39371;
  assign n39373 = pi17 ? n32 : ~n2653;
  assign n39374 = pi16 ? n32 : n39373;
  assign n39375 = pi15 ? n39372 : n39374;
  assign n39376 = pi14 ? n39370 : n39375;
  assign n39377 = pi13 ? n39368 : n39376;
  assign n39378 = pi12 ? n39362 : n39377;
  assign n39379 = pi11 ? n39358 : n39378;
  assign n39380 = pi10 ? n39314 : n39379;
  assign n39381 = pi09 ? n32 : n39380;
  assign n39382 = pi08 ? n39351 : n39381;
  assign n39383 = pi07 ? n39309 : n39382;
  assign n39384 = pi06 ? n39226 : n39383;
  assign n39385 = pi05 ? n39079 : n39384;
  assign n39386 = pi14 ? n25377 : n17039;
  assign n39387 = pi13 ? n39230 : n39386;
  assign n39388 = pi15 ? n17039 : n26322;
  assign n39389 = pi14 ? n39388 : n38628;
  assign n39390 = pi13 ? n39389 : n16837;
  assign n39391 = pi12 ? n39387 : n39390;
  assign n39392 = pi11 ? n39288 : n39391;
  assign n39393 = pi14 ? n39042 : n16452;
  assign n39394 = pi15 ? n16293 : n16105;
  assign n39395 = pi14 ? n39045 : n39394;
  assign n39396 = pi13 ? n39393 : n39395;
  assign n39397 = pi15 ? n14917 : n15244;
  assign n39398 = pi14 ? n24504 : n39397;
  assign n39399 = pi13 ? n39398 : n24742;
  assign n39400 = pi12 ? n39396 : n39399;
  assign n39401 = pi19 ? n1818 : ~n2614;
  assign n39402 = pi18 ? n32 : n39401;
  assign n39403 = pi17 ? n32 : n39402;
  assign n39404 = pi16 ? n32 : n39403;
  assign n39405 = pi15 ? n24742 : n39404;
  assign n39406 = pi15 ? n26663 : n22437;
  assign n39407 = pi14 ? n39405 : n39406;
  assign n39408 = pi15 ? n22434 : n24543;
  assign n39409 = pi15 ? n24543 : n13913;
  assign n39410 = pi14 ? n39408 : n39409;
  assign n39411 = pi13 ? n39407 : n39410;
  assign n39412 = pi15 ? n14152 : n32685;
  assign n39413 = pi18 ? n289 : ~n323;
  assign n39414 = pi17 ? n32 : n39413;
  assign n39415 = pi16 ? n32 : n39414;
  assign n39416 = pi15 ? n10247 : n39415;
  assign n39417 = pi14 ? n39412 : n39416;
  assign n39418 = pi18 ? n237 : ~n532;
  assign n39419 = pi17 ? n32 : n39418;
  assign n39420 = pi16 ? n32 : n39419;
  assign n39421 = pi18 ? n1813 : ~n532;
  assign n39422 = pi17 ? n32 : n39421;
  assign n39423 = pi16 ? n32 : n39422;
  assign n39424 = pi15 ? n39420 : n39423;
  assign n39425 = pi14 ? n39424 : n39423;
  assign n39426 = pi13 ? n39417 : n39425;
  assign n39427 = pi12 ? n39411 : n39426;
  assign n39428 = pi11 ? n39400 : n39427;
  assign n39429 = pi10 ? n39392 : n39428;
  assign n39430 = pi09 ? n32 : n39429;
  assign n39431 = pi14 ? n17273 : n39229;
  assign n39432 = pi13 ? n39431 : n39386;
  assign n39433 = pi12 ? n39432 : n39390;
  assign n39434 = pi11 ? n39288 : n39433;
  assign n39435 = pi15 ? n24742 : n23169;
  assign n39436 = pi15 ? n23443 : n22437;
  assign n39437 = pi14 ? n39435 : n39436;
  assign n39438 = pi13 ? n39437 : n39410;
  assign n39439 = pi15 ? n14156 : n32685;
  assign n39440 = pi18 ? n350 : ~n323;
  assign n39441 = pi17 ? n32 : n39440;
  assign n39442 = pi16 ? n32 : n39441;
  assign n39443 = pi18 ? n2318 : ~n323;
  assign n39444 = pi17 ? n32 : n39443;
  assign n39445 = pi16 ? n32 : n39444;
  assign n39446 = pi15 ? n39442 : n39445;
  assign n39447 = pi14 ? n39439 : n39446;
  assign n39448 = pi17 ? n32 : n32624;
  assign n39449 = pi16 ? n32 : n39448;
  assign n39450 = pi18 ? n2318 : ~n532;
  assign n39451 = pi17 ? n32 : n39450;
  assign n39452 = pi16 ? n32 : n39451;
  assign n39453 = pi15 ? n39449 : n39452;
  assign n39454 = pi14 ? n39449 : n39453;
  assign n39455 = pi13 ? n39447 : n39454;
  assign n39456 = pi12 ? n39438 : n39455;
  assign n39457 = pi11 ? n39400 : n39456;
  assign n39458 = pi10 ? n39434 : n39457;
  assign n39459 = pi09 ? n32 : n39458;
  assign n39460 = pi08 ? n39430 : n39459;
  assign n39461 = pi15 ? n17061 : n32;
  assign n39462 = pi14 ? n39388 : n39461;
  assign n39463 = pi15 ? n16837 : n16392;
  assign n39464 = pi14 ? n16837 : n39463;
  assign n39465 = pi13 ? n39462 : n39464;
  assign n39466 = pi12 ? n39432 : n39465;
  assign n39467 = pi11 ? n39288 : n39466;
  assign n39468 = pi15 ? n16204 : n16105;
  assign n39469 = pi14 ? n16298 : n39468;
  assign n39470 = pi13 ? n39393 : n39469;
  assign n39471 = pi19 ? n32 : ~n11590;
  assign n39472 = pi18 ? n32 : n39471;
  assign n39473 = pi17 ? n32 : n39472;
  assign n39474 = pi16 ? n32 : n39473;
  assign n39475 = pi15 ? n15700 : n39474;
  assign n39476 = pi15 ? n14917 : n24838;
  assign n39477 = pi14 ? n39475 : n39476;
  assign n39478 = pi14 ? n24838 : n24742;
  assign n39479 = pi13 ? n39477 : n39478;
  assign n39480 = pi12 ? n39470 : n39479;
  assign n39481 = pi15 ? n23443 : n21853;
  assign n39482 = pi15 ? n21853 : n14967;
  assign n39483 = pi14 ? n39481 : n39482;
  assign n39484 = pi19 ? n6727 : n32;
  assign n39485 = pi18 ? n32 : n39484;
  assign n39486 = pi17 ? n32 : n39485;
  assign n39487 = pi16 ? n32 : n39486;
  assign n39488 = pi15 ? n39487 : n24543;
  assign n39489 = pi14 ? n39488 : n39439;
  assign n39490 = pi13 ? n39483 : n39489;
  assign n39491 = pi18 ? n39007 : ~n323;
  assign n39492 = pi17 ? n32 : n39491;
  assign n39493 = pi16 ? n32 : n39492;
  assign n39494 = pi18 ? n532 : ~n22159;
  assign n39495 = pi17 ? n32 : n39494;
  assign n39496 = pi16 ? n32 : n39495;
  assign n39497 = pi15 ? n39493 : n39496;
  assign n39498 = pi14 ? n39439 : n39497;
  assign n39499 = pi18 ? n532 : ~n418;
  assign n39500 = pi17 ? n32 : n39499;
  assign n39501 = pi16 ? n32 : n39500;
  assign n39502 = pi15 ? n32709 : n39501;
  assign n39503 = pi14 ? n32709 : n39502;
  assign n39504 = pi13 ? n39498 : n39503;
  assign n39505 = pi12 ? n39490 : n39504;
  assign n39506 = pi11 ? n39480 : n39505;
  assign n39507 = pi10 ? n39467 : n39506;
  assign n39508 = pi09 ? n32 : n39507;
  assign n39509 = pi13 ? n17239 : n39386;
  assign n39510 = pi12 ? n39509 : n39465;
  assign n39511 = pi11 ? n39288 : n39510;
  assign n39512 = pi15 ? n16298 : n16204;
  assign n39513 = pi15 ? n16204 : n15700;
  assign n39514 = pi14 ? n39512 : n39513;
  assign n39515 = pi13 ? n39393 : n39514;
  assign n39516 = pi15 ? n23569 : n24097;
  assign n39517 = pi19 ? n322 : ~n2848;
  assign n39518 = pi18 ? n32 : n39517;
  assign n39519 = pi17 ? n32 : n39518;
  assign n39520 = pi16 ? n32 : n39519;
  assign n39521 = pi15 ? n39520 : n25657;
  assign n39522 = pi14 ? n39516 : n39521;
  assign n39523 = pi13 ? n39522 : n24742;
  assign n39524 = pi12 ? n39515 : n39523;
  assign n39525 = pi20 ? n32 : ~n2180;
  assign n39526 = pi19 ? n39525 : n32;
  assign n39527 = pi18 ? n32 : n39526;
  assign n39528 = pi17 ? n32 : n39527;
  assign n39529 = pi16 ? n32 : n39528;
  assign n39530 = pi15 ? n39529 : n14147;
  assign n39531 = pi14 ? n39530 : n39439;
  assign n39532 = pi13 ? n39483 : n39531;
  assign n39533 = pi18 ? n605 : ~n22159;
  assign n39534 = pi17 ? n32 : n39533;
  assign n39535 = pi16 ? n32 : n39534;
  assign n39536 = pi15 ? n10958 : n39535;
  assign n39537 = pi14 ? n39439 : n39536;
  assign n39538 = pi18 ? n605 : ~n532;
  assign n39539 = pi17 ? n32 : n39538;
  assign n39540 = pi16 ? n32 : n39539;
  assign n39541 = pi18 ? n2291 : ~n418;
  assign n39542 = pi17 ? n32 : n39541;
  assign n39543 = pi16 ? n32 : n39542;
  assign n39544 = pi15 ? n39540 : n39543;
  assign n39545 = pi14 ? n39540 : n39544;
  assign n39546 = pi13 ? n39537 : n39545;
  assign n39547 = pi12 ? n39532 : n39546;
  assign n39548 = pi11 ? n39524 : n39547;
  assign n39549 = pi10 ? n39511 : n39548;
  assign n39550 = pi09 ? n32 : n39549;
  assign n39551 = pi08 ? n39508 : n39550;
  assign n39552 = pi07 ? n39460 : n39551;
  assign n39553 = pi15 ? n17286 : n16850;
  assign n39554 = pi14 ? n32 : n39553;
  assign n39555 = pi13 ? n39554 : n39386;
  assign n39556 = pi15 ? n17056 : n26322;
  assign n39557 = pi14 ? n39556 : n39461;
  assign n39558 = pi15 ? n25814 : n16546;
  assign n39559 = pi14 ? n16837 : n39558;
  assign n39560 = pi13 ? n39557 : n39559;
  assign n39561 = pi12 ? n39555 : n39560;
  assign n39562 = pi11 ? n39288 : n39561;
  assign n39563 = pi15 ? n16606 : n16452;
  assign n39564 = pi14 ? n38634 : n39563;
  assign n39565 = pi20 ? n27235 : n32;
  assign n39566 = pi19 ? n32 : n39565;
  assign n39567 = pi18 ? n32 : n39566;
  assign n39568 = pi17 ? n32 : n39567;
  assign n39569 = pi16 ? n32 : n39568;
  assign n39570 = pi15 ? n39569 : n15700;
  assign n39571 = pi14 ? n39570 : n15700;
  assign n39572 = pi13 ? n39564 : n39571;
  assign n39573 = pi15 ? n26837 : n24511;
  assign n39574 = pi14 ? n39573 : n24659;
  assign n39575 = pi15 ? n25466 : n27229;
  assign n39576 = pi14 ? n24659 : n39575;
  assign n39577 = pi13 ? n39574 : n39576;
  assign n39578 = pi12 ? n39572 : n39577;
  assign n39579 = pi19 ? n18865 : n32;
  assign n39580 = pi18 ? n32 : n39579;
  assign n39581 = pi17 ? n32 : n39580;
  assign n39582 = pi16 ? n32 : n39581;
  assign n39583 = pi15 ? n23443 : n39582;
  assign n39584 = pi15 ? n21928 : n39487;
  assign n39585 = pi14 ? n39583 : n39584;
  assign n39586 = pi21 ? n174 : n6898;
  assign n39587 = pi20 ? n321 : ~n39586;
  assign n39588 = pi19 ? n39587 : n32;
  assign n39589 = pi18 ? n32 : n39588;
  assign n39590 = pi17 ? n32 : n39589;
  assign n39591 = pi16 ? n32 : n39590;
  assign n39592 = pi15 ? n39591 : n13629;
  assign n39593 = pi17 ? n32 : n34131;
  assign n39594 = pi16 ? n32 : n39593;
  assign n39595 = pi14 ? n39592 : n39594;
  assign n39596 = pi13 ? n39585 : n39595;
  assign n39597 = pi20 ? n32 : ~n160;
  assign n39598 = pi19 ? n39597 : ~n32;
  assign n39599 = pi18 ? n323 : ~n39598;
  assign n39600 = pi17 ? n32 : n39599;
  assign n39601 = pi16 ? n32 : n39600;
  assign n39602 = pi18 ? n1326 : ~n22159;
  assign n39603 = pi17 ? n32 : n39602;
  assign n39604 = pi16 ? n32 : n39603;
  assign n39605 = pi15 ? n39601 : n39604;
  assign n39606 = pi14 ? n39594 : n39605;
  assign n39607 = pi18 ? n508 : ~n532;
  assign n39608 = pi17 ? n32 : n39607;
  assign n39609 = pi16 ? n32 : n39608;
  assign n39610 = pi15 ? n39609 : n33130;
  assign n39611 = pi18 ? n508 : ~n418;
  assign n39612 = pi17 ? n32 : n39611;
  assign n39613 = pi16 ? n32 : n39612;
  assign n39614 = pi15 ? n39609 : n39613;
  assign n39615 = pi14 ? n39610 : n39614;
  assign n39616 = pi13 ? n39606 : n39615;
  assign n39617 = pi12 ? n39596 : n39616;
  assign n39618 = pi11 ? n39578 : n39617;
  assign n39619 = pi10 ? n39562 : n39618;
  assign n39620 = pi09 ? n32 : n39619;
  assign n39621 = pi14 ? n17278 : n26537;
  assign n39622 = pi13 ? n32 : n39621;
  assign n39623 = pi12 ? n32 : n39622;
  assign n39624 = pi11 ? n39623 : n39561;
  assign n39625 = pi21 ? n1939 : ~n100;
  assign n39626 = pi20 ? n39625 : n32;
  assign n39627 = pi19 ? n32 : n39626;
  assign n39628 = pi18 ? n32 : n39627;
  assign n39629 = pi17 ? n32 : n39628;
  assign n39630 = pi16 ? n32 : n39629;
  assign n39631 = pi15 ? n39630 : n15700;
  assign n39632 = pi14 ? n39631 : n15700;
  assign n39633 = pi13 ? n39564 : n39632;
  assign n39634 = pi15 ? n25466 : n37644;
  assign n39635 = pi14 ? n24659 : n39634;
  assign n39636 = pi13 ? n39574 : n39635;
  assign n39637 = pi12 ? n39633 : n39636;
  assign n39638 = pi22 ? n50 : n84;
  assign n39639 = pi21 ? n206 : ~n39638;
  assign n39640 = pi20 ? n32 : ~n39639;
  assign n39641 = pi19 ? n39640 : n32;
  assign n39642 = pi18 ? n32 : n39641;
  assign n39643 = pi17 ? n32 : n39642;
  assign n39644 = pi16 ? n32 : n39643;
  assign n39645 = pi15 ? n21853 : n39644;
  assign n39646 = pi14 ? n39481 : n39645;
  assign n39647 = pi15 ? n39591 : n13626;
  assign n39648 = pi14 ? n39647 : n33939;
  assign n39649 = pi13 ? n39646 : n39648;
  assign n39650 = pi15 ? n33939 : n39594;
  assign n39651 = pi15 ? n39609 : n33135;
  assign n39652 = pi14 ? n39650 : n39651;
  assign n39653 = pi15 ? n33135 : n11429;
  assign n39654 = pi14 ? n33135 : n39653;
  assign n39655 = pi13 ? n39652 : n39654;
  assign n39656 = pi12 ? n39649 : n39655;
  assign n39657 = pi11 ? n39637 : n39656;
  assign n39658 = pi10 ? n39624 : n39657;
  assign n39659 = pi09 ? n32 : n39658;
  assign n39660 = pi08 ? n39620 : n39659;
  assign n39661 = pi13 ? n39554 : n17039;
  assign n39662 = pi15 ? n25814 : n16467;
  assign n39663 = pi14 ? n16837 : n39662;
  assign n39664 = pi13 ? n39557 : n39663;
  assign n39665 = pi12 ? n39661 : n39664;
  assign n39666 = pi11 ? n39623 : n39665;
  assign n39667 = pi19 ? n32 : n21369;
  assign n39668 = pi18 ? n32 : n39667;
  assign n39669 = pi17 ? n32 : n39668;
  assign n39670 = pi16 ? n32 : n39669;
  assign n39671 = pi15 ? n39670 : n24495;
  assign n39672 = pi15 ? n24495 : n25384;
  assign n39673 = pi14 ? n39671 : n39672;
  assign n39674 = pi15 ? n27304 : n15700;
  assign n39675 = pi14 ? n39674 : n26837;
  assign n39676 = pi13 ? n39673 : n39675;
  assign n39677 = pi18 ? n16834 : n21287;
  assign n39678 = pi17 ? n32 : n39677;
  assign n39679 = pi16 ? n32 : n39678;
  assign n39680 = pi15 ? n39679 : n24247;
  assign n39681 = pi14 ? n39680 : n24659;
  assign n39682 = pi13 ? n39681 : n39635;
  assign n39683 = pi12 ? n39676 : n39682;
  assign n39684 = pi20 ? n32 : ~n23668;
  assign n39685 = pi19 ? n39684 : n32;
  assign n39686 = pi18 ? n32 : n39685;
  assign n39687 = pi17 ? n32 : n39686;
  assign n39688 = pi16 ? n32 : n39687;
  assign n39689 = pi15 ? n14397 : n39688;
  assign n39690 = pi14 ? n39481 : n39689;
  assign n39691 = pi20 ? n321 : ~n7108;
  assign n39692 = pi19 ? n39691 : n32;
  assign n39693 = pi18 ? n32 : n39692;
  assign n39694 = pi17 ? n32 : n39693;
  assign n39695 = pi16 ? n32 : n39694;
  assign n39696 = pi20 ? n321 : ~n18610;
  assign n39697 = pi19 ? n39696 : n32;
  assign n39698 = pi18 ? n32 : n39697;
  assign n39699 = pi17 ? n32 : n39698;
  assign n39700 = pi16 ? n32 : n39699;
  assign n39701 = pi15 ? n39695 : n39700;
  assign n39702 = pi14 ? n39701 : n33939;
  assign n39703 = pi13 ? n39690 : n39702;
  assign n39704 = pi20 ? n321 : ~n7013;
  assign n39705 = pi19 ? n39704 : n32;
  assign n39706 = pi18 ? n32 : n39705;
  assign n39707 = pi17 ? n32 : n39706;
  assign n39708 = pi16 ? n32 : n39707;
  assign n39709 = pi15 ? n33939 : n39708;
  assign n39710 = pi14 ? n39709 : n33618;
  assign n39711 = pi18 ? n697 : ~n35365;
  assign n39712 = pi17 ? n32 : n39711;
  assign n39713 = pi16 ? n32 : n39712;
  assign n39714 = pi15 ? n11657 : n39713;
  assign n39715 = pi14 ? n33618 : n39714;
  assign n39716 = pi13 ? n39710 : n39715;
  assign n39717 = pi12 ? n39703 : n39716;
  assign n39718 = pi11 ? n39683 : n39717;
  assign n39719 = pi10 ? n39666 : n39718;
  assign n39720 = pi09 ? n32 : n39719;
  assign n39721 = pi12 ? n39661 : n39560;
  assign n39722 = pi11 ? n39623 : n39721;
  assign n39723 = pi15 ? n16601 : n25384;
  assign n39724 = pi14 ? n16601 : n39723;
  assign n39725 = pi15 ? n25211 : n15700;
  assign n39726 = pi14 ? n39725 : n26837;
  assign n39727 = pi13 ? n39724 : n39726;
  assign n39728 = pi19 ? n236 : ~n9724;
  assign n39729 = pi18 ? n16896 : ~n39728;
  assign n39730 = pi17 ? n32 : n39729;
  assign n39731 = pi16 ? n32 : n39730;
  assign n39732 = pi15 ? n39731 : n24247;
  assign n39733 = pi14 ? n39732 : n24659;
  assign n39734 = pi15 ? n14765 : n37644;
  assign n39735 = pi14 ? n36816 : n39734;
  assign n39736 = pi13 ? n39733 : n39735;
  assign n39737 = pi12 ? n39727 : n39736;
  assign n39738 = pi20 ? n321 : ~n1324;
  assign n39739 = pi19 ? n39738 : n32;
  assign n39740 = pi18 ? n32 : n39739;
  assign n39741 = pi17 ? n32 : n39740;
  assign n39742 = pi16 ? n32 : n39741;
  assign n39743 = pi15 ? n39742 : n23874;
  assign n39744 = pi14 ? n39743 : n33939;
  assign n39745 = pi13 ? n39690 : n39744;
  assign n39746 = pi14 ? n39709 : n33448;
  assign n39747 = pi15 ? n11863 : n20151;
  assign n39748 = pi14 ? n33448 : n39747;
  assign n39749 = pi13 ? n39746 : n39748;
  assign n39750 = pi12 ? n39745 : n39749;
  assign n39751 = pi11 ? n39737 : n39750;
  assign n39752 = pi10 ? n39722 : n39751;
  assign n39753 = pi09 ? n32 : n39752;
  assign n39754 = pi08 ? n39720 : n39753;
  assign n39755 = pi07 ? n39660 : n39754;
  assign n39756 = pi06 ? n39552 : n39755;
  assign n39757 = pi14 ? n17278 : n37565;
  assign n39758 = pi13 ? n32 : n39757;
  assign n39759 = pi12 ? n32 : n39758;
  assign n39760 = pi14 ? n32 : n16852;
  assign n39761 = pi13 ? n39760 : n17039;
  assign n39762 = pi15 ? n17056 : n38750;
  assign n39763 = pi14 ? n39762 : n32;
  assign n39764 = pi21 ? n32 : ~n11567;
  assign n39765 = pi20 ? n39764 : n32;
  assign n39766 = pi19 ? n32 : n39765;
  assign n39767 = pi18 ? n32 : n39766;
  assign n39768 = pi17 ? n32 : n39767;
  assign n39769 = pi16 ? n32 : n39768;
  assign n39770 = pi15 ? n16452 : n39769;
  assign n39771 = pi20 ? n321 : n481;
  assign n39772 = pi19 ? n32 : n39771;
  assign n39773 = pi18 ? n32 : n39772;
  assign n39774 = pi17 ? n32 : n39773;
  assign n39775 = pi16 ? n32 : n39774;
  assign n39776 = pi15 ? n39775 : n15847;
  assign n39777 = pi14 ? n39770 : n39776;
  assign n39778 = pi13 ? n39763 : n39777;
  assign n39779 = pi12 ? n39761 : n39778;
  assign n39780 = pi11 ? n39759 : n39779;
  assign n39781 = pi19 ? n32 : n20508;
  assign n39782 = pi18 ? n32 : n39781;
  assign n39783 = pi17 ? n32 : n39782;
  assign n39784 = pi16 ? n32 : n39783;
  assign n39785 = pi15 ? n25044 : n39784;
  assign n39786 = pi14 ? n16452 : n39785;
  assign n39787 = pi15 ? n15867 : n15700;
  assign n39788 = pi21 ? n51 : n259;
  assign n39789 = pi20 ? n39788 : ~n32;
  assign n39790 = pi19 ? n322 : ~n39789;
  assign n39791 = pi18 ? n32 : n39790;
  assign n39792 = pi17 ? n32 : n39791;
  assign n39793 = pi16 ? n32 : n39792;
  assign n39794 = pi15 ? n15700 : n39793;
  assign n39795 = pi14 ? n39787 : n39794;
  assign n39796 = pi13 ? n39786 : n39795;
  assign n39797 = pi15 ? n37501 : n14917;
  assign n39798 = pi15 ? n25466 : n24659;
  assign n39799 = pi14 ? n39797 : n39798;
  assign n39800 = pi19 ? n322 : ~n10447;
  assign n39801 = pi18 ? n32 : n39800;
  assign n39802 = pi17 ? n32 : n39801;
  assign n39803 = pi16 ? n32 : n39802;
  assign n39804 = pi15 ? n23443 : n39803;
  assign n39805 = pi19 ? n322 : n53;
  assign n39806 = pi18 ? n32 : n39805;
  assign n39807 = pi17 ? n32 : n39806;
  assign n39808 = pi16 ? n32 : n39807;
  assign n39809 = pi19 ? n1464 : n358;
  assign n39810 = pi18 ? n32 : n39809;
  assign n39811 = pi17 ? n32 : n39810;
  assign n39812 = pi16 ? n32 : n39811;
  assign n39813 = pi15 ? n39808 : n39812;
  assign n39814 = pi14 ? n39804 : n39813;
  assign n39815 = pi13 ? n39799 : n39814;
  assign n39816 = pi12 ? n39796 : n39815;
  assign n39817 = pi21 ? n206 : n1009;
  assign n39818 = pi20 ? n32 : n39817;
  assign n39819 = pi19 ? n39818 : n32;
  assign n39820 = pi18 ? n32 : n39819;
  assign n39821 = pi17 ? n32 : n39820;
  assign n39822 = pi16 ? n32 : n39821;
  assign n39823 = pi21 ? n206 : ~n7478;
  assign n39824 = pi20 ? n342 : n39823;
  assign n39825 = pi19 ? n39824 : n32;
  assign n39826 = pi18 ? n32 : n39825;
  assign n39827 = pi17 ? n32 : n39826;
  assign n39828 = pi16 ? n32 : n39827;
  assign n39829 = pi15 ? n39822 : n39828;
  assign n39830 = pi14 ? n34408 : n39829;
  assign n39831 = pi20 ? n342 : n1685;
  assign n39832 = pi19 ? n39831 : n32;
  assign n39833 = pi18 ? n32 : n39832;
  assign n39834 = pi17 ? n32 : n39833;
  assign n39835 = pi16 ? n32 : n39834;
  assign n39836 = pi15 ? n39835 : n13920;
  assign n39837 = pi19 ? n15983 : n32;
  assign n39838 = pi18 ? n32 : n39837;
  assign n39839 = pi17 ? n32 : n39838;
  assign n39840 = pi16 ? n32 : n39839;
  assign n39841 = pi15 ? n39840 : n32685;
  assign n39842 = pi14 ? n39836 : n39841;
  assign n39843 = pi13 ? n39830 : n39842;
  assign n39844 = pi15 ? n33939 : n13369;
  assign n39845 = pi18 ? n1741 : ~n605;
  assign n39846 = pi17 ? n32 : n39845;
  assign n39847 = pi16 ? n32 : n39846;
  assign n39848 = pi16 ? n32 : n810;
  assign n39849 = pi15 ? n39847 : n39848;
  assign n39850 = pi14 ? n39844 : n39849;
  assign n39851 = pi15 ? n11863 : n20883;
  assign n39852 = pi14 ? n39851 : n20319;
  assign n39853 = pi13 ? n39850 : n39852;
  assign n39854 = pi12 ? n39843 : n39853;
  assign n39855 = pi11 ? n39816 : n39854;
  assign n39856 = pi10 ? n39780 : n39855;
  assign n39857 = pi09 ? n32 : n39856;
  assign n39858 = pi14 ? n17278 : n32;
  assign n39859 = pi13 ? n32 : n39858;
  assign n39860 = pi12 ? n32 : n39859;
  assign n39861 = pi15 ? n26322 : n38750;
  assign n39862 = pi14 ? n39861 : n24962;
  assign n39863 = pi15 ? n16452 : n39775;
  assign n39864 = pi14 ? n39863 : n15847;
  assign n39865 = pi13 ? n39862 : n39864;
  assign n39866 = pi12 ? n39761 : n39865;
  assign n39867 = pi11 ? n39860 : n39866;
  assign n39868 = pi15 ? n27304 : n39784;
  assign n39869 = pi14 ? n16452 : n39868;
  assign n39870 = pi20 ? n111 : n321;
  assign n39871 = pi19 ? n39870 : ~n589;
  assign n39872 = pi18 ? n32 : n39871;
  assign n39873 = pi17 ? n32 : n39872;
  assign n39874 = pi16 ? n32 : n39873;
  assign n39875 = pi15 ? n15700 : n39874;
  assign n39876 = pi14 ? n39787 : n39875;
  assign n39877 = pi13 ? n39869 : n39876;
  assign n39878 = pi15 ? n23443 : n25247;
  assign n39879 = pi14 ? n39878 : n39481;
  assign n39880 = pi13 ? n39799 : n39879;
  assign n39881 = pi12 ? n39877 : n39880;
  assign n39882 = pi21 ? n206 : ~n1392;
  assign n39883 = pi20 ? n32 : n39882;
  assign n39884 = pi19 ? n39883 : n32;
  assign n39885 = pi18 ? n32 : n39884;
  assign n39886 = pi17 ? n32 : n39885;
  assign n39887 = pi16 ? n32 : n39886;
  assign n39888 = pi15 ? n39887 : n39828;
  assign n39889 = pi14 ? n34408 : n39888;
  assign n39890 = pi20 ? n342 : n7388;
  assign n39891 = pi19 ? n39890 : n32;
  assign n39892 = pi18 ? n32 : n39891;
  assign n39893 = pi17 ? n32 : n39892;
  assign n39894 = pi16 ? n32 : n39893;
  assign n39895 = pi15 ? n39894 : n13642;
  assign n39896 = pi15 ? n24213 : n39840;
  assign n39897 = pi14 ? n39895 : n39896;
  assign n39898 = pi13 ? n39889 : n39897;
  assign n39899 = pi18 ? n209 : ~n2298;
  assign n39900 = pi17 ? n32 : n39899;
  assign n39901 = pi16 ? n32 : n39900;
  assign n39902 = pi15 ? n12304 : n39901;
  assign n39903 = pi14 ? n39844 : n39902;
  assign n39904 = pi18 ? n209 : ~n418;
  assign n39905 = pi17 ? n32 : n39904;
  assign n39906 = pi16 ? n32 : n39905;
  assign n39907 = pi15 ? n39906 : n39901;
  assign n39908 = pi17 ? n32 : n20899;
  assign n39909 = pi16 ? n32 : n39908;
  assign n39910 = pi14 ? n39907 : n39909;
  assign n39911 = pi13 ? n39903 : n39910;
  assign n39912 = pi12 ? n39898 : n39911;
  assign n39913 = pi11 ? n39881 : n39912;
  assign n39914 = pi10 ? n39867 : n39913;
  assign n39915 = pi09 ? n32 : n39914;
  assign n39916 = pi08 ? n39857 : n39915;
  assign n39917 = pi15 ? n26322 : n32;
  assign n39918 = pi14 ? n39917 : n32;
  assign n39919 = pi15 ? n24874 : n25708;
  assign n39920 = pi14 ? n39919 : n26831;
  assign n39921 = pi13 ? n39918 : n39920;
  assign n39922 = pi12 ? n39761 : n39921;
  assign n39923 = pi11 ? n39860 : n39922;
  assign n39924 = pi15 ? n25211 : n16105;
  assign n39925 = pi14 ? n16452 : n39924;
  assign n39926 = pi15 ? n16105 : n24659;
  assign n39927 = pi14 ? n16105 : n39926;
  assign n39928 = pi13 ? n39925 : n39927;
  assign n39929 = pi15 ? n35030 : n14580;
  assign n39930 = pi15 ? n22825 : n27471;
  assign n39931 = pi14 ? n39929 : n39930;
  assign n39932 = pi13 ? n24659 : n39931;
  assign n39933 = pi12 ? n39928 : n39932;
  assign n39934 = pi15 ? n27471 : n14397;
  assign n39935 = pi21 ? n35 : n206;
  assign n39936 = pi20 ? n32 : ~n39935;
  assign n39937 = pi19 ? n39936 : n32;
  assign n39938 = pi18 ? n32 : n39937;
  assign n39939 = pi17 ? n32 : n39938;
  assign n39940 = pi16 ? n32 : n39939;
  assign n39941 = pi15 ? n39940 : n32685;
  assign n39942 = pi14 ? n39934 : n39941;
  assign n39943 = pi15 ? n13660 : n21346;
  assign n39944 = pi14 ? n32685 : n39943;
  assign n39945 = pi13 ? n39942 : n39944;
  assign n39946 = pi14 ? n13369 : n20997;
  assign n39947 = pi18 ? n940 : ~n344;
  assign n39948 = pi17 ? n32 : n39947;
  assign n39949 = pi16 ? n32 : n39948;
  assign n39950 = pi18 ? n863 : ~n1548;
  assign n39951 = pi17 ? n32 : n39950;
  assign n39952 = pi16 ? n32 : n39951;
  assign n39953 = pi15 ? n23240 : n39952;
  assign n39954 = pi14 ? n39949 : n39953;
  assign n39955 = pi13 ? n39946 : n39954;
  assign n39956 = pi12 ? n39945 : n39955;
  assign n39957 = pi11 ? n39933 : n39956;
  assign n39958 = pi10 ? n39923 : n39957;
  assign n39959 = pi09 ? n32 : n39958;
  assign n39960 = pi14 ? n32 : n16736;
  assign n39961 = pi13 ? n39960 : n17039;
  assign n39962 = pi12 ? n39961 : n39921;
  assign n39963 = pi11 ? n39860 : n39962;
  assign n39964 = pi19 ? n2359 : ~n236;
  assign n39965 = pi18 ? n32 : n39964;
  assign n39966 = pi17 ? n32 : n39965;
  assign n39967 = pi16 ? n32 : n39966;
  assign n39968 = pi15 ? n24659 : n39967;
  assign n39969 = pi14 ? n24659 : n39968;
  assign n39970 = pi19 ? n340 : ~n236;
  assign n39971 = pi18 ? n32 : n39970;
  assign n39972 = pi17 ? n32 : n39971;
  assign n39973 = pi16 ? n32 : n39972;
  assign n39974 = pi15 ? n39973 : n14580;
  assign n39975 = pi14 ? n39974 : n39930;
  assign n39976 = pi13 ? n39969 : n39975;
  assign n39977 = pi12 ? n39928 : n39976;
  assign n39978 = pi15 ? n27471 : n21954;
  assign n39979 = pi19 ? n261 : n32;
  assign n39980 = pi18 ? n32 : n39979;
  assign n39981 = pi17 ? n32 : n39980;
  assign n39982 = pi16 ? n32 : n39981;
  assign n39983 = pi15 ? n39982 : n32685;
  assign n39984 = pi14 ? n39978 : n39983;
  assign n39985 = pi13 ? n39984 : n39944;
  assign n39986 = pi14 ? n13369 : n12542;
  assign n39987 = pi15 ? n20072 : n20089;
  assign n39988 = pi14 ? n20072 : n39987;
  assign n39989 = pi13 ? n39986 : n39988;
  assign n39990 = pi12 ? n39985 : n39989;
  assign n39991 = pi11 ? n39977 : n39990;
  assign n39992 = pi10 ? n39963 : n39991;
  assign n39993 = pi09 ? n32 : n39992;
  assign n39994 = pi08 ? n39959 : n39993;
  assign n39995 = pi07 ? n39916 : n39994;
  assign n39996 = pi15 ? n16397 : n17039;
  assign n39997 = pi14 ? n32 : n39996;
  assign n39998 = pi15 ? n17039 : n17056;
  assign n39999 = pi14 ? n17039 : n39998;
  assign n40000 = pi13 ? n39997 : n39999;
  assign n40001 = pi15 ? n38071 : n24874;
  assign n40002 = pi14 ? n40001 : n24874;
  assign n40003 = pi13 ? n25133 : n40002;
  assign n40004 = pi12 ? n40000 : n40003;
  assign n40005 = pi11 ? n39860 : n40004;
  assign n40006 = pi15 ? n16606 : n27304;
  assign n40007 = pi14 ? n40006 : n39924;
  assign n40008 = pi15 ? n24504 : n15834;
  assign n40009 = pi19 ? n32 : n29918;
  assign n40010 = pi18 ? n32 : n40009;
  assign n40011 = pi17 ? n32 : n40010;
  assign n40012 = pi16 ? n32 : n40011;
  assign n40013 = pi15 ? n40012 : n23484;
  assign n40014 = pi14 ? n40008 : n40013;
  assign n40015 = pi13 ? n40007 : n40014;
  assign n40016 = pi19 ? n4721 : ~n236;
  assign n40017 = pi18 ? n32 : n40016;
  assign n40018 = pi17 ? n32 : n40017;
  assign n40019 = pi16 ? n32 : n40018;
  assign n40020 = pi15 ? n40019 : n14138;
  assign n40021 = pi14 ? n24660 : n40020;
  assign n40022 = pi19 ? n340 : n32;
  assign n40023 = pi18 ? n32 : n40022;
  assign n40024 = pi17 ? n32 : n40023;
  assign n40025 = pi16 ? n32 : n40024;
  assign n40026 = pi15 ? n40025 : n22825;
  assign n40027 = pi15 ? n22825 : n33970;
  assign n40028 = pi14 ? n40026 : n40027;
  assign n40029 = pi13 ? n40021 : n40028;
  assign n40030 = pi12 ? n40015 : n40029;
  assign n40031 = pi15 ? n20660 : n13660;
  assign n40032 = pi14 ? n32 : n40031;
  assign n40033 = pi15 ? n32685 : n13360;
  assign n40034 = pi15 ? n32698 : n13369;
  assign n40035 = pi14 ? n40033 : n40034;
  assign n40036 = pi13 ? n40032 : n40035;
  assign n40037 = pi14 ? n13381 : n13083;
  assign n40038 = pi15 ? n20323 : n20067;
  assign n40039 = pi14 ? n40038 : n19814;
  assign n40040 = pi13 ? n40037 : n40039;
  assign n40041 = pi12 ? n40036 : n40040;
  assign n40042 = pi11 ? n40030 : n40041;
  assign n40043 = pi10 ? n40005 : n40042;
  assign n40044 = pi09 ? n32 : n40043;
  assign n40045 = pi14 ? n17273 : n39996;
  assign n40046 = pi14 ? n17039 : n39388;
  assign n40047 = pi13 ? n40045 : n40046;
  assign n40048 = pi15 ? n25708 : n24874;
  assign n40049 = pi14 ? n40048 : n24874;
  assign n40050 = pi13 ? n25133 : n40049;
  assign n40051 = pi12 ? n40047 : n40050;
  assign n40052 = pi11 ? n39860 : n40051;
  assign n40053 = pi20 ? n17389 : n32;
  assign n40054 = pi19 ? n32 : n40053;
  assign n40055 = pi18 ? n32 : n40054;
  assign n40056 = pi17 ? n32 : n40055;
  assign n40057 = pi16 ? n32 : n40056;
  assign n40058 = pi15 ? n40057 : n23484;
  assign n40059 = pi14 ? n40008 : n40058;
  assign n40060 = pi13 ? n40007 : n40059;
  assign n40061 = pi18 ? n32 : n6623;
  assign n40062 = pi17 ? n32 : n40061;
  assign n40063 = pi16 ? n32 : n40062;
  assign n40064 = pi15 ? n22825 : n40063;
  assign n40065 = pi14 ? n40026 : n40064;
  assign n40066 = pi13 ? n40021 : n40065;
  assign n40067 = pi12 ? n40060 : n40066;
  assign n40068 = pi15 ? n13948 : n13660;
  assign n40069 = pi14 ? n32 : n40068;
  assign n40070 = pi20 ? n749 : n357;
  assign n40071 = pi19 ? n40070 : n32;
  assign n40072 = pi18 ? n32 : n40071;
  assign n40073 = pi17 ? n32 : n40072;
  assign n40074 = pi16 ? n32 : n40073;
  assign n40075 = pi15 ? n32698 : n40074;
  assign n40076 = pi14 ? n21636 : n40075;
  assign n40077 = pi13 ? n40069 : n40076;
  assign n40078 = pi19 ? n15674 : n32;
  assign n40079 = pi18 ? n32 : n40078;
  assign n40080 = pi17 ? n32 : n40079;
  assign n40081 = pi16 ? n32 : n40080;
  assign n40082 = pi15 ? n40081 : n20692;
  assign n40083 = pi19 ? n16247 : n32;
  assign n40084 = pi18 ? n32 : n40083;
  assign n40085 = pi17 ? n32 : n40084;
  assign n40086 = pi16 ? n32 : n40085;
  assign n40087 = pi15 ? n40086 : n20692;
  assign n40088 = pi14 ? n40082 : n40087;
  assign n40089 = pi15 ? n19805 : n19235;
  assign n40090 = pi14 ? n40089 : n32;
  assign n40091 = pi13 ? n40088 : n40090;
  assign n40092 = pi12 ? n40077 : n40091;
  assign n40093 = pi11 ? n40067 : n40092;
  assign n40094 = pi10 ? n40052 : n40093;
  assign n40095 = pi09 ? n32 : n40094;
  assign n40096 = pi08 ? n40044 : n40095;
  assign n40097 = pi15 ? n16397 : n32;
  assign n40098 = pi14 ? n17273 : n40097;
  assign n40099 = pi14 ? n25133 : n39388;
  assign n40100 = pi13 ? n40098 : n40099;
  assign n40101 = pi15 ? n17039 : n16837;
  assign n40102 = pi14 ? n25133 : n40101;
  assign n40103 = pi15 ? n25704 : n26009;
  assign n40104 = pi15 ? n24874 : n26009;
  assign n40105 = pi14 ? n40103 : n40104;
  assign n40106 = pi13 ? n40102 : n40105;
  assign n40107 = pi12 ? n40100 : n40106;
  assign n40108 = pi11 ? n39860 : n40107;
  assign n40109 = pi15 ? n16452 : n25211;
  assign n40110 = pi19 ? n2092 : ~n236;
  assign n40111 = pi18 ? n32 : n40110;
  assign n40112 = pi17 ? n32 : n40111;
  assign n40113 = pi16 ? n32 : n40112;
  assign n40114 = pi15 ? n24504 : n40113;
  assign n40115 = pi14 ? n40109 : n40114;
  assign n40116 = pi15 ? n23250 : n15834;
  assign n40117 = pi19 ? n4491 : n15651;
  assign n40118 = pi18 ? n32 : n40117;
  assign n40119 = pi17 ? n32 : n40118;
  assign n40120 = pi16 ? n32 : n40119;
  assign n40121 = pi15 ? n40120 : n39354;
  assign n40122 = pi14 ? n40116 : n40121;
  assign n40123 = pi13 ? n40115 : n40122;
  assign n40124 = pi15 ? n25657 : n24659;
  assign n40125 = pi15 ? n36631 : n14138;
  assign n40126 = pi14 ? n40124 : n40125;
  assign n40127 = pi15 ? n40025 : n39982;
  assign n40128 = pi15 ? n14379 : n14156;
  assign n40129 = pi14 ? n40127 : n40128;
  assign n40130 = pi13 ? n40126 : n40129;
  assign n40131 = pi12 ? n40123 : n40130;
  assign n40132 = pi14 ? n33931 : n40068;
  assign n40133 = pi15 ? n13360 : n13369;
  assign n40134 = pi19 ? n25700 : n32;
  assign n40135 = pi18 ? n32 : n40134;
  assign n40136 = pi17 ? n32 : n40135;
  assign n40137 = pi16 ? n32 : n40136;
  assign n40138 = pi15 ? n40137 : n20618;
  assign n40139 = pi14 ? n40133 : n40138;
  assign n40140 = pi13 ? n40132 : n40139;
  assign n40141 = pi15 ? n13386 : n19972;
  assign n40142 = pi14 ? n19755 : n32;
  assign n40143 = pi13 ? n40141 : n40142;
  assign n40144 = pi12 ? n40140 : n40143;
  assign n40145 = pi11 ? n40131 : n40144;
  assign n40146 = pi10 ? n40108 : n40145;
  assign n40147 = pi09 ? n32 : n40146;
  assign n40148 = pi14 ? n16985 : n40097;
  assign n40149 = pi20 ? n428 : n6229;
  assign n40150 = pi19 ? n32 : n40149;
  assign n40151 = pi18 ? n32 : n40150;
  assign n40152 = pi17 ? n32 : n40151;
  assign n40153 = pi16 ? n32 : n40152;
  assign n40154 = pi15 ? n40153 : n26322;
  assign n40155 = pi14 ? n25133 : n40154;
  assign n40156 = pi13 ? n40148 : n40155;
  assign n40157 = pi20 ? n13785 : n481;
  assign n40158 = pi19 ? n32 : n40157;
  assign n40159 = pi18 ? n32 : n40158;
  assign n40160 = pi17 ? n32 : n40159;
  assign n40161 = pi16 ? n32 : n40160;
  assign n40162 = pi15 ? n17039 : n40161;
  assign n40163 = pi14 ? n25133 : n40162;
  assign n40164 = pi14 ? n40103 : n24874;
  assign n40165 = pi13 ? n40163 : n40164;
  assign n40166 = pi12 ? n40156 : n40165;
  assign n40167 = pi11 ? n39860 : n40166;
  assign n40168 = pi15 ? n24504 : n23484;
  assign n40169 = pi14 ? n40109 : n40168;
  assign n40170 = pi19 ? n857 : ~n349;
  assign n40171 = pi18 ? n32 : n40170;
  assign n40172 = pi17 ? n32 : n40171;
  assign n40173 = pi16 ? n32 : n40172;
  assign n40174 = pi15 ? n23250 : n40173;
  assign n40175 = pi20 ? n32 : n9013;
  assign n40176 = pi19 ? n40175 : ~n236;
  assign n40177 = pi18 ? n32 : n40176;
  assign n40178 = pi17 ? n32 : n40177;
  assign n40179 = pi16 ? n32 : n40178;
  assign n40180 = pi15 ? n40179 : n24742;
  assign n40181 = pi14 ? n40174 : n40180;
  assign n40182 = pi13 ? n40169 : n40181;
  assign n40183 = pi19 ? n355 : n32;
  assign n40184 = pi18 ? n32 : n40183;
  assign n40185 = pi17 ? n32 : n40184;
  assign n40186 = pi16 ? n32 : n40185;
  assign n40187 = pi15 ? n40186 : n39982;
  assign n40188 = pi15 ? n39982 : n21954;
  assign n40189 = pi14 ? n40187 : n40188;
  assign n40190 = pi13 ? n40126 : n40189;
  assign n40191 = pi12 ? n40182 : n40190;
  assign n40192 = pi15 ? n20660 : n14156;
  assign n40193 = pi19 ? n1011 : n32;
  assign n40194 = pi18 ? n32 : n40193;
  assign n40195 = pi17 ? n32 : n40194;
  assign n40196 = pi16 ? n32 : n40195;
  assign n40197 = pi15 ? n40196 : n13660;
  assign n40198 = pi14 ? n40192 : n40197;
  assign n40199 = pi15 ? n20301 : n20048;
  assign n40200 = pi14 ? n21346 : n40199;
  assign n40201 = pi13 ? n40198 : n40200;
  assign n40202 = pi12 ? n40201 : n32;
  assign n40203 = pi11 ? n40191 : n40202;
  assign n40204 = pi10 ? n40167 : n40203;
  assign n40205 = pi09 ? n32 : n40204;
  assign n40206 = pi08 ? n40147 : n40205;
  assign n40207 = pi07 ? n40096 : n40206;
  assign n40208 = pi06 ? n39995 : n40207;
  assign n40209 = pi05 ? n39756 : n40208;
  assign n40210 = pi04 ? n39385 : n40209;
  assign n40211 = pi15 ? n32 : n17286;
  assign n40212 = pi14 ? n40211 : n40097;
  assign n40213 = pi15 ? n17056 : n26479;
  assign n40214 = pi14 ? n26163 : n40213;
  assign n40215 = pi13 ? n40212 : n40214;
  assign n40216 = pi20 ? n1319 : ~n243;
  assign n40217 = pi19 ? n32 : n40216;
  assign n40218 = pi18 ? n32 : n40217;
  assign n40219 = pi17 ? n32 : n40218;
  assign n40220 = pi16 ? n32 : n40219;
  assign n40221 = pi15 ? n17039 : n40220;
  assign n40222 = pi14 ? n25133 : n40221;
  assign n40223 = pi15 ? n26009 : n24874;
  assign n40224 = pi14 ? n40103 : n40223;
  assign n40225 = pi13 ? n40222 : n40224;
  assign n40226 = pi12 ? n40215 : n40225;
  assign n40227 = pi11 ? n39860 : n40226;
  assign n40228 = pi19 ? n32 : ~n20517;
  assign n40229 = pi18 ? n32 : n40228;
  assign n40230 = pi17 ? n32 : n40229;
  assign n40231 = pi16 ? n32 : n40230;
  assign n40232 = pi15 ? n40231 : n24700;
  assign n40233 = pi15 ? n24511 : n24247;
  assign n40234 = pi14 ? n40232 : n40233;
  assign n40235 = pi15 ? n24572 : n15123;
  assign n40236 = pi15 ? n23484 : n35030;
  assign n40237 = pi14 ? n40235 : n40236;
  assign n40238 = pi13 ? n40234 : n40237;
  assign n40239 = pi15 ? n14358 : n40025;
  assign n40240 = pi14 ? n39929 : n40239;
  assign n40241 = pi15 ? n40025 : n14363;
  assign n40242 = pi14 ? n40241 : n14156;
  assign n40243 = pi13 ? n40240 : n40242;
  assign n40244 = pi12 ? n40238 : n40243;
  assign n40245 = pi15 ? n14156 : n13948;
  assign n40246 = pi14 ? n40245 : n13948;
  assign n40247 = pi14 ? n13953 : n32;
  assign n40248 = pi13 ? n40246 : n40247;
  assign n40249 = pi12 ? n40248 : n32;
  assign n40250 = pi11 ? n40244 : n40249;
  assign n40251 = pi10 ? n40227 : n40250;
  assign n40252 = pi09 ? n32 : n40251;
  assign n40253 = pi15 ? n16392 : n40220;
  assign n40254 = pi14 ? n25133 : n40253;
  assign n40255 = pi15 ? n25704 : n39670;
  assign n40256 = pi14 ? n40255 : n24874;
  assign n40257 = pi13 ? n40254 : n40256;
  assign n40258 = pi12 ? n40215 : n40257;
  assign n40259 = pi11 ? n39860 : n40258;
  assign n40260 = pi19 ? n126 : ~n20517;
  assign n40261 = pi18 ? n32 : n40260;
  assign n40262 = pi17 ? n32 : n40261;
  assign n40263 = pi16 ? n32 : n40262;
  assign n40264 = pi15 ? n40263 : n24700;
  assign n40265 = pi15 ? n24640 : n24247;
  assign n40266 = pi14 ? n40264 : n40265;
  assign n40267 = pi15 ? n24572 : n32;
  assign n40268 = pi20 ? n1393 : ~n32;
  assign n40269 = pi19 ? n208 : ~n40268;
  assign n40270 = pi18 ? n32 : n40269;
  assign n40271 = pi17 ? n32 : n40270;
  assign n40272 = pi16 ? n32 : n40271;
  assign n40273 = pi15 ? n23484 : n40272;
  assign n40274 = pi14 ? n40267 : n40273;
  assign n40275 = pi13 ? n40266 : n40274;
  assign n40276 = pi15 ? n40272 : n14580;
  assign n40277 = pi14 ? n40276 : n40239;
  assign n40278 = pi19 ? n365 : n32;
  assign n40279 = pi18 ? n32 : n40278;
  assign n40280 = pi17 ? n32 : n40279;
  assign n40281 = pi16 ? n32 : n40280;
  assign n40282 = pi15 ? n40281 : n14363;
  assign n40283 = pi14 ? n40282 : n21954;
  assign n40284 = pi13 ? n40277 : n40283;
  assign n40285 = pi12 ? n40275 : n40284;
  assign n40286 = pi20 ? n32 : n15961;
  assign n40287 = pi19 ? n40286 : n32;
  assign n40288 = pi18 ? n32 : n40287;
  assign n40289 = pi17 ? n32 : n40288;
  assign n40290 = pi16 ? n32 : n40289;
  assign n40291 = pi15 ? n40290 : n20660;
  assign n40292 = pi15 ? n666 : n32;
  assign n40293 = pi14 ? n40291 : n40292;
  assign n40294 = pi13 ? n40293 : n32;
  assign n40295 = pi12 ? n40294 : n32;
  assign n40296 = pi11 ? n40285 : n40295;
  assign n40297 = pi10 ? n40259 : n40296;
  assign n40298 = pi09 ? n32 : n40297;
  assign n40299 = pi08 ? n40252 : n40298;
  assign n40300 = pi15 ? n16824 : n26479;
  assign n40301 = pi14 ? n16393 : n40300;
  assign n40302 = pi13 ? n40212 : n40301;
  assign n40303 = pi15 ? n32 : n40220;
  assign n40304 = pi14 ? n16392 : n40303;
  assign n40305 = pi15 ? n26009 : n39670;
  assign n40306 = pi14 ? n40305 : n24874;
  assign n40307 = pi13 ? n40304 : n40306;
  assign n40308 = pi12 ? n40302 : n40307;
  assign n40309 = pi11 ? n39860 : n40308;
  assign n40310 = pi19 ? n32 : ~n12020;
  assign n40311 = pi18 ? n32 : n40310;
  assign n40312 = pi17 ? n32 : n40311;
  assign n40313 = pi16 ? n32 : n40312;
  assign n40314 = pi19 ? n1818 : ~n343;
  assign n40315 = pi18 ? n32 : n40314;
  assign n40316 = pi17 ? n32 : n40315;
  assign n40317 = pi16 ? n32 : n40316;
  assign n40318 = pi15 ? n40313 : n40317;
  assign n40319 = pi21 ? n35 : ~n259;
  assign n40320 = pi20 ? n32 : n40319;
  assign n40321 = pi19 ? n40320 : ~n2317;
  assign n40322 = pi18 ? n32 : n40321;
  assign n40323 = pi17 ? n32 : n40322;
  assign n40324 = pi16 ? n32 : n40323;
  assign n40325 = pi19 ? n662 : ~n589;
  assign n40326 = pi18 ? n32 : n40325;
  assign n40327 = pi17 ? n32 : n40326;
  assign n40328 = pi16 ? n32 : n40327;
  assign n40329 = pi15 ? n40324 : n40328;
  assign n40330 = pi14 ? n40318 : n40329;
  assign n40331 = pi15 ? n26623 : n24659;
  assign n40332 = pi14 ? n32 : n40331;
  assign n40333 = pi13 ? n40330 : n40332;
  assign n40334 = pi19 ? n1165 : n32;
  assign n40335 = pi18 ? n32 : n40334;
  assign n40336 = pi17 ? n32 : n40335;
  assign n40337 = pi16 ? n32 : n40336;
  assign n40338 = pi19 ? n750 : ~n617;
  assign n40339 = pi18 ? n32 : n40338;
  assign n40340 = pi17 ? n32 : n40339;
  assign n40341 = pi16 ? n32 : n40340;
  assign n40342 = pi15 ? n40337 : n40341;
  assign n40343 = pi15 ? n40341 : n25247;
  assign n40344 = pi14 ? n40342 : n40343;
  assign n40345 = pi19 ? n24204 : n32;
  assign n40346 = pi18 ? n32 : n40345;
  assign n40347 = pi17 ? n32 : n40346;
  assign n40348 = pi16 ? n32 : n40347;
  assign n40349 = pi15 ? n40348 : n40063;
  assign n40350 = pi15 ? n14397 : n21141;
  assign n40351 = pi14 ? n40349 : n40350;
  assign n40352 = pi13 ? n40344 : n40351;
  assign n40353 = pi12 ? n40333 : n40352;
  assign n40354 = pi14 ? n40350 : n32128;
  assign n40355 = pi13 ? n40354 : n32;
  assign n40356 = pi12 ? n40355 : n32;
  assign n40357 = pi11 ? n40353 : n40356;
  assign n40358 = pi10 ? n40309 : n40357;
  assign n40359 = pi09 ? n32 : n40358;
  assign n40360 = pi15 ? n39670 : n26009;
  assign n40361 = pi14 ? n40360 : n24874;
  assign n40362 = pi13 ? n40304 : n40361;
  assign n40363 = pi12 ? n40302 : n40362;
  assign n40364 = pi11 ? n39860 : n40363;
  assign n40365 = pi15 ? n24640 : n24511;
  assign n40366 = pi14 ? n24700 : n40365;
  assign n40367 = pi19 ? n38400 : n32;
  assign n40368 = pi18 ? n32 : n40367;
  assign n40369 = pi17 ? n32 : n40368;
  assign n40370 = pi16 ? n32 : n40369;
  assign n40371 = pi15 ? n32 : n40370;
  assign n40372 = pi14 ? n40371 : n40331;
  assign n40373 = pi13 ? n40366 : n40372;
  assign n40374 = pi21 ? n66 : ~n309;
  assign n40375 = pi20 ? n32 : n40374;
  assign n40376 = pi19 ? n40375 : n32;
  assign n40377 = pi18 ? n32 : n40376;
  assign n40378 = pi17 ? n32 : n40377;
  assign n40379 = pi16 ? n32 : n40378;
  assign n40380 = pi15 ? n40379 : n40341;
  assign n40381 = pi14 ? n40380 : n40343;
  assign n40382 = pi21 ? n100 : n174;
  assign n40383 = pi20 ? n32 : n40382;
  assign n40384 = pi19 ? n40383 : n32;
  assign n40385 = pi18 ? n32 : n40384;
  assign n40386 = pi17 ? n32 : n40385;
  assign n40387 = pi16 ? n32 : n40386;
  assign n40388 = pi15 ? n26663 : n40387;
  assign n40389 = pi21 ? n100 : n51;
  assign n40390 = pi20 ? n32 : n40389;
  assign n40391 = pi19 ? n40390 : n32;
  assign n40392 = pi18 ? n32 : n40391;
  assign n40393 = pi17 ? n32 : n40392;
  assign n40394 = pi16 ? n32 : n40393;
  assign n40395 = pi15 ? n40394 : n648;
  assign n40396 = pi14 ? n40388 : n40395;
  assign n40397 = pi13 ? n40381 : n40396;
  assign n40398 = pi12 ? n40373 : n40397;
  assign n40399 = pi15 ? n658 : n32;
  assign n40400 = pi14 ? n40399 : n32;
  assign n40401 = pi13 ? n40400 : n32;
  assign n40402 = pi12 ? n40401 : n32;
  assign n40403 = pi11 ? n40398 : n40402;
  assign n40404 = pi10 ? n40364 : n40403;
  assign n40405 = pi09 ? n32 : n40404;
  assign n40406 = pi08 ? n40359 : n40405;
  assign n40407 = pi07 ? n40299 : n40406;
  assign n40408 = pi19 ? n32 : n40175;
  assign n40409 = pi18 ? n32 : n40408;
  assign n40410 = pi17 ? n32 : n40409;
  assign n40411 = pi16 ? n32 : n40410;
  assign n40412 = pi15 ? n17278 : n40411;
  assign n40413 = pi14 ? n40412 : n32;
  assign n40414 = pi13 ? n32 : n40413;
  assign n40415 = pi12 ? n32 : n40414;
  assign n40416 = pi15 ? n16984 : n16392;
  assign n40417 = pi14 ? n16851 : n40416;
  assign n40418 = pi20 ? n342 : n7487;
  assign n40419 = pi19 ? n32 : n40418;
  assign n40420 = pi18 ? n32 : n40419;
  assign n40421 = pi17 ? n32 : n40420;
  assign n40422 = pi16 ? n32 : n40421;
  assign n40423 = pi19 ? n32 : n17641;
  assign n40424 = pi18 ? n32 : n40423;
  assign n40425 = pi17 ? n32 : n40424;
  assign n40426 = pi16 ? n32 : n40425;
  assign n40427 = pi15 ? n40422 : n40426;
  assign n40428 = pi14 ? n16392 : n40427;
  assign n40429 = pi13 ? n40417 : n40428;
  assign n40430 = pi20 ? n151 : ~n243;
  assign n40431 = pi19 ? n32 : n40430;
  assign n40432 = pi18 ? n32 : n40431;
  assign n40433 = pi17 ? n32 : n40432;
  assign n40434 = pi16 ? n32 : n40433;
  assign n40435 = pi15 ? n32 : n40434;
  assign n40436 = pi14 ? n16392 : n40435;
  assign n40437 = pi15 ? n24874 : n37998;
  assign n40438 = pi14 ? n37774 : n40437;
  assign n40439 = pi13 ? n40436 : n40438;
  assign n40440 = pi12 ? n40429 : n40439;
  assign n40441 = pi11 ? n40415 : n40440;
  assign n40442 = pi19 ? n507 : n3692;
  assign n40443 = pi18 ? n32 : n40442;
  assign n40444 = pi17 ? n32 : n40443;
  assign n40445 = pi16 ? n32 : n40444;
  assign n40446 = pi15 ? n40445 : n24700;
  assign n40447 = pi15 ? n32 : n15244;
  assign n40448 = pi14 ? n40446 : n40447;
  assign n40449 = pi15 ? n15362 : n22540;
  assign n40450 = pi15 ? n26623 : n15263;
  assign n40451 = pi14 ? n40449 : n40450;
  assign n40452 = pi13 ? n40448 : n40451;
  assign n40453 = pi21 ? n100 : ~n7500;
  assign n40454 = pi20 ? n32 : n40453;
  assign n40455 = pi19 ? n40454 : n32;
  assign n40456 = pi18 ? n32 : n40455;
  assign n40457 = pi17 ? n32 : n40456;
  assign n40458 = pi16 ? n32 : n40457;
  assign n40459 = pi15 ? n40458 : n14785;
  assign n40460 = pi15 ? n25247 : n14798;
  assign n40461 = pi14 ? n40459 : n40460;
  assign n40462 = pi15 ? n21928 : n14798;
  assign n40463 = pi14 ? n21928 : n40462;
  assign n40464 = pi13 ? n40461 : n40463;
  assign n40465 = pi12 ? n40452 : n40464;
  assign n40466 = pi11 ? n40465 : n32;
  assign n40467 = pi10 ? n40441 : n40466;
  assign n40468 = pi09 ? n32 : n40467;
  assign n40469 = pi14 ? n17279 : n32;
  assign n40470 = pi13 ? n32 : n40469;
  assign n40471 = pi12 ? n32 : n40470;
  assign n40472 = pi14 ? n16851 : n25498;
  assign n40473 = pi13 ? n40472 : n40428;
  assign n40474 = pi20 ? n3523 : ~n243;
  assign n40475 = pi19 ? n32 : n40474;
  assign n40476 = pi18 ? n32 : n40475;
  assign n40477 = pi17 ? n32 : n40476;
  assign n40478 = pi16 ? n32 : n40477;
  assign n40479 = pi15 ? n32 : n40478;
  assign n40480 = pi14 ? n16392 : n40479;
  assign n40481 = pi19 ? n23123 : ~n429;
  assign n40482 = pi18 ? n32 : n40481;
  assign n40483 = pi17 ? n32 : n40482;
  assign n40484 = pi16 ? n32 : n40483;
  assign n40485 = pi15 ? n24874 : n40484;
  assign n40486 = pi14 ? n37774 : n40485;
  assign n40487 = pi13 ? n40480 : n40486;
  assign n40488 = pi12 ? n40473 : n40487;
  assign n40489 = pi11 ? n40471 : n40488;
  assign n40490 = pi15 ? n26623 : n15123;
  assign n40491 = pi14 ? n40449 : n40490;
  assign n40492 = pi13 ? n40448 : n40491;
  assign n40493 = pi15 ? n23447 : n14967;
  assign n40494 = pi15 ? n14951 : n14967;
  assign n40495 = pi14 ? n40493 : n40494;
  assign n40496 = pi13 ? n40495 : n32;
  assign n40497 = pi12 ? n40492 : n40496;
  assign n40498 = pi11 ? n40497 : n32;
  assign n40499 = pi10 ? n40489 : n40498;
  assign n40500 = pi09 ? n32 : n40499;
  assign n40501 = pi08 ? n40468 : n40500;
  assign n40502 = pi14 ? n39229 : n25498;
  assign n40503 = pi13 ? n40502 : n16392;
  assign n40504 = pi14 ? n16392 : n39563;
  assign n40505 = pi19 ? n472 : ~n343;
  assign n40506 = pi18 ? n32 : n40505;
  assign n40507 = pi17 ? n32 : n40506;
  assign n40508 = pi16 ? n32 : n40507;
  assign n40509 = pi15 ? n16101 : n40508;
  assign n40510 = pi14 ? n16452 : n40509;
  assign n40511 = pi13 ? n40504 : n40510;
  assign n40512 = pi12 ? n40503 : n40511;
  assign n40513 = pi11 ? n40471 : n40512;
  assign n40514 = pi19 ? n472 : n3692;
  assign n40515 = pi18 ? n32 : n40514;
  assign n40516 = pi17 ? n32 : n40515;
  assign n40517 = pi16 ? n32 : n40516;
  assign n40518 = pi15 ? n40517 : n24511;
  assign n40519 = pi15 ? n22817 : n15244;
  assign n40520 = pi14 ? n40518 : n40519;
  assign n40521 = pi14 ? n36865 : n22252;
  assign n40522 = pi13 ? n40520 : n40521;
  assign n40523 = pi14 ? n22817 : n15267;
  assign n40524 = pi13 ? n40523 : n32;
  assign n40525 = pi12 ? n40522 : n40524;
  assign n40526 = pi11 ? n40525 : n32;
  assign n40527 = pi10 ? n40513 : n40526;
  assign n40528 = pi09 ? n32 : n40527;
  assign n40529 = pi15 ? n16101 : n24700;
  assign n40530 = pi14 ? n16452 : n40529;
  assign n40531 = pi13 ? n40504 : n40530;
  assign n40532 = pi12 ? n40503 : n40531;
  assign n40533 = pi11 ? n40471 : n40532;
  assign n40534 = pi15 ? n16101 : n24511;
  assign n40535 = pi19 ? n2141 : ~n349;
  assign n40536 = pi18 ? n32 : n40535;
  assign n40537 = pi17 ? n32 : n40536;
  assign n40538 = pi16 ? n32 : n40537;
  assign n40539 = pi15 ? n22540 : n40538;
  assign n40540 = pi14 ? n40534 : n40539;
  assign n40541 = pi15 ? n40538 : n32;
  assign n40542 = pi14 ? n40541 : n22205;
  assign n40543 = pi13 ? n40540 : n40542;
  assign n40544 = pi14 ? n15263 : n32;
  assign n40545 = pi13 ? n40544 : n32;
  assign n40546 = pi12 ? n40543 : n40545;
  assign n40547 = pi11 ? n40546 : n32;
  assign n40548 = pi10 ? n40533 : n40547;
  assign n40549 = pi09 ? n32 : n40548;
  assign n40550 = pi08 ? n40528 : n40549;
  assign n40551 = pi07 ? n40501 : n40550;
  assign n40552 = pi06 ? n40407 : n40551;
  assign n40553 = pi14 ? n17188 : n16832;
  assign n40554 = pi20 ? n342 : n6229;
  assign n40555 = pi19 ? n32 : n40554;
  assign n40556 = pi18 ? n32 : n40555;
  assign n40557 = pi17 ? n32 : n40556;
  assign n40558 = pi16 ? n32 : n40557;
  assign n40559 = pi15 ? n16392 : n40558;
  assign n40560 = pi14 ? n40559 : n16392;
  assign n40561 = pi13 ? n40553 : n40560;
  assign n40562 = pi15 ? n16392 : n32;
  assign n40563 = pi14 ? n40562 : n39563;
  assign n40564 = pi19 ? n594 : ~n343;
  assign n40565 = pi18 ? n32 : n40564;
  assign n40566 = pi17 ? n32 : n40565;
  assign n40567 = pi16 ? n32 : n40566;
  assign n40568 = pi15 ? n40567 : n24700;
  assign n40569 = pi14 ? n16452 : n40568;
  assign n40570 = pi13 ? n40563 : n40569;
  assign n40571 = pi12 ? n40561 : n40570;
  assign n40572 = pi11 ? n40471 : n40571;
  assign n40573 = pi15 ? n24504 : n24511;
  assign n40574 = pi19 ? n1574 : ~n236;
  assign n40575 = pi18 ? n32 : n40574;
  assign n40576 = pi17 ? n32 : n40575;
  assign n40577 = pi16 ? n32 : n40576;
  assign n40578 = pi15 ? n40577 : n24528;
  assign n40579 = pi14 ? n40573 : n40578;
  assign n40580 = pi15 ? n24528 : n22923;
  assign n40581 = pi14 ? n40580 : n22923;
  assign n40582 = pi13 ? n40579 : n40581;
  assign n40583 = pi12 ? n40582 : n32;
  assign n40584 = pi11 ? n40583 : n32;
  assign n40585 = pi10 ? n40572 : n40584;
  assign n40586 = pi09 ? n32 : n40585;
  assign n40587 = pi14 ? n17273 : n16832;
  assign n40588 = pi13 ? n40587 : n16392;
  assign n40589 = pi14 ? n16452 : n15501;
  assign n40590 = pi13 ? n40563 : n40589;
  assign n40591 = pi12 ? n40588 : n40590;
  assign n40592 = pi11 ? n40471 : n40591;
  assign n40593 = pi15 ? n23484 : n24274;
  assign n40594 = pi14 ? n25779 : n40593;
  assign n40595 = pi15 ? n24274 : n15665;
  assign n40596 = pi14 ? n24274 : n40595;
  assign n40597 = pi13 ? n40594 : n40596;
  assign n40598 = pi12 ? n40597 : n32;
  assign n40599 = pi11 ? n40598 : n32;
  assign n40600 = pi10 ? n40592 : n40599;
  assign n40601 = pi09 ? n32 : n40600;
  assign n40602 = pi08 ? n40586 : n40601;
  assign n40603 = pi14 ? n27678 : n16452;
  assign n40604 = pi21 ? n1939 : ~n405;
  assign n40605 = pi20 ? n40604 : n32;
  assign n40606 = pi19 ? n32 : n40605;
  assign n40607 = pi18 ? n32 : n40606;
  assign n40608 = pi17 ? n32 : n40607;
  assign n40609 = pi16 ? n32 : n40608;
  assign n40610 = pi15 ? n40609 : n16101;
  assign n40611 = pi15 ? n16101 : n15834;
  assign n40612 = pi14 ? n40610 : n40611;
  assign n40613 = pi13 ? n40603 : n40612;
  assign n40614 = pi12 ? n40588 : n40613;
  assign n40615 = pi11 ? n40471 : n40614;
  assign n40616 = pi15 ? n16319 : n15650;
  assign n40617 = pi15 ? n15650 : n16108;
  assign n40618 = pi14 ? n40616 : n40617;
  assign n40619 = pi13 ? n40618 : n32;
  assign n40620 = pi12 ? n40619 : n32;
  assign n40621 = pi11 ? n40620 : n32;
  assign n40622 = pi10 ? n40615 : n40621;
  assign n40623 = pi09 ? n32 : n40622;
  assign n40624 = pi15 ? n17111 : n17188;
  assign n40625 = pi14 ? n40624 : n16832;
  assign n40626 = pi13 ? n40625 : n16392;
  assign n40627 = pi21 ? n66 : ~n206;
  assign n40628 = pi20 ? n40627 : n32;
  assign n40629 = pi19 ? n32 : n40628;
  assign n40630 = pi18 ? n32 : n40629;
  assign n40631 = pi17 ? n32 : n40630;
  assign n40632 = pi16 ? n32 : n40631;
  assign n40633 = pi15 ? n16392 : n40632;
  assign n40634 = pi14 ? n40633 : n16452;
  assign n40635 = pi15 ? n16101 : n15966;
  assign n40636 = pi14 ? n40610 : n40635;
  assign n40637 = pi13 ? n40634 : n40636;
  assign n40638 = pi12 ? n40626 : n40637;
  assign n40639 = pi11 ? n40471 : n40638;
  assign n40640 = pi21 ? n7659 : n32;
  assign n40641 = pi20 ? n40640 : n32;
  assign n40642 = pi19 ? n32 : n40641;
  assign n40643 = pi18 ? n32 : n40642;
  assign n40644 = pi17 ? n32 : n40643;
  assign n40645 = pi16 ? n32 : n40644;
  assign n40646 = pi15 ? n40645 : n15966;
  assign n40647 = pi15 ? n15966 : n23741;
  assign n40648 = pi14 ? n40646 : n40647;
  assign n40649 = pi13 ? n40648 : n23327;
  assign n40650 = pi12 ? n40649 : n32;
  assign n40651 = pi11 ? n40650 : n32;
  assign n40652 = pi10 ? n40639 : n40651;
  assign n40653 = pi09 ? n32 : n40652;
  assign n40654 = pi08 ? n40623 : n40653;
  assign n40655 = pi07 ? n40602 : n40654;
  assign n40656 = pi20 ? n321 : n564;
  assign n40657 = pi19 ? n32 : n40656;
  assign n40658 = pi18 ? n32 : n40657;
  assign n40659 = pi17 ? n32 : n40658;
  assign n40660 = pi16 ? n32 : n40659;
  assign n40661 = pi15 ? n40660 : n16485;
  assign n40662 = pi14 ? n40661 : n16485;
  assign n40663 = pi15 ? n16352 : n15847;
  assign n40664 = pi14 ? n40663 : n15847;
  assign n40665 = pi13 ? n40662 : n40664;
  assign n40666 = pi15 ? n15847 : n23569;
  assign n40667 = pi14 ? n40666 : n37774;
  assign n40668 = pi15 ? n16204 : n16101;
  assign n40669 = pi14 ? n40668 : n40635;
  assign n40670 = pi13 ? n40667 : n40669;
  assign n40671 = pi12 ? n40665 : n40670;
  assign n40672 = pi11 ? n40471 : n40671;
  assign n40673 = pi15 ? n40645 : n16105;
  assign n40674 = pi14 ? n40673 : n23421;
  assign n40675 = pi13 ? n40674 : n32;
  assign n40676 = pi12 ? n40675 : n32;
  assign n40677 = pi11 ? n40676 : n32;
  assign n40678 = pi10 ? n40672 : n40677;
  assign n40679 = pi09 ? n32 : n40678;
  assign n40680 = pi15 ? n15852 : n16485;
  assign n40681 = pi14 ? n40680 : n16485;
  assign n40682 = pi13 ? n40681 : n40664;
  assign n40683 = pi15 ? n16452 : n40609;
  assign n40684 = pi14 ? n25818 : n40683;
  assign n40685 = pi21 ? n11567 : ~n206;
  assign n40686 = pi20 ? n40685 : n32;
  assign n40687 = pi19 ? n32 : n40686;
  assign n40688 = pi18 ? n32 : n40687;
  assign n40689 = pi17 ? n32 : n40688;
  assign n40690 = pi16 ? n32 : n40689;
  assign n40691 = pi15 ? n40690 : n15700;
  assign n40692 = pi14 ? n40668 : n40691;
  assign n40693 = pi13 ? n40684 : n40692;
  assign n40694 = pi12 ? n40682 : n40693;
  assign n40695 = pi11 ? n40471 : n40694;
  assign n40696 = pi14 ? n15700 : n32;
  assign n40697 = pi13 ? n40696 : n32;
  assign n40698 = pi12 ? n40697 : n32;
  assign n40699 = pi11 ? n40698 : n32;
  assign n40700 = pi10 ? n40695 : n40699;
  assign n40701 = pi09 ? n32 : n40700;
  assign n40702 = pi08 ? n40679 : n40701;
  assign n40703 = pi15 ? n24874 : n16298;
  assign n40704 = pi14 ? n24633 : n40703;
  assign n40705 = pi15 ? n16293 : n16319;
  assign n40706 = pi14 ? n16298 : n40705;
  assign n40707 = pi13 ? n40704 : n40706;
  assign n40708 = pi12 ? n40682 : n40707;
  assign n40709 = pi11 ? n40471 : n40708;
  assign n40710 = pi13 ? n37047 : n32;
  assign n40711 = pi12 ? n40710 : n32;
  assign n40712 = pi11 ? n40711 : n32;
  assign n40713 = pi10 ? n40709 : n40712;
  assign n40714 = pi09 ? n32 : n40713;
  assign n40715 = pi14 ? n24633 : n38362;
  assign n40716 = pi15 ? n16452 : n16293;
  assign n40717 = pi14 ? n40716 : n25070;
  assign n40718 = pi13 ? n40715 : n40717;
  assign n40719 = pi12 ? n40682 : n40718;
  assign n40720 = pi11 ? n40471 : n40719;
  assign n40721 = pi10 ? n40720 : n32;
  assign n40722 = pi09 ? n32 : n40721;
  assign n40723 = pi08 ? n40714 : n40722;
  assign n40724 = pi07 ? n40702 : n40723;
  assign n40725 = pi06 ? n40655 : n40724;
  assign n40726 = pi05 ? n40552 : n40725;
  assign n40727 = pi14 ? n17388 : n32;
  assign n40728 = pi13 ? n32 : n40727;
  assign n40729 = pi12 ? n32 : n40728;
  assign n40730 = pi20 ? n342 : n1010;
  assign n40731 = pi19 ? n32 : n40730;
  assign n40732 = pi18 ? n32 : n40731;
  assign n40733 = pi17 ? n32 : n40732;
  assign n40734 = pi16 ? n32 : n40733;
  assign n40735 = pi15 ? n40734 : n16832;
  assign n40736 = pi14 ? n40735 : n16832;
  assign n40737 = pi15 ? n40426 : n16392;
  assign n40738 = pi14 ? n40737 : n25502;
  assign n40739 = pi13 ? n40736 : n40738;
  assign n40740 = pi14 ? n38635 : n16377;
  assign n40741 = pi13 ? n16515 : n40740;
  assign n40742 = pi12 ? n40739 : n40741;
  assign n40743 = pi11 ? n40729 : n40742;
  assign n40744 = pi10 ? n40743 : n32;
  assign n40745 = pi09 ? n32 : n40744;
  assign n40746 = pi14 ? n16833 : n16832;
  assign n40747 = pi15 ? n16392 : n16333;
  assign n40748 = pi14 ? n40737 : n40747;
  assign n40749 = pi13 ? n40746 : n40748;
  assign n40750 = pi14 ? n16515 : n16378;
  assign n40751 = pi13 ? n16515 : n40750;
  assign n40752 = pi12 ? n40749 : n40751;
  assign n40753 = pi11 ? n40729 : n40752;
  assign n40754 = pi10 ? n40753 : n32;
  assign n40755 = pi09 ? n32 : n40754;
  assign n40756 = pi08 ? n40745 : n40755;
  assign n40757 = pi14 ? n16832 : n25633;
  assign n40758 = pi15 ? n16392 : n16546;
  assign n40759 = pi14 ? n40758 : n38511;
  assign n40760 = pi13 ? n40757 : n40759;
  assign n40761 = pi13 ? n16606 : n32;
  assign n40762 = pi12 ? n40760 : n40761;
  assign n40763 = pi11 ? n32 : n40762;
  assign n40764 = pi10 ? n40763 : n32;
  assign n40765 = pi09 ? n32 : n40764;
  assign n40766 = pi07 ? n40756 : n40765;
  assign n40767 = pi12 ? n32 : n25289;
  assign n40768 = pi14 ? n37225 : n25633;
  assign n40769 = pi15 ? n16392 : n16467;
  assign n40770 = pi14 ? n40769 : n16467;
  assign n40771 = pi13 ? n40768 : n40770;
  assign n40772 = pi15 ? n24495 : n32;
  assign n40773 = pi14 ? n39671 : n40772;
  assign n40774 = pi13 ? n40773 : n32;
  assign n40775 = pi12 ? n40771 : n40774;
  assign n40776 = pi11 ? n40767 : n40775;
  assign n40777 = pi10 ? n40776 : n32;
  assign n40778 = pi09 ? n32 : n40777;
  assign n40779 = pi13 ? n40768 : n16467;
  assign n40780 = pi14 ? n39671 : n32;
  assign n40781 = pi13 ? n40780 : n32;
  assign n40782 = pi12 ? n40779 : n40781;
  assign n40783 = pi11 ? n40767 : n40782;
  assign n40784 = pi10 ? n40783 : n32;
  assign n40785 = pi09 ? n32 : n40784;
  assign n40786 = pi08 ? n40778 : n40785;
  assign n40787 = pi14 ? n16392 : n26250;
  assign n40788 = pi13 ? n40757 : n40787;
  assign n40789 = pi12 ? n40788 : n32;
  assign n40790 = pi11 ? n40767 : n40789;
  assign n40791 = pi10 ? n40790 : n32;
  assign n40792 = pi09 ? n32 : n40791;
  assign n40793 = pi07 ? n40786 : n40792;
  assign n40794 = pi06 ? n40766 : n40793;
  assign n40795 = pi15 ? n16953 : n16965;
  assign n40796 = pi14 ? n17036 : n40795;
  assign n40797 = pi15 ? n16965 : n36851;
  assign n40798 = pi14 ? n16965 : n40797;
  assign n40799 = pi13 ? n40796 : n40798;
  assign n40800 = pi15 ? n36851 : n32;
  assign n40801 = pi14 ? n40800 : n32;
  assign n40802 = pi13 ? n40801 : n32;
  assign n40803 = pi12 ? n40799 : n40802;
  assign n40804 = pi11 ? n40767 : n40803;
  assign n40805 = pi10 ? n40804 : n32;
  assign n40806 = pi09 ? n32 : n40805;
  assign n40807 = pi14 ? n16953 : n40795;
  assign n40808 = pi15 ? n16965 : n32;
  assign n40809 = pi14 ? n16965 : n40808;
  assign n40810 = pi13 ? n40807 : n40809;
  assign n40811 = pi12 ? n40810 : n32;
  assign n40812 = pi11 ? n40767 : n40811;
  assign n40813 = pi10 ? n40812 : n32;
  assign n40814 = pi09 ? n32 : n40813;
  assign n40815 = pi08 ? n40806 : n40814;
  assign n40816 = pi14 ? n32 : n37568;
  assign n40817 = pi13 ? n32 : n40816;
  assign n40818 = pi12 ? n32 : n40817;
  assign n40819 = pi14 ? n17036 : n27858;
  assign n40820 = pi14 ? n17039 : n32;
  assign n40821 = pi13 ? n40819 : n40820;
  assign n40822 = pi12 ? n40821 : n32;
  assign n40823 = pi11 ? n40818 : n40822;
  assign n40824 = pi10 ? n40823 : n32;
  assign n40825 = pi09 ? n32 : n40824;
  assign n40826 = pi13 ? n17036 : n40820;
  assign n40827 = pi12 ? n40826 : n32;
  assign n40828 = pi11 ? n40818 : n40827;
  assign n40829 = pi10 ? n40828 : n32;
  assign n40830 = pi09 ? n32 : n40829;
  assign n40831 = pi08 ? n40825 : n40830;
  assign n40832 = pi07 ? n40815 : n40831;
  assign n40833 = pi14 ? n16914 : n25492;
  assign n40834 = pi13 ? n32 : n40833;
  assign n40835 = pi12 ? n32 : n40834;
  assign n40836 = pi14 ? n17091 : n17036;
  assign n40837 = pi14 ? n16913 : n32;
  assign n40838 = pi13 ? n40836 : n40837;
  assign n40839 = pi12 ? n40838 : n32;
  assign n40840 = pi11 ? n40835 : n40839;
  assign n40841 = pi10 ? n40840 : n32;
  assign n40842 = pi09 ? n32 : n40841;
  assign n40843 = pi14 ? n32 : n17188;
  assign n40844 = pi13 ? n32 : n40843;
  assign n40845 = pi12 ? n32 : n40844;
  assign n40846 = pi14 ? n17090 : n17133;
  assign n40847 = pi15 ? n16913 : n32;
  assign n40848 = pi14 ? n40847 : n32;
  assign n40849 = pi13 ? n40846 : n40848;
  assign n40850 = pi12 ? n40849 : n32;
  assign n40851 = pi11 ? n40845 : n40850;
  assign n40852 = pi10 ? n40851 : n32;
  assign n40853 = pi09 ? n32 : n40852;
  assign n40854 = pi08 ? n40842 : n40853;
  assign n40855 = pi14 ? n32 : n17189;
  assign n40856 = pi13 ? n32 : n40855;
  assign n40857 = pi12 ? n32 : n40856;
  assign n40858 = pi13 ? n40846 : n32;
  assign n40859 = pi12 ? n40858 : n32;
  assign n40860 = pi11 ? n40857 : n40859;
  assign n40861 = pi10 ? n40860 : n32;
  assign n40862 = pi09 ? n32 : n40861;
  assign n40863 = pi14 ? n17188 : n17100;
  assign n40864 = pi13 ? n40863 : n32;
  assign n40865 = pi12 ? n40864 : n32;
  assign n40866 = pi11 ? n32 : n40865;
  assign n40867 = pi10 ? n40866 : n32;
  assign n40868 = pi09 ? n32 : n40867;
  assign n40869 = pi08 ? n40862 : n40868;
  assign n40870 = pi07 ? n40854 : n40869;
  assign n40871 = pi06 ? n40832 : n40870;
  assign n40872 = pi05 ? n40794 : n40871;
  assign n40873 = pi04 ? n40726 : n40872;
  assign n40874 = pi03 ? n40210 : n40873;
  assign n40875 = pi14 ? n17273 : n17189;
  assign n40876 = pi13 ? n40875 : n32;
  assign n40877 = pi12 ? n40876 : n32;
  assign n40878 = pi11 ? n32 : n40877;
  assign n40879 = pi10 ? n40878 : n32;
  assign n40880 = pi09 ? n32 : n40879;
  assign n40881 = pi13 ? n40855 : n32;
  assign n40882 = pi12 ? n40881 : n32;
  assign n40883 = pi11 ? n32 : n40882;
  assign n40884 = pi10 ? n40883 : n32;
  assign n40885 = pi09 ? n32 : n40884;
  assign n40886 = pi08 ? n40880 : n40885;
  assign n40887 = pi07 ? n40886 : n40885;
  assign n40888 = pi07 ? n40885 : n32;
  assign n40889 = pi06 ? n40887 : n40888;
  assign n40890 = pi05 ? n40889 : n32;
  assign n40891 = pi04 ? n40890 : n17568;
  assign n40892 = pi03 ? n40891 : n17568;
  assign n40893 = pi02 ? n40874 : n40892;
  assign n40894 = pi06 ? n32 : n17601;
  assign n40895 = pi05 ? n17572 : n40894;
  assign n40896 = pi08 ? n17601 : n17625;
  assign n40897 = pi07 ? n40896 : n32;
  assign n40898 = pi06 ? n17601 : n40897;
  assign n40899 = pi05 ? n40898 : n32;
  assign n40900 = pi04 ? n40895 : n40899;
  assign n40901 = pi03 ? n17568 : n40900;
  assign n40902 = pi02 ? n40901 : n32;
  assign n40903 = pi01 ? n40893 : n40902;
  assign n40904 = pi00 ? n38613 : n40903;
  assign n40905 = pi14 ? n28051 : n32;
  assign n40906 = pi13 ? n32 : n40905;
  assign n40907 = pi12 ? n32 : n40906;
  assign n40908 = pi20 ? n342 : n111;
  assign n40909 = pi19 ? n9007 : n40908;
  assign n40910 = pi18 ? n40909 : n32;
  assign n40911 = pi17 ? n28031 : n40910;
  assign n40912 = pi16 ? n19171 : n40911;
  assign n40913 = pi19 ? n266 : ~n236;
  assign n40914 = pi18 ? n17118 : n40913;
  assign n40915 = pi20 ? n220 : ~n111;
  assign n40916 = pi19 ? n9007 : ~n40915;
  assign n40917 = pi18 ? n40916 : n32;
  assign n40918 = pi17 ? n40914 : n40917;
  assign n40919 = pi16 ? n19171 : n40918;
  assign n40920 = pi15 ? n40912 : n40919;
  assign n40921 = pi14 ? n28022 : n40920;
  assign n40922 = pi18 ? n2387 : ~n32;
  assign n40923 = pi17 ? n32 : n40922;
  assign n40924 = pi16 ? n40923 : ~n2144;
  assign n40925 = pi16 ? n1705 : ~n1581;
  assign n40926 = pi15 ? n40924 : n40925;
  assign n40927 = pi14 ? n40926 : n29240;
  assign n40928 = pi13 ? n40921 : n40927;
  assign n40929 = pi19 ? n17644 : ~n15751;
  assign n40930 = pi18 ? n40929 : ~n32;
  assign n40931 = pi17 ? n17643 : n40930;
  assign n40932 = pi16 ? n1214 : ~n40931;
  assign n40933 = pi15 ? n40932 : n28098;
  assign n40934 = pi14 ? n40933 : n28051;
  assign n40935 = pi20 ? n439 : n18834;
  assign n40936 = pi19 ? n40935 : n36826;
  assign n40937 = pi18 ? n4127 : ~n40936;
  assign n40938 = pi17 ? n32 : n40937;
  assign n40939 = pi20 ? n11107 : ~n7939;
  assign n40940 = pi20 ? n246 : n439;
  assign n40941 = pi19 ? n40939 : n40940;
  assign n40942 = pi20 ? n439 : ~n206;
  assign n40943 = pi19 ? n40942 : n439;
  assign n40944 = pi18 ? n40941 : n40943;
  assign n40945 = pi20 ? n439 : ~n260;
  assign n40946 = pi20 ? n6621 : n206;
  assign n40947 = pi19 ? n40945 : n40946;
  assign n40948 = pi18 ? n40947 : ~n32;
  assign n40949 = pi17 ? n40944 : n40948;
  assign n40950 = pi16 ? n40938 : ~n40949;
  assign n40951 = pi20 ? n18261 : n18408;
  assign n40952 = pi19 ? n40951 : ~n18782;
  assign n40953 = pi18 ? n28071 : ~n40952;
  assign n40954 = pi17 ? n32 : n40953;
  assign n40955 = pi21 ? n173 : ~n1939;
  assign n40956 = pi20 ? n18832 : n40955;
  assign n40957 = pi19 ? n28081 : ~n40956;
  assign n40958 = pi18 ? n40957 : ~n32;
  assign n40959 = pi17 ? n28080 : ~n40958;
  assign n40960 = pi16 ? n40954 : n40959;
  assign n40961 = pi15 ? n40950 : n40960;
  assign n40962 = pi20 ? n9488 : n40955;
  assign n40963 = pi19 ? n28092 : ~n40962;
  assign n40964 = pi18 ? n40963 : ~n32;
  assign n40965 = pi17 ? n28091 : ~n40964;
  assign n40966 = pi16 ? n28075 : n40965;
  assign n40967 = pi18 ? n268 : n9170;
  assign n40968 = pi17 ? n32 : n40967;
  assign n40969 = pi20 ? n2358 : ~n220;
  assign n40970 = pi19 ? n32 : ~n40969;
  assign n40971 = pi19 ? n23307 : n321;
  assign n40972 = pi18 ? n40970 : n40971;
  assign n40973 = pi20 ? n220 : ~n1324;
  assign n40974 = pi20 ? n18129 : n14601;
  assign n40975 = pi19 ? n40973 : n40974;
  assign n40976 = pi18 ? n40975 : n32;
  assign n40977 = pi17 ? n40972 : n40976;
  assign n40978 = pi16 ? n40968 : n40977;
  assign n40979 = pi15 ? n40966 : n40978;
  assign n40980 = pi14 ? n40961 : n40979;
  assign n40981 = pi13 ? n40934 : n40980;
  assign n40982 = pi12 ? n40928 : n40981;
  assign n40983 = pi11 ? n40907 : n40982;
  assign n40984 = pi18 ? n209 : n28362;
  assign n40985 = pi17 ? n32 : n40984;
  assign n40986 = pi19 ? n4670 : n9007;
  assign n40987 = pi19 ? n9345 : n207;
  assign n40988 = pi18 ? n40986 : ~n40987;
  assign n40989 = pi20 ? n246 : n2140;
  assign n40990 = pi19 ? n30849 : ~n40989;
  assign n40991 = pi18 ? n40990 : n32;
  assign n40992 = pi17 ? n40988 : ~n40991;
  assign n40993 = pi16 ? n40985 : ~n40992;
  assign n40994 = pi18 ? n268 : n4689;
  assign n40995 = pi17 ? n32 : n40994;
  assign n40996 = pi19 ? n17766 : n9007;
  assign n40997 = pi18 ? n29140 : n40996;
  assign n40998 = pi20 ? n342 : n7880;
  assign n40999 = pi19 ? n18390 : ~n40998;
  assign n41000 = pi18 ? n40999 : ~n32;
  assign n41001 = pi17 ? n40997 : ~n41000;
  assign n41002 = pi16 ? n40995 : n41001;
  assign n41003 = pi15 ? n41002 : n17702;
  assign n41004 = pi14 ? n40993 : n41003;
  assign n41005 = pi14 ? n28106 : n18170;
  assign n41006 = pi13 ? n41004 : n41005;
  assign n41007 = pi14 ? n17698 : n32;
  assign n41008 = pi21 ? n405 : n85;
  assign n41009 = pi20 ? n32 : n41008;
  assign n41010 = pi19 ? n32 : n41009;
  assign n41011 = pi18 ? n41010 : n32;
  assign n41012 = pi17 ? n32 : n41011;
  assign n41013 = pi16 ? n32 : n41012;
  assign n41014 = pi15 ? n17856 : n41013;
  assign n41015 = pi14 ? n32 : n41014;
  assign n41016 = pi13 ? n41007 : n41015;
  assign n41017 = pi12 ? n41006 : n41016;
  assign n41018 = pi18 ? n19082 : n32;
  assign n41019 = pi17 ? n32 : n41018;
  assign n41020 = pi16 ? n32 : n41019;
  assign n41021 = pi15 ? n41020 : n32;
  assign n41022 = pi14 ? n41021 : n32;
  assign n41023 = pi20 ? n220 : ~n12884;
  assign n41024 = pi20 ? n13171 : n17652;
  assign n41025 = pi19 ? n41023 : ~n41024;
  assign n41026 = pi18 ? n28053 : ~n41025;
  assign n41027 = pi17 ? n32 : n41026;
  assign n41028 = pi20 ? n310 : ~n220;
  assign n41029 = pi19 ? n41028 : n32;
  assign n41030 = pi19 ? n32 : n17649;
  assign n41031 = pi18 ? n41029 : n41030;
  assign n41032 = pi17 ? n41031 : n32;
  assign n41033 = pi16 ? n41027 : n41032;
  assign n41034 = pi15 ? n32 : n41033;
  assign n41035 = pi18 ? n28178 : ~n28141;
  assign n41036 = pi17 ? n32 : n41035;
  assign n41037 = pi19 ? n9037 : ~n9345;
  assign n41038 = pi18 ? n41037 : n32;
  assign n41039 = pi17 ? n28147 : n41038;
  assign n41040 = pi16 ? n41036 : n41039;
  assign n41041 = pi19 ? n41023 : n22698;
  assign n41042 = pi18 ? n28178 : ~n41041;
  assign n41043 = pi17 ? n32 : n41042;
  assign n41044 = pi20 ? n266 : ~n357;
  assign n41045 = pi19 ? n9037 : ~n41044;
  assign n41046 = pi18 ? n41045 : n32;
  assign n41047 = pi17 ? n28147 : n41046;
  assign n41048 = pi16 ? n41043 : n41047;
  assign n41049 = pi15 ? n41040 : n41048;
  assign n41050 = pi14 ? n41034 : n41049;
  assign n41051 = pi13 ? n41022 : n41050;
  assign n41052 = pi19 ? n1464 : n5004;
  assign n41053 = pi18 ? n1613 : ~n41052;
  assign n41054 = pi17 ? n32 : n41053;
  assign n41055 = pi19 ? n28041 : ~n32;
  assign n41056 = pi18 ? n41055 : ~n16234;
  assign n41057 = pi18 ? n8203 : ~n32;
  assign n41058 = pi17 ? n41056 : ~n41057;
  assign n41059 = pi16 ? n41054 : n41058;
  assign n41060 = pi15 ? n29780 : n41059;
  assign n41061 = pi18 ? n366 : ~n20020;
  assign n41062 = pi17 ? n32 : n41061;
  assign n41063 = pi16 ? n41062 : ~n1214;
  assign n41064 = pi17 ? n17743 : n1697;
  assign n41065 = pi16 ? n41062 : ~n41064;
  assign n41066 = pi15 ? n41063 : n41065;
  assign n41067 = pi14 ? n41060 : n41066;
  assign n41068 = pi19 ? n22185 : ~n9822;
  assign n41069 = pi18 ? n940 : n41068;
  assign n41070 = pi17 ? n32 : n41069;
  assign n41071 = pi19 ? n9345 : ~n349;
  assign n41072 = pi19 ? n17749 : n33796;
  assign n41073 = pi18 ? n41071 : n41072;
  assign n41074 = pi19 ? n28134 : ~n6298;
  assign n41075 = pi18 ? n41074 : n32;
  assign n41076 = pi17 ? n41073 : n41075;
  assign n41077 = pi16 ? n41070 : n41076;
  assign n41078 = pi19 ? n221 : n21349;
  assign n41079 = pi18 ? n41078 : ~n32;
  assign n41080 = pi17 ? n17759 : n41079;
  assign n41081 = pi16 ? n1214 : ~n41080;
  assign n41082 = pi15 ? n41077 : n41081;
  assign n41083 = pi20 ? n1331 : n785;
  assign n41084 = pi20 ? n206 : n357;
  assign n41085 = pi19 ? n41083 : n41084;
  assign n41086 = pi18 ? n209 : ~n41085;
  assign n41087 = pi17 ? n32 : n41086;
  assign n41088 = pi19 ? n34314 : ~n17766;
  assign n41089 = pi18 ? n41088 : ~n28185;
  assign n41090 = pi17 ? n41089 : ~n28188;
  assign n41091 = pi16 ? n41087 : n41090;
  assign n41092 = pi17 ? n17768 : n1213;
  assign n41093 = pi16 ? n1214 : ~n41092;
  assign n41094 = pi15 ? n41091 : n41093;
  assign n41095 = pi14 ? n41082 : n41094;
  assign n41096 = pi13 ? n41067 : n41095;
  assign n41097 = pi12 ? n41051 : n41096;
  assign n41098 = pi11 ? n41017 : n41097;
  assign n41099 = pi10 ? n40983 : n41098;
  assign n41100 = pi09 ? n32 : n41099;
  assign n41101 = pi14 ? n17637 : n32;
  assign n41102 = pi13 ? n32 : n41101;
  assign n41103 = pi12 ? n32 : n41102;
  assign n41104 = pi15 ? n17813 : n32;
  assign n41105 = pi19 ? n9007 : n34159;
  assign n41106 = pi18 ? n41105 : n32;
  assign n41107 = pi17 ? n28031 : n41106;
  assign n41108 = pi16 ? n19171 : n41107;
  assign n41109 = pi20 ? n220 : ~n175;
  assign n41110 = pi19 ? n9007 : ~n41109;
  assign n41111 = pi18 ? n41110 : n32;
  assign n41112 = pi17 ? n40914 : n41111;
  assign n41113 = pi16 ? n19171 : n41112;
  assign n41114 = pi15 ? n41108 : n41113;
  assign n41115 = pi14 ? n41104 : n41114;
  assign n41116 = pi19 ? n32 : n30521;
  assign n41117 = pi18 ? n41116 : ~n32;
  assign n41118 = pi17 ? n32 : n41117;
  assign n41119 = pi16 ? n41118 : ~n1577;
  assign n41120 = pi16 ? n1705 : ~n1577;
  assign n41121 = pi15 ? n41119 : n41120;
  assign n41122 = pi16 ? n1214 : ~n1577;
  assign n41123 = pi16 ? n1214 : ~n18985;
  assign n41124 = pi15 ? n41122 : n41123;
  assign n41125 = pi14 ? n41121 : n41124;
  assign n41126 = pi13 ? n41115 : n41125;
  assign n41127 = pi16 ? n18561 : n17812;
  assign n41128 = pi15 ? n40932 : n41127;
  assign n41129 = pi14 ? n41128 : n17813;
  assign n41130 = pi20 ? n274 : n17671;
  assign n41131 = pi19 ? n41130 : n28481;
  assign n41132 = pi18 ? n37954 : ~n41131;
  assign n41133 = pi17 ? n32 : n41132;
  assign n41134 = pi20 ? n1331 : ~n18173;
  assign n41135 = pi20 ? n3523 : n274;
  assign n41136 = pi19 ? n41134 : n41135;
  assign n41137 = pi20 ? n274 : ~n785;
  assign n41138 = pi19 ? n41137 : n274;
  assign n41139 = pi18 ? n41136 : n41138;
  assign n41140 = pi20 ? n274 : ~n260;
  assign n41141 = pi20 ? n18129 : n2385;
  assign n41142 = pi19 ? n41140 : n41141;
  assign n41143 = pi18 ? n41142 : ~n32;
  assign n41144 = pi17 ? n41139 : n41143;
  assign n41145 = pi16 ? n41133 : ~n41144;
  assign n41146 = pi20 ? n7939 : n18173;
  assign n41147 = pi19 ? n41146 : ~n28243;
  assign n41148 = pi18 ? n19082 : ~n41147;
  assign n41149 = pi17 ? n32 : n41148;
  assign n41150 = pi20 ? n9491 : n3695;
  assign n41151 = pi19 ? n18621 : ~n41150;
  assign n41152 = pi18 ? n41151 : ~n32;
  assign n41153 = pi17 ? n28251 : ~n41152;
  assign n41154 = pi16 ? n41149 : n41153;
  assign n41155 = pi15 ? n41145 : n41154;
  assign n41156 = pi21 ? n173 : ~n14513;
  assign n41157 = pi20 ? n9488 : n41156;
  assign n41158 = pi19 ? n28092 : ~n41157;
  assign n41159 = pi18 ? n41158 : ~n32;
  assign n41160 = pi17 ? n28091 : ~n41159;
  assign n41161 = pi16 ? n28075 : n41160;
  assign n41162 = pi20 ? n18129 : n10878;
  assign n41163 = pi19 ? n40973 : n41162;
  assign n41164 = pi18 ? n41163 : n32;
  assign n41165 = pi17 ? n40972 : n41164;
  assign n41166 = pi16 ? n40968 : n41165;
  assign n41167 = pi15 ? n41161 : n41166;
  assign n41168 = pi14 ? n41155 : n41167;
  assign n41169 = pi13 ? n41129 : n41168;
  assign n41170 = pi12 ? n41126 : n41169;
  assign n41171 = pi11 ? n41103 : n41170;
  assign n41172 = pi19 ? n30849 : ~n22106;
  assign n41173 = pi18 ? n41172 : n32;
  assign n41174 = pi17 ? n40988 : ~n41173;
  assign n41175 = pi16 ? n40985 : ~n41174;
  assign n41176 = pi19 ? n18390 : ~n18396;
  assign n41177 = pi18 ? n41176 : ~n32;
  assign n41178 = pi17 ? n40997 : ~n41177;
  assign n41179 = pi16 ? n40995 : n41178;
  assign n41180 = pi15 ? n41179 : n18326;
  assign n41181 = pi14 ? n41175 : n41180;
  assign n41182 = pi15 ? n17825 : n17822;
  assign n41183 = pi14 ? n28269 : n41182;
  assign n41184 = pi13 ? n41181 : n41183;
  assign n41185 = pi15 ? n17822 : n32;
  assign n41186 = pi14 ? n41185 : n32;
  assign n41187 = pi14 ? n32 : n17851;
  assign n41188 = pi13 ? n41186 : n41187;
  assign n41189 = pi12 ? n41184 : n41188;
  assign n41190 = pi15 ? n32 : n17856;
  assign n41191 = pi14 ? n32 : n41190;
  assign n41192 = pi21 ? n10182 : n174;
  assign n41193 = pi20 ? n32 : n41192;
  assign n41194 = pi19 ? n32 : n41193;
  assign n41195 = pi18 ? n41194 : ~n41025;
  assign n41196 = pi17 ? n32 : n41195;
  assign n41197 = pi16 ? n41196 : n41032;
  assign n41198 = pi15 ? n32 : n41197;
  assign n41199 = pi20 ? n32 : n17140;
  assign n41200 = pi19 ? n32 : n41199;
  assign n41201 = pi18 ? n41200 : ~n28141;
  assign n41202 = pi17 ? n32 : n41201;
  assign n41203 = pi16 ? n41202 : n41039;
  assign n41204 = pi15 ? n41203 : n41048;
  assign n41205 = pi14 ? n41198 : n41204;
  assign n41206 = pi13 ? n41191 : n41205;
  assign n41207 = pi18 ? n341 : ~n20020;
  assign n41208 = pi17 ? n32 : n41207;
  assign n41209 = pi16 ? n41208 : ~n1214;
  assign n41210 = pi15 ? n41209 : n41065;
  assign n41211 = pi14 ? n41060 : n41210;
  assign n41212 = pi18 ? n29325 : n41068;
  assign n41213 = pi17 ? n32 : n41212;
  assign n41214 = pi16 ? n41213 : n41076;
  assign n41215 = pi16 ? n19652 : ~n41080;
  assign n41216 = pi15 ? n41214 : n41215;
  assign n41217 = pi16 ? n28182 : n41090;
  assign n41218 = pi17 ? n17768 : n1971;
  assign n41219 = pi16 ? n19652 : ~n41218;
  assign n41220 = pi15 ? n41217 : n41219;
  assign n41221 = pi14 ? n41216 : n41220;
  assign n41222 = pi13 ? n41211 : n41221;
  assign n41223 = pi12 ? n41206 : n41222;
  assign n41224 = pi11 ? n41189 : n41223;
  assign n41225 = pi10 ? n41171 : n41224;
  assign n41226 = pi09 ? n32 : n41225;
  assign n41227 = pi08 ? n41100 : n41226;
  assign n41228 = pi07 ? n32 : n41227;
  assign n41229 = pi06 ? n32 : n41228;
  assign n41230 = pi14 ? n17885 : n32;
  assign n41231 = pi13 ? n32 : n41230;
  assign n41232 = pi12 ? n32 : n41231;
  assign n41233 = pi20 ? n9491 : n9194;
  assign n41234 = pi19 ? n41233 : n18404;
  assign n41235 = pi18 ? n863 : n41234;
  assign n41236 = pi17 ? n32 : n41235;
  assign n41237 = pi20 ? n18253 : n820;
  assign n41238 = pi19 ? n18409 : ~n41237;
  assign n41239 = pi20 ? n820 : ~n3843;
  assign n41240 = pi20 ? n18832 : ~n333;
  assign n41241 = pi19 ? n41239 : n41240;
  assign n41242 = pi18 ? n41238 : ~n41241;
  assign n41243 = pi21 ? n173 : ~n6898;
  assign n41244 = pi20 ? n2019 : n41243;
  assign n41245 = pi19 ? n5614 : n41244;
  assign n41246 = pi18 ? n41245 : ~n32;
  assign n41247 = pi17 ? n41242 : n41246;
  assign n41248 = pi16 ? n41236 : ~n41247;
  assign n41249 = pi15 ? n17876 : n41248;
  assign n41250 = pi18 ? n1862 : n28073;
  assign n41251 = pi17 ? n32 : n41250;
  assign n41252 = pi19 ? n18404 : ~n41237;
  assign n41253 = pi18 ? n41252 : ~n41241;
  assign n41254 = pi21 ? n173 : n9326;
  assign n41255 = pi20 ? n448 : n41254;
  assign n41256 = pi19 ? n5614 : n41255;
  assign n41257 = pi18 ? n41256 : ~n32;
  assign n41258 = pi17 ? n41253 : n41257;
  assign n41259 = pi16 ? n41251 : ~n41258;
  assign n41260 = pi20 ? n820 : ~n310;
  assign n41261 = pi19 ? n41260 : n41240;
  assign n41262 = pi18 ? n41252 : ~n41261;
  assign n41263 = pi20 ? n501 : ~n41254;
  assign n41264 = pi19 ? n5614 : ~n41263;
  assign n41265 = pi18 ? n41264 : ~n32;
  assign n41266 = pi17 ? n41262 : n41265;
  assign n41267 = pi16 ? n41251 : ~n41266;
  assign n41268 = pi15 ? n41259 : n41267;
  assign n41269 = pi14 ? n41249 : n41268;
  assign n41270 = pi17 ? n32 : n5671;
  assign n41271 = pi16 ? n1471 : ~n41270;
  assign n41272 = pi16 ? n1214 : ~n1834;
  assign n41273 = pi15 ? n41271 : n41272;
  assign n41274 = pi18 ? n209 : ~n4671;
  assign n41275 = pi17 ? n32 : n41274;
  assign n41276 = pi19 ? n247 : n342;
  assign n41277 = pi18 ? n29140 : n41276;
  assign n41278 = pi18 ? n41105 : ~n32;
  assign n41279 = pi17 ? n41277 : n41278;
  assign n41280 = pi16 ? n41275 : ~n41279;
  assign n41281 = pi15 ? n30304 : n41280;
  assign n41282 = pi14 ? n41273 : n41281;
  assign n41283 = pi13 ? n41269 : n41282;
  assign n41284 = pi20 ? n32 : n18255;
  assign n41285 = pi19 ? n32 : n41284;
  assign n41286 = pi19 ? n18282 : n28058;
  assign n41287 = pi18 ? n41285 : ~n41286;
  assign n41288 = pi17 ? n32 : n41287;
  assign n41289 = pi20 ? n6822 : n17652;
  assign n41290 = pi19 ? n18778 : ~n41289;
  assign n41291 = pi20 ? n17652 : n6822;
  assign n41292 = pi19 ? n41291 : n18282;
  assign n41293 = pi18 ? n41290 : ~n41292;
  assign n41294 = pi20 ? n18253 : n18415;
  assign n41295 = pi19 ? n29877 : ~n41294;
  assign n41296 = pi18 ? n41295 : ~n32;
  assign n41297 = pi17 ? n41293 : ~n41296;
  assign n41298 = pi16 ? n41288 : n41297;
  assign n41299 = pi15 ? n29240 : n41298;
  assign n41300 = pi20 ? n18415 : n17652;
  assign n41301 = pi19 ? n41300 : n18253;
  assign n41302 = pi18 ? n28060 : ~n41301;
  assign n41303 = pi20 ? n18415 : n310;
  assign n41304 = pi20 ? n9491 : n18073;
  assign n41305 = pi19 ? n41303 : ~n41304;
  assign n41306 = pi18 ? n41305 : ~n32;
  assign n41307 = pi17 ? n41302 : ~n41306;
  assign n41308 = pi16 ? n28057 : n41307;
  assign n41309 = pi15 ? n41308 : n28349;
  assign n41310 = pi14 ? n41299 : n41309;
  assign n41311 = pi20 ? n357 : n1817;
  assign n41312 = pi19 ? n32 : n41311;
  assign n41313 = pi20 ? n175 : ~n354;
  assign n41314 = pi19 ? n3495 : n41313;
  assign n41315 = pi18 ? n41312 : n41314;
  assign n41316 = pi19 ? n4476 : ~n1574;
  assign n41317 = pi18 ? n41316 : n32;
  assign n41318 = pi17 ? n41315 : ~n41317;
  assign n41319 = pi16 ? n1214 : ~n41318;
  assign n41320 = pi20 ? n32 : n29457;
  assign n41321 = pi19 ? n32 : n41320;
  assign n41322 = pi19 ? n18129 : ~n18246;
  assign n41323 = pi18 ? n41321 : ~n41322;
  assign n41324 = pi17 ? n32 : n41323;
  assign n41325 = pi20 ? n6303 : n9194;
  assign n41326 = pi20 ? n1368 : n1817;
  assign n41327 = pi19 ? n41325 : n41326;
  assign n41328 = pi20 ? n1817 : n1368;
  assign n41329 = pi19 ? n41328 : n1331;
  assign n41330 = pi18 ? n41327 : n41329;
  assign n41331 = pi20 ? n274 : n23668;
  assign n41332 = pi19 ? n3495 : n41331;
  assign n41333 = pi18 ? n41332 : ~n32;
  assign n41334 = pi17 ? n41330 : n41333;
  assign n41335 = pi16 ? n41324 : ~n41334;
  assign n41336 = pi15 ? n41319 : n41335;
  assign n41337 = pi19 ? n28365 : n30044;
  assign n41338 = pi18 ? n41321 : n41337;
  assign n41339 = pi17 ? n32 : n41338;
  assign n41340 = pi20 ? n29457 : n17652;
  assign n41341 = pi19 ? n36181 : ~n41340;
  assign n41342 = pi20 ? n5854 : ~n9194;
  assign n41343 = pi19 ? n41342 : n17652;
  assign n41344 = pi18 ? n41341 : ~n41343;
  assign n41345 = pi20 ? n17652 : n20501;
  assign n41346 = pi19 ? n28140 : ~n41345;
  assign n41347 = pi18 ? n41346 : n32;
  assign n41348 = pi17 ? n41344 : ~n41347;
  assign n41349 = pi16 ? n41339 : ~n41348;
  assign n41350 = pi15 ? n41349 : n41122;
  assign n41351 = pi14 ? n41336 : n41350;
  assign n41352 = pi13 ? n41310 : n41351;
  assign n41353 = pi12 ? n41283 : n41352;
  assign n41354 = pi11 ? n41232 : n41353;
  assign n41355 = pi18 ? n268 : n248;
  assign n41356 = pi17 ? n32 : n41355;
  assign n41357 = pi19 ? n32 : ~n5004;
  assign n41358 = pi19 ? n18211 : n321;
  assign n41359 = pi18 ? n41357 : n41358;
  assign n41360 = pi19 ? n18396 : n247;
  assign n41361 = pi18 ? n41360 : ~n32;
  assign n41362 = pi17 ? n41359 : ~n41361;
  assign n41363 = pi16 ? n41356 : n41362;
  assign n41364 = pi19 ? n32 : ~n4964;
  assign n41365 = pi18 ? n41364 : n36115;
  assign n41366 = pi19 ? n4342 : n1464;
  assign n41367 = pi18 ? n41366 : ~n32;
  assign n41368 = pi17 ? n41365 : ~n41367;
  assign n41369 = pi16 ? n32 : n41368;
  assign n41370 = pi15 ? n41363 : n41369;
  assign n41371 = pi19 ? n17766 : n321;
  assign n41372 = pi18 ? n29140 : n41371;
  assign n41373 = pi19 ? n4342 : ~n23688;
  assign n41374 = pi18 ? n41373 : ~n32;
  assign n41375 = pi17 ? n41372 : ~n41374;
  assign n41376 = pi16 ? n32 : n41375;
  assign n41377 = pi15 ? n41376 : n28385;
  assign n41378 = pi14 ? n41370 : n41377;
  assign n41379 = pi19 ? n11374 : n17685;
  assign n41380 = pi18 ? n41379 : n32;
  assign n41381 = pi17 ? n3282 : n41380;
  assign n41382 = pi16 ? n32 : n41381;
  assign n41383 = pi15 ? n32 : n41382;
  assign n41384 = pi14 ? n17903 : n41383;
  assign n41385 = pi13 ? n41378 : n41384;
  assign n41386 = pi15 ? n17910 : n32;
  assign n41387 = pi14 ? n41386 : n32;
  assign n41388 = pi13 ? n41387 : n32;
  assign n41389 = pi12 ? n41385 : n41388;
  assign n41390 = pi18 ? n341 : ~n248;
  assign n41391 = pi17 ? n32 : n41390;
  assign n41392 = pi17 ? n28422 : n1227;
  assign n41393 = pi16 ? n41391 : ~n41392;
  assign n41394 = pi15 ? n32 : n41393;
  assign n41395 = pi19 ? n208 : ~n17194;
  assign n41396 = pi18 ? n41395 : ~n32;
  assign n41397 = pi17 ? n28428 : n41396;
  assign n41398 = pi16 ? n1233 : ~n41397;
  assign n41399 = pi18 ? n366 : ~n6145;
  assign n41400 = pi17 ? n32 : n41399;
  assign n41401 = pi16 ? n41400 : ~n1135;
  assign n41402 = pi15 ? n41398 : n41401;
  assign n41403 = pi14 ? n41394 : n41402;
  assign n41404 = pi13 ? n32 : n41403;
  assign n41405 = pi16 ? n1135 : ~n4729;
  assign n41406 = pi18 ? n341 : ~n34006;
  assign n41407 = pi17 ? n32 : n41406;
  assign n41408 = pi16 ? n41407 : ~n4060;
  assign n41409 = pi15 ? n41405 : n41408;
  assign n41410 = pi17 ? n17951 : n1978;
  assign n41411 = pi16 ? n1135 : ~n41410;
  assign n41412 = pi18 ? n6071 : n248;
  assign n41413 = pi19 ? n322 : n207;
  assign n41414 = pi18 ? n41413 : ~n32;
  assign n41415 = pi17 ? n41412 : n41414;
  assign n41416 = pi16 ? n1135 : ~n41415;
  assign n41417 = pi15 ? n41411 : n41416;
  assign n41418 = pi14 ? n41409 : n41417;
  assign n41419 = pi20 ? n175 : n246;
  assign n41420 = pi19 ? n41419 : ~n207;
  assign n41421 = pi18 ? n18710 : ~n41420;
  assign n41422 = pi17 ? n32 : n41421;
  assign n41423 = pi19 ? n4406 : n28184;
  assign n41424 = pi18 ? n38793 : ~n41423;
  assign n41425 = pi19 ? n322 : ~n5004;
  assign n41426 = pi18 ? n41425 : ~n32;
  assign n41427 = pi17 ? n41424 : n41426;
  assign n41428 = pi16 ? n41422 : ~n41427;
  assign n41429 = pi19 ? n208 : ~n5004;
  assign n41430 = pi18 ? n41429 : ~n32;
  assign n41431 = pi17 ? n32 : n41430;
  assign n41432 = pi16 ? n1233 : ~n41431;
  assign n41433 = pi15 ? n41428 : n41432;
  assign n41434 = pi17 ? n17976 : n28453;
  assign n41435 = pi16 ? n28449 : ~n41434;
  assign n41436 = pi19 ? n1818 : n208;
  assign n41437 = pi18 ? n41436 : ~n32;
  assign n41438 = pi17 ? n32 : n41437;
  assign n41439 = pi16 ? n1233 : ~n41438;
  assign n41440 = pi15 ? n41435 : n41439;
  assign n41441 = pi14 ? n41433 : n41440;
  assign n41442 = pi13 ? n41418 : n41441;
  assign n41443 = pi12 ? n41404 : n41442;
  assign n41444 = pi11 ? n41389 : n41443;
  assign n41445 = pi10 ? n41354 : n41444;
  assign n41446 = pi09 ? n32 : n41445;
  assign n41447 = pi20 ? n32 : n17159;
  assign n41448 = pi19 ? n32 : n41447;
  assign n41449 = pi18 ? n41448 : ~n32;
  assign n41450 = pi17 ? n32 : n41449;
  assign n41451 = pi16 ? n41450 : ~n1683;
  assign n41452 = pi15 ? n32 : n41451;
  assign n41453 = pi21 ? n10182 : ~n309;
  assign n41454 = pi20 ? n32 : n41453;
  assign n41455 = pi19 ? n32 : n41454;
  assign n41456 = pi18 ? n41455 : ~n41131;
  assign n41457 = pi17 ? n32 : n41456;
  assign n41458 = pi20 ? n274 : n3523;
  assign n41459 = pi19 ? n41458 : n274;
  assign n41460 = pi18 ? n41136 : n41459;
  assign n41461 = pi19 ? n5614 : n20933;
  assign n41462 = pi18 ? n41461 : ~n32;
  assign n41463 = pi17 ? n41460 : n41462;
  assign n41464 = pi16 ? n41457 : ~n41463;
  assign n41465 = pi18 ? n41116 : ~n41131;
  assign n41466 = pi17 ? n32 : n41465;
  assign n41467 = pi19 ? n21107 : n274;
  assign n41468 = pi18 ? n41136 : n41467;
  assign n41469 = pi19 ? n5614 : ~n18333;
  assign n41470 = pi18 ? n41469 : ~n32;
  assign n41471 = pi17 ? n41468 : n41470;
  assign n41472 = pi16 ? n41466 : ~n41471;
  assign n41473 = pi15 ? n41464 : n41472;
  assign n41474 = pi14 ? n41452 : n41473;
  assign n41475 = pi19 ? n507 : n857;
  assign n41476 = pi18 ? n41475 : n1676;
  assign n41477 = pi17 ? n32 : n41476;
  assign n41478 = pi16 ? n1471 : ~n41477;
  assign n41479 = pi16 ? n1214 : ~n1678;
  assign n41480 = pi15 ? n41478 : n41479;
  assign n41481 = pi16 ? n1214 : ~n3356;
  assign n41482 = pi18 ? n41105 : n618;
  assign n41483 = pi17 ? n41277 : n41482;
  assign n41484 = pi16 ? n41275 : ~n41483;
  assign n41485 = pi15 ? n41481 : n41484;
  assign n41486 = pi14 ? n41480 : n41485;
  assign n41487 = pi13 ? n41474 : n41486;
  assign n41488 = pi18 ? n863 : n618;
  assign n41489 = pi17 ? n32 : n41488;
  assign n41490 = pi16 ? n1214 : ~n41489;
  assign n41491 = pi18 ? n41285 : n18779;
  assign n41492 = pi17 ? n32 : n41491;
  assign n41493 = pi20 ? n18408 : n9488;
  assign n41494 = pi19 ? n18782 : n41493;
  assign n41495 = pi20 ? n9488 : ~n29457;
  assign n41496 = pi20 ? n9488 : ~n17652;
  assign n41497 = pi19 ? n41495 : n41496;
  assign n41498 = pi18 ? n41494 : n41497;
  assign n41499 = pi20 ? n2180 : n17652;
  assign n41500 = pi19 ? n29877 : ~n41499;
  assign n41501 = pi18 ? n41500 : n618;
  assign n41502 = pi17 ? n41498 : ~n41501;
  assign n41503 = pi16 ? n41492 : n41502;
  assign n41504 = pi15 ? n41490 : n41503;
  assign n41505 = pi18 ? n28053 : n28478;
  assign n41506 = pi17 ? n32 : n41505;
  assign n41507 = pi19 ? n28481 : n18129;
  assign n41508 = pi20 ? n1331 : ~n314;
  assign n41509 = pi19 ? n29912 : n41508;
  assign n41510 = pi18 ? n41507 : n41509;
  assign n41511 = pi20 ? n1076 : n9641;
  assign n41512 = pi19 ? n41303 : ~n41511;
  assign n41513 = pi18 ? n41512 : ~n32;
  assign n41514 = pi17 ? n41510 : ~n41513;
  assign n41515 = pi16 ? n41506 : n41514;
  assign n41516 = pi15 ? n41515 : n28349;
  assign n41517 = pi14 ? n41504 : n41516;
  assign n41518 = pi19 ? n4476 : ~n32;
  assign n41519 = pi18 ? n41518 : n32;
  assign n41520 = pi17 ? n41315 : ~n41519;
  assign n41521 = pi16 ? n1214 : ~n41520;
  assign n41522 = pi19 ? n3495 : n274;
  assign n41523 = pi18 ? n41522 : ~n32;
  assign n41524 = pi17 ? n41330 : n41523;
  assign n41525 = pi16 ? n41324 : ~n41524;
  assign n41526 = pi15 ? n41521 : n41525;
  assign n41527 = pi19 ? n28140 : ~n31309;
  assign n41528 = pi18 ? n41527 : n32;
  assign n41529 = pi17 ? n41344 : ~n41528;
  assign n41530 = pi16 ? n41339 : ~n41529;
  assign n41531 = pi15 ? n41530 : n30304;
  assign n41532 = pi14 ? n41526 : n41531;
  assign n41533 = pi13 ? n41517 : n41532;
  assign n41534 = pi12 ? n41487 : n41533;
  assign n41535 = pi11 ? n41232 : n41534;
  assign n41536 = pi18 ? n41360 : n1676;
  assign n41537 = pi17 ? n41359 : ~n41536;
  assign n41538 = pi16 ? n41356 : n41537;
  assign n41539 = pi18 ? n41366 : n1676;
  assign n41540 = pi17 ? n41365 : ~n41539;
  assign n41541 = pi16 ? n32 : n41540;
  assign n41542 = pi15 ? n41538 : n41541;
  assign n41543 = pi18 ? n41373 : n1676;
  assign n41544 = pi17 ? n41372 : ~n41543;
  assign n41545 = pi16 ? n32 : n41544;
  assign n41546 = pi15 ? n41545 : n28516;
  assign n41547 = pi14 ? n41542 : n41546;
  assign n41548 = pi19 ? n11374 : n507;
  assign n41549 = pi18 ? n41548 : n32;
  assign n41550 = pi17 ? n3282 : n41549;
  assign n41551 = pi16 ? n32 : n41550;
  assign n41552 = pi15 ? n32 : n41551;
  assign n41553 = pi14 ? n17891 : n41552;
  assign n41554 = pi13 ? n41547 : n41553;
  assign n41555 = pi14 ? n18005 : n32;
  assign n41556 = pi13 ? n41555 : n32;
  assign n41557 = pi12 ? n41554 : n41556;
  assign n41558 = pi19 ? n208 : ~n9007;
  assign n41559 = pi18 ? n41558 : ~n32;
  assign n41560 = pi17 ? n28428 : n41559;
  assign n41561 = pi16 ? n1135 : ~n41560;
  assign n41562 = pi16 ? n28949 : ~n1135;
  assign n41563 = pi15 ? n41561 : n41562;
  assign n41564 = pi14 ? n41394 : n41563;
  assign n41565 = pi13 ? n32 : n41564;
  assign n41566 = pi20 ? n32 : ~n86;
  assign n41567 = pi19 ? n32 : n41566;
  assign n41568 = pi18 ? n41567 : ~n32;
  assign n41569 = pi17 ? n32 : n41568;
  assign n41570 = pi16 ? n1233 : ~n41569;
  assign n41571 = pi18 ? n366 : ~n34006;
  assign n41572 = pi17 ? n32 : n41571;
  assign n41573 = pi20 ? n321 : ~n86;
  assign n41574 = pi19 ? n594 : n41573;
  assign n41575 = pi18 ? n41574 : ~n32;
  assign n41576 = pi17 ? n32 : n41575;
  assign n41577 = pi16 ? n41572 : ~n41576;
  assign n41578 = pi15 ? n41570 : n41577;
  assign n41579 = pi16 ? n1233 : ~n41410;
  assign n41580 = pi16 ? n1233 : ~n41415;
  assign n41581 = pi15 ? n41579 : n41580;
  assign n41582 = pi14 ? n41578 : n41581;
  assign n41583 = pi19 ? n32 : n22154;
  assign n41584 = pi18 ? n41583 : ~n41423;
  assign n41585 = pi17 ? n41584 : n41426;
  assign n41586 = pi16 ? n41422 : ~n41585;
  assign n41587 = pi16 ? n1135 : ~n41431;
  assign n41588 = pi15 ? n41586 : n41587;
  assign n41589 = pi17 ? n32234 : n28550;
  assign n41590 = pi16 ? n28449 : ~n41589;
  assign n41591 = pi15 ? n41590 : n29780;
  assign n41592 = pi14 ? n41588 : n41591;
  assign n41593 = pi13 ? n41582 : n41592;
  assign n41594 = pi12 ? n41565 : n41593;
  assign n41595 = pi11 ? n41557 : n41594;
  assign n41596 = pi10 ? n41535 : n41595;
  assign n41597 = pi09 ? n32 : n41596;
  assign n41598 = pi08 ? n41446 : n41597;
  assign n41599 = pi14 ? n32 : n18008;
  assign n41600 = pi13 ? n32 : n41599;
  assign n41601 = pi12 ? n32 : n41600;
  assign n41602 = pi18 ? n18391 : n618;
  assign n41603 = pi17 ? n18389 : ~n41602;
  assign n41604 = pi16 ? n18109 : n41603;
  assign n41605 = pi15 ? n18008 : n41604;
  assign n41606 = pi19 ? n4670 : ~n18502;
  assign n41607 = pi18 ? n863 : n41606;
  assign n41608 = pi17 ? n32 : n41607;
  assign n41609 = pi19 ? n18678 : n1490;
  assign n41610 = pi19 ? n9822 : n7089;
  assign n41611 = pi18 ? n41609 : n41610;
  assign n41612 = pi19 ? n9345 : ~n18390;
  assign n41613 = pi18 ? n41612 : ~n32;
  assign n41614 = pi17 ? n41611 : ~n41613;
  assign n41615 = pi16 ? n41608 : n41614;
  assign n41616 = pi16 ? n29327 : ~n1678;
  assign n41617 = pi15 ? n41615 : n41616;
  assign n41618 = pi14 ? n41605 : n41617;
  assign n41619 = pi16 ? n1471 : ~n1678;
  assign n41620 = pi15 ? n41619 : n41479;
  assign n41621 = pi16 ? n1214 : ~n3352;
  assign n41622 = pi17 ? n32 : n6394;
  assign n41623 = pi18 ? n18088 : n3350;
  assign n41624 = pi17 ? n18087 : n41623;
  assign n41625 = pi16 ? n41622 : ~n41624;
  assign n41626 = pi15 ? n41621 : n41625;
  assign n41627 = pi14 ? n41620 : n41626;
  assign n41628 = pi13 ? n41618 : n41627;
  assign n41629 = pi18 ? n19350 : n18096;
  assign n41630 = pi17 ? n32 : n41629;
  assign n41631 = pi18 ? n18102 : n32;
  assign n41632 = pi17 ? n18101 : ~n41631;
  assign n41633 = pi16 ? n41630 : ~n41632;
  assign n41634 = pi20 ? n309 : n1611;
  assign n41635 = pi19 ? n41634 : n18095;
  assign n41636 = pi18 ? n19350 : n41635;
  assign n41637 = pi17 ? n32 : n41636;
  assign n41638 = pi20 ? n7942 : n9491;
  assign n41639 = pi19 ? n18099 : n41638;
  assign n41640 = pi20 ? n9491 : n12884;
  assign n41641 = pi20 ? n6085 : ~n6050;
  assign n41642 = pi19 ? n41640 : n41641;
  assign n41643 = pi18 ? n41639 : n41642;
  assign n41644 = pi20 ? n206 : ~n18415;
  assign n41645 = pi19 ? n41644 : ~n11107;
  assign n41646 = pi18 ? n41645 : ~n32;
  assign n41647 = pi17 ? n41643 : ~n41646;
  assign n41648 = pi16 ? n41637 : n41647;
  assign n41649 = pi15 ? n41633 : n41648;
  assign n41650 = pi18 ? n19082 : n248;
  assign n41651 = pi17 ? n32 : n41650;
  assign n41652 = pi19 ? n32 : n18113;
  assign n41653 = pi19 ? n17649 : n9007;
  assign n41654 = pi18 ? n41652 : n41653;
  assign n41655 = pi20 ? n32 : ~n17669;
  assign n41656 = pi19 ? n41655 : ~n428;
  assign n41657 = pi18 ? n41656 : n3350;
  assign n41658 = pi17 ? n41654 : ~n41657;
  assign n41659 = pi16 ? n41651 : n41658;
  assign n41660 = pi15 ? n32 : n41659;
  assign n41661 = pi14 ? n41649 : n41660;
  assign n41662 = pi17 ? n36573 : n2123;
  assign n41663 = pi16 ? n1214 : ~n41662;
  assign n41664 = pi19 ? n246 : n4670;
  assign n41665 = pi18 ? n32 : n41664;
  assign n41666 = pi17 ? n32 : n41665;
  assign n41667 = pi19 ? n267 : n246;
  assign n41668 = pi18 ? n33239 : ~n41667;
  assign n41669 = pi18 ? n36402 : ~n618;
  assign n41670 = pi17 ? n41668 : ~n41669;
  assign n41671 = pi16 ? n41666 : ~n41670;
  assign n41672 = pi15 ? n41663 : n41671;
  assign n41673 = pi18 ? n18397 : n618;
  assign n41674 = pi17 ? n18395 : n41673;
  assign n41675 = pi16 ? n1471 : ~n41674;
  assign n41676 = pi19 ? n266 : n246;
  assign n41677 = pi18 ? n18503 : ~n41676;
  assign n41678 = pi19 ? n11879 : ~n16002;
  assign n41679 = pi18 ? n41678 : n32;
  assign n41680 = pi17 ? n41677 : ~n41679;
  assign n41681 = pi16 ? n16391 : ~n41680;
  assign n41682 = pi15 ? n41675 : n41681;
  assign n41683 = pi14 ? n41672 : n41682;
  assign n41684 = pi13 ? n41661 : n41683;
  assign n41685 = pi12 ? n41628 : n41684;
  assign n41686 = pi11 ? n41601 : n41685;
  assign n41687 = pi19 ? n32 : n5688;
  assign n41688 = pi19 ? n34188 : n246;
  assign n41689 = pi18 ? n41687 : n41688;
  assign n41690 = pi19 ? n32302 : n246;
  assign n41691 = pi18 ? n41690 : ~n32;
  assign n41692 = pi17 ? n41689 : ~n41691;
  assign n41693 = pi16 ? n32 : n41692;
  assign n41694 = pi15 ? n41693 : n41369;
  assign n41695 = pi19 ? n4342 : ~n4342;
  assign n41696 = pi18 ? n41695 : n1676;
  assign n41697 = pi17 ? n8193 : ~n41696;
  assign n41698 = pi16 ? n32 : n41697;
  assign n41699 = pi15 ? n41698 : n28620;
  assign n41700 = pi14 ? n41694 : n41699;
  assign n41701 = pi13 ? n41700 : n28629;
  assign n41702 = pi12 ? n41701 : n32;
  assign n41703 = pi15 ? n32 : n17707;
  assign n41704 = pi18 ? n38424 : n32;
  assign n41705 = pi17 ? n32 : n41704;
  assign n41706 = pi16 ? n32 : n41705;
  assign n41707 = pi15 ? n32 : n41706;
  assign n41708 = pi14 ? n41703 : n41707;
  assign n41709 = pi19 ? n9864 : n462;
  assign n41710 = pi18 ? n41709 : n32;
  assign n41711 = pi17 ? n32 : n41710;
  assign n41712 = pi16 ? n32 : n41711;
  assign n41713 = pi20 ? n333 : n3523;
  assign n41714 = pi19 ? n275 : n41713;
  assign n41715 = pi18 ? n17927 : ~n41714;
  assign n41716 = pi17 ? n32 : n41715;
  assign n41717 = pi20 ? n18415 : ~n1331;
  assign n41718 = pi19 ? n41717 : ~n32;
  assign n41719 = pi18 ? n41718 : ~n334;
  assign n41720 = pi19 ? n6327 : ~n32;
  assign n41721 = pi18 ? n41720 : ~n32;
  assign n41722 = pi17 ? n41719 : ~n41721;
  assign n41723 = pi16 ? n41716 : n41722;
  assign n41724 = pi15 ? n41712 : n41723;
  assign n41725 = pi20 ? n274 : n3843;
  assign n41726 = pi19 ? n41135 : n41725;
  assign n41727 = pi18 ? n341 : ~n41726;
  assign n41728 = pi17 ? n32 : n41727;
  assign n41729 = pi20 ? n175 : n333;
  assign n41730 = pi19 ? n6057 : n41729;
  assign n41731 = pi19 ? n21588 : n4491;
  assign n41732 = pi18 ? n41730 : n41731;
  assign n41733 = pi20 ? n174 : n207;
  assign n41734 = pi19 ? n41733 : ~n32;
  assign n41735 = pi18 ? n41734 : ~n32;
  assign n41736 = pi17 ? n41732 : n41735;
  assign n41737 = pi16 ? n41728 : ~n41736;
  assign n41738 = pi20 ? n1324 : n17671;
  assign n41739 = pi20 ? n274 : n310;
  assign n41740 = pi19 ? n41738 : n41739;
  assign n41741 = pi18 ? n356 : ~n41740;
  assign n41742 = pi17 ? n32 : n41741;
  assign n41743 = pi20 ? n175 : n13171;
  assign n41744 = pi19 ? n267 : n41743;
  assign n41745 = pi20 ? n405 : n32;
  assign n41746 = pi19 ? n21588 : n41745;
  assign n41747 = pi18 ? n41744 : n41746;
  assign n41748 = pi19 ? n17974 : n208;
  assign n41749 = pi18 ? n41748 : ~n32;
  assign n41750 = pi17 ? n41747 : n41749;
  assign n41751 = pi16 ? n41742 : ~n41750;
  assign n41752 = pi15 ? n41737 : n41751;
  assign n41753 = pi14 ? n41724 : n41752;
  assign n41754 = pi13 ? n41708 : n41753;
  assign n41755 = pi20 ? n1324 : ~n10878;
  assign n41756 = pi19 ? n41755 : n22652;
  assign n41757 = pi18 ? n222 : ~n41756;
  assign n41758 = pi17 ? n32 : n41757;
  assign n41759 = pi20 ? n28761 : n18415;
  assign n41760 = pi19 ? n35706 : n41759;
  assign n41761 = pi20 ? n8644 : n12884;
  assign n41762 = pi19 ? n41761 : n21108;
  assign n41763 = pi18 ? n41760 : n41762;
  assign n41764 = pi20 ? n18173 : n32;
  assign n41765 = pi19 ? n17974 : ~n41764;
  assign n41766 = pi18 ? n41765 : ~n32;
  assign n41767 = pi17 ? n41763 : n41766;
  assign n41768 = pi16 ? n41758 : ~n41767;
  assign n41769 = pi18 ? n209 : ~n13949;
  assign n41770 = pi17 ? n32 : n41769;
  assign n41771 = pi16 ? n41770 : ~n4064;
  assign n41772 = pi15 ? n41768 : n41771;
  assign n41773 = pi16 ? n1135 : ~n4060;
  assign n41774 = pi20 ? n2358 : ~n2385;
  assign n41775 = pi19 ? n18332 : n41774;
  assign n41776 = pi18 ? n19350 : n41775;
  assign n41777 = pi17 ? n32 : n41776;
  assign n41778 = pi20 ? n1368 : n3523;
  assign n41779 = pi19 ? n6171 : n41778;
  assign n41780 = pi20 ? n6303 : n2385;
  assign n41781 = pi20 ? n17665 : n2385;
  assign n41782 = pi19 ? n41780 : n41781;
  assign n41783 = pi18 ? n41779 : n41782;
  assign n41784 = pi17 ? n41783 : n41414;
  assign n41785 = pi16 ? n41777 : ~n41784;
  assign n41786 = pi15 ? n41773 : n41785;
  assign n41787 = pi14 ? n41772 : n41786;
  assign n41788 = pi20 ? n623 : n207;
  assign n41789 = pi20 ? n321 : n5854;
  assign n41790 = pi19 ? n41788 : n41789;
  assign n41791 = pi18 ? n19350 : n41790;
  assign n41792 = pi17 ? n32 : n41791;
  assign n41793 = pi21 ? n405 : ~n313;
  assign n41794 = pi20 ? n1324 : n41793;
  assign n41795 = pi20 ? n19554 : ~n310;
  assign n41796 = pi19 ? n41794 : ~n41795;
  assign n41797 = pi20 ? n13171 : n2385;
  assign n41798 = pi20 ? n12884 : n2385;
  assign n41799 = pi19 ? n41797 : n41798;
  assign n41800 = pi18 ? n41796 : n41799;
  assign n41801 = pi17 ? n41800 : n41426;
  assign n41802 = pi16 ? n41792 : ~n41801;
  assign n41803 = pi18 ? n4380 : n29440;
  assign n41804 = pi17 ? n32 : n41803;
  assign n41805 = pi17 ? n1028 : ~n28286;
  assign n41806 = pi16 ? n41804 : ~n41805;
  assign n41807 = pi15 ? n41802 : n41806;
  assign n41808 = pi18 ? n1395 : ~n9012;
  assign n41809 = pi17 ? n32 : n41808;
  assign n41810 = pi19 ? n1464 : n750;
  assign n41811 = pi18 ? n41810 : ~n32;
  assign n41812 = pi17 ? n32 : n41811;
  assign n41813 = pi16 ? n41809 : ~n41812;
  assign n41814 = pi15 ? n28681 : n41813;
  assign n41815 = pi14 ? n41807 : n41814;
  assign n41816 = pi13 ? n41787 : n41815;
  assign n41817 = pi12 ? n41754 : n41816;
  assign n41818 = pi11 ? n41702 : n41817;
  assign n41819 = pi10 ? n41686 : n41818;
  assign n41820 = pi09 ? n32 : n41819;
  assign n41821 = pi18 ? n18556 : n618;
  assign n41822 = pi17 ? n18554 : ~n41821;
  assign n41823 = pi16 ? n18260 : n41822;
  assign n41824 = pi15 ? n18008 : n41823;
  assign n41825 = pi17 ? n32 : n3100;
  assign n41826 = pi16 ? n1471 : ~n41825;
  assign n41827 = pi15 ? n41615 : n41826;
  assign n41828 = pi14 ? n41824 : n41827;
  assign n41829 = pi16 ? n1214 : ~n41825;
  assign n41830 = pi15 ? n41826 : n41829;
  assign n41831 = pi18 ? n18088 : n618;
  assign n41832 = pi17 ? n18087 : n41831;
  assign n41833 = pi16 ? n41622 : ~n41832;
  assign n41834 = pi15 ? n19711 : n41833;
  assign n41835 = pi14 ? n41830 : n41834;
  assign n41836 = pi13 ? n41828 : n41835;
  assign n41837 = pi20 ? n357 : n1611;
  assign n41838 = pi19 ? n41837 : n18095;
  assign n41839 = pi18 ? n19350 : n41838;
  assign n41840 = pi17 ? n32 : n41839;
  assign n41841 = pi16 ? n41840 : n41647;
  assign n41842 = pi15 ? n28600 : n41841;
  assign n41843 = pi18 ? n41656 : n237;
  assign n41844 = pi17 ? n41654 : ~n41843;
  assign n41845 = pi16 ? n41651 : n41844;
  assign n41846 = pi15 ? n32 : n41845;
  assign n41847 = pi14 ? n41842 : n41846;
  assign n41848 = pi18 ? n18397 : n3350;
  assign n41849 = pi17 ? n18395 : n41848;
  assign n41850 = pi16 ? n1471 : ~n41849;
  assign n41851 = pi15 ? n41850 : n41681;
  assign n41852 = pi14 ? n41672 : n41851;
  assign n41853 = pi13 ? n41847 : n41852;
  assign n41854 = pi12 ? n41836 : n41853;
  assign n41855 = pi11 ? n41601 : n41854;
  assign n41856 = pi18 ? n41366 : n618;
  assign n41857 = pi17 ? n41365 : ~n41856;
  assign n41858 = pi16 ? n32 : n41857;
  assign n41859 = pi15 ? n41693 : n41858;
  assign n41860 = pi18 ? n41695 : n618;
  assign n41861 = pi17 ? n8193 : ~n41860;
  assign n41862 = pi16 ? n32 : n41861;
  assign n41863 = pi15 ? n41862 : n28727;
  assign n41864 = pi14 ? n41859 : n41863;
  assign n41865 = pi13 ? n41864 : n28734;
  assign n41866 = pi12 ? n41865 : n32;
  assign n41867 = pi14 ? n41703 : n28104;
  assign n41868 = pi20 ? n333 : ~n18173;
  assign n41869 = pi19 ? n41868 : ~n41294;
  assign n41870 = pi18 ? n30697 : n41869;
  assign n41871 = pi17 ? n32 : n41870;
  assign n41872 = pi20 ? n333 : ~n7939;
  assign n41873 = pi20 ? n18624 : n19554;
  assign n41874 = pi19 ? n41872 : ~n41873;
  assign n41875 = pi20 ? n18624 : n18073;
  assign n41876 = pi19 ? n28777 : n41875;
  assign n41877 = pi18 ? n41874 : n41876;
  assign n41878 = pi20 ? n41793 : ~n623;
  assign n41879 = pi19 ? n41878 : ~n462;
  assign n41880 = pi18 ? n41879 : ~n32;
  assign n41881 = pi17 ? n41877 : n41880;
  assign n41882 = pi16 ? n41871 : ~n41881;
  assign n41883 = pi19 ? n32 : n6139;
  assign n41884 = pi18 ? n41883 : ~n28751;
  assign n41885 = pi17 ? n32 : n41884;
  assign n41886 = pi19 ? n28762 : n32;
  assign n41887 = pi18 ? n41886 : n32;
  assign n41888 = pi17 ? n28760 : n41887;
  assign n41889 = pi16 ? n41885 : n41888;
  assign n41890 = pi15 ? n41882 : n41889;
  assign n41891 = pi20 ? n310 : n6085;
  assign n41892 = pi19 ? n28774 : ~n41891;
  assign n41893 = pi20 ? n501 : n18073;
  assign n41894 = pi20 ? n206 : n18073;
  assign n41895 = pi19 ? n41893 : n41894;
  assign n41896 = pi18 ? n41892 : n41895;
  assign n41897 = pi20 ? n785 : ~n357;
  assign n41898 = pi19 ? n41897 : ~n32;
  assign n41899 = pi18 ? n41898 : ~n32;
  assign n41900 = pi17 ? n41896 : n41899;
  assign n41901 = pi16 ? n41742 : ~n41900;
  assign n41902 = pi19 ? n9169 : n6057;
  assign n41903 = pi18 ? n366 : ~n41902;
  assign n41904 = pi17 ? n32 : n41903;
  assign n41905 = pi20 ? n175 : n19554;
  assign n41906 = pi19 ? n275 : n41905;
  assign n41907 = pi18 ? n41906 : n41731;
  assign n41908 = pi19 ? n176 : n208;
  assign n41909 = pi18 ? n41908 : ~n32;
  assign n41910 = pi17 ? n41907 : n41909;
  assign n41911 = pi16 ? n41904 : ~n41910;
  assign n41912 = pi15 ? n41901 : n41911;
  assign n41913 = pi14 ? n41890 : n41912;
  assign n41914 = pi13 ? n41867 : n41913;
  assign n41915 = pi21 ? n1392 : ~n405;
  assign n41916 = pi20 ? n32 : n41915;
  assign n41917 = pi19 ? n32 : n41916;
  assign n41918 = pi20 ? n3523 : ~n749;
  assign n41919 = pi20 ? n1331 : n9863;
  assign n41920 = pi19 ? n41918 : n41919;
  assign n41921 = pi18 ? n41917 : ~n41920;
  assign n41922 = pi17 ? n32 : n41921;
  assign n41923 = pi20 ? n1331 : n274;
  assign n41924 = pi20 ? n14286 : n19554;
  assign n41925 = pi19 ? n41923 : n41924;
  assign n41926 = pi20 ? n41793 : n3523;
  assign n41927 = pi20 ? n428 : n3523;
  assign n41928 = pi19 ? n41926 : n41927;
  assign n41929 = pi18 ? n41925 : n41928;
  assign n41930 = pi19 ? n176 : ~n41764;
  assign n41931 = pi18 ? n41930 : ~n32;
  assign n41932 = pi17 ? n41929 : n41931;
  assign n41933 = pi16 ? n41922 : ~n41932;
  assign n41934 = pi18 ? n1395 : ~n13949;
  assign n41935 = pi17 ? n32 : n41934;
  assign n41936 = pi16 ? n41935 : ~n4064;
  assign n41937 = pi15 ? n41933 : n41936;
  assign n41938 = pi20 ? n1324 : n18337;
  assign n41939 = pi20 ? n20396 : n12884;
  assign n41940 = pi19 ? n41938 : n41939;
  assign n41941 = pi20 ? n28761 : ~n206;
  assign n41942 = pi20 ? n18073 : n206;
  assign n41943 = pi19 ? n41941 : ~n41942;
  assign n41944 = pi18 ? n41940 : ~n41943;
  assign n41945 = pi19 ? n18345 : n207;
  assign n41946 = pi18 ? n41945 : ~n32;
  assign n41947 = pi17 ? n41944 : n41946;
  assign n41948 = pi16 ? n41777 : ~n41947;
  assign n41949 = pi15 ? n41773 : n41948;
  assign n41950 = pi14 ? n41937 : n41949;
  assign n41951 = pi19 ? n8230 : ~n11929;
  assign n41952 = pi20 ? n175 : ~n206;
  assign n41953 = pi19 ? n41952 : ~n31675;
  assign n41954 = pi18 ? n41951 : ~n41953;
  assign n41955 = pi19 ? n18345 : ~n5004;
  assign n41956 = pi18 ? n41955 : ~n32;
  assign n41957 = pi17 ? n41954 : n41956;
  assign n41958 = pi16 ? n41792 : ~n41957;
  assign n41959 = pi16 ? n41804 : ~n1029;
  assign n41960 = pi15 ? n41958 : n41959;
  assign n41961 = pi18 ? n209 : ~n9012;
  assign n41962 = pi17 ? n32 : n41961;
  assign n41963 = pi16 ? n41962 : ~n41812;
  assign n41964 = pi15 ? n28805 : n41963;
  assign n41965 = pi14 ? n41960 : n41964;
  assign n41966 = pi13 ? n41950 : n41965;
  assign n41967 = pi12 ? n41914 : n41966;
  assign n41968 = pi11 ? n41866 : n41967;
  assign n41969 = pi10 ? n41855 : n41968;
  assign n41970 = pi09 ? n32 : n41969;
  assign n41971 = pi08 ? n41820 : n41970;
  assign n41972 = pi07 ? n41598 : n41971;
  assign n41973 = pi13 ? n32 : n18953;
  assign n41974 = pi12 ? n32 : n41973;
  assign n41975 = pi21 ? n1009 : n405;
  assign n41976 = pi20 ? n32 : n41975;
  assign n41977 = pi19 ? n32 : n41976;
  assign n41978 = pi20 ? n9491 : n18129;
  assign n41979 = pi19 ? n5854 : n41978;
  assign n41980 = pi18 ? n41977 : n41979;
  assign n41981 = pi17 ? n32 : n41980;
  assign n41982 = pi20 ? n785 : n3695;
  assign n41983 = pi20 ? n11107 : n274;
  assign n41984 = pi19 ? n41982 : ~n41983;
  assign n41985 = pi20 ? n274 : ~n1385;
  assign n41986 = pi19 ? n41985 : n5854;
  assign n41987 = pi18 ? n41984 : ~n41986;
  assign n41988 = pi18 ? n28855 : ~n237;
  assign n41989 = pi17 ? n41987 : ~n41988;
  assign n41990 = pi16 ? n41981 : ~n41989;
  assign n41991 = pi15 ? n32 : n41990;
  assign n41992 = pi21 ? n124 : ~n174;
  assign n41993 = pi20 ? n32 : n41992;
  assign n41994 = pi19 ? n32 : n41993;
  assign n41995 = pi20 ? n9491 : ~n17652;
  assign n41996 = pi19 ? n501 : n41995;
  assign n41997 = pi18 ? n41994 : n41996;
  assign n41998 = pi17 ? n32 : n41997;
  assign n41999 = pi20 ? n1076 : n6085;
  assign n42000 = pi19 ? n41999 : ~n19115;
  assign n42001 = pi20 ? n501 : ~n175;
  assign n42002 = pi19 ? n42001 : n30682;
  assign n42003 = pi18 ? n42000 : ~n42002;
  assign n42004 = pi19 ? n1844 : n1817;
  assign n42005 = pi18 ? n42004 : n237;
  assign n42006 = pi17 ? n42003 : n42005;
  assign n42007 = pi16 ? n41998 : ~n42006;
  assign n42008 = pi20 ? n274 : n1817;
  assign n42009 = pi19 ? n339 : ~n42008;
  assign n42010 = pi18 ? n940 : n42009;
  assign n42011 = pi17 ? n32 : n42010;
  assign n42012 = pi20 ? n314 : n339;
  assign n42013 = pi19 ? n176 : ~n42012;
  assign n42014 = pi20 ? n339 : ~n1331;
  assign n42015 = pi19 ? n42014 : n339;
  assign n42016 = pi18 ? n42013 : ~n42015;
  assign n42017 = pi19 ? n617 : ~n357;
  assign n42018 = pi18 ? n42017 : ~n1942;
  assign n42019 = pi17 ? n42016 : ~n42018;
  assign n42020 = pi16 ? n42011 : ~n42019;
  assign n42021 = pi15 ? n42007 : n42020;
  assign n42022 = pi14 ? n41991 : n42021;
  assign n42023 = pi16 ? n1705 : ~n1944;
  assign n42024 = pi16 ? n1471 : ~n1944;
  assign n42025 = pi15 ? n42023 : n42024;
  assign n42026 = pi18 ? n4380 : n18096;
  assign n42027 = pi17 ? n32 : n42026;
  assign n42028 = pi18 ? n18378 : n54;
  assign n42029 = pi17 ? n18376 : ~n42028;
  assign n42030 = pi16 ? n42027 : ~n42029;
  assign n42031 = pi15 ? n42024 : n42030;
  assign n42032 = pi14 ? n42025 : n42031;
  assign n42033 = pi13 ? n42022 : n42032;
  assign n42034 = pi19 ? n9007 : n32082;
  assign n42035 = pi19 ? n9169 : n8622;
  assign n42036 = pi18 ? n42034 : n42035;
  assign n42037 = pi19 ? n339 : ~n175;
  assign n42038 = pi18 ? n42037 : ~n237;
  assign n42039 = pi17 ? n42036 : ~n42038;
  assign n42040 = pi16 ? n28888 : ~n42039;
  assign n42041 = pi20 ? n9488 : ~n1091;
  assign n42042 = pi19 ? n32 : n42041;
  assign n42043 = pi18 ? n32 : n42042;
  assign n42044 = pi17 ? n32 : n42043;
  assign n42045 = pi18 ? n36866 : n42035;
  assign n42046 = pi18 ? n42037 : ~n3350;
  assign n42047 = pi17 ? n42045 : ~n42046;
  assign n42048 = pi16 ? n42044 : ~n42047;
  assign n42049 = pi15 ? n42040 : n42048;
  assign n42050 = pi19 ? n32 : n35462;
  assign n42051 = pi18 ? n32 : n42050;
  assign n42052 = pi17 ? n32 : n42051;
  assign n42053 = pi16 ? n42052 : n19473;
  assign n42054 = pi20 ? n9194 : n18261;
  assign n42055 = pi19 ? n42054 : ~n5855;
  assign n42056 = pi18 ? n42055 : ~n32;
  assign n42057 = pi17 ? n42056 : ~n2123;
  assign n42058 = pi16 ? n32 : n42057;
  assign n42059 = pi15 ? n42053 : n42058;
  assign n42060 = pi14 ? n42049 : n42059;
  assign n42061 = pi13 ? n28885 : n42060;
  assign n42062 = pi12 ? n42033 : n42061;
  assign n42063 = pi11 ? n41974 : n42062;
  assign n42064 = pi20 ? n18415 : n18281;
  assign n42065 = pi19 ? n857 : ~n42064;
  assign n42066 = pi19 ? n18761 : n29918;
  assign n42067 = pi18 ? n42065 : ~n42066;
  assign n42068 = pi18 ? n248 : n618;
  assign n42069 = pi17 ? n42067 : ~n42068;
  assign n42070 = pi16 ? n32 : n42069;
  assign n42071 = pi20 ? n14286 : ~n428;
  assign n42072 = pi19 ? n32 : n42071;
  assign n42073 = pi18 ? n32 : n42072;
  assign n42074 = pi20 ? n1324 : n333;
  assign n42075 = pi20 ? n310 : n3523;
  assign n42076 = pi19 ? n42074 : n42075;
  assign n42077 = pi18 ? n42076 : n618;
  assign n42078 = pi17 ? n42073 : ~n42077;
  assign n42079 = pi16 ? n32 : n42078;
  assign n42080 = pi15 ? n42070 : n42079;
  assign n42081 = pi19 ? n18722 : n1757;
  assign n42082 = pi18 ? n42081 : n618;
  assign n42083 = pi17 ? n17119 : ~n42082;
  assign n42084 = pi16 ? n32 : n42083;
  assign n42085 = pi15 ? n42084 : n18008;
  assign n42086 = pi14 ? n42080 : n42085;
  assign n42087 = pi13 ? n42086 : n28932;
  assign n42088 = pi15 ? n17894 : n17885;
  assign n42089 = pi14 ? n42088 : n28507;
  assign n42090 = pi13 ? n42089 : n32;
  assign n42091 = pi12 ? n42087 : n42090;
  assign n42092 = pi19 ? n32 : ~n8818;
  assign n42093 = pi18 ? n42092 : n32;
  assign n42094 = pi17 ? n32 : n42093;
  assign n42095 = pi16 ? n22816 : n42094;
  assign n42096 = pi15 ? n130 : n42095;
  assign n42097 = pi18 ? n3776 : ~n32;
  assign n42098 = pi17 ? n32 : n42097;
  assign n42099 = pi16 ? n1135 : ~n42098;
  assign n42100 = pi15 ? n41405 : n42099;
  assign n42101 = pi14 ? n42096 : n42100;
  assign n42102 = pi13 ? n32 : n42101;
  assign n42103 = pi19 ? n267 : ~n1757;
  assign n42104 = pi18 ? n42103 : ~n32;
  assign n42105 = pi17 ? n32 : n42104;
  assign n42106 = pi16 ? n28949 : ~n42105;
  assign n42107 = pi20 ? n32 : n18261;
  assign n42108 = pi19 ? n32 : n42107;
  assign n42109 = pi20 ? n12884 : ~n314;
  assign n42110 = pi20 ? n501 : ~n6621;
  assign n42111 = pi19 ? n42109 : ~n42110;
  assign n42112 = pi18 ? n42108 : n42111;
  assign n42113 = pi17 ? n32 : n42112;
  assign n42114 = pi20 ? n19731 : ~n274;
  assign n42115 = pi20 ? n6617 : ~n428;
  assign n42116 = pi19 ? n42114 : n42115;
  assign n42117 = pi20 ? n1091 : n18129;
  assign n42118 = pi20 ? n6085 : ~n17652;
  assign n42119 = pi19 ? n42117 : n42118;
  assign n42120 = pi18 ? n42116 : ~n42119;
  assign n42121 = pi19 ? n38705 : ~n32;
  assign n42122 = pi18 ? n42121 : ~n32;
  assign n42123 = pi17 ? n42120 : ~n42122;
  assign n42124 = pi16 ? n42113 : n42123;
  assign n42125 = pi15 ? n42106 : n42124;
  assign n42126 = pi18 ? n463 : n18474;
  assign n42127 = pi17 ? n32 : n42126;
  assign n42128 = pi16 ? n42127 : n32;
  assign n42129 = pi19 ? n322 : ~n18478;
  assign n42130 = pi18 ? n863 : n42129;
  assign n42131 = pi17 ? n32 : n42130;
  assign n42132 = pi16 ? n42131 : n29937;
  assign n42133 = pi15 ? n42128 : n42132;
  assign n42134 = pi14 ? n42125 : n42133;
  assign n42135 = pi18 ? n1395 : n350;
  assign n42136 = pi17 ? n32 : n42135;
  assign n42137 = pi17 ? n18491 : n1500;
  assign n42138 = pi16 ? n42136 : ~n42137;
  assign n42139 = pi19 ? n9007 : ~n18497;
  assign n42140 = pi18 ? n32 : n42139;
  assign n42141 = pi17 ? n32 : n42140;
  assign n42142 = pi16 ? n42141 : n28989;
  assign n42143 = pi15 ? n42138 : n42142;
  assign n42144 = pi16 ? n19652 : ~n1471;
  assign n42145 = pi15 ? n42144 : n29519;
  assign n42146 = pi14 ? n42143 : n42145;
  assign n42147 = pi13 ? n42134 : n42146;
  assign n42148 = pi12 ? n42102 : n42147;
  assign n42149 = pi11 ? n42091 : n42148;
  assign n42150 = pi10 ? n42063 : n42149;
  assign n42151 = pi09 ? n32 : n42150;
  assign n42152 = pi13 ? n32 : n19163;
  assign n42153 = pi12 ? n32 : n42152;
  assign n42154 = pi18 ? n936 : n41979;
  assign n42155 = pi17 ? n32 : n42154;
  assign n42156 = pi16 ? n42155 : ~n41989;
  assign n42157 = pi15 ? n32 : n42156;
  assign n42158 = pi18 ? n18402 : n41996;
  assign n42159 = pi17 ? n32 : n42158;
  assign n42160 = pi16 ? n42159 : ~n42006;
  assign n42161 = pi20 ? n18832 : ~n18282;
  assign n42162 = pi19 ? n314 : n42161;
  assign n42163 = pi18 ? n18402 : n42162;
  assign n42164 = pi17 ? n32 : n42163;
  assign n42165 = pi20 ? n1368 : n6085;
  assign n42166 = pi19 ? n42165 : ~n18253;
  assign n42167 = pi20 ? n18253 : ~n18129;
  assign n42168 = pi20 ? n314 : n820;
  assign n42169 = pi19 ? n42167 : n42168;
  assign n42170 = pi18 ? n42166 : ~n42169;
  assign n42171 = pi20 ? n18832 : n339;
  assign n42172 = pi19 ? n42171 : ~n9194;
  assign n42173 = pi22 ? n84 : n50;
  assign n42174 = pi21 ? n42173 : ~n32;
  assign n42175 = pi20 ? n42174 : ~n32;
  assign n42176 = pi19 ? n42175 : ~n32;
  assign n42177 = pi18 ? n42172 : ~n42176;
  assign n42178 = pi17 ? n42170 : ~n42177;
  assign n42179 = pi16 ? n42164 : ~n42178;
  assign n42180 = pi15 ? n42160 : n42179;
  assign n42181 = pi14 ? n42157 : n42180;
  assign n42182 = pi16 ? n1471 : ~n2326;
  assign n42183 = pi15 ? n42023 : n42182;
  assign n42184 = pi18 ? n18542 : n32;
  assign n42185 = pi17 ? n18539 : ~n42184;
  assign n42186 = pi16 ? n28597 : ~n42185;
  assign n42187 = pi15 ? n42182 : n42186;
  assign n42188 = pi14 ? n42183 : n42187;
  assign n42189 = pi13 ? n42181 : n42188;
  assign n42190 = pi16 ? n29060 : ~n42039;
  assign n42191 = pi19 ? n32 : n13747;
  assign n42192 = pi18 ? n32 : n42191;
  assign n42193 = pi17 ? n32 : n42192;
  assign n42194 = pi17 ? n42045 : ~n42038;
  assign n42195 = pi16 ? n42193 : ~n42194;
  assign n42196 = pi15 ? n42190 : n42195;
  assign n42197 = pi17 ? n32 : n4319;
  assign n42198 = pi17 ? n2008 : ~n2325;
  assign n42199 = pi16 ? n42197 : n42198;
  assign n42200 = pi20 ? n175 : n2385;
  assign n42201 = pi19 ? n42200 : ~n5855;
  assign n42202 = pi18 ? n42201 : ~n32;
  assign n42203 = pi17 ? n42202 : ~n2123;
  assign n42204 = pi16 ? n32 : n42203;
  assign n42205 = pi15 ? n42199 : n42204;
  assign n42206 = pi14 ? n42196 : n42205;
  assign n42207 = pi13 ? n29056 : n42206;
  assign n42208 = pi12 ? n42189 : n42207;
  assign n42209 = pi11 ? n42153 : n42208;
  assign n42210 = pi19 ? n32 : ~n29918;
  assign n42211 = pi18 ? n32 : n42210;
  assign n42212 = pi18 ? n248 : n3350;
  assign n42213 = pi17 ? n42211 : ~n42212;
  assign n42214 = pi16 ? n32 : n42213;
  assign n42215 = pi18 ? n42076 : n3350;
  assign n42216 = pi17 ? n42073 : ~n42215;
  assign n42217 = pi16 ? n32 : n42216;
  assign n42218 = pi15 ? n42214 : n42217;
  assign n42219 = pi15 ? n42084 : n18297;
  assign n42220 = pi14 ? n42218 : n42219;
  assign n42221 = pi13 ? n42220 : n29080;
  assign n42222 = pi15 ? n32 : n17885;
  assign n42223 = pi14 ? n42222 : n28507;
  assign n42224 = pi13 ? n42223 : n32;
  assign n42225 = pi12 ? n42221 : n42224;
  assign n42226 = pi15 ? n32 : n42095;
  assign n42227 = pi16 ? n1233 : ~n42098;
  assign n42228 = pi15 ? n41405 : n42227;
  assign n42229 = pi14 ? n42226 : n42228;
  assign n42230 = pi13 ? n32 : n42229;
  assign n42231 = pi19 ? n267 : ~n32082;
  assign n42232 = pi18 ? n42231 : ~n32;
  assign n42233 = pi17 ? n32 : n42232;
  assign n42234 = pi16 ? n28949 : ~n42233;
  assign n42235 = pi19 ? n12885 : ~n18502;
  assign n42236 = pi18 ? n42108 : n42235;
  assign n42237 = pi17 ? n32 : n42236;
  assign n42238 = pi20 ? n19731 : ~n333;
  assign n42239 = pi19 ? n42238 : n18622;
  assign n42240 = pi20 ? n3523 : ~n18624;
  assign n42241 = pi20 ? n9491 : ~n9641;
  assign n42242 = pi19 ? n42240 : ~n42241;
  assign n42243 = pi18 ? n42239 : n42242;
  assign n42244 = pi20 ? n18073 : ~n28761;
  assign n42245 = pi19 ? n42244 : ~n32;
  assign n42246 = pi18 ? n42245 : ~n32;
  assign n42247 = pi17 ? n42243 : ~n42246;
  assign n42248 = pi16 ? n42237 : n42247;
  assign n42249 = pi15 ? n42234 : n42248;
  assign n42250 = pi14 ? n42249 : n42133;
  assign n42251 = pi18 ? n209 : n350;
  assign n42252 = pi17 ? n32 : n42251;
  assign n42253 = pi16 ? n42252 : ~n42137;
  assign n42254 = pi15 ? n42253 : n42142;
  assign n42255 = pi15 ? n28992 : n29676;
  assign n42256 = pi14 ? n42254 : n42255;
  assign n42257 = pi13 ? n42250 : n42256;
  assign n42258 = pi12 ? n42230 : n42257;
  assign n42259 = pi11 ? n42225 : n42258;
  assign n42260 = pi10 ? n42209 : n42259;
  assign n42261 = pi09 ? n32 : n42260;
  assign n42262 = pi08 ? n42151 : n42261;
  assign n42263 = pi13 ? n29128 : n29865;
  assign n42264 = pi12 ? n32 : n42263;
  assign n42265 = pi17 ? n13946 : n20200;
  assign n42266 = pi16 ? n32 : n42265;
  assign n42267 = pi15 ? n32 : n42266;
  assign n42268 = pi15 ? n18676 : n18672;
  assign n42269 = pi14 ? n42267 : n42268;
  assign n42270 = pi19 ? n21105 : n41134;
  assign n42271 = pi18 ? n940 : ~n42270;
  assign n42272 = pi17 ? n32 : n42271;
  assign n42273 = pi19 ? n28243 : n357;
  assign n42274 = pi20 ? n6085 : n174;
  assign n42275 = pi19 ? n18665 : n42274;
  assign n42276 = pi18 ? n42273 : n42275;
  assign n42277 = pi19 ? n5614 : n266;
  assign n42278 = pi18 ? n42277 : n237;
  assign n42279 = pi17 ? n42276 : n42278;
  assign n42280 = pi16 ? n42272 : ~n42279;
  assign n42281 = pi15 ? n42280 : n32;
  assign n42282 = pi14 ? n18676 : n42281;
  assign n42283 = pi13 ? n42269 : n42282;
  assign n42284 = pi19 ? n29173 : n18332;
  assign n42285 = pi18 ? n42284 : ~n16981;
  assign n42286 = pi18 ? n618 : ~n237;
  assign n42287 = pi17 ? n42285 : n42286;
  assign n42288 = pi16 ? n32 : n42287;
  assign n42289 = pi20 ? n32 : n6085;
  assign n42290 = pi20 ? n18408 : n29452;
  assign n42291 = pi19 ? n42289 : n42290;
  assign n42292 = pi20 ? n1324 : n266;
  assign n42293 = pi19 ? n42292 : n1324;
  assign n42294 = pi18 ? n42291 : ~n42293;
  assign n42295 = pi20 ? n428 : n310;
  assign n42296 = pi20 ? n785 : n2180;
  assign n42297 = pi19 ? n42295 : ~n42296;
  assign n42298 = pi18 ? n42297 : n237;
  assign n42299 = pi17 ? n42294 : ~n42298;
  assign n42300 = pi16 ? n32 : n42299;
  assign n42301 = pi15 ? n42288 : n42300;
  assign n42302 = pi20 ? n32 : ~n1611;
  assign n42303 = pi19 ? n28833 : n42302;
  assign n42304 = pi18 ? n32 : n42303;
  assign n42305 = pi20 ? n321 : n310;
  assign n42306 = pi19 ? n42305 : ~n28036;
  assign n42307 = pi18 ? n42306 : n237;
  assign n42308 = pi17 ? n42304 : ~n42307;
  assign n42309 = pi16 ? n32 : n42308;
  assign n42310 = pi19 ? n349 : ~n22525;
  assign n42311 = pi18 ? n42310 : n618;
  assign n42312 = pi17 ? n17346 : ~n42311;
  assign n42313 = pi16 ? n32 : n42312;
  assign n42314 = pi15 ? n42309 : n42313;
  assign n42315 = pi14 ? n42301 : n42314;
  assign n42316 = pi13 ? n29172 : n42315;
  assign n42317 = pi12 ? n42283 : n42316;
  assign n42318 = pi11 ? n42264 : n42317;
  assign n42319 = pi19 ? n349 : ~n1077;
  assign n42320 = pi18 ? n42319 : n618;
  assign n42321 = pi17 ? n23052 : ~n42320;
  assign n42322 = pi16 ? n32 : n42321;
  assign n42323 = pi18 ? n13182 : n618;
  assign n42324 = pi17 ? n23052 : ~n42323;
  assign n42325 = pi16 ? n32 : n42324;
  assign n42326 = pi15 ? n42322 : n42325;
  assign n42327 = pi18 ? n29192 : n18076;
  assign n42328 = pi17 ? n3282 : n42327;
  assign n42329 = pi16 ? n32 : n42328;
  assign n42330 = pi15 ? n42329 : n18142;
  assign n42331 = pi14 ? n42326 : n42330;
  assign n42332 = pi13 ? n42331 : n29199;
  assign n42333 = pi14 ? n32 : n28507;
  assign n42334 = pi13 ? n42333 : n32;
  assign n42335 = pi12 ? n42332 : n42334;
  assign n42336 = pi15 ? n466 : n29676;
  assign n42337 = pi20 ? n32 : n314;
  assign n42338 = pi19 ? n32 : n42337;
  assign n42339 = pi19 ? n594 : n274;
  assign n42340 = pi18 ? n42338 : ~n42339;
  assign n42341 = pi17 ? n32 : n42340;
  assign n42342 = pi19 ? n9169 : n41745;
  assign n42343 = pi18 ? n42342 : n18532;
  assign n42344 = pi18 ? n8612 : ~n32;
  assign n42345 = pi17 ? n42343 : n42344;
  assign n42346 = pi16 ? n42341 : ~n42345;
  assign n42347 = pi15 ? n41405 : n42346;
  assign n42348 = pi14 ? n42336 : n42347;
  assign n42349 = pi13 ? n32 : n42348;
  assign n42350 = pi19 ? n18722 : n5688;
  assign n42351 = pi18 ? n222 : n42350;
  assign n42352 = pi17 ? n32 : n42351;
  assign n42353 = pi17 ? n18718 : n32;
  assign n42354 = pi16 ? n42352 : n42353;
  assign n42355 = pi19 ? n22891 : ~n29269;
  assign n42356 = pi18 ? n18727 : ~n42355;
  assign n42357 = pi18 ? n5436 : ~n32;
  assign n42358 = pi17 ? n42356 : n42357;
  assign n42359 = pi16 ? n1135 : ~n42358;
  assign n42360 = pi15 ? n42354 : n42359;
  assign n42361 = pi14 ? n32 : n42360;
  assign n42362 = pi21 ? n10182 : n259;
  assign n42363 = pi20 ? n32 : n42362;
  assign n42364 = pi19 ? n32 : n42363;
  assign n42365 = pi20 ? n274 : ~n339;
  assign n42366 = pi19 ? n42365 : ~n42001;
  assign n42367 = pi18 ? n42364 : ~n42366;
  assign n42368 = pi17 ? n32 : n42367;
  assign n42369 = pi18 ? n177 : n32;
  assign n42370 = pi17 ? n42369 : n2355;
  assign n42371 = pi16 ? n42368 : ~n42370;
  assign n42372 = pi19 ? n9345 : ~n23644;
  assign n42373 = pi18 ? n209 : n42372;
  assign n42374 = pi17 ? n32 : n42373;
  assign n42375 = pi19 ? n18741 : n24204;
  assign n42376 = pi18 ? n42375 : ~n32;
  assign n42377 = pi17 ? n32 : n42376;
  assign n42378 = pi16 ? n42374 : ~n42377;
  assign n42379 = pi15 ? n42371 : n42378;
  assign n42380 = pi14 ? n42379 : n42144;
  assign n42381 = pi13 ? n42361 : n42380;
  assign n42382 = pi12 ? n42349 : n42381;
  assign n42383 = pi11 ? n42335 : n42382;
  assign n42384 = pi10 ? n42318 : n42383;
  assign n42385 = pi09 ? n32 : n42384;
  assign n42386 = pi14 ? n32 : n20583;
  assign n42387 = pi14 ? n20583 : n32;
  assign n42388 = pi13 ? n42386 : n42387;
  assign n42389 = pi14 ? n19531 : n32;
  assign n42390 = pi13 ? n29314 : n42389;
  assign n42391 = pi12 ? n42388 : n42390;
  assign n42392 = pi18 ? n18402 : ~n18779;
  assign n42393 = pi17 ? n32 : n42392;
  assign n42394 = pi20 ? n9488 : n6621;
  assign n42395 = pi19 ? n18785 : n42394;
  assign n42396 = pi18 ? n18784 : n42395;
  assign n42397 = pi19 ? n7435 : n1685;
  assign n42398 = pi18 ? n42397 : n237;
  assign n42399 = pi17 ? n42396 : n42398;
  assign n42400 = pi16 ? n42393 : ~n42399;
  assign n42401 = pi15 ? n42400 : n32;
  assign n42402 = pi14 ? n18676 : n42401;
  assign n42403 = pi13 ? n42269 : n42402;
  assign n42404 = pi19 ? n29340 : n18332;
  assign n42405 = pi18 ? n42404 : ~n16981;
  assign n42406 = pi18 ? n618 : ~n1942;
  assign n42407 = pi17 ? n42405 : n42406;
  assign n42408 = pi16 ? n32 : n42407;
  assign n42409 = pi20 ? n1331 : n6621;
  assign n42410 = pi19 ? n32 : n42409;
  assign n42411 = pi18 ? n42410 : ~n42293;
  assign n42412 = pi18 ? n42297 : n1942;
  assign n42413 = pi17 ? n42411 : ~n42412;
  assign n42414 = pi16 ? n32 : n42413;
  assign n42415 = pi15 ? n42408 : n42414;
  assign n42416 = pi19 ? n32 : n42302;
  assign n42417 = pi18 ? n32 : n42416;
  assign n42418 = pi18 ? n42306 : n1942;
  assign n42419 = pi17 ? n42417 : ~n42418;
  assign n42420 = pi16 ? n32 : n42419;
  assign n42421 = pi15 ? n42420 : n42313;
  assign n42422 = pi14 ? n42415 : n42421;
  assign n42423 = pi13 ? n29339 : n42422;
  assign n42424 = pi12 ? n42403 : n42423;
  assign n42425 = pi11 ? n42391 : n42424;
  assign n42426 = pi18 ? n29192 : n359;
  assign n42427 = pi17 ? n3282 : n42426;
  assign n42428 = pi16 ? n32 : n42427;
  assign n42429 = pi15 ? n42428 : n18294;
  assign n42430 = pi14 ? n42326 : n42429;
  assign n42431 = pi13 ? n42430 : n29360;
  assign n42432 = pi12 ? n42431 : n42334;
  assign n42433 = pi20 ? n32 : n18253;
  assign n42434 = pi19 ? n32 : n42433;
  assign n42435 = pi18 ? n42434 : n18836;
  assign n42436 = pi17 ? n32 : n42435;
  assign n42437 = pi19 ? n18847 : ~n1686;
  assign n42438 = pi18 ? n42437 : n32;
  assign n42439 = pi17 ? n18846 : ~n42438;
  assign n42440 = pi16 ? n42436 : ~n42439;
  assign n42441 = pi15 ? n41405 : n42440;
  assign n42442 = pi14 ? n42336 : n42441;
  assign n42443 = pi13 ? n32 : n42442;
  assign n42444 = pi21 ? n173 : ~n174;
  assign n42445 = pi20 ? n42444 : n339;
  assign n42446 = pi20 ? n501 : ~n1368;
  assign n42447 = pi19 ? n42445 : n42446;
  assign n42448 = pi18 ? n2387 : n42447;
  assign n42449 = pi17 ? n32 : n42448;
  assign n42450 = pi20 ? n342 : n333;
  assign n42451 = pi20 ? n339 : ~n1817;
  assign n42452 = pi19 ? n42450 : ~n42451;
  assign n42453 = pi20 ? n18073 : n32;
  assign n42454 = pi19 ? n275 : n42453;
  assign n42455 = pi18 ? n42452 : n42454;
  assign n42456 = pi20 ? n18073 : n207;
  assign n42457 = pi19 ? n42456 : ~n32;
  assign n42458 = pi18 ? n42457 : ~n32;
  assign n42459 = pi17 ? n42455 : n42458;
  assign n42460 = pi16 ? n42449 : ~n42459;
  assign n42461 = pi19 ? n18741 : n519;
  assign n42462 = pi18 ? n42461 : ~n32;
  assign n42463 = pi17 ? n32 : n42462;
  assign n42464 = pi16 ? n42374 : ~n42463;
  assign n42465 = pi15 ? n42460 : n42464;
  assign n42466 = pi14 ? n42465 : n29403;
  assign n42467 = pi13 ? n42361 : n42466;
  assign n42468 = pi12 ? n42443 : n42467;
  assign n42469 = pi11 ? n42432 : n42468;
  assign n42470 = pi10 ? n42425 : n42469;
  assign n42471 = pi09 ? n32 : n42470;
  assign n42472 = pi08 ? n42385 : n42471;
  assign n42473 = pi07 ? n42262 : n42472;
  assign n42474 = pi06 ? n41972 : n42473;
  assign n42475 = pi05 ? n41229 : n42474;
  assign n42476 = pi04 ? n32 : n42475;
  assign n42477 = pi14 ? n32 : n34363;
  assign n42478 = pi14 ? n18906 : n32;
  assign n42479 = pi13 ? n42477 : n42478;
  assign n42480 = pi14 ? n32 : n18890;
  assign n42481 = pi13 ? n42480 : n42478;
  assign n42482 = pi12 ? n42479 : n42481;
  assign n42483 = pi16 ? n1705 : ~n2326;
  assign n42484 = pi15 ? n32 : n42483;
  assign n42485 = pi18 ? n8106 : n814;
  assign n42486 = pi17 ? n13950 : n42485;
  assign n42487 = pi16 ? n1471 : ~n42486;
  assign n42488 = pi15 ? n42487 : n18798;
  assign n42489 = pi14 ? n42484 : n42488;
  assign n42490 = pi16 ? n1214 : ~n1815;
  assign n42491 = pi18 ? n940 : ~n20020;
  assign n42492 = pi17 ? n32 : n42491;
  assign n42493 = pi16 ? n42492 : ~n1815;
  assign n42494 = pi15 ? n42490 : n42493;
  assign n42495 = pi18 ? n18920 : ~n19893;
  assign n42496 = pi17 ? n18917 : ~n42495;
  assign n42497 = pi16 ? n32 : n42496;
  assign n42498 = pi17 ? n18929 : n18482;
  assign n42499 = pi16 ? n17038 : n42498;
  assign n42500 = pi15 ? n42497 : n42499;
  assign n42501 = pi14 ? n42494 : n42500;
  assign n42502 = pi13 ? n42489 : n42501;
  assign n42503 = pi19 ? n32 : n42289;
  assign n42504 = pi18 ? n32 : n42503;
  assign n42505 = pi17 ? n32 : n42504;
  assign n42506 = pi18 ? n18941 : n32;
  assign n42507 = pi17 ? n18929 : n42506;
  assign n42508 = pi16 ? n42505 : n42507;
  assign n42509 = pi20 ? n5854 : n1076;
  assign n42510 = pi19 ? n32 : n42509;
  assign n42511 = pi20 ? n1076 : n266;
  assign n42512 = pi19 ? n42511 : n19598;
  assign n42513 = pi18 ? n42510 : n42512;
  assign n42514 = pi19 ? n19601 : ~n41146;
  assign n42515 = pi18 ? n42514 : ~n1813;
  assign n42516 = pi17 ? n42513 : n42515;
  assign n42517 = pi16 ? n32 : n42516;
  assign n42518 = pi15 ? n42508 : n42517;
  assign n42519 = pi20 ? n18073 : ~n310;
  assign n42520 = pi19 ? n29363 : n42519;
  assign n42521 = pi18 ? n42520 : ~n6059;
  assign n42522 = pi17 ? n42521 : ~n1814;
  assign n42523 = pi16 ? n32 : n42522;
  assign n42524 = pi15 ? n42523 : n29487;
  assign n42525 = pi14 ? n42518 : n42524;
  assign n42526 = pi20 ? n3523 : ~n28553;
  assign n42527 = pi20 ? n18282 : n406;
  assign n42528 = pi19 ? n42526 : ~n42527;
  assign n42529 = pi18 ? n32 : n42528;
  assign n42530 = pi20 ? n18253 : ~n32;
  assign n42531 = pi19 ? n42074 : ~n42530;
  assign n42532 = pi18 ? n42531 : n814;
  assign n42533 = pi17 ? n42529 : ~n42532;
  assign n42534 = pi16 ? n32 : n42533;
  assign n42535 = pi20 ? n342 : n9491;
  assign n42536 = pi19 ? n617 : ~n42535;
  assign n42537 = pi18 ? n42536 : n237;
  assign n42538 = pi17 ? n32 : ~n42537;
  assign n42539 = pi16 ? n32 : n42538;
  assign n42540 = pi15 ? n42534 : n42539;
  assign n42541 = pi15 ? n19061 : n19073;
  assign n42542 = pi14 ? n42540 : n42541;
  assign n42543 = pi13 ? n42525 : n42542;
  assign n42544 = pi12 ? n42502 : n42543;
  assign n42545 = pi11 ? n42482 : n42544;
  assign n42546 = pi18 ? n11884 : n237;
  assign n42547 = pi17 ? n32 : ~n42546;
  assign n42548 = pi16 ? n32 : n42547;
  assign n42549 = pi15 ? n42548 : n29496;
  assign n42550 = pi14 ? n42549 : n29499;
  assign n42551 = pi14 ? n29504 : n32;
  assign n42552 = pi13 ? n42550 : n42551;
  assign n42553 = pi13 ? n18008 : n32;
  assign n42554 = pi12 ? n42552 : n42553;
  assign n42555 = pi16 ? n1233 : ~n3726;
  assign n42556 = pi15 ? n32 : n42555;
  assign n42557 = pi14 ? n32 : n42556;
  assign n42558 = pi19 ? n322 : n507;
  assign n42559 = pi18 ? n42558 : ~n32;
  assign n42560 = pi17 ? n32 : n42559;
  assign n42561 = pi16 ? n1233 : ~n42560;
  assign n42562 = pi18 ? n366 : ~n18249;
  assign n42563 = pi17 ? n32 : n42562;
  assign n42564 = pi19 ? n8622 : n176;
  assign n42565 = pi18 ? n42564 : n32;
  assign n42566 = pi17 ? n42565 : n2555;
  assign n42567 = pi16 ? n42563 : ~n42566;
  assign n42568 = pi15 ? n42561 : n42567;
  assign n42569 = pi16 ? n16391 : n17636;
  assign n42570 = pi15 ? n32 : n42569;
  assign n42571 = pi14 ? n42568 : n42570;
  assign n42572 = pi13 ? n42557 : n42571;
  assign n42573 = pi16 ? n1135 : ~n4066;
  assign n42574 = pi20 ? n32 : n13426;
  assign n42575 = pi19 ? n32 : n42574;
  assign n42576 = pi18 ? n42575 : ~n16449;
  assign n42577 = pi17 ? n32 : n42576;
  assign n42578 = pi16 ? n42577 : ~n4733;
  assign n42579 = pi15 ? n42573 : n42578;
  assign n42580 = pi14 ? n29566 : n42579;
  assign n42581 = pi18 ? n22865 : ~n32;
  assign n42582 = pi17 ? n32 : n42581;
  assign n42583 = pi16 ? n1135 : ~n42582;
  assign n42584 = pi15 ? n42583 : n29519;
  assign n42585 = pi16 ? n1233 : ~n1594;
  assign n42586 = pi15 ? n42585 : n29875;
  assign n42587 = pi14 ? n42584 : n42586;
  assign n42588 = pi13 ? n42580 : n42587;
  assign n42589 = pi12 ? n42572 : n42588;
  assign n42590 = pi11 ? n42554 : n42589;
  assign n42591 = pi10 ? n42545 : n42590;
  assign n42592 = pi09 ? n32 : n42591;
  assign n42593 = pi15 ? n18657 : n19628;
  assign n42594 = pi14 ? n166 : n42593;
  assign n42595 = pi13 ? n42594 : n42478;
  assign n42596 = pi14 ? n32 : n165;
  assign n42597 = pi14 ? n19147 : n32;
  assign n42598 = pi13 ? n42596 : n42597;
  assign n42599 = pi12 ? n42595 : n42598;
  assign n42600 = pi18 ? n32 : n20023;
  assign n42601 = pi17 ? n32 : n42600;
  assign n42602 = pi16 ? n1705 : ~n42601;
  assign n42603 = pi15 ? n32 : n42602;
  assign n42604 = pi18 ? n8106 : n1813;
  assign n42605 = pi17 ? n13950 : n42604;
  assign n42606 = pi16 ? n5262 : ~n42605;
  assign n42607 = pi16 ? n5262 : ~n1815;
  assign n42608 = pi15 ? n42606 : n42607;
  assign n42609 = pi14 ? n42603 : n42608;
  assign n42610 = pi18 ? n41448 : ~n20020;
  assign n42611 = pi17 ? n32 : n42610;
  assign n42612 = pi16 ? n42611 : ~n1815;
  assign n42613 = pi15 ? n20104 : n42612;
  assign n42614 = pi18 ? n18920 : ~n441;
  assign n42615 = pi17 ? n18917 : ~n42614;
  assign n42616 = pi16 ? n32 : n42615;
  assign n42617 = pi19 ? n18919 : n4491;
  assign n42618 = pi18 ? n1819 : n42617;
  assign n42619 = pi17 ? n32 : n42618;
  assign n42620 = pi18 ? n6059 : n18658;
  assign n42621 = pi17 ? n18929 : n42620;
  assign n42622 = pi16 ? n42619 : n42621;
  assign n42623 = pi15 ? n42616 : n42622;
  assign n42624 = pi14 ? n42613 : n42623;
  assign n42625 = pi13 ? n42609 : n42624;
  assign n42626 = pi16 ? n32 : n42507;
  assign n42627 = pi15 ? n42626 : n42517;
  assign n42628 = pi20 ? n17665 : ~n310;
  assign n42629 = pi19 ? n1818 : n42628;
  assign n42630 = pi18 ? n42629 : ~n6059;
  assign n42631 = pi17 ? n42630 : ~n1814;
  assign n42632 = pi16 ? n32 : n42631;
  assign n42633 = pi15 ? n42632 : n29633;
  assign n42634 = pi14 ? n42627 : n42633;
  assign n42635 = pi20 ? n321 : n18415;
  assign n42636 = pi19 ? n42635 : ~n19612;
  assign n42637 = pi18 ? n42636 : n814;
  assign n42638 = pi17 ? n23052 : ~n42637;
  assign n42639 = pi16 ? n32 : n42638;
  assign n42640 = pi20 ? n175 : n9491;
  assign n42641 = pi19 ? n617 : ~n42640;
  assign n42642 = pi18 ? n42641 : n237;
  assign n42643 = pi17 ? n32 : ~n42642;
  assign n42644 = pi16 ? n32 : n42643;
  assign n42645 = pi15 ? n42639 : n42644;
  assign n42646 = pi15 ? n18814 : n19073;
  assign n42647 = pi14 ? n42645 : n42646;
  assign n42648 = pi13 ? n42634 : n42647;
  assign n42649 = pi12 ? n42625 : n42648;
  assign n42650 = pi11 ? n42599 : n42649;
  assign n42651 = pi18 ? n11884 : n1942;
  assign n42652 = pi17 ? n32 : ~n42651;
  assign n42653 = pi16 ? n32 : n42652;
  assign n42654 = pi15 ? n42653 : n29642;
  assign n42655 = pi14 ? n42654 : n29647;
  assign n42656 = pi14 ? n29652 : n32;
  assign n42657 = pi13 ? n42655 : n42656;
  assign n42658 = pi14 ? n32 : n18148;
  assign n42659 = pi13 ? n42658 : n32;
  assign n42660 = pi12 ? n42657 : n42659;
  assign n42661 = pi16 ? n1135 : ~n3726;
  assign n42662 = pi15 ? n32 : n42661;
  assign n42663 = pi14 ? n32 : n42662;
  assign n42664 = pi16 ? n1135 : ~n42560;
  assign n42665 = pi18 ? n42338 : ~n19084;
  assign n42666 = pi17 ? n32 : n42665;
  assign n42667 = pi18 ? n19095 : ~n32;
  assign n42668 = pi17 ? n19093 : n42667;
  assign n42669 = pi16 ? n42666 : ~n42668;
  assign n42670 = pi15 ? n42664 : n42669;
  assign n42671 = pi18 ? n127 : n16389;
  assign n42672 = pi17 ? n32 : n42671;
  assign n42673 = pi16 ? n42672 : n17909;
  assign n42674 = pi15 ? n32 : n42673;
  assign n42675 = pi14 ? n42670 : n42674;
  assign n42676 = pi13 ? n42663 : n42675;
  assign n42677 = pi20 ? n32 : n7939;
  assign n42678 = pi19 ? n32 : n42677;
  assign n42679 = pi18 ? n42678 : ~n16449;
  assign n42680 = pi17 ? n32 : n42679;
  assign n42681 = pi16 ? n42680 : ~n4733;
  assign n42682 = pi15 ? n42573 : n42681;
  assign n42683 = pi14 ? n29566 : n42682;
  assign n42684 = pi15 ? n42583 : n29676;
  assign n42685 = pi16 ? n1135 : ~n1594;
  assign n42686 = pi15 ? n42685 : n29780;
  assign n42687 = pi14 ? n42684 : n42686;
  assign n42688 = pi13 ? n42683 : n42687;
  assign n42689 = pi12 ? n42676 : n42688;
  assign n42690 = pi11 ? n42660 : n42689;
  assign n42691 = pi10 ? n42650 : n42690;
  assign n42692 = pi09 ? n32 : n42691;
  assign n42693 = pi08 ? n42592 : n42692;
  assign n42694 = pi15 ? n165 : n19694;
  assign n42695 = pi14 ? n19236 : n42694;
  assign n42696 = pi14 ? n20746 : n32;
  assign n42697 = pi13 ? n42695 : n42696;
  assign n42698 = pi14 ? n21124 : n32;
  assign n42699 = pi13 ? n42596 : n42698;
  assign n42700 = pi12 ? n42697 : n42699;
  assign n42701 = pi20 ? n1611 : n448;
  assign n42702 = pi19 ? n1464 : n42701;
  assign n42703 = pi18 ? n32 : n42702;
  assign n42704 = pi17 ? n32 : n42703;
  assign n42705 = pi20 ? n2180 : ~n29457;
  assign n42706 = pi20 ? n17652 : n1324;
  assign n42707 = pi19 ? n42705 : ~n42706;
  assign n42708 = pi20 ? n1324 : n17669;
  assign n42709 = pi19 ? n41738 : n42708;
  assign n42710 = pi18 ? n42707 : ~n42709;
  assign n42711 = pi20 ? n18173 : n18253;
  assign n42712 = pi19 ? n18578 : ~n42711;
  assign n42713 = pi18 ? n42712 : ~n618;
  assign n42714 = pi17 ? n42710 : ~n42713;
  assign n42715 = pi16 ? n42704 : ~n42714;
  assign n42716 = pi19 ? n38323 : n236;
  assign n42717 = pi18 ? n858 : n42716;
  assign n42718 = pi17 ? n32 : n42717;
  assign n42719 = pi18 ? n19142 : n814;
  assign n42720 = pi17 ? n13950 : n42719;
  assign n42721 = pi16 ? n42718 : ~n42720;
  assign n42722 = pi15 ? n42715 : n42721;
  assign n42723 = pi20 ? n9863 : ~n207;
  assign n42724 = pi19 ? n28070 : ~n42723;
  assign n42725 = pi18 ? n32 : n42724;
  assign n42726 = pi17 ? n32 : n42725;
  assign n42727 = pi19 ? n1464 : n267;
  assign n42728 = pi18 ? n42727 : n814;
  assign n42729 = pi17 ? n36651 : n42728;
  assign n42730 = pi16 ? n42726 : ~n42729;
  assign n42731 = pi20 ? n18282 : n18253;
  assign n42732 = pi19 ? n594 : n42731;
  assign n42733 = pi18 ? n32 : n42732;
  assign n42734 = pi17 ? n32 : n42733;
  assign n42735 = pi16 ? n42734 : ~n1808;
  assign n42736 = pi15 ? n42730 : n42735;
  assign n42737 = pi14 ? n42722 : n42736;
  assign n42738 = pi18 ? n32 : n28821;
  assign n42739 = pi17 ? n32 : n42738;
  assign n42740 = pi17 ? n932 : ~n1807;
  assign n42741 = pi16 ? n42739 : n42740;
  assign n42742 = pi15 ? n42741 : n5050;
  assign n42743 = pi20 ? n974 : ~n448;
  assign n42744 = pi19 ? n42743 : ~n32;
  assign n42745 = pi18 ? n42744 : ~n32;
  assign n42746 = pi17 ? n42745 : ~n2136;
  assign n42747 = pi16 ? n32 : n42746;
  assign n42748 = pi20 ? n1091 : ~n518;
  assign n42749 = pi19 ? n6139 : n42748;
  assign n42750 = pi18 ? n42749 : ~n342;
  assign n42751 = pi18 ? n19152 : n237;
  assign n42752 = pi17 ? n42750 : ~n42751;
  assign n42753 = pi16 ? n32 : n42752;
  assign n42754 = pi15 ? n42747 : n42753;
  assign n42755 = pi14 ? n42742 : n42754;
  assign n42756 = pi13 ? n42737 : n42755;
  assign n42757 = pi20 ? n9641 : n9491;
  assign n42758 = pi19 ? n594 : n42757;
  assign n42759 = pi20 ? n310 : ~n314;
  assign n42760 = pi19 ? n42759 : n32;
  assign n42761 = pi18 ? n42758 : ~n42760;
  assign n42762 = pi17 ? n42761 : ~n1807;
  assign n42763 = pi16 ? n32 : n42762;
  assign n42764 = pi19 ? n32 : n29473;
  assign n42765 = pi18 ? n32 : n42764;
  assign n42766 = pi20 ? n266 : ~n18415;
  assign n42767 = pi20 ? n29452 : n9488;
  assign n42768 = pi19 ? n42766 : n42767;
  assign n42769 = pi18 ? n42768 : n350;
  assign n42770 = pi17 ? n42765 : ~n42769;
  assign n42771 = pi16 ? n32 : n42770;
  assign n42772 = pi15 ? n42763 : n42771;
  assign n42773 = pi19 ? n857 : n9488;
  assign n42774 = pi18 ? n32 : n42773;
  assign n42775 = pi20 ? n18408 : n18073;
  assign n42776 = pi20 ? n18282 : n321;
  assign n42777 = pi19 ? n42775 : n42776;
  assign n42778 = pi18 ? n42777 : ~n350;
  assign n42779 = pi17 ? n42774 : n42778;
  assign n42780 = pi16 ? n32 : n42779;
  assign n42781 = pi15 ? n42780 : n19628;
  assign n42782 = pi14 ? n42772 : n42781;
  assign n42783 = pi18 ? n751 : ~n814;
  assign n42784 = pi17 ? n32 : n42783;
  assign n42785 = pi16 ? n32 : n42784;
  assign n42786 = pi18 ? n2387 : ~n814;
  assign n42787 = pi17 ? n32 : n42786;
  assign n42788 = pi16 ? n32 : n42787;
  assign n42789 = pi15 ? n42785 : n42788;
  assign n42790 = pi18 ? n2387 : ~n237;
  assign n42791 = pi17 ? n32 : n42790;
  assign n42792 = pi16 ? n32 : n42791;
  assign n42793 = pi19 ? n207 : n18211;
  assign n42794 = pi18 ? n127 : ~n42793;
  assign n42795 = pi17 ? n32 : n42794;
  assign n42796 = pi19 ? n28686 : n220;
  assign n42797 = pi19 ? n5675 : n9007;
  assign n42798 = pi18 ? n42796 : ~n42797;
  assign n42799 = pi19 ? n5741 : n322;
  assign n42800 = pi18 ? n42799 : ~n237;
  assign n42801 = pi17 ? n42798 : n42800;
  assign n42802 = pi16 ? n42795 : n42801;
  assign n42803 = pi15 ? n42792 : n42802;
  assign n42804 = pi14 ? n42789 : n42803;
  assign n42805 = pi13 ? n42782 : n42804;
  assign n42806 = pi12 ? n42756 : n42805;
  assign n42807 = pi11 ? n42700 : n42806;
  assign n42808 = pi19 ? n207 : n28957;
  assign n42809 = pi18 ? n32 : ~n42808;
  assign n42810 = pi17 ? n32 : n42809;
  assign n42811 = pi19 ? n6018 : n17749;
  assign n42812 = pi18 ? n42811 : n16449;
  assign n42813 = pi18 ? n23504 : n237;
  assign n42814 = pi17 ? n42812 : n42813;
  assign n42815 = pi16 ? n42810 : ~n42814;
  assign n42816 = pi15 ? n42815 : n18814;
  assign n42817 = pi15 ? n19073 : n19172;
  assign n42818 = pi14 ? n42816 : n42817;
  assign n42819 = pi14 ? n19461 : n32;
  assign n42820 = pi13 ? n42818 : n42819;
  assign n42821 = pi12 ? n42820 : n32;
  assign n42822 = pi15 ? n32 : n33111;
  assign n42823 = pi14 ? n32 : n42822;
  assign n42824 = pi18 ? n356 : ~n19188;
  assign n42825 = pi17 ? n32 : n42824;
  assign n42826 = pi18 ? n19194 : n32;
  assign n42827 = pi17 ? n19193 : n42826;
  assign n42828 = pi16 ? n42825 : n42827;
  assign n42829 = pi15 ? n28947 : n42828;
  assign n42830 = pi16 ? n17120 : n32;
  assign n42831 = pi18 ? n463 : n19202;
  assign n42832 = pi17 ? n32 : n42831;
  assign n42833 = pi16 ? n42832 : n32;
  assign n42834 = pi15 ? n42830 : n42833;
  assign n42835 = pi14 ? n42829 : n42834;
  assign n42836 = pi13 ? n42823 : n42835;
  assign n42837 = pi18 ? n268 : n24647;
  assign n42838 = pi17 ? n32 : n42837;
  assign n42839 = pi16 ? n42838 : n32;
  assign n42840 = pi15 ? n32 : n42839;
  assign n42841 = pi20 ? n7839 : n12882;
  assign n42842 = pi19 ? n42841 : ~n5748;
  assign n42843 = pi18 ? n19350 : n42842;
  assign n42844 = pi17 ? n32 : n42843;
  assign n42845 = pi20 ? n1685 : n9863;
  assign n42846 = pi19 ? n42845 : n358;
  assign n42847 = pi18 ? n42846 : n19082;
  assign n42848 = pi19 ? n6057 : n4406;
  assign n42849 = pi18 ? n42848 : ~n32;
  assign n42850 = pi17 ? n42847 : n42849;
  assign n42851 = pi16 ? n42844 : ~n42850;
  assign n42852 = pi15 ? n41405 : n42851;
  assign n42853 = pi14 ? n42840 : n42852;
  assign n42854 = pi18 ? n209 : ~n6071;
  assign n42855 = pi17 ? n32 : n42854;
  assign n42856 = pi16 ? n42855 : ~n1581;
  assign n42857 = pi16 ? n1214 : ~n1594;
  assign n42858 = pi15 ? n42856 : n42857;
  assign n42859 = pi18 ? n209 : ~n17118;
  assign n42860 = pi17 ? n32 : n42859;
  assign n42861 = pi16 ? n42860 : ~n1594;
  assign n42862 = pi14 ? n42858 : n42861;
  assign n42863 = pi13 ? n42853 : n42862;
  assign n42864 = pi12 ? n42836 : n42863;
  assign n42865 = pi11 ? n42821 : n42864;
  assign n42866 = pi10 ? n42807 : n42865;
  assign n42867 = pi09 ? n32 : n42866;
  assign n42868 = pi15 ? n19235 : n19240;
  assign n42869 = pi14 ? n19236 : n42868;
  assign n42870 = pi14 ? n30369 : n32;
  assign n42871 = pi13 ? n42869 : n42870;
  assign n42872 = pi12 ? n42697 : n42871;
  assign n42873 = pi20 ? n32 : n3695;
  assign n42874 = pi20 ? n18261 : ~n2180;
  assign n42875 = pi19 ? n42873 : n42874;
  assign n42876 = pi18 ? n32 : n42875;
  assign n42877 = pi17 ? n32 : n42876;
  assign n42878 = pi20 ? n1368 : ~n6050;
  assign n42879 = pi20 ? n18415 : n2358;
  assign n42880 = pi19 ? n42878 : ~n42879;
  assign n42881 = pi20 ? n2358 : n18281;
  assign n42882 = pi19 ? n42881 : n2358;
  assign n42883 = pi18 ? n42880 : ~n42882;
  assign n42884 = pi20 ? n18408 : n9194;
  assign n42885 = pi19 ? n18416 : ~n42884;
  assign n42886 = pi18 ? n42885 : ~n822;
  assign n42887 = pi17 ? n42883 : ~n42886;
  assign n42888 = pi16 ? n42877 : ~n42887;
  assign n42889 = pi18 ? n32 : n8975;
  assign n42890 = pi17 ? n32 : n42889;
  assign n42891 = pi16 ? n42890 : ~n42720;
  assign n42892 = pi15 ? n42888 : n42891;
  assign n42893 = pi20 ? n7839 : ~n207;
  assign n42894 = pi19 ? n32 : ~n42893;
  assign n42895 = pi18 ? n32 : n42894;
  assign n42896 = pi17 ? n32 : n42895;
  assign n42897 = pi16 ? n42896 : ~n42729;
  assign n42898 = pi20 ? n1817 : n9194;
  assign n42899 = pi19 ? n32 : n42898;
  assign n42900 = pi18 ? n32 : n42899;
  assign n42901 = pi17 ? n32 : n42900;
  assign n42902 = pi16 ? n42901 : ~n1808;
  assign n42903 = pi15 ? n42897 : n42902;
  assign n42904 = pi14 ? n42892 : n42903;
  assign n42905 = pi19 ? n35462 : ~n32;
  assign n42906 = pi18 ? n42905 : ~n32;
  assign n42907 = pi17 ? n42906 : ~n2136;
  assign n42908 = pi16 ? n32 : n42907;
  assign n42909 = pi20 ? n17665 : ~n518;
  assign n42910 = pi19 ? n1818 : n42909;
  assign n42911 = pi18 ? n42910 : ~n342;
  assign n42912 = pi17 ? n42911 : ~n42751;
  assign n42913 = pi16 ? n32 : n42912;
  assign n42914 = pi15 ? n42908 : n42913;
  assign n42915 = pi14 ? n5050 : n42914;
  assign n42916 = pi13 ? n42904 : n42915;
  assign n42917 = pi20 ? n6050 : ~n2358;
  assign n42918 = pi19 ? n42917 : n32;
  assign n42919 = pi18 ? n858 : ~n42918;
  assign n42920 = pi17 ? n42919 : ~n1807;
  assign n42921 = pi16 ? n32 : n42920;
  assign n42922 = pi15 ? n42921 : n42771;
  assign n42923 = pi18 ? n940 : ~n350;
  assign n42924 = pi17 ? n32 : n42923;
  assign n42925 = pi16 ? n32 : n42924;
  assign n42926 = pi15 ? n42925 : n19628;
  assign n42927 = pi14 ? n42922 : n42926;
  assign n42928 = pi18 ? n751 : ~n1813;
  assign n42929 = pi17 ? n32 : n42928;
  assign n42930 = pi16 ? n32 : n42929;
  assign n42931 = pi18 ? n2387 : ~n1813;
  assign n42932 = pi17 ? n32 : n42931;
  assign n42933 = pi16 ? n32 : n42932;
  assign n42934 = pi15 ? n42930 : n42933;
  assign n42935 = pi18 ? n32 : ~n42793;
  assign n42936 = pi17 ? n32 : n42935;
  assign n42937 = pi16 ? n42936 : n42801;
  assign n42938 = pi15 ? n18814 : n42937;
  assign n42939 = pi14 ? n42934 : n42938;
  assign n42940 = pi13 ? n42927 : n42939;
  assign n42941 = pi12 ? n42916 : n42940;
  assign n42942 = pi11 ? n42872 : n42941;
  assign n42943 = pi18 ? n23504 : n814;
  assign n42944 = pi17 ? n42812 : n42943;
  assign n42945 = pi16 ? n42810 : ~n42944;
  assign n42946 = pi15 ? n42945 : n19536;
  assign n42947 = pi14 ? n42946 : n29869;
  assign n42948 = pi14 ? n29871 : n32;
  assign n42949 = pi13 ? n42947 : n42948;
  assign n42950 = pi12 ? n42949 : n32;
  assign n42951 = pi15 ? n17894 : n33111;
  assign n42952 = pi14 ? n32 : n42951;
  assign n42953 = pi18 ? n356 : ~n19281;
  assign n42954 = pi17 ? n32 : n42953;
  assign n42955 = pi16 ? n42954 : n42827;
  assign n42956 = pi15 ? n28947 : n42955;
  assign n42957 = pi16 ? n17434 : n32;
  assign n42958 = pi15 ? n42957 : n42833;
  assign n42959 = pi14 ? n42956 : n42958;
  assign n42960 = pi13 ? n42952 : n42959;
  assign n42961 = pi16 ? n1233 : ~n4729;
  assign n42962 = pi20 ? n246 : n12882;
  assign n42963 = pi19 ? n42962 : ~n5748;
  assign n42964 = pi18 ? n4380 : n42963;
  assign n42965 = pi17 ? n32 : n42964;
  assign n42966 = pi20 ? n1685 : n7839;
  assign n42967 = pi20 ? n17652 : ~n32;
  assign n42968 = pi19 ? n42966 : ~n42967;
  assign n42969 = pi20 ? n831 : ~n310;
  assign n42970 = pi19 ? n5614 : ~n42969;
  assign n42971 = pi18 ? n42968 : n42970;
  assign n42972 = pi19 ? n42295 : n12801;
  assign n42973 = pi18 ? n42972 : ~n32;
  assign n42974 = pi17 ? n42971 : n42973;
  assign n42975 = pi16 ? n42965 : ~n42974;
  assign n42976 = pi15 ? n42961 : n42975;
  assign n42977 = pi14 ? n42840 : n42976;
  assign n42978 = pi13 ? n42977 : n42862;
  assign n42979 = pi12 ? n42960 : n42978;
  assign n42980 = pi11 ? n42950 : n42979;
  assign n42981 = pi10 ? n42942 : n42980;
  assign n42982 = pi09 ? n32 : n42981;
  assign n42983 = pi08 ? n42867 : n42982;
  assign n42984 = pi07 ? n42693 : n42983;
  assign n42985 = pi14 ? n92 : n19235;
  assign n42986 = pi15 ? n19240 : n32;
  assign n42987 = pi14 ? n42986 : n32;
  assign n42988 = pi13 ? n42985 : n42987;
  assign n42989 = pi14 ? n19236 : n19235;
  assign n42990 = pi14 ? n19326 : n32;
  assign n42991 = pi13 ? n42989 : n42990;
  assign n42992 = pi12 ? n42988 : n42991;
  assign n42993 = pi18 ? n237 : ~n13949;
  assign n42994 = pi18 ? n19316 : n350;
  assign n42995 = pi17 ? n42993 : ~n42994;
  assign n42996 = pi16 ? n4578 : n42995;
  assign n42997 = pi18 ? n350 : ~n13949;
  assign n42998 = pi17 ? n42997 : ~n42994;
  assign n42999 = pi16 ? n32 : n42998;
  assign n43000 = pi15 ? n42996 : n42999;
  assign n43001 = pi18 ? n29919 : n32;
  assign n43002 = pi17 ? n43001 : n1807;
  assign n43003 = pi16 ? n32 : ~n43002;
  assign n43004 = pi17 ? n1219 : ~n3337;
  assign n43005 = pi16 ? n32 : n43004;
  assign n43006 = pi15 ? n43003 : n43005;
  assign n43007 = pi14 ? n43000 : n43006;
  assign n43008 = pi17 ? n4408 : ~n3337;
  assign n43009 = pi16 ? n32 : n43008;
  assign n43010 = pi17 ? n2519 : ~n3337;
  assign n43011 = pi16 ? n32 : n43010;
  assign n43012 = pi15 ? n43009 : n43011;
  assign n43013 = pi17 ? n2512 : ~n3337;
  assign n43014 = pi16 ? n32 : n43013;
  assign n43015 = pi19 ? n9668 : ~n32;
  assign n43016 = pi18 ? n32 : n43015;
  assign n43017 = pi17 ? n2855 : ~n43016;
  assign n43018 = pi16 ? n32 : n43017;
  assign n43019 = pi15 ? n43014 : n43018;
  assign n43020 = pi14 ? n43012 : n43019;
  assign n43021 = pi13 ? n43007 : n43020;
  assign n43022 = pi17 ? n2750 : ~n3337;
  assign n43023 = pi16 ? n32 : n43022;
  assign n43024 = pi15 ? n43023 : n19691;
  assign n43025 = pi14 ? n43024 : n29955;
  assign n43026 = pi13 ? n43025 : n19264;
  assign n43027 = pi12 ? n43021 : n43026;
  assign n43028 = pi11 ? n42992 : n43027;
  assign n43029 = pi20 ? n3523 : n357;
  assign n43030 = pi19 ? n43029 : n3495;
  assign n43031 = pi18 ? n32 : n43030;
  assign n43032 = pi18 ? n33807 : ~n237;
  assign n43033 = pi17 ? n43031 : n43032;
  assign n43034 = pi16 ? n32 : n43033;
  assign n43035 = pi15 ? n43034 : n32;
  assign n43036 = pi14 ? n43035 : n19334;
  assign n43037 = pi13 ? n43036 : n29636;
  assign n43038 = pi13 ? n30215 : n32;
  assign n43039 = pi12 ? n43037 : n43038;
  assign n43040 = pi18 ? n36761 : ~n32;
  assign n43041 = pi17 ? n32 : n43040;
  assign n43042 = pi16 ? n19652 : ~n43041;
  assign n43043 = pi15 ? n33111 : n43042;
  assign n43044 = pi14 ? n32 : n43043;
  assign n43045 = pi18 ? n1395 : ~n268;
  assign n43046 = pi17 ? n32 : n43045;
  assign n43047 = pi16 ? n43046 : ~n1581;
  assign n43048 = pi18 ? n127 : n4380;
  assign n43049 = pi17 ? n32 : n43048;
  assign n43050 = pi16 ? n43049 : n32;
  assign n43051 = pi15 ? n43047 : n43050;
  assign n43052 = pi18 ? n32 : n19350;
  assign n43053 = pi17 ? n32 : n43052;
  assign n43054 = pi16 ? n43053 : n32;
  assign n43055 = pi15 ? n32 : n43054;
  assign n43056 = pi14 ? n43051 : n43055;
  assign n43057 = pi13 ? n43044 : n43056;
  assign n43058 = pi18 ? n917 : n880;
  assign n43059 = pi17 ? n32 : n43058;
  assign n43060 = pi16 ? n43059 : ~n1501;
  assign n43061 = pi15 ? n271 : n43060;
  assign n43062 = pi18 ? n19364 : ~n32;
  assign n43063 = pi17 ? n32 : n43062;
  assign n43064 = pi16 ? n1214 : ~n43063;
  assign n43065 = pi15 ? n29676 : n43064;
  assign n43066 = pi14 ? n43061 : n43065;
  assign n43067 = pi18 ? n341 : ~n1819;
  assign n43068 = pi17 ? n32 : n43067;
  assign n43069 = pi16 ? n43068 : ~n2144;
  assign n43070 = pi15 ? n43069 : n29240;
  assign n43071 = pi14 ? n43070 : n29240;
  assign n43072 = pi13 ? n43066 : n43071;
  assign n43073 = pi12 ? n43057 : n43072;
  assign n43074 = pi11 ? n43039 : n43073;
  assign n43075 = pi10 ? n43028 : n43074;
  assign n43076 = pi09 ? n32 : n43075;
  assign n43077 = pi13 ? n42985 : n42990;
  assign n43078 = pi14 ? n92 : n19384;
  assign n43079 = pi14 ? n30011 : n32;
  assign n43080 = pi13 ? n43078 : n43079;
  assign n43081 = pi12 ? n43077 : n43080;
  assign n43082 = pi17 ? n2519 : ~n1807;
  assign n43083 = pi16 ? n32 : n43082;
  assign n43084 = pi15 ? n43009 : n43083;
  assign n43085 = pi19 ? n32 : n314;
  assign n43086 = pi18 ? n32 : n43085;
  assign n43087 = pi19 ? n36253 : ~n1817;
  assign n43088 = pi18 ? n43087 : ~n43015;
  assign n43089 = pi17 ? n43086 : n43088;
  assign n43090 = pi16 ? n32 : n43089;
  assign n43091 = pi15 ? n43014 : n43090;
  assign n43092 = pi14 ? n43084 : n43091;
  assign n43093 = pi13 ? n43007 : n43092;
  assign n43094 = pi14 ? n43024 : n19691;
  assign n43095 = pi14 ? n19628 : n19264;
  assign n43096 = pi13 ? n43094 : n43095;
  assign n43097 = pi12 ? n43093 : n43096;
  assign n43098 = pi11 ? n43081 : n43097;
  assign n43099 = pi17 ? n18560 : n19170;
  assign n43100 = pi16 ? n32 : n43099;
  assign n43101 = pi15 ? n43100 : n32;
  assign n43102 = pi14 ? n43101 : n19399;
  assign n43103 = pi15 ? n18531 : n32;
  assign n43104 = pi14 ? n43103 : n32;
  assign n43105 = pi13 ? n43102 : n43104;
  assign n43106 = pi15 ? n19172 : n41;
  assign n43107 = pi14 ? n43106 : n32;
  assign n43108 = pi13 ? n43107 : n32;
  assign n43109 = pi12 ? n43105 : n43108;
  assign n43110 = pi16 ? n1214 : ~n43041;
  assign n43111 = pi15 ? n33111 : n43110;
  assign n43112 = pi14 ? n32 : n43111;
  assign n43113 = pi18 ? n209 : ~n268;
  assign n43114 = pi17 ? n32 : n43113;
  assign n43115 = pi16 ? n43114 : ~n1581;
  assign n43116 = pi16 ? n26461 : n32;
  assign n43117 = pi15 ? n43115 : n43116;
  assign n43118 = pi14 ? n43117 : n43055;
  assign n43119 = pi13 ? n43112 : n43118;
  assign n43120 = pi16 ? n19652 : ~n43063;
  assign n43121 = pi15 ? n29519 : n43120;
  assign n43122 = pi14 ? n43061 : n43121;
  assign n43123 = pi16 ? n43068 : ~n1581;
  assign n43124 = pi15 ? n43123 : n29240;
  assign n43125 = pi14 ? n43124 : n29240;
  assign n43126 = pi13 ? n43122 : n43125;
  assign n43127 = pi12 ? n43119 : n43126;
  assign n43128 = pi11 ? n43109 : n43127;
  assign n43129 = pi10 ? n43098 : n43128;
  assign n43130 = pi09 ? n32 : n43129;
  assign n43131 = pi08 ? n43076 : n43130;
  assign n43132 = pi14 ? n19925 : n91;
  assign n43133 = pi14 ? n19447 : n32;
  assign n43134 = pi13 ? n43132 : n43133;
  assign n43135 = pi14 ? n92 : n91;
  assign n43136 = pi13 ? n43135 : n43133;
  assign n43137 = pi12 ? n43134 : n43136;
  assign n43138 = pi18 ? n237 : ~n4492;
  assign n43139 = pi18 ? n19439 : n350;
  assign n43140 = pi17 ? n43138 : ~n43139;
  assign n43141 = pi16 ? n32 : n43140;
  assign n43142 = pi18 ? n6063 : ~n5749;
  assign n43143 = pi17 ? n43142 : ~n43139;
  assign n43144 = pi16 ? n32 : n43143;
  assign n43145 = pi15 ? n43141 : n43144;
  assign n43146 = pi20 ? n342 : n501;
  assign n43147 = pi19 ? n43146 : ~n32;
  assign n43148 = pi18 ? n43147 : ~n32;
  assign n43149 = pi17 ? n43148 : ~n2537;
  assign n43150 = pi16 ? n32 : n43149;
  assign n43151 = pi18 ? n25110 : ~n32;
  assign n43152 = pi17 ? n43151 : ~n2537;
  assign n43153 = pi16 ? n32 : n43152;
  assign n43154 = pi15 ? n43150 : n43153;
  assign n43155 = pi14 ? n43145 : n43154;
  assign n43156 = pi17 ? n2119 : ~n2537;
  assign n43157 = pi16 ? n32 : n43156;
  assign n43158 = pi17 ? n2519 : ~n2537;
  assign n43159 = pi16 ? n32 : n43158;
  assign n43160 = pi15 ? n43157 : n43159;
  assign n43161 = pi17 ? n6236 : ~n2537;
  assign n43162 = pi16 ? n32 : n43161;
  assign n43163 = pi19 ? n32 : n23026;
  assign n43164 = pi18 ? n32 : n43163;
  assign n43165 = pi19 ? n6398 : n37542;
  assign n43166 = pi18 ? n43165 : n1548;
  assign n43167 = pi17 ? n43164 : ~n43166;
  assign n43168 = pi16 ? n32 : n43167;
  assign n43169 = pi15 ? n43162 : n43168;
  assign n43170 = pi14 ? n43160 : n43169;
  assign n43171 = pi13 ? n43155 : n43170;
  assign n43172 = pi17 ? n3067 : ~n2880;
  assign n43173 = pi16 ? n32 : n43172;
  assign n43174 = pi15 ? n43173 : n19235;
  assign n43175 = pi14 ? n43174 : n20646;
  assign n43176 = pi14 ? n20960 : n19399;
  assign n43177 = pi13 ? n43175 : n43176;
  assign n43178 = pi12 ? n43171 : n43177;
  assign n43179 = pi11 ? n43137 : n43178;
  assign n43180 = pi14 ? n19333 : n18535;
  assign n43181 = pi13 ? n43180 : n19261;
  assign n43182 = pi14 ? n30211 : n32;
  assign n43183 = pi14 ? n32 : n18016;
  assign n43184 = pi13 ? n43182 : n43183;
  assign n43185 = pi12 ? n43181 : n43184;
  assign n43186 = pi15 ? n33111 : n30025;
  assign n43187 = pi14 ? n18005 : n43186;
  assign n43188 = pi20 ? n32 : n15732;
  assign n43189 = pi19 ? n32 : n43188;
  assign n43190 = pi20 ? n274 : ~n17652;
  assign n43191 = pi19 ? n1817 : n43190;
  assign n43192 = pi18 ? n43189 : ~n43191;
  assign n43193 = pi17 ? n32 : n43192;
  assign n43194 = pi20 ? n18129 : n342;
  assign n43195 = pi19 ? n43194 : n6049;
  assign n43196 = pi20 ? n32 : n18337;
  assign n43197 = pi19 ? n43196 : ~n29914;
  assign n43198 = pi18 ? n43195 : n43197;
  assign n43199 = pi20 ? n428 : n1331;
  assign n43200 = pi19 ? n43199 : n507;
  assign n43201 = pi18 ? n43200 : ~n32;
  assign n43202 = pi17 ? n43198 : n43201;
  assign n43203 = pi16 ? n43193 : ~n43202;
  assign n43204 = pi18 ? n127 : n936;
  assign n43205 = pi17 ? n32 : n43204;
  assign n43206 = pi16 ? n43205 : ~n2009;
  assign n43207 = pi15 ? n43203 : n43206;
  assign n43208 = pi18 ? n463 : n863;
  assign n43209 = pi17 ? n32 : n43208;
  assign n43210 = pi16 ? n43209 : ~n2009;
  assign n43211 = pi15 ? n32 : n43210;
  assign n43212 = pi14 ? n43207 : n43211;
  assign n43213 = pi13 ? n43187 : n43212;
  assign n43214 = pi17 ? n32 : n268;
  assign n43215 = pi16 ? n43214 : ~n1029;
  assign n43216 = pi18 ? n268 : n880;
  assign n43217 = pi17 ? n32 : n43216;
  assign n43218 = pi16 ? n43217 : ~n1501;
  assign n43219 = pi15 ? n43215 : n43218;
  assign n43220 = pi20 ? n32 : n18173;
  assign n43221 = pi19 ? n32 : n43220;
  assign n43222 = pi20 ? n1331 : n246;
  assign n43223 = pi19 ? n3523 : n43222;
  assign n43224 = pi18 ? n43221 : ~n43223;
  assign n43225 = pi17 ? n32 : n43224;
  assign n43226 = pi20 ? n274 : ~n266;
  assign n43227 = pi19 ? n5614 : n43226;
  assign n43228 = pi18 ? n43227 : ~n32;
  assign n43229 = pi17 ? n28638 : n43228;
  assign n43230 = pi16 ? n43225 : ~n43229;
  assign n43231 = pi15 ? n43230 : n29240;
  assign n43232 = pi14 ? n43219 : n43231;
  assign n43233 = pi16 ? n1046 : ~n1834;
  assign n43234 = pi15 ? n43233 : n42685;
  assign n43235 = pi14 ? n43234 : n28947;
  assign n43236 = pi13 ? n43232 : n43235;
  assign n43237 = pi12 ? n43213 : n43236;
  assign n43238 = pi11 ? n43185 : n43237;
  assign n43239 = pi10 ? n43179 : n43238;
  assign n43240 = pi09 ? n32 : n43239;
  assign n43241 = pi14 ? n19504 : n19503;
  assign n43242 = pi14 ? n19618 : n32;
  assign n43243 = pi13 ? n43241 : n43242;
  assign n43244 = pi12 ? n43134 : n43243;
  assign n43245 = pi18 ? n19439 : n1548;
  assign n43246 = pi17 ? n43138 : ~n43245;
  assign n43247 = pi16 ? n32 : n43246;
  assign n43248 = pi17 ? n43142 : ~n43245;
  assign n43249 = pi16 ? n32 : n43248;
  assign n43250 = pi15 ? n43247 : n43249;
  assign n43251 = pi14 ? n43250 : n43154;
  assign n43252 = pi13 ? n43251 : n43170;
  assign n43253 = pi15 ? n43173 : n30155;
  assign n43254 = pi14 ? n43253 : n30155;
  assign n43255 = pi15 ? n18657 : n19691;
  assign n43256 = pi14 ? n43255 : n19698;
  assign n43257 = pi13 ? n43254 : n43256;
  assign n43258 = pi12 ? n43252 : n43257;
  assign n43259 = pi11 ? n43244 : n43258;
  assign n43260 = pi14 ? n20960 : n30199;
  assign n43261 = pi13 ? n43260 : n32;
  assign n43262 = pi12 ? n43261 : n43184;
  assign n43263 = pi15 ? n33111 : n28947;
  assign n43264 = pi14 ? n18005 : n43263;
  assign n43265 = pi18 ? n35362 : ~n43191;
  assign n43266 = pi17 ? n32 : n43265;
  assign n43267 = pi20 ? n6085 : n9491;
  assign n43268 = pi19 ? n43194 : n43267;
  assign n43269 = pi20 ? n17652 : n1076;
  assign n43270 = pi19 ? n41084 : n43269;
  assign n43271 = pi18 ? n43268 : ~n43270;
  assign n43272 = pi20 ? n13171 : ~n310;
  assign n43273 = pi19 ? n43272 : n19559;
  assign n43274 = pi18 ? n43273 : n32;
  assign n43275 = pi17 ? n43271 : ~n43274;
  assign n43276 = pi16 ? n43266 : ~n43275;
  assign n43277 = pi16 ? n3283 : ~n2009;
  assign n43278 = pi15 ? n43276 : n43277;
  assign n43279 = pi14 ? n43278 : n43211;
  assign n43280 = pi13 ? n43264 : n43279;
  assign n43281 = pi20 ? n17671 : ~n266;
  assign n43282 = pi19 ? n5614 : n43281;
  assign n43283 = pi18 ? n43282 : ~n32;
  assign n43284 = pi17 ? n28638 : n43283;
  assign n43285 = pi16 ? n43225 : ~n43284;
  assign n43286 = pi15 ? n43285 : n29240;
  assign n43287 = pi14 ? n43219 : n43286;
  assign n43288 = pi13 ? n43287 : n43235;
  assign n43289 = pi12 ? n43280 : n43288;
  assign n43290 = pi11 ? n43262 : n43289;
  assign n43291 = pi10 ? n43259 : n43290;
  assign n43292 = pi09 ? n32 : n43291;
  assign n43293 = pi08 ? n43240 : n43292;
  assign n43294 = pi07 ? n43131 : n43293;
  assign n43295 = pi06 ? n42984 : n43294;
  assign n43296 = pi14 ? n19869 : n19805;
  assign n43297 = pi13 ? n43296 : n43242;
  assign n43298 = pi14 ? n157 : n19503;
  assign n43299 = pi13 ? n43298 : n43242;
  assign n43300 = pi12 ? n43297 : n43299;
  assign n43301 = pi18 ? n32 : ~n20361;
  assign n43302 = pi20 ? n915 : n342;
  assign n43303 = pi19 ? n34314 : ~n43302;
  assign n43304 = pi18 ? n43303 : ~n19232;
  assign n43305 = pi17 ? n43301 : ~n43304;
  assign n43306 = pi16 ? n32 : n43305;
  assign n43307 = pi15 ? n43306 : n19235;
  assign n43308 = pi18 ? n8192 : ~n20164;
  assign n43309 = pi17 ? n43308 : ~n2537;
  assign n43310 = pi16 ? n32 : n43309;
  assign n43311 = pi19 ? n247 : ~n349;
  assign n43312 = pi18 ? n8192 : ~n43311;
  assign n43313 = pi17 ? n43312 : ~n2319;
  assign n43314 = pi16 ? n32 : n43313;
  assign n43315 = pi15 ? n43310 : n43314;
  assign n43316 = pi14 ? n43307 : n43315;
  assign n43317 = pi17 ? n2750 : ~n2319;
  assign n43318 = pi16 ? n32 : n43317;
  assign n43319 = pi20 ? n9641 : n18415;
  assign n43320 = pi19 ? n32 : n43319;
  assign n43321 = pi18 ? n32 : n43320;
  assign n43322 = pi20 ? n18282 : n1091;
  assign n43323 = pi19 ? n20938 : n43322;
  assign n43324 = pi21 ? n173 : ~n242;
  assign n43325 = pi20 ? n43324 : n32;
  assign n43326 = pi19 ? n43325 : n32;
  assign n43327 = pi18 ? n43323 : ~n43326;
  assign n43328 = pi17 ? n43321 : ~n43327;
  assign n43329 = pi16 ? n32 : n43328;
  assign n43330 = pi15 ? n43329 : n19999;
  assign n43331 = pi14 ? n43318 : n43330;
  assign n43332 = pi13 ? n43316 : n43331;
  assign n43333 = pi18 ? n35798 : n2318;
  assign n43334 = pi17 ? n32 : ~n43333;
  assign n43335 = pi16 ? n32 : n43334;
  assign n43336 = pi15 ? n43335 : n19936;
  assign n43337 = pi14 ? n43336 : n19936;
  assign n43338 = pi15 ? n19531 : n30199;
  assign n43339 = pi20 ? n32 : n18840;
  assign n43340 = pi19 ? n43339 : n462;
  assign n43341 = pi18 ? n32 : n43340;
  assign n43342 = pi17 ? n43341 : n19529;
  assign n43343 = pi16 ? n32 : n43342;
  assign n43344 = pi15 ? n30199 : n43343;
  assign n43345 = pi14 ? n43338 : n43344;
  assign n43346 = pi13 ? n43337 : n43345;
  assign n43347 = pi12 ? n43332 : n43346;
  assign n43348 = pi11 ? n43300 : n43347;
  assign n43349 = pi13 ? n30210 : n32;
  assign n43350 = pi12 ? n43349 : n32;
  assign n43351 = pi19 ? n7939 : n29682;
  assign n43352 = pi18 ? n4380 : ~n43351;
  assign n43353 = pi17 ? n32 : n43352;
  assign n43354 = pi20 ? n4279 : n5854;
  assign n43355 = pi19 ? n1076 : n43354;
  assign n43356 = pi19 ? n28970 : n28973;
  assign n43357 = pi18 ? n43355 : ~n43356;
  assign n43358 = pi20 ? n310 : n17669;
  assign n43359 = pi20 ? n310 : n11107;
  assign n43360 = pi19 ? n43358 : n43359;
  assign n43361 = pi18 ? n43360 : ~n32;
  assign n43362 = pi17 ? n43357 : ~n43361;
  assign n43363 = pi16 ? n43353 : n43362;
  assign n43364 = pi15 ? n32 : n43363;
  assign n43365 = pi15 ? n41405 : n18979;
  assign n43366 = pi14 ? n43364 : n43365;
  assign n43367 = pi16 ? n465 : n29937;
  assign n43368 = pi17 ? n19655 : n32;
  assign n43369 = pi16 ? n129 : n43368;
  assign n43370 = pi15 ? n32 : n43369;
  assign n43371 = pi14 ? n43367 : n43370;
  assign n43372 = pi13 ? n43366 : n43371;
  assign n43373 = pi16 ? n1214 : ~n4729;
  assign n43374 = pi16 ? n1214 : ~n1214;
  assign n43375 = pi15 ? n43373 : n43374;
  assign n43376 = pi17 ? n1500 : ~n1682;
  assign n43377 = pi16 ? n1471 : n43376;
  assign n43378 = pi16 ? n1471 : ~n1834;
  assign n43379 = pi15 ? n43377 : n43378;
  assign n43380 = pi14 ? n43375 : n43379;
  assign n43381 = pi17 ? n2005 : ~n2899;
  assign n43382 = pi16 ? n1471 : n43381;
  assign n43383 = pi16 ? n1214 : ~n5259;
  assign n43384 = pi15 ? n43382 : n43383;
  assign n43385 = pi16 ? n1471 : ~n5259;
  assign n43386 = pi15 ? n43385 : n41272;
  assign n43387 = pi14 ? n43384 : n43386;
  assign n43388 = pi13 ? n43380 : n43387;
  assign n43389 = pi12 ? n43372 : n43388;
  assign n43390 = pi11 ? n43350 : n43389;
  assign n43391 = pi10 ? n43348 : n43390;
  assign n43392 = pi09 ? n32 : n43391;
  assign n43393 = pi14 ? n19932 : n32;
  assign n43394 = pi13 ? n43296 : n43393;
  assign n43395 = pi15 ? n116 : n19874;
  assign n43396 = pi14 ? n117 : n43395;
  assign n43397 = pi15 ? n19874 : n32;
  assign n43398 = pi18 ? n6114 : n32;
  assign n43399 = pi17 ? n32 : n43398;
  assign n43400 = pi16 ? n32 : n43399;
  assign n43401 = pi15 ? n32 : n43400;
  assign n43402 = pi14 ? n43397 : n43401;
  assign n43403 = pi13 ? n43396 : n43402;
  assign n43404 = pi12 ? n43394 : n43403;
  assign n43405 = pi17 ? n2750 : ~n2537;
  assign n43406 = pi16 ? n32 : n43405;
  assign n43407 = pi20 ? n9641 : n333;
  assign n43408 = pi19 ? n32 : n43407;
  assign n43409 = pi18 ? n32 : n43408;
  assign n43410 = pi20 ? n18073 : n17652;
  assign n43411 = pi20 ? n17652 : n13171;
  assign n43412 = pi19 ? n43410 : n43411;
  assign n43413 = pi18 ? n43412 : ~n29919;
  assign n43414 = pi17 ? n43409 : ~n43413;
  assign n43415 = pi16 ? n32 : n43414;
  assign n43416 = pi15 ? n43415 : n20089;
  assign n43417 = pi14 ? n43406 : n43416;
  assign n43418 = pi13 ? n43316 : n43417;
  assign n43419 = pi15 ? n19936 : n20067;
  assign n43420 = pi14 ? n43336 : n43419;
  assign n43421 = pi15 ? n19814 : n30199;
  assign n43422 = pi19 ? n21412 : n462;
  assign n43423 = pi18 ? n32 : n43422;
  assign n43424 = pi17 ? n43423 : n19529;
  assign n43425 = pi16 ? n32 : n43424;
  assign n43426 = pi15 ? n30199 : n43425;
  assign n43427 = pi14 ? n43421 : n43426;
  assign n43428 = pi13 ? n43420 : n43427;
  assign n43429 = pi12 ? n43418 : n43428;
  assign n43430 = pi11 ? n43404 : n43429;
  assign n43431 = pi13 ? n30264 : n28705;
  assign n43432 = pi12 ? n43431 : n32;
  assign n43433 = pi21 ? n10182 : ~n405;
  assign n43434 = pi20 ? n32 : n43433;
  assign n43435 = pi19 ? n32 : n43434;
  assign n43436 = pi21 ? n309 : n173;
  assign n43437 = pi20 ? n43436 : n310;
  assign n43438 = pi19 ? n406 : n43437;
  assign n43439 = pi18 ? n43435 : ~n43438;
  assign n43440 = pi17 ? n32 : n43439;
  assign n43441 = pi20 ? n1076 : n2180;
  assign n43442 = pi20 ? n10889 : ~n18762;
  assign n43443 = pi19 ? n43441 : n43442;
  assign n43444 = pi19 ? n29291 : n29293;
  assign n43445 = pi18 ? n43443 : ~n43444;
  assign n43446 = pi20 ? n1331 : n11107;
  assign n43447 = pi19 ? n29537 : n43446;
  assign n43448 = pi18 ? n43447 : ~n32;
  assign n43449 = pi17 ? n43445 : ~n43448;
  assign n43450 = pi16 ? n43440 : n43449;
  assign n43451 = pi15 ? n32 : n43450;
  assign n43452 = pi15 ? n42961 : n18979;
  assign n43453 = pi14 ? n43451 : n43452;
  assign n43454 = pi16 ? n32 : n43368;
  assign n43455 = pi15 ? n32 : n43454;
  assign n43456 = pi14 ? n43367 : n43455;
  assign n43457 = pi13 ? n43453 : n43456;
  assign n43458 = pi12 ? n43457 : n43388;
  assign n43459 = pi11 ? n43432 : n43458;
  assign n43460 = pi10 ? n43430 : n43459;
  assign n43461 = pi09 ? n32 : n43460;
  assign n43462 = pi08 ? n43392 : n43461;
  assign n43463 = pi15 ? n32 : n20531;
  assign n43464 = pi14 ? n43463 : n19868;
  assign n43465 = pi13 ? n43464 : n40142;
  assign n43466 = pi15 ? n116 : n20538;
  assign n43467 = pi14 ? n117 : n43466;
  assign n43468 = pi15 ? n20538 : n31854;
  assign n43469 = pi19 ? n594 : n4491;
  assign n43470 = pi18 ? n32 : n43469;
  assign n43471 = pi17 ? n43470 : n41018;
  assign n43472 = pi16 ? n32 : n43471;
  assign n43473 = pi15 ? n43472 : n32;
  assign n43474 = pi14 ? n43468 : n43473;
  assign n43475 = pi13 ? n43467 : n43474;
  assign n43476 = pi12 ? n43465 : n43475;
  assign n43477 = pi17 ? n23052 : n18482;
  assign n43478 = pi16 ? n32 : n43477;
  assign n43479 = pi15 ? n43478 : n19805;
  assign n43480 = pi17 ? n43308 : ~n1933;
  assign n43481 = pi16 ? n32 : n43480;
  assign n43482 = pi17 ? n43312 : ~n1933;
  assign n43483 = pi16 ? n32 : n43482;
  assign n43484 = pi15 ? n43481 : n43483;
  assign n43485 = pi14 ? n43479 : n43484;
  assign n43486 = pi17 ? n2750 : ~n1933;
  assign n43487 = pi16 ? n32 : n43486;
  assign n43488 = pi15 ? n30286 : n20072;
  assign n43489 = pi14 ? n43487 : n43488;
  assign n43490 = pi13 ? n43485 : n43489;
  assign n43491 = pi18 ? n35798 : n344;
  assign n43492 = pi17 ? n32 : ~n43491;
  assign n43493 = pi16 ? n32 : n43492;
  assign n43494 = pi15 ? n43493 : n20067;
  assign n43495 = pi14 ? n43494 : n20067;
  assign n43496 = pi18 ? n17848 : n19811;
  assign n43497 = pi17 ? n32 : n43496;
  assign n43498 = pi16 ? n32 : n43497;
  assign n43499 = pi15 ? n43498 : n19942;
  assign n43500 = pi14 ? n43499 : n30290;
  assign n43501 = pi13 ? n43495 : n43500;
  assign n43502 = pi12 ? n43490 : n43501;
  assign n43503 = pi11 ? n43476 : n43502;
  assign n43504 = pi13 ? n30301 : n32;
  assign n43505 = pi12 ? n43504 : n32;
  assign n43506 = pi15 ? n32 : n18979;
  assign n43507 = pi14 ? n43506 : n18979;
  assign n43508 = pi17 ? n19775 : n32;
  assign n43509 = pi16 ? n32 : n43508;
  assign n43510 = pi17 ? n19779 : n32;
  assign n43511 = pi16 ? n465 : n43510;
  assign n43512 = pi15 ? n32 : n43511;
  assign n43513 = pi14 ? n43509 : n43512;
  assign n43514 = pi13 ? n43507 : n43513;
  assign n43515 = pi16 ? n19652 : ~n4729;
  assign n43516 = pi16 ? n19652 : ~n3356;
  assign n43517 = pi15 ? n43515 : n43516;
  assign n43518 = pi18 ? n4689 : n32;
  assign n43519 = pi17 ? n43518 : n1682;
  assign n43520 = pi16 ? n29318 : ~n43519;
  assign n43521 = pi16 ? n20208 : ~n1683;
  assign n43522 = pi15 ? n43520 : n43521;
  assign n43523 = pi14 ? n43517 : n43522;
  assign n43524 = pi17 ? n1227 : ~n1682;
  assign n43525 = pi16 ? n20208 : n43524;
  assign n43526 = pi16 ? n1135 : ~n1834;
  assign n43527 = pi15 ? n43525 : n43526;
  assign n43528 = pi16 ? n20208 : ~n1834;
  assign n43529 = pi16 ? n1233 : ~n1834;
  assign n43530 = pi15 ? n43528 : n43529;
  assign n43531 = pi14 ? n43527 : n43530;
  assign n43532 = pi13 ? n43523 : n43531;
  assign n43533 = pi12 ? n43514 : n43532;
  assign n43534 = pi11 ? n43505 : n43533;
  assign n43535 = pi10 ? n43503 : n43534;
  assign n43536 = pi09 ? n32 : n43535;
  assign n43537 = pi14 ? n32 : n30345;
  assign n43538 = pi17 ? n32 : n2650;
  assign n43539 = pi16 ? n1233 : ~n43538;
  assign n43540 = pi15 ? n20315 : n43539;
  assign n43541 = pi20 ? n428 : n9641;
  assign n43542 = pi19 ? n594 : n43541;
  assign n43543 = pi18 ? n28876 : n43542;
  assign n43544 = pi19 ? n6398 : n6057;
  assign n43545 = pi18 ? n43544 : n32;
  assign n43546 = pi17 ? n43543 : n43545;
  assign n43547 = pi16 ? n32 : n43546;
  assign n43548 = pi15 ? n43547 : n32;
  assign n43549 = pi14 ? n43540 : n43548;
  assign n43550 = pi13 ? n43537 : n43549;
  assign n43551 = pi12 ? n43465 : n43550;
  assign n43552 = pi15 ? n30355 : n20072;
  assign n43553 = pi14 ? n43487 : n43552;
  assign n43554 = pi13 ? n43485 : n43553;
  assign n43555 = pi15 ? n20067 : n20252;
  assign n43556 = pi14 ? n43494 : n43555;
  assign n43557 = pi18 ? n17848 : n19933;
  assign n43558 = pi17 ? n32 : n43557;
  assign n43559 = pi16 ? n32 : n43558;
  assign n43560 = pi15 ? n43559 : n19942;
  assign n43561 = pi14 ? n43560 : n30290;
  assign n43562 = pi13 ? n43556 : n43561;
  assign n43563 = pi12 ? n43554 : n43562;
  assign n43564 = pi11 ? n43551 : n43563;
  assign n43565 = pi13 ? n30370 : n32;
  assign n43566 = pi12 ? n43565 : n32;
  assign n43567 = pi15 ? n32 : n19100;
  assign n43568 = pi14 ? n43567 : n19100;
  assign n43569 = pi13 ? n43568 : n43513;
  assign n43570 = pi15 ? n43373 : n41481;
  assign n43571 = pi16 ? n20208 : ~n43519;
  assign n43572 = pi15 ? n43571 : n43521;
  assign n43573 = pi14 ? n43570 : n43572;
  assign n43574 = pi16 ? n1135 : ~n1577;
  assign n43575 = pi15 ? n43525 : n43574;
  assign n43576 = pi16 ? n20208 : ~n1577;
  assign n43577 = pi16 ? n1233 : ~n1577;
  assign n43578 = pi15 ? n43576 : n43577;
  assign n43579 = pi14 ? n43575 : n43578;
  assign n43580 = pi13 ? n43573 : n43579;
  assign n43581 = pi12 ? n43569 : n43580;
  assign n43582 = pi11 ? n43566 : n43581;
  assign n43583 = pi10 ? n43564 : n43582;
  assign n43584 = pi09 ? n32 : n43583;
  assign n43585 = pi08 ? n43536 : n43584;
  assign n43586 = pi07 ? n43462 : n43585;
  assign n43587 = pi14 ? n19970 : n180;
  assign n43588 = pi13 ? n43587 : n30395;
  assign n43589 = pi14 ? n32 : n180;
  assign n43590 = pi18 ? n18710 : ~n6641;
  assign n43591 = pi17 ? n32 : n43590;
  assign n43592 = pi18 ? n34283 : n430;
  assign n43593 = pi17 ? n18487 : ~n43592;
  assign n43594 = pi16 ? n43591 : n43593;
  assign n43595 = pi15 ? n180 : n43594;
  assign n43596 = pi19 ? n507 : n6303;
  assign n43597 = pi20 ? n1324 : n2180;
  assign n43598 = pi19 ? n43597 : n1076;
  assign n43599 = pi18 ? n43596 : n43598;
  assign n43600 = pi19 ? n6398 : n267;
  assign n43601 = pi18 ? n43600 : ~n289;
  assign n43602 = pi17 ? n43599 : n43601;
  assign n43603 = pi16 ? n32 : n43602;
  assign n43604 = pi15 ? n17885 : n43603;
  assign n43605 = pi14 ? n43595 : n43604;
  assign n43606 = pi13 ? n43589 : n43605;
  assign n43607 = pi12 ? n43588 : n43606;
  assign n43608 = pi20 ? n17665 : ~n287;
  assign n43609 = pi19 ? n32 : n43608;
  assign n43610 = pi20 ? n1076 : n9194;
  assign n43611 = pi20 ? n1368 : n1076;
  assign n43612 = pi19 ? n43610 : n43611;
  assign n43613 = pi18 ? n43609 : n43612;
  assign n43614 = pi19 ? n1464 : n275;
  assign n43615 = pi18 ? n43614 : n19811;
  assign n43616 = pi17 ? n43613 : n43615;
  assign n43617 = pi16 ? n32 : n43616;
  assign n43618 = pi18 ? n30775 : n248;
  assign n43619 = pi17 ? n23052 : n43618;
  assign n43620 = pi16 ? n32 : n43619;
  assign n43621 = pi15 ? n43617 : n43620;
  assign n43622 = pi19 ? n342 : n18396;
  assign n43623 = pi18 ? n10078 : n43622;
  assign n43624 = pi19 ? n11879 : ~n30681;
  assign n43625 = pi18 ? n43624 : n4689;
  assign n43626 = pi17 ? n43623 : n43625;
  assign n43627 = pi16 ? n32 : n43626;
  assign n43628 = pi19 ? n617 : n247;
  assign n43629 = pi18 ? n32 : ~n43628;
  assign n43630 = pi18 ? n9012 : n2304;
  assign n43631 = pi17 ? n43629 : ~n43630;
  assign n43632 = pi16 ? n32 : n43631;
  assign n43633 = pi15 ? n43627 : n43632;
  assign n43634 = pi14 ? n43621 : n43633;
  assign n43635 = pi17 ? n2733 : ~n2305;
  assign n43636 = pi16 ? n32 : n43635;
  assign n43637 = pi20 ? n2385 : n339;
  assign n43638 = pi19 ? n32 : n43637;
  assign n43639 = pi18 ? n32 : n43638;
  assign n43640 = pi19 ? n32 : n18575;
  assign n43641 = pi21 ? n174 : n1939;
  assign n43642 = pi20 ? n43641 : ~n32;
  assign n43643 = pi19 ? n43642 : ~n32;
  assign n43644 = pi18 ? n43640 : n43643;
  assign n43645 = pi17 ? n43639 : ~n43644;
  assign n43646 = pi16 ? n32 : n43645;
  assign n43647 = pi15 ? n43636 : n43646;
  assign n43648 = pi20 ? n2385 : n915;
  assign n43649 = pi19 ? n43648 : n30400;
  assign n43650 = pi18 ? n43649 : n20249;
  assign n43651 = pi17 ? n32 : n43650;
  assign n43652 = pi16 ? n32 : n43651;
  assign n43653 = pi20 ? n175 : n18832;
  assign n43654 = pi19 ? n32 : n43653;
  assign n43655 = pi18 ? n32 : n43654;
  assign n43656 = pi20 ? n339 : ~n18129;
  assign n43657 = pi20 ? n1368 : n9194;
  assign n43658 = pi19 ? n43656 : ~n43657;
  assign n43659 = pi18 ? n43658 : ~n43643;
  assign n43660 = pi17 ? n43655 : n43659;
  assign n43661 = pi16 ? n32 : n43660;
  assign n43662 = pi15 ? n43652 : n43661;
  assign n43663 = pi14 ? n43647 : n43662;
  assign n43664 = pi13 ? n43634 : n43663;
  assign n43665 = pi18 ? n32 : n1054;
  assign n43666 = pi18 ? n858 : n2304;
  assign n43667 = pi17 ? n43665 : ~n43666;
  assign n43668 = pi16 ? n32 : n43667;
  assign n43669 = pi15 ? n43668 : n19531;
  assign n43670 = pi19 ? n1325 : n311;
  assign n43671 = pi19 ? n10863 : n32;
  assign n43672 = pi18 ? n43670 : n43671;
  assign n43673 = pi17 ? n32 : n43672;
  assign n43674 = pi16 ? n32 : n43673;
  assign n43675 = pi15 ? n20636 : n43674;
  assign n43676 = pi14 ? n43669 : n43675;
  assign n43677 = pi19 ? n1325 : n23193;
  assign n43678 = pi18 ? n43677 : n19933;
  assign n43679 = pi17 ? n32 : n43678;
  assign n43680 = pi16 ? n32 : n43679;
  assign n43681 = pi19 ? n30521 : n28356;
  assign n43682 = pi18 ? n43681 : n6059;
  assign n43683 = pi17 ? n32 : n43682;
  assign n43684 = pi16 ? n32 : n43683;
  assign n43685 = pi15 ? n43680 : n43684;
  assign n43686 = pi15 ? n19235 : n19942;
  assign n43687 = pi14 ? n43685 : n43686;
  assign n43688 = pi13 ? n43676 : n43687;
  assign n43689 = pi12 ? n43664 : n43688;
  assign n43690 = pi11 ? n43607 : n43689;
  assign n43691 = pi13 ? n30440 : n32;
  assign n43692 = pi12 ? n43691 : n32;
  assign n43693 = pi15 ? n43526 : n28947;
  assign n43694 = pi15 ? n18979 : n31707;
  assign n43695 = pi14 ? n43693 : n43694;
  assign n43696 = pi16 ? n32 : n29752;
  assign n43697 = pi17 ? n19907 : n32;
  assign n43698 = pi16 ? n568 : n43697;
  assign n43699 = pi15 ? n32 : n43698;
  assign n43700 = pi14 ? n43696 : n43699;
  assign n43701 = pi13 ? n43695 : n43700;
  assign n43702 = pi15 ? n43516 : n30473;
  assign n43703 = pi15 ? n30477 : n18979;
  assign n43704 = pi14 ? n43702 : n43703;
  assign n43705 = pi17 ? n30475 : n2133;
  assign n43706 = pi16 ? n1135 : ~n43705;
  assign n43707 = pi17 ? n32 : n2133;
  assign n43708 = pi16 ? n1135 : ~n43707;
  assign n43709 = pi15 ? n43706 : n43708;
  assign n43710 = pi15 ? n18979 : n19100;
  assign n43711 = pi14 ? n43709 : n43710;
  assign n43712 = pi13 ? n43704 : n43711;
  assign n43713 = pi12 ? n43701 : n43712;
  assign n43714 = pi11 ? n43692 : n43713;
  assign n43715 = pi10 ? n43690 : n43714;
  assign n43716 = pi09 ? n32 : n43715;
  assign n43717 = pi14 ? n32 : n13392;
  assign n43718 = pi18 ? n34283 : n2298;
  assign n43719 = pi17 ? n18487 : ~n43718;
  assign n43720 = pi16 ? n43591 : n43719;
  assign n43721 = pi15 ? n13392 : n43720;
  assign n43722 = pi18 ? n30406 : n32;
  assign n43723 = pi17 ? n18006 : n43722;
  assign n43724 = pi16 ? n32 : n43723;
  assign n43725 = pi15 ? n43724 : n43603;
  assign n43726 = pi14 ? n43721 : n43725;
  assign n43727 = pi13 ? n43717 : n43726;
  assign n43728 = pi12 ? n43588 : n43727;
  assign n43729 = pi19 ? n16289 : n32;
  assign n43730 = pi18 ? n30775 : n43729;
  assign n43731 = pi17 ? n23052 : n43730;
  assign n43732 = pi16 ? n32 : n43731;
  assign n43733 = pi15 ? n43617 : n43732;
  assign n43734 = pi18 ? n9012 : n344;
  assign n43735 = pi17 ? n43629 : ~n43734;
  assign n43736 = pi16 ? n32 : n43735;
  assign n43737 = pi15 ? n43627 : n43736;
  assign n43738 = pi14 ? n43733 : n43737;
  assign n43739 = pi20 ? n342 : n18415;
  assign n43740 = pi19 ? n32 : n43739;
  assign n43741 = pi18 ? n32 : n43740;
  assign n43742 = pi20 ? n18073 : n18282;
  assign n43743 = pi20 ? n18282 : n17665;
  assign n43744 = pi19 ? n43742 : n43743;
  assign n43745 = pi18 ? n43744 : ~n30130;
  assign n43746 = pi17 ? n43741 : ~n43745;
  assign n43747 = pi16 ? n32 : n43746;
  assign n43748 = pi15 ? n43636 : n43747;
  assign n43749 = pi20 ? n13171 : ~n29452;
  assign n43750 = pi19 ? n43749 : ~n30501;
  assign n43751 = pi18 ? n43750 : ~n20249;
  assign n43752 = pi17 ? n30499 : ~n43751;
  assign n43753 = pi16 ? n32 : n43752;
  assign n43754 = pi20 ? n1368 : n17665;
  assign n43755 = pi19 ? n43656 : ~n43754;
  assign n43756 = pi19 ? n4558 : ~n32;
  assign n43757 = pi18 ? n43755 : ~n43756;
  assign n43758 = pi17 ? n43655 : n43757;
  assign n43759 = pi16 ? n32 : n43758;
  assign n43760 = pi15 ? n43753 : n43759;
  assign n43761 = pi14 ? n43748 : n43760;
  assign n43762 = pi13 ? n43738 : n43761;
  assign n43763 = pi17 ? n43665 : ~n2305;
  assign n43764 = pi16 ? n32 : n43763;
  assign n43765 = pi19 ? n7449 : n32;
  assign n43766 = pi18 ? n32 : n43765;
  assign n43767 = pi17 ? n32 : n43766;
  assign n43768 = pi16 ? n32 : n43767;
  assign n43769 = pi15 ? n43764 : n43768;
  assign n43770 = pi18 ? n43670 : n30514;
  assign n43771 = pi17 ? n32 : n43770;
  assign n43772 = pi16 ? n32 : n43771;
  assign n43773 = pi15 ? n20636 : n43772;
  assign n43774 = pi14 ? n43769 : n43773;
  assign n43775 = pi18 ? n43677 : n4689;
  assign n43776 = pi17 ? n32 : n43775;
  assign n43777 = pi16 ? n32 : n43776;
  assign n43778 = pi15 ? n43777 : n43684;
  assign n43779 = pi15 ? n19384 : n20157;
  assign n43780 = pi14 ? n43778 : n43779;
  assign n43781 = pi13 ? n43774 : n43780;
  assign n43782 = pi12 ? n43762 : n43781;
  assign n43783 = pi11 ? n43728 : n43782;
  assign n43784 = pi13 ? n30545 : n32;
  assign n43785 = pi12 ? n43784 : n32;
  assign n43786 = pi15 ? n43529 : n30025;
  assign n43787 = pi16 ? n1233 : ~n2326;
  assign n43788 = pi15 ? n19100 : n43787;
  assign n43789 = pi14 ? n43786 : n43788;
  assign n43790 = pi16 ? n919 : n43697;
  assign n43791 = pi15 ? n32 : n43790;
  assign n43792 = pi14 ? n43696 : n43791;
  assign n43793 = pi13 ? n43789 : n43792;
  assign n43794 = pi15 ? n41621 : n30556;
  assign n43795 = pi14 ? n43794 : n43703;
  assign n43796 = pi13 ? n43795 : n43711;
  assign n43797 = pi12 ? n43793 : n43796;
  assign n43798 = pi11 ? n43785 : n43797;
  assign n43799 = pi10 ? n43783 : n43798;
  assign n43800 = pi09 ? n32 : n43799;
  assign n43801 = pi08 ? n43716 : n43800;
  assign n43802 = pi14 ? n32926 : n19976;
  assign n43803 = pi14 ? n19969 : n32;
  assign n43804 = pi13 ? n43802 : n43803;
  assign n43805 = pi15 ? n19969 : n20236;
  assign n43806 = pi14 ? n32 : n43805;
  assign n43807 = pi18 ? n940 : ~n6641;
  assign n43808 = pi17 ? n32 : n43807;
  assign n43809 = pi18 ? n34283 : n2304;
  assign n43810 = pi17 ? n18487 : ~n43809;
  assign n43811 = pi16 ? n43808 : n43810;
  assign n43812 = pi15 ? n20236 : n43811;
  assign n43813 = pi19 ? n857 : n41313;
  assign n43814 = pi20 ? n2358 : n17669;
  assign n43815 = pi19 ? n502 : n43814;
  assign n43816 = pi18 ? n43813 : ~n43815;
  assign n43817 = pi19 ? n28774 : ~n28076;
  assign n43818 = pi18 ? n43817 : n3508;
  assign n43819 = pi17 ? n43816 : ~n43818;
  assign n43820 = pi16 ? n32 : n43819;
  assign n43821 = pi15 ? n19805 : n43820;
  assign n43822 = pi14 ? n43812 : n43821;
  assign n43823 = pi13 ? n43806 : n43822;
  assign n43824 = pi12 ? n43804 : n43823;
  assign n43825 = pi20 ? n820 : n18261;
  assign n43826 = pi19 ? n6683 : n43825;
  assign n43827 = pi18 ? n37005 : ~n43826;
  assign n43828 = pi20 ? n17669 : n6050;
  assign n43829 = pi19 ? n43828 : n30984;
  assign n43830 = pi18 ? n43829 : ~n5856;
  assign n43831 = pi17 ? n43827 : ~n43830;
  assign n43832 = pi16 ? n32 : n43831;
  assign n43833 = pi20 ? n18073 : n18281;
  assign n43834 = pi19 ? n594 : n43833;
  assign n43835 = pi20 ? n17652 : n314;
  assign n43836 = pi19 ? n43835 : ~n20933;
  assign n43837 = pi18 ? n43834 : n43836;
  assign n43838 = pi20 ? n17671 : n32;
  assign n43839 = pi19 ? n43742 : n43838;
  assign n43840 = pi18 ? n43839 : n430;
  assign n43841 = pi17 ? n43837 : ~n43840;
  assign n43842 = pi16 ? n32 : n43841;
  assign n43843 = pi15 ? n43832 : n43842;
  assign n43844 = pi19 ? n32 : n1076;
  assign n43845 = pi20 ? n342 : n18253;
  assign n43846 = pi19 ? n43845 : n41294;
  assign n43847 = pi18 ? n43844 : n43846;
  assign n43848 = pi20 ? n18245 : n32;
  assign n43849 = pi19 ? n43848 : n32;
  assign n43850 = pi18 ? n43744 : ~n43849;
  assign n43851 = pi17 ? n43847 : ~n43850;
  assign n43852 = pi16 ? n32 : n43851;
  assign n43853 = pi19 ? n1369 : ~n9169;
  assign n43854 = pi18 ? n32 : n43853;
  assign n43855 = pi18 ? n9012 : n430;
  assign n43856 = pi17 ? n43854 : ~n43855;
  assign n43857 = pi16 ? n32 : n43856;
  assign n43858 = pi15 ? n43852 : n43857;
  assign n43859 = pi14 ? n43843 : n43858;
  assign n43860 = pi17 ? n2726 : ~n2410;
  assign n43861 = pi16 ? n32 : n43860;
  assign n43862 = pi19 ? n43742 : n31309;
  assign n43863 = pi18 ? n43862 : n20525;
  assign n43864 = pi17 ? n30283 : ~n43863;
  assign n43865 = pi16 ? n32 : n43864;
  assign n43866 = pi15 ? n43861 : n43865;
  assign n43867 = pi19 ? n1817 : n5854;
  assign n43868 = pi18 ? n43867 : n20525;
  assign n43869 = pi17 ? n30283 : ~n43868;
  assign n43870 = pi16 ? n32 : n43869;
  assign n43871 = pi20 ? n2180 : n17665;
  assign n43872 = pi19 ? n30593 : ~n43871;
  assign n43873 = pi18 ? n43872 : n43849;
  assign n43874 = pi17 ? n3282 : n43873;
  assign n43875 = pi16 ? n32 : n43874;
  assign n43876 = pi15 ? n43870 : n43875;
  assign n43877 = pi14 ? n43866 : n43876;
  assign n43878 = pi13 ? n43859 : n43877;
  assign n43879 = pi17 ? n3164 : ~n33153;
  assign n43880 = pi16 ? n32 : n43879;
  assign n43881 = pi19 ? n7435 : n32;
  assign n43882 = pi18 ? n32 : n43881;
  assign n43883 = pi17 ? n32 : n43882;
  assign n43884 = pi16 ? n32 : n43883;
  assign n43885 = pi15 ? n43880 : n43884;
  assign n43886 = pi19 ? n1464 : n462;
  assign n43887 = pi18 ? n43886 : n4689;
  assign n43888 = pi17 ? n32 : n43887;
  assign n43889 = pi16 ? n32 : n43888;
  assign n43890 = pi15 ? n43777 : n43889;
  assign n43891 = pi14 ? n43885 : n43890;
  assign n43892 = pi19 ? n6057 : n23193;
  assign n43893 = pi18 ? n43892 : n4689;
  assign n43894 = pi17 ? n32 : n43893;
  assign n43895 = pi16 ? n32 : n43894;
  assign n43896 = pi19 ? n2386 : ~n247;
  assign n43897 = pi18 ? n43896 : ~n350;
  assign n43898 = pi17 ? n32 : n43897;
  assign n43899 = pi16 ? n32 : n43898;
  assign n43900 = pi15 ? n43895 : n43899;
  assign n43901 = pi15 ? n17637 : n30610;
  assign n43902 = pi14 ? n43900 : n43901;
  assign n43903 = pi13 ? n43891 : n43902;
  assign n43904 = pi12 ? n43878 : n43903;
  assign n43905 = pi11 ? n43824 : n43904;
  assign n43906 = pi14 ? n30620 : n32;
  assign n43907 = pi13 ? n43906 : n32;
  assign n43908 = pi12 ? n43907 : n32;
  assign n43909 = pi18 ? n32 : ~n18532;
  assign n43910 = pi17 ? n20021 : n43909;
  assign n43911 = pi16 ? n1135 : ~n43910;
  assign n43912 = pi17 ? n20021 : n2325;
  assign n43913 = pi16 ? n1135 : ~n43912;
  assign n43914 = pi15 ? n43911 : n43913;
  assign n43915 = pi14 ? n18979 : n43914;
  assign n43916 = pi17 ? n20031 : n32;
  assign n43917 = pi16 ? n465 : n43916;
  assign n43918 = pi16 ? n919 : n30736;
  assign n43919 = pi15 ? n32 : n43918;
  assign n43920 = pi14 ? n43917 : n43919;
  assign n43921 = pi13 ? n43915 : n43920;
  assign n43922 = pi15 ? n19711 : n30657;
  assign n43923 = pi18 ? n936 : n3350;
  assign n43924 = pi17 ? n32 : n43923;
  assign n43925 = pi16 ? n1214 : ~n43924;
  assign n43926 = pi15 ? n30663 : n43925;
  assign n43927 = pi14 ? n43922 : n43926;
  assign n43928 = pi17 ? n32752 : n43923;
  assign n43929 = pi16 ? n1214 : ~n43928;
  assign n43930 = pi17 ? n32 : n2433;
  assign n43931 = pi16 ? n1135 : ~n43930;
  assign n43932 = pi15 ? n43929 : n43931;
  assign n43933 = pi16 ? n1233 : ~n3356;
  assign n43934 = pi15 ? n41490 : n43933;
  assign n43935 = pi14 ? n43932 : n43934;
  assign n43936 = pi13 ? n43927 : n43935;
  assign n43937 = pi12 ? n43921 : n43936;
  assign n43938 = pi11 ? n43908 : n43937;
  assign n43939 = pi10 ? n43905 : n43938;
  assign n43940 = pi09 ? n32 : n43939;
  assign n43941 = pi15 ? n106 : n20048;
  assign n43942 = pi14 ? n32 : n43941;
  assign n43943 = pi16 ? n43808 : n43593;
  assign n43944 = pi15 ? n19972 : n43943;
  assign n43945 = pi18 ? n43817 : n19740;
  assign n43946 = pi17 ? n43816 : ~n43945;
  assign n43947 = pi16 ? n32 : n43946;
  assign n43948 = pi15 ? n20531 : n43947;
  assign n43949 = pi14 ? n43944 : n43948;
  assign n43950 = pi13 ? n43942 : n43949;
  assign n43951 = pi12 ? n43804 : n43950;
  assign n43952 = pi18 ? n43829 : ~n22411;
  assign n43953 = pi17 ? n43827 : ~n43952;
  assign n43954 = pi16 ? n32 : n43953;
  assign n43955 = pi20 ? n9641 : n18282;
  assign n43956 = pi19 ? n594 : n43955;
  assign n43957 = pi19 ? n41289 : ~n9488;
  assign n43958 = pi18 ? n43956 : n43957;
  assign n43959 = pi19 ? n43742 : n28750;
  assign n43960 = pi18 ? n43959 : n19740;
  assign n43961 = pi17 ? n43958 : ~n43960;
  assign n43962 = pi16 ? n32 : n43961;
  assign n43963 = pi15 ? n43954 : n43962;
  assign n43964 = pi14 ? n43963 : n43858;
  assign n43965 = pi19 ? n43742 : n31183;
  assign n43966 = pi18 ? n43965 : n30702;
  assign n43967 = pi17 ? n30698 : ~n43966;
  assign n43968 = pi16 ? n32 : n43967;
  assign n43969 = pi15 ? n43861 : n43968;
  assign n43970 = pi20 ? n6303 : n1817;
  assign n43971 = pi19 ? n1817 : n43970;
  assign n43972 = pi18 ? n43971 : n30702;
  assign n43973 = pi17 ? n30283 : ~n43972;
  assign n43974 = pi16 ? n32 : n43973;
  assign n43975 = pi20 ? n354 : ~n18129;
  assign n43976 = pi19 ? n43975 : ~n43754;
  assign n43977 = pi18 ? n43976 : ~n30702;
  assign n43978 = pi17 ? n36054 : n43977;
  assign n43979 = pi16 ? n32 : n43978;
  assign n43980 = pi15 ? n43974 : n43979;
  assign n43981 = pi14 ? n43969 : n43980;
  assign n43982 = pi13 ? n43964 : n43981;
  assign n43983 = pi18 ? n43886 : n20320;
  assign n43984 = pi17 ? n32 : n43983;
  assign n43985 = pi16 ? n32 : n43984;
  assign n43986 = pi15 ? n43777 : n43985;
  assign n43987 = pi14 ? n43885 : n43986;
  assign n43988 = pi18 ? n43892 : n20249;
  assign n43989 = pi17 ? n32 : n43988;
  assign n43990 = pi16 ? n32 : n43989;
  assign n43991 = pi15 ? n43990 : n43899;
  assign n43992 = pi14 ? n43991 : n43901;
  assign n43993 = pi13 ? n43987 : n43992;
  assign n43994 = pi12 ? n43982 : n43993;
  assign n43995 = pi11 ? n43951 : n43994;
  assign n43996 = pi14 ? n30727 : n32;
  assign n43997 = pi13 ? n43996 : n32;
  assign n43998 = pi12 ? n43997 : n32;
  assign n43999 = pi16 ? n1233 : ~n43912;
  assign n44000 = pi15 ? n43911 : n43999;
  assign n44001 = pi14 ? n18979 : n44000;
  assign n44002 = pi16 ? n1014 : n43916;
  assign n44003 = pi14 ? n44002 : n43919;
  assign n44004 = pi13 ? n44001 : n44003;
  assign n44005 = pi16 ? n1214 : ~n43930;
  assign n44006 = pi15 ? n30743 : n44005;
  assign n44007 = pi14 ? n43922 : n44006;
  assign n44008 = pi17 ? n32752 : n2433;
  assign n44009 = pi16 ? n1214 : ~n44008;
  assign n44010 = pi15 ? n44009 : n43931;
  assign n44011 = pi14 ? n44010 : n43934;
  assign n44012 = pi13 ? n44007 : n44011;
  assign n44013 = pi12 ? n44004 : n44012;
  assign n44014 = pi11 ? n43998 : n44013;
  assign n44015 = pi10 ? n43995 : n44014;
  assign n44016 = pi09 ? n32 : n44015;
  assign n44017 = pi08 ? n43940 : n44016;
  assign n44018 = pi07 ? n43801 : n44017;
  assign n44019 = pi06 ? n43586 : n44018;
  assign n44020 = pi05 ? n43295 : n44019;
  assign n44021 = pi15 ? n13380 : n20692;
  assign n44022 = pi14 ? n20297 : n44021;
  assign n44023 = pi14 ? n30981 : n32;
  assign n44024 = pi13 ? n44022 : n44023;
  assign n44025 = pi14 ? n32 : n20048;
  assign n44026 = pi20 ? n17652 : ~n448;
  assign n44027 = pi19 ? n32 : n44026;
  assign n44028 = pi18 ? n127 : n44027;
  assign n44029 = pi17 ? n32 : n44028;
  assign n44030 = pi16 ? n44029 : ~n3625;
  assign n44031 = pi18 ? n276 : n1758;
  assign n44032 = pi17 ? n32 : n44031;
  assign n44033 = pi16 ? n44032 : ~n2530;
  assign n44034 = pi15 ? n44030 : n44033;
  assign n44035 = pi20 ? n17652 : ~n6085;
  assign n44036 = pi19 ? n594 : n44035;
  assign n44037 = pi19 ? n28823 : n28826;
  assign n44038 = pi18 ? n44036 : ~n44037;
  assign n44039 = pi19 ? n32 : n31723;
  assign n44040 = pi18 ? n44039 : n19740;
  assign n44041 = pi17 ? n44038 : ~n44040;
  assign n44042 = pi16 ? n32 : n44041;
  assign n44043 = pi20 ? n1076 : n785;
  assign n44044 = pi19 ? n32 : n44043;
  assign n44045 = pi20 ? n6050 : n207;
  assign n44046 = pi19 ? n44045 : ~n32;
  assign n44047 = pi18 ? n44044 : n44046;
  assign n44048 = pi17 ? n44047 : ~n2410;
  assign n44049 = pi16 ? n32 : n44048;
  assign n44050 = pi15 ? n44042 : n44049;
  assign n44051 = pi14 ? n44034 : n44050;
  assign n44052 = pi13 ? n44025 : n44051;
  assign n44053 = pi12 ? n44024 : n44052;
  assign n44054 = pi18 ? n17118 : n2360;
  assign n44055 = pi17 ? n44054 : ~n1933;
  assign n44056 = pi16 ? n32 : n44055;
  assign n44057 = pi19 ? n246 : ~n207;
  assign n44058 = pi18 ? n32 : n44057;
  assign n44059 = pi17 ? n32 : n44058;
  assign n44060 = pi19 ? n22501 : ~n17749;
  assign n44061 = pi19 ? n37542 : ~n236;
  assign n44062 = pi18 ? n44060 : n44061;
  assign n44063 = pi17 ? n44062 : n2410;
  assign n44064 = pi16 ? n44059 : ~n44063;
  assign n44065 = pi15 ? n44056 : n44064;
  assign n44066 = pi17 ? n3067 : ~n2410;
  assign n44067 = pi16 ? n32 : n44066;
  assign n44068 = pi19 ? n17757 : n342;
  assign n44069 = pi18 ? n32 : n44068;
  assign n44070 = pi17 ? n32 : n44069;
  assign n44071 = pi19 ? n18396 : n28685;
  assign n44072 = pi19 ? n18478 : n247;
  assign n44073 = pi18 ? n44071 : ~n44072;
  assign n44074 = pi17 ? n44073 : ~n2299;
  assign n44075 = pi16 ? n44070 : n44074;
  assign n44076 = pi15 ? n44067 : n44075;
  assign n44077 = pi14 ? n44065 : n44076;
  assign n44078 = pi20 ? n354 : ~n175;
  assign n44079 = pi19 ? n44078 : ~n176;
  assign n44080 = pi18 ? n44079 : ~n2298;
  assign n44081 = pi17 ? n36054 : n44080;
  assign n44082 = pi16 ? n32 : n44081;
  assign n44083 = pi17 ? n2954 : ~n2410;
  assign n44084 = pi16 ? n32 : n44083;
  assign n44085 = pi15 ? n44082 : n44084;
  assign n44086 = pi17 ? n32 : n33062;
  assign n44087 = pi16 ? n32 : n44086;
  assign n44088 = pi18 ? n344 : ~n344;
  assign n44089 = pi17 ? n32 : n44088;
  assign n44090 = pi16 ? n32 : n44089;
  assign n44091 = pi15 ? n44087 : n44090;
  assign n44092 = pi14 ? n44085 : n44091;
  assign n44093 = pi13 ? n44077 : n44092;
  assign n44094 = pi18 ? n858 : n19853;
  assign n44095 = pi17 ? n32 : n44094;
  assign n44096 = pi16 ? n32 : n44095;
  assign n44097 = pi15 ? n33042 : n44096;
  assign n44098 = pi20 ? n2358 : ~n18624;
  assign n44099 = pi19 ? n32 : ~n44098;
  assign n44100 = pi18 ? n44099 : ~n20267;
  assign n44101 = pi17 ? n32 : n44100;
  assign n44102 = pi16 ? n32 : n44101;
  assign n44103 = pi15 ? n44096 : n44102;
  assign n44104 = pi14 ? n44097 : n44103;
  assign n44105 = pi19 ? n594 : n246;
  assign n44106 = pi18 ? n44105 : n20366;
  assign n44107 = pi17 ? n16450 : n44106;
  assign n44108 = pi16 ? n32 : n44107;
  assign n44109 = pi20 ? n18282 : n5854;
  assign n44110 = pi19 ? n594 : n44109;
  assign n44111 = pi20 ? n18834 : ~n32;
  assign n44112 = pi19 ? n44111 : ~n32;
  assign n44113 = pi18 ? n44110 : ~n44112;
  assign n44114 = pi17 ? n16317 : n44113;
  assign n44115 = pi16 ? n32 : n44114;
  assign n44116 = pi15 ? n44108 : n44115;
  assign n44117 = pi18 ? n4127 : n4689;
  assign n44118 = pi17 ? n32 : n44117;
  assign n44119 = pi16 ? n32 : n44118;
  assign n44120 = pi15 ? n44119 : n30799;
  assign n44121 = pi14 ? n44116 : n44120;
  assign n44122 = pi13 ? n44104 : n44121;
  assign n44123 = pi12 ? n44093 : n44122;
  assign n44124 = pi11 ? n44053 : n44123;
  assign n44125 = pi18 ? n4392 : ~n31385;
  assign n44126 = pi17 ? n32 : n44125;
  assign n44127 = pi16 ? n32 : n44126;
  assign n44128 = pi15 ? n44127 : n32;
  assign n44129 = pi14 ? n44128 : n32;
  assign n44130 = pi13 ? n44129 : n32;
  assign n44131 = pi18 ? n1819 : n274;
  assign n44132 = pi17 ? n32 : n44131;
  assign n44133 = pi19 ? n339 : n44078;
  assign n44134 = pi20 ? n1817 : n174;
  assign n44135 = pi20 ? n174 : n246;
  assign n44136 = pi19 ? n44134 : n44135;
  assign n44137 = pi18 ? n44133 : ~n44136;
  assign n44138 = pi20 ? n259 : ~n6621;
  assign n44139 = pi20 ? n1817 : n6621;
  assign n44140 = pi19 ? n44138 : ~n44139;
  assign n44141 = pi18 ? n44140 : ~n32;
  assign n44142 = pi17 ? n44137 : n44141;
  assign n44143 = pi16 ? n44132 : ~n44142;
  assign n44144 = pi15 ? n18890 : n44143;
  assign n44145 = pi14 ? n32 : n44144;
  assign n44146 = pi13 ? n32 : n44145;
  assign n44147 = pi12 ? n44130 : n44146;
  assign n44148 = pi17 ? n20173 : n2325;
  assign n44149 = pi16 ? n1135 : ~n44148;
  assign n44150 = pi18 ? n19350 : ~n32;
  assign n44151 = pi17 ? n20183 : n44150;
  assign n44152 = pi16 ? n1135 : ~n44151;
  assign n44153 = pi15 ? n44149 : n44152;
  assign n44154 = pi18 ? n20189 : ~n32;
  assign n44155 = pi17 ? n20188 : n44154;
  assign n44156 = pi16 ? n1135 : ~n44155;
  assign n44157 = pi18 ? n20193 : n18532;
  assign n44158 = pi17 ? n10245 : n44157;
  assign n44159 = pi16 ? n1135 : n44158;
  assign n44160 = pi15 ? n44156 : n44159;
  assign n44161 = pi14 ? n44153 : n44160;
  assign n44162 = pi17 ? n20200 : n32;
  assign n44163 = pi16 ? n465 : n44162;
  assign n44164 = pi17 ? n20200 : n19170;
  assign n44165 = pi16 ? n465 : n44164;
  assign n44166 = pi15 ? n44163 : n44165;
  assign n44167 = pi17 ? n20209 : n17901;
  assign n44168 = pi16 ? n270 : n44167;
  assign n44169 = pi15 ? n44168 : n31707;
  assign n44170 = pi14 ? n44166 : n44169;
  assign n44171 = pi13 ? n44161 : n44170;
  assign n44172 = pi16 ? n1214 : ~n30875;
  assign n44173 = pi15 ? n44172 : n19711;
  assign n44174 = pi14 ? n44173 : n19711;
  assign n44175 = pi15 ? n44005 : n41481;
  assign n44176 = pi16 ? n1471 : ~n3356;
  assign n44177 = pi15 ? n44176 : n43933;
  assign n44178 = pi14 ? n44175 : n44177;
  assign n44179 = pi13 ? n44174 : n44178;
  assign n44180 = pi12 ? n44171 : n44179;
  assign n44181 = pi11 ? n44147 : n44180;
  assign n44182 = pi10 ? n44124 : n44181;
  assign n44183 = pi09 ? n32 : n44182;
  assign n44184 = pi14 ? n20297 : n13684;
  assign n44185 = pi20 ? n17652 : n501;
  assign n44186 = pi19 ? n32 : n44185;
  assign n44187 = pi18 ? n32 : n44186;
  assign n44188 = pi17 ? n32 : n44187;
  assign n44189 = pi16 ? n44188 : ~n3788;
  assign n44190 = pi17 ? n32 : n7396;
  assign n44191 = pi16 ? n44190 : ~n2530;
  assign n44192 = pi15 ? n44189 : n44191;
  assign n44193 = pi20 ? n333 : ~n9491;
  assign n44194 = pi19 ? n32 : n44193;
  assign n44195 = pi20 ? n18253 : n9194;
  assign n44196 = pi20 ? n9194 : n18073;
  assign n44197 = pi19 ? n44195 : n44196;
  assign n44198 = pi18 ? n44194 : ~n44197;
  assign n44199 = pi20 ? n333 : ~n18253;
  assign n44200 = pi20 ? n18253 : n18832;
  assign n44201 = pi19 ? n44199 : ~n44200;
  assign n44202 = pi18 ? n44201 : n19740;
  assign n44203 = pi17 ? n44198 : ~n44202;
  assign n44204 = pi16 ? n32 : n44203;
  assign n44205 = pi15 ? n44204 : n44049;
  assign n44206 = pi14 ? n44192 : n44205;
  assign n44207 = pi13 ? n44184 : n44206;
  assign n44208 = pi12 ? n44024 : n44207;
  assign n44209 = pi17 ? n3067 : ~n2299;
  assign n44210 = pi16 ? n32 : n44209;
  assign n44211 = pi15 ? n44210 : n44075;
  assign n44212 = pi14 ? n44065 : n44211;
  assign n44213 = pi19 ? n44078 : ~n43754;
  assign n44214 = pi20 ? n23668 : ~n32;
  assign n44215 = pi19 ? n44214 : ~n32;
  assign n44216 = pi18 ? n44213 : ~n44215;
  assign n44217 = pi17 ? n36054 : n44216;
  assign n44218 = pi16 ? n32 : n44217;
  assign n44219 = pi17 ? n2954 : ~n2299;
  assign n44220 = pi16 ? n32 : n44219;
  assign n44221 = pi15 ? n44218 : n44220;
  assign n44222 = pi18 ? n344 : ~n30575;
  assign n44223 = pi17 ? n32 : n44222;
  assign n44224 = pi16 ? n32 : n44223;
  assign n44225 = pi15 ? n44087 : n44224;
  assign n44226 = pi14 ? n44221 : n44225;
  assign n44227 = pi13 ? n44212 : n44226;
  assign n44228 = pi18 ? n858 : n20615;
  assign n44229 = pi17 ? n32 : n44228;
  assign n44230 = pi16 ? n32 : n44229;
  assign n44231 = pi18 ? n44099 : ~n31385;
  assign n44232 = pi17 ? n32 : n44231;
  assign n44233 = pi16 ? n32 : n44232;
  assign n44234 = pi15 ? n44230 : n44233;
  assign n44235 = pi14 ? n44097 : n44234;
  assign n44236 = pi19 ? n594 : n30539;
  assign n44237 = pi21 ? n313 : n1939;
  assign n44238 = pi20 ? n44237 : ~n32;
  assign n44239 = pi19 ? n44238 : ~n32;
  assign n44240 = pi18 ? n44236 : ~n44239;
  assign n44241 = pi17 ? n16317 : n44240;
  assign n44242 = pi16 ? n32 : n44241;
  assign n44243 = pi15 ? n44108 : n44242;
  assign n44244 = pi18 ? n4127 : n20249;
  assign n44245 = pi17 ? n32 : n44244;
  assign n44246 = pi16 ? n32 : n44245;
  assign n44247 = pi15 ? n44246 : n30929;
  assign n44248 = pi14 ? n44243 : n44247;
  assign n44249 = pi13 ? n44235 : n44248;
  assign n44250 = pi12 ? n44227 : n44249;
  assign n44251 = pi11 ? n44208 : n44250;
  assign n44252 = pi18 ? n4392 : ~n22194;
  assign n44253 = pi17 ? n32 : n44252;
  assign n44254 = pi16 ? n32 : n44253;
  assign n44255 = pi15 ? n44254 : n32;
  assign n44256 = pi14 ? n44255 : n32;
  assign n44257 = pi13 ? n44256 : n32;
  assign n44258 = pi20 ? n32 : n6303;
  assign n44259 = pi19 ? n32 : n44258;
  assign n44260 = pi18 ? n44259 : n333;
  assign n44261 = pi17 ? n32 : n44260;
  assign n44262 = pi20 ? n18415 : n287;
  assign n44263 = pi20 ? n29457 : ~n9491;
  assign n44264 = pi19 ? n44262 : n44263;
  assign n44265 = pi20 ? n6621 : n21111;
  assign n44266 = pi19 ? n44134 : n44265;
  assign n44267 = pi18 ? n44264 : ~n44266;
  assign n44268 = pi20 ? n287 : n17669;
  assign n44269 = pi20 ? n246 : ~n17669;
  assign n44270 = pi19 ? n44268 : ~n44269;
  assign n44271 = pi18 ? n44270 : ~n32;
  assign n44272 = pi17 ? n44267 : n44271;
  assign n44273 = pi16 ? n44261 : ~n44272;
  assign n44274 = pi15 ? n32 : n44273;
  assign n44275 = pi14 ? n32 : n44274;
  assign n44276 = pi13 ? n32 : n44275;
  assign n44277 = pi12 ? n44257 : n44276;
  assign n44278 = pi16 ? n30460 : n44167;
  assign n44279 = pi15 ? n44278 : n19778;
  assign n44280 = pi14 ? n44166 : n44279;
  assign n44281 = pi13 ? n44161 : n44280;
  assign n44282 = pi16 ? n1214 : ~n30951;
  assign n44283 = pi16 ? n1214 : ~n1944;
  assign n44284 = pi15 ? n44282 : n44283;
  assign n44285 = pi17 ? n1542 : n2325;
  assign n44286 = pi16 ? n1214 : ~n44285;
  assign n44287 = pi15 ? n44286 : n19711;
  assign n44288 = pi14 ? n44284 : n44287;
  assign n44289 = pi16 ? n1233 : ~n3352;
  assign n44290 = pi15 ? n44176 : n44289;
  assign n44291 = pi14 ? n44175 : n44290;
  assign n44292 = pi13 ? n44288 : n44291;
  assign n44293 = pi12 ? n44281 : n44292;
  assign n44294 = pi11 ? n44277 : n44293;
  assign n44295 = pi10 ? n44251 : n44294;
  assign n44296 = pi09 ? n32 : n44295;
  assign n44297 = pi08 ? n44183 : n44296;
  assign n44298 = pi14 ? n20416 : n13381;
  assign n44299 = pi14 ? n146 : n32;
  assign n44300 = pi13 ? n44298 : n44299;
  assign n44301 = pi15 ? n146 : n20779;
  assign n44302 = pi14 ? n20297 : n44301;
  assign n44303 = pi20 ? n246 : ~n448;
  assign n44304 = pi19 ? n44303 : ~n358;
  assign n44305 = pi18 ? n44304 : ~n32;
  assign n44306 = pi17 ? n44305 : ~n3787;
  assign n44307 = pi16 ? n32 : n44306;
  assign n44308 = pi17 ? n1582 : ~n2299;
  assign n44309 = pi16 ? n32 : n44308;
  assign n44310 = pi15 ? n44307 : n44309;
  assign n44311 = pi20 ? n1076 : n207;
  assign n44312 = pi19 ? n507 : n44311;
  assign n44313 = pi18 ? n32 : n44312;
  assign n44314 = pi19 ? n5350 : n246;
  assign n44315 = pi18 ? n44314 : n20525;
  assign n44316 = pi17 ? n44313 : ~n44315;
  assign n44317 = pi16 ? n32 : n44316;
  assign n44318 = pi20 ? n11107 : n310;
  assign n44319 = pi19 ? n23944 : n44318;
  assign n44320 = pi18 ? n268 : n44319;
  assign n44321 = pi20 ? n5854 : ~n1611;
  assign n44322 = pi20 ? n9491 : n18832;
  assign n44323 = pi19 ? n44321 : ~n44322;
  assign n44324 = pi18 ? n44323 : ~n30986;
  assign n44325 = pi17 ? n44320 : ~n44324;
  assign n44326 = pi16 ? n32 : n44325;
  assign n44327 = pi15 ? n44317 : n44326;
  assign n44328 = pi14 ? n44310 : n44327;
  assign n44329 = pi13 ? n44302 : n44328;
  assign n44330 = pi12 ? n44300 : n44329;
  assign n44331 = pi19 ? n1464 : n31668;
  assign n44332 = pi18 ? n32 : n44331;
  assign n44333 = pi20 ? n501 : n5854;
  assign n44334 = pi19 ? n30587 : ~n44333;
  assign n44335 = pi18 ? n44334 : n33338;
  assign n44336 = pi17 ? n44332 : n44335;
  assign n44337 = pi16 ? n32 : n44336;
  assign n44338 = pi17 ? n3067 : ~n2531;
  assign n44339 = pi16 ? n32 : n44338;
  assign n44340 = pi15 ? n44337 : n44339;
  assign n44341 = pi17 ? n3164 : ~n2531;
  assign n44342 = pi16 ? n32 : n44341;
  assign n44343 = pi14 ? n44340 : n44342;
  assign n44344 = pi20 ? n175 : ~n428;
  assign n44345 = pi20 ? n974 : n3523;
  assign n44346 = pi19 ? n44344 : ~n44345;
  assign n44347 = pi19 ? n3775 : ~n32;
  assign n44348 = pi18 ? n44346 : ~n44347;
  assign n44349 = pi17 ? n32 : n44348;
  assign n44350 = pi16 ? n32 : n44349;
  assign n44351 = pi15 ? n30989 : n44350;
  assign n44352 = pi18 ? n22159 : ~n532;
  assign n44353 = pi17 ? n32 : n44352;
  assign n44354 = pi16 ? n32 : n44353;
  assign n44355 = pi15 ? n44354 : n39609;
  assign n44356 = pi14 ? n44351 : n44355;
  assign n44357 = pi13 ? n44343 : n44356;
  assign n44358 = pi18 ? n4428 : ~n423;
  assign n44359 = pi17 ? n32 : n44358;
  assign n44360 = pi16 ? n32 : n44359;
  assign n44361 = pi20 ? n29457 : n18624;
  assign n44362 = pi19 ? n594 : n44361;
  assign n44363 = pi20 ? n174 : ~n32;
  assign n44364 = pi19 ? n44363 : ~n32;
  assign n44365 = pi18 ? n44362 : ~n44364;
  assign n44366 = pi17 ? n32 : n44365;
  assign n44367 = pi16 ? n32 : n44366;
  assign n44368 = pi15 ? n44360 : n44367;
  assign n44369 = pi19 ? n32 : n44361;
  assign n44370 = pi18 ? n44369 : ~n31102;
  assign n44371 = pi17 ? n32 : n44370;
  assign n44372 = pi16 ? n32 : n44371;
  assign n44373 = pi20 ? n29457 : n287;
  assign n44374 = pi19 ? n32 : n44373;
  assign n44375 = pi18 ? n44374 : ~n30702;
  assign n44376 = pi17 ? n32 : n44375;
  assign n44377 = pi16 ? n32 : n44376;
  assign n44378 = pi15 ? n44372 : n44377;
  assign n44379 = pi14 ? n44368 : n44378;
  assign n44380 = pi18 ? n697 : ~n430;
  assign n44381 = pi17 ? n32 : n44380;
  assign n44382 = pi16 ? n32 : n44381;
  assign n44383 = pi18 ? n4127 : n19750;
  assign n44384 = pi17 ? n32 : n44383;
  assign n44385 = pi16 ? n32 : n44384;
  assign n44386 = pi15 ? n44382 : n44385;
  assign n44387 = pi15 ? n30999 : n31014;
  assign n44388 = pi14 ? n44386 : n44387;
  assign n44389 = pi13 ? n44379 : n44388;
  assign n44390 = pi12 ? n44357 : n44389;
  assign n44391 = pi11 ? n44330 : n44390;
  assign n44392 = pi15 ? n20315 : n32;
  assign n44393 = pi14 ? n44392 : n32;
  assign n44394 = pi13 ? n44393 : n32;
  assign n44395 = pi18 ? n728 : ~n342;
  assign n44396 = pi17 ? n32 : n44395;
  assign n44397 = pi19 ? n18728 : ~n5371;
  assign n44398 = pi19 ? n30849 : ~n32090;
  assign n44399 = pi18 ? n44397 : ~n44398;
  assign n44400 = pi19 ? n7642 : ~n30849;
  assign n44401 = pi18 ? n44400 : ~n19232;
  assign n44402 = pi17 ? n44399 : n44401;
  assign n44403 = pi16 ? n44396 : ~n44402;
  assign n44404 = pi15 ? n19235 : n44403;
  assign n44405 = pi14 ? n32 : n44404;
  assign n44406 = pi13 ? n32 : n44405;
  assign n44407 = pi12 ? n44394 : n44406;
  assign n44408 = pi17 ? n16103 : n2123;
  assign n44409 = pi16 ? n1233 : ~n44408;
  assign n44410 = pi18 ? n20361 : n32;
  assign n44411 = pi17 ? n20360 : ~n44410;
  assign n44412 = pi16 ? n1233 : ~n44411;
  assign n44413 = pi15 ? n44409 : n44412;
  assign n44414 = pi18 ? n20369 : n32;
  assign n44415 = pi17 ? n20367 : ~n44414;
  assign n44416 = pi16 ? n1233 : ~n44415;
  assign n44417 = pi17 ? n20373 : ~n44157;
  assign n44418 = pi16 ? n1135 : ~n44417;
  assign n44419 = pi15 ? n44416 : n44418;
  assign n44420 = pi14 ? n44413 : n44419;
  assign n44421 = pi17 ? n20381 : n32;
  assign n44422 = pi16 ? n465 : n44421;
  assign n44423 = pi17 ? n20385 : n19262;
  assign n44424 = pi16 ? n465 : n44423;
  assign n44425 = pi15 ? n44422 : n44424;
  assign n44426 = pi18 ? n209 : ~n20392;
  assign n44427 = pi17 ? n32 : n44426;
  assign n44428 = pi18 ? n20402 : n814;
  assign n44429 = pi17 ? n20399 : n44428;
  assign n44430 = pi16 ? n44427 : ~n44429;
  assign n44431 = pi15 ? n44430 : n20034;
  assign n44432 = pi14 ? n44425 : n44431;
  assign n44433 = pi13 ? n44420 : n44432;
  assign n44434 = pi17 ? n20385 : n2136;
  assign n44435 = pi16 ? n1135 : ~n44434;
  assign n44436 = pi15 ? n44435 : n20034;
  assign n44437 = pi17 ? n29699 : n2325;
  assign n44438 = pi16 ? n19652 : ~n44437;
  assign n44439 = pi15 ? n20034 : n44438;
  assign n44440 = pi14 ? n44436 : n44439;
  assign n44441 = pi15 ? n44438 : n43787;
  assign n44442 = pi16 ? n29318 : ~n2326;
  assign n44443 = pi15 ? n44442 : n43787;
  assign n44444 = pi14 ? n44441 : n44443;
  assign n44445 = pi13 ? n44440 : n44444;
  assign n44446 = pi12 ? n44433 : n44445;
  assign n44447 = pi11 ? n44407 : n44446;
  assign n44448 = pi10 ? n44391 : n44447;
  assign n44449 = pi09 ? n32 : n44448;
  assign n44450 = pi20 ? n1611 : ~n339;
  assign n44451 = pi19 ? n44450 : n32;
  assign n44452 = pi18 ? n32 : n44451;
  assign n44453 = pi17 ? n32 : n44452;
  assign n44454 = pi16 ? n32 : n44453;
  assign n44455 = pi15 ? n13952 : n44454;
  assign n44456 = pi14 ? n20416 : n44455;
  assign n44457 = pi20 ? n246 : n501;
  assign n44458 = pi19 ? n44457 : n236;
  assign n44459 = pi18 ? n44458 : ~n32;
  assign n44460 = pi17 ? n44459 : ~n2653;
  assign n44461 = pi16 ? n32 : n44460;
  assign n44462 = pi17 ? n4917 : ~n2531;
  assign n44463 = pi16 ? n32 : n44462;
  assign n44464 = pi15 ? n44461 : n44463;
  assign n44465 = pi18 ? n44314 : n20788;
  assign n44466 = pi17 ? n44313 : ~n44465;
  assign n44467 = pi16 ? n32 : n44466;
  assign n44468 = pi20 ? n18256 : n6050;
  assign n44469 = pi19 ? n23944 : n44468;
  assign n44470 = pi18 ? n268 : n44469;
  assign n44471 = pi20 ? n1817 : n6303;
  assign n44472 = pi19 ? n44471 : n333;
  assign n44473 = pi20 ? n314 : n32;
  assign n44474 = pi19 ? n44473 : n32;
  assign n44475 = pi18 ? n44472 : ~n44474;
  assign n44476 = pi17 ? n44470 : ~n44475;
  assign n44477 = pi16 ? n32 : n44476;
  assign n44478 = pi15 ? n44467 : n44477;
  assign n44479 = pi14 ? n44464 : n44478;
  assign n44480 = pi13 ? n44456 : n44479;
  assign n44481 = pi12 ? n44300 : n44480;
  assign n44482 = pi20 ? n1385 : n17669;
  assign n44483 = pi19 ? n1464 : n44482;
  assign n44484 = pi18 ? n32 : n44483;
  assign n44485 = pi20 ? n2180 : n1817;
  assign n44486 = pi19 ? n30587 : ~n44485;
  assign n44487 = pi20 ? n820 : n32;
  assign n44488 = pi19 ? n44487 : n32;
  assign n44489 = pi18 ? n44486 : n44488;
  assign n44490 = pi17 ? n44484 : n44489;
  assign n44491 = pi16 ? n32 : n44490;
  assign n44492 = pi15 ? n44491 : n44339;
  assign n44493 = pi14 ? n44492 : n44342;
  assign n44494 = pi13 ? n44493 : n44356;
  assign n44495 = pi18 ? n4428 : ~n532;
  assign n44496 = pi17 ? n32 : n44495;
  assign n44497 = pi16 ? n32 : n44496;
  assign n44498 = pi18 ? n44362 : ~n31102;
  assign n44499 = pi17 ? n32 : n44498;
  assign n44500 = pi16 ? n32 : n44499;
  assign n44501 = pi15 ? n44497 : n44500;
  assign n44502 = pi20 ? n274 : n141;
  assign n44503 = pi19 ? n44502 : ~n32;
  assign n44504 = pi18 ? n44369 : ~n44503;
  assign n44505 = pi17 ? n32 : n44504;
  assign n44506 = pi16 ? n32 : n44505;
  assign n44507 = pi15 ? n44506 : n44377;
  assign n44508 = pi14 ? n44501 : n44507;
  assign n44509 = pi18 ? n4127 : n19848;
  assign n44510 = pi17 ? n32 : n44509;
  assign n44511 = pi16 ? n32 : n44510;
  assign n44512 = pi15 ? n44382 : n44511;
  assign n44513 = pi15 ? n30999 : n31135;
  assign n44514 = pi14 ? n44512 : n44513;
  assign n44515 = pi13 ? n44508 : n44514;
  assign n44516 = pi12 ? n44494 : n44515;
  assign n44517 = pi11 ? n44481 : n44516;
  assign n44518 = pi13 ? n43242 : n32;
  assign n44519 = pi18 ? n262 : ~n342;
  assign n44520 = pi17 ? n32 : n44519;
  assign n44521 = pi18 ? n44400 : ~n19318;
  assign n44522 = pi17 ? n44399 : n44521;
  assign n44523 = pi16 ? n44520 : ~n44522;
  assign n44524 = pi15 ? n19235 : n44523;
  assign n44525 = pi14 ? n32 : n44524;
  assign n44526 = pi13 ? n32 : n44525;
  assign n44527 = pi12 ? n44518 : n44526;
  assign n44528 = pi16 ? n1135 : ~n44408;
  assign n44529 = pi16 ? n1135 : ~n44411;
  assign n44530 = pi15 ? n44528 : n44529;
  assign n44531 = pi16 ? n1135 : ~n44415;
  assign n44532 = pi15 ? n44531 : n44418;
  assign n44533 = pi14 ? n44530 : n44532;
  assign n44534 = pi18 ? n1395 : ~n20392;
  assign n44535 = pi17 ? n32 : n44534;
  assign n44536 = pi16 ? n44535 : ~n44429;
  assign n44537 = pi16 ? n1233 : ~n1815;
  assign n44538 = pi15 ? n44536 : n44537;
  assign n44539 = pi14 ? n44425 : n44538;
  assign n44540 = pi13 ? n44533 : n44539;
  assign n44541 = pi16 ? n1214 : ~n44437;
  assign n44542 = pi15 ? n20034 : n44541;
  assign n44543 = pi14 ? n44436 : n44542;
  assign n44544 = pi15 ? n44541 : n31707;
  assign n44545 = pi16 ? n20208 : ~n2326;
  assign n44546 = pi15 ? n44545 : n43787;
  assign n44547 = pi14 ? n44544 : n44546;
  assign n44548 = pi13 ? n44543 : n44547;
  assign n44549 = pi12 ? n44540 : n44548;
  assign n44550 = pi11 ? n44527 : n44549;
  assign n44551 = pi10 ? n44517 : n44550;
  assign n44552 = pi09 ? n32 : n44551;
  assign n44553 = pi08 ? n44449 : n44552;
  assign n44554 = pi07 ? n44297 : n44553;
  assign n44555 = pi14 ? n487 : n21357;
  assign n44556 = pi13 ? n44555 : n31121;
  assign n44557 = pi16 ? n3438 : ~n2654;
  assign n44558 = pi15 ? n13952 : n44557;
  assign n44559 = pi14 ? n20416 : n44558;
  assign n44560 = pi19 ? n28416 : ~n32;
  assign n44561 = pi18 ? n44560 : ~n32;
  assign n44562 = pi17 ? n44561 : ~n2653;
  assign n44563 = pi16 ? n32 : n44562;
  assign n44564 = pi19 ? n32 : n14260;
  assign n44565 = pi18 ? n44564 : ~n19121;
  assign n44566 = pi17 ? n44565 : ~n2531;
  assign n44567 = pi16 ? n32 : n44566;
  assign n44568 = pi15 ? n44563 : n44567;
  assign n44569 = pi19 ? n594 : n44318;
  assign n44570 = pi18 ? n32 : n44569;
  assign n44571 = pi20 ? n342 : n2385;
  assign n44572 = pi19 ? n6308 : ~n44571;
  assign n44573 = pi18 ? n44572 : ~n4343;
  assign n44574 = pi17 ? n44570 : ~n44573;
  assign n44575 = pi16 ? n32 : n44574;
  assign n44576 = pi18 ? n2387 : n4343;
  assign n44577 = pi17 ? n17037 : n44576;
  assign n44578 = pi16 ? n32 : n44577;
  assign n44579 = pi15 ? n44575 : n44578;
  assign n44580 = pi14 ? n44568 : n44579;
  assign n44581 = pi13 ? n44559 : n44580;
  assign n44582 = pi12 ? n44556 : n44581;
  assign n44583 = pi20 ? n2358 : ~n141;
  assign n44584 = pi19 ? n44583 : n32;
  assign n44585 = pi18 ? n44334 : n44584;
  assign n44586 = pi17 ? n30283 : n44585;
  assign n44587 = pi16 ? n32 : n44586;
  assign n44588 = pi17 ? n3164 : ~n3787;
  assign n44589 = pi16 ? n32 : n44588;
  assign n44590 = pi15 ? n44587 : n44589;
  assign n44591 = pi18 ? n237 : ~n21068;
  assign n44592 = pi17 ? n32 : n44591;
  assign n44593 = pi16 ? n32 : n44592;
  assign n44594 = pi20 ? n18337 : ~n17652;
  assign n44595 = pi19 ? n44594 : ~n28750;
  assign n44596 = pi20 ? n28553 : ~n141;
  assign n44597 = pi19 ? n44596 : n32;
  assign n44598 = pi18 ? n44595 : n44597;
  assign n44599 = pi17 ? n32 : n44598;
  assign n44600 = pi16 ? n32 : n44599;
  assign n44601 = pi15 ? n44593 : n44600;
  assign n44602 = pi14 ? n44590 : n44601;
  assign n44603 = pi19 ? n31182 : ~n43838;
  assign n44604 = pi18 ? n44603 : n33554;
  assign n44605 = pi17 ? n32 : n44604;
  assign n44606 = pi16 ? n32 : n44605;
  assign n44607 = pi20 ? n32 : ~n1091;
  assign n44608 = pi19 ? n44607 : ~n5614;
  assign n44609 = pi20 ? n339 : ~n141;
  assign n44610 = pi19 ? n44609 : n32;
  assign n44611 = pi18 ? n44608 : n44610;
  assign n44612 = pi17 ? n32 : n44611;
  assign n44613 = pi16 ? n32 : n44612;
  assign n44614 = pi15 ? n44606 : n44613;
  assign n44615 = pi19 ? n792 : ~n43970;
  assign n44616 = pi18 ? n44615 : n44488;
  assign n44617 = pi17 ? n32 : n44616;
  assign n44618 = pi16 ? n32 : n44617;
  assign n44619 = pi18 ? n32194 : ~n3786;
  assign n44620 = pi17 ? n32 : n44619;
  assign n44621 = pi16 ? n32 : n44620;
  assign n44622 = pi15 ? n44618 : n44621;
  assign n44623 = pi14 ? n44614 : n44622;
  assign n44624 = pi13 ? n44602 : n44623;
  assign n44625 = pi20 ? n1324 : n141;
  assign n44626 = pi19 ? n44625 : ~n32;
  assign n44627 = pi18 ? n880 : ~n44626;
  assign n44628 = pi17 ? n32 : n44627;
  assign n44629 = pi16 ? n32 : n44628;
  assign n44630 = pi15 ? n33451 : n44629;
  assign n44631 = pi18 ? n4127 : n43765;
  assign n44632 = pi17 ? n32 : n44631;
  assign n44633 = pi16 ? n32 : n44632;
  assign n44634 = pi15 ? n31515 : n44633;
  assign n44635 = pi14 ? n44630 : n44634;
  assign n44636 = pi19 ? n25514 : n32;
  assign n44637 = pi18 ? n463 : n44636;
  assign n44638 = pi17 ? n32 : n44637;
  assign n44639 = pi16 ? n32 : n44638;
  assign n44640 = pi15 ? n44639 : n32;
  assign n44641 = pi21 ? n405 : n7107;
  assign n44642 = pi20 ? n44641 : n32;
  assign n44643 = pi19 ? n44642 : n32;
  assign n44644 = pi18 ? n268 : n44643;
  assign n44645 = pi17 ? n32 : n44644;
  assign n44646 = pi16 ? n32 : n44645;
  assign n44647 = pi15 ? n44646 : n31229;
  assign n44648 = pi14 ? n44640 : n44647;
  assign n44649 = pi13 ? n44635 : n44648;
  assign n44650 = pi12 ? n44624 : n44649;
  assign n44651 = pi11 ? n44582 : n44650;
  assign n44652 = pi18 ? n21287 : n496;
  assign n44653 = pi18 ? n20547 : ~n32;
  assign n44654 = pi17 ? n44652 : n44653;
  assign n44655 = pi16 ? n1214 : ~n44654;
  assign n44656 = pi15 ? n31262 : n44655;
  assign n44657 = pi14 ? n32 : n44656;
  assign n44658 = pi13 ? n32 : n44657;
  assign n44659 = pi12 ? n32 : n44658;
  assign n44660 = pi18 ? n20556 : n32;
  assign n44661 = pi17 ? n3067 : ~n44660;
  assign n44662 = pi16 ? n19652 : ~n44661;
  assign n44663 = pi17 ? n20560 : ~n30107;
  assign n44664 = pi16 ? n19652 : ~n44663;
  assign n44665 = pi15 ? n44662 : n44664;
  assign n44666 = pi17 ? n20570 : n32;
  assign n44667 = pi16 ? n919 : n44666;
  assign n44668 = pi15 ? n30109 : n44667;
  assign n44669 = pi14 ? n44665 : n44668;
  assign n44670 = pi18 ? n268 : n237;
  assign n44671 = pi17 ? n32 : n44670;
  assign n44672 = pi16 ? n1471 : ~n44671;
  assign n44673 = pi15 ? n44667 : n44672;
  assign n44674 = pi15 ? n20034 : n18798;
  assign n44675 = pi14 ? n44673 : n44674;
  assign n44676 = pi13 ? n44669 : n44675;
  assign n44677 = pi17 ? n33128 : n1814;
  assign n44678 = pi16 ? n3283 : ~n44677;
  assign n44679 = pi18 ? n4343 : n323;
  assign n44680 = pi17 ? n44679 : ~n1814;
  assign n44681 = pi16 ? n32 : n44680;
  assign n44682 = pi15 ? n44678 : n44681;
  assign n44683 = pi19 ? n4964 : ~n9822;
  assign n44684 = pi18 ? n44683 : n1813;
  assign n44685 = pi17 ? n2736 : ~n44684;
  assign n44686 = pi16 ? n32 : n44685;
  assign n44687 = pi19 ? n4982 : ~n1490;
  assign n44688 = pi18 ? n268 : ~n44687;
  assign n44689 = pi17 ? n32 : n44688;
  assign n44690 = pi17 ? n21288 : n2136;
  assign n44691 = pi16 ? n44689 : ~n44690;
  assign n44692 = pi15 ? n44686 : n44691;
  assign n44693 = pi14 ? n44682 : n44692;
  assign n44694 = pi20 ? n6621 : n342;
  assign n44695 = pi19 ? n44694 : n342;
  assign n44696 = pi18 ? n19082 : n44695;
  assign n44697 = pi17 ? n32 : n44696;
  assign n44698 = pi19 ? n32 : ~n3524;
  assign n44699 = pi18 ? n44698 : n32;
  assign n44700 = pi17 ? n44699 : n2325;
  assign n44701 = pi16 ? n44697 : ~n44700;
  assign n44702 = pi15 ? n44701 : n19653;
  assign n44703 = pi17 ? n29510 : n2325;
  assign n44704 = pi16 ? n1233 : ~n44703;
  assign n44705 = pi15 ? n44283 : n44704;
  assign n44706 = pi14 ? n44702 : n44705;
  assign n44707 = pi13 ? n44693 : n44706;
  assign n44708 = pi12 ? n44676 : n44707;
  assign n44709 = pi11 ? n44659 : n44708;
  assign n44710 = pi10 ? n44651 : n44709;
  assign n44711 = pi09 ? n32 : n44710;
  assign n44712 = pi15 ? n20486 : n13952;
  assign n44713 = pi14 ? n487 : n44712;
  assign n44714 = pi14 ? n672 : n32;
  assign n44715 = pi13 ? n44713 : n44714;
  assign n44716 = pi16 ? n3438 : ~n2426;
  assign n44717 = pi15 ? n486 : n44716;
  assign n44718 = pi14 ? n487 : n44717;
  assign n44719 = pi19 ? n29298 : ~n32;
  assign n44720 = pi18 ? n44719 : ~n32;
  assign n44721 = pi17 ? n44720 : ~n2425;
  assign n44722 = pi16 ? n32 : n44721;
  assign n44723 = pi18 ? n8231 : ~n19137;
  assign n44724 = pi17 ? n44723 : ~n2531;
  assign n44725 = pi16 ? n32 : n44724;
  assign n44726 = pi15 ? n44722 : n44725;
  assign n44727 = pi19 ? n594 : n44468;
  assign n44728 = pi18 ? n32 : n44727;
  assign n44729 = pi20 ? n9863 : n1091;
  assign n44730 = pi19 ? n44729 : n13171;
  assign n44731 = pi18 ? n44730 : ~n33338;
  assign n44732 = pi17 ? n44728 : ~n44731;
  assign n44733 = pi16 ? n32 : n44732;
  assign n44734 = pi19 ? n32 : n43541;
  assign n44735 = pi18 ? n32 : n44734;
  assign n44736 = pi19 ? n6398 : n2386;
  assign n44737 = pi18 ? n44736 : n4343;
  assign n44738 = pi17 ? n44735 : n44737;
  assign n44739 = pi16 ? n32 : n44738;
  assign n44740 = pi15 ? n44733 : n44739;
  assign n44741 = pi14 ? n44726 : n44740;
  assign n44742 = pi13 ? n44718 : n44741;
  assign n44743 = pi12 ? n44715 : n44742;
  assign n44744 = pi17 ? n30283 : n44489;
  assign n44745 = pi16 ? n32 : n44744;
  assign n44746 = pi17 ? n3164 : ~n2653;
  assign n44747 = pi16 ? n32 : n44746;
  assign n44748 = pi15 ? n44745 : n44747;
  assign n44749 = pi18 ? n237 : ~n21180;
  assign n44750 = pi17 ? n32 : n44749;
  assign n44751 = pi16 ? n32 : n44750;
  assign n44752 = pi20 ? n175 : n6085;
  assign n44753 = pi20 ? n9194 : n9491;
  assign n44754 = pi19 ? n44752 : n44753;
  assign n44755 = pi20 ? n6822 : ~n339;
  assign n44756 = pi19 ? n44755 : n32;
  assign n44757 = pi18 ? n44754 : n44756;
  assign n44758 = pi17 ? n32 : n44757;
  assign n44759 = pi16 ? n32 : n44758;
  assign n44760 = pi15 ? n44751 : n44759;
  assign n44761 = pi14 ? n44748 : n44760;
  assign n44762 = pi19 ? n31182 : ~n28750;
  assign n44763 = pi20 ? n18415 : ~n339;
  assign n44764 = pi19 ? n44763 : n32;
  assign n44765 = pi18 ? n44762 : n44764;
  assign n44766 = pi17 ? n32 : n44765;
  assign n44767 = pi16 ? n32 : n44766;
  assign n44768 = pi19 ? n44607 : ~n333;
  assign n44769 = pi18 ? n44768 : n44764;
  assign n44770 = pi17 ? n32 : n44769;
  assign n44771 = pi16 ? n32 : n44770;
  assign n44772 = pi15 ? n44767 : n44771;
  assign n44773 = pi19 ? n792 : ~n5854;
  assign n44774 = pi20 ? n2358 : ~n339;
  assign n44775 = pi19 ? n44774 : n32;
  assign n44776 = pi18 ? n44773 : n44775;
  assign n44777 = pi17 ? n32 : n44776;
  assign n44778 = pi16 ? n32 : n44777;
  assign n44779 = pi19 ? n6398 : ~n31723;
  assign n44780 = pi20 ? n1331 : n339;
  assign n44781 = pi19 ? n44780 : ~n32;
  assign n44782 = pi18 ? n44779 : ~n44781;
  assign n44783 = pi17 ? n32 : n44782;
  assign n44784 = pi16 ? n32 : n44783;
  assign n44785 = pi15 ? n44778 : n44784;
  assign n44786 = pi14 ? n44772 : n44785;
  assign n44787 = pi13 ? n44761 : n44786;
  assign n44788 = pi19 ? n7622 : ~n32;
  assign n44789 = pi18 ? n880 : ~n44788;
  assign n44790 = pi17 ? n32 : n44789;
  assign n44791 = pi16 ? n32 : n44790;
  assign n44792 = pi15 ? n11429 : n44791;
  assign n44793 = pi18 ? n4127 : n43881;
  assign n44794 = pi17 ? n32 : n44793;
  assign n44795 = pi16 ? n32 : n44794;
  assign n44796 = pi15 ? n20982 : n44795;
  assign n44797 = pi14 ? n44792 : n44796;
  assign n44798 = pi14 ? n18906 : n31347;
  assign n44799 = pi13 ? n44797 : n44798;
  assign n44800 = pi12 ? n44787 : n44799;
  assign n44801 = pi11 ? n44743 : n44800;
  assign n44802 = pi16 ? n1214 : ~n44661;
  assign n44803 = pi16 ? n1214 : ~n44663;
  assign n44804 = pi15 ? n44802 : n44803;
  assign n44805 = pi14 ? n44804 : n44668;
  assign n44806 = pi15 ? n20034 : n29729;
  assign n44807 = pi14 ? n44673 : n44806;
  assign n44808 = pi13 ? n44805 : n44807;
  assign n44809 = pi17 ? n33128 : n2136;
  assign n44810 = pi16 ? n3283 : ~n44809;
  assign n44811 = pi17 ? n44679 : ~n2136;
  assign n44812 = pi16 ? n32 : n44811;
  assign n44813 = pi15 ? n44810 : n44812;
  assign n44814 = pi18 ? n44683 : n814;
  assign n44815 = pi17 ? n2736 : ~n44814;
  assign n44816 = pi16 ? n32 : n44815;
  assign n44817 = pi15 ? n44816 : n44691;
  assign n44818 = pi14 ? n44813 : n44817;
  assign n44819 = pi15 ? n44701 : n19711;
  assign n44820 = pi15 ? n19711 : n44704;
  assign n44821 = pi14 ? n44819 : n44820;
  assign n44822 = pi13 ? n44818 : n44821;
  assign n44823 = pi12 ? n44808 : n44822;
  assign n44824 = pi11 ? n44659 : n44823;
  assign n44825 = pi10 ? n44801 : n44824;
  assign n44826 = pi09 ? n32 : n44825;
  assign n44827 = pi08 ? n44711 : n44826;
  assign n44828 = pi15 ? n13948 : n486;
  assign n44829 = pi14 ? n20844 : n44828;
  assign n44830 = pi13 ? n44829 : n31305;
  assign n44831 = pi15 ? n32 : n44716;
  assign n44832 = pi14 ? n32 : n44831;
  assign n44833 = pi18 ? n6926 : ~n32;
  assign n44834 = pi17 ? n44833 : ~n2425;
  assign n44835 = pi16 ? n32 : n44834;
  assign n44836 = pi20 ? n3843 : ~n32;
  assign n44837 = pi19 ? n44836 : ~n32;
  assign n44838 = pi18 ? n312 : n44837;
  assign n44839 = pi17 ? n44838 : ~n2653;
  assign n44840 = pi16 ? n32 : n44839;
  assign n44841 = pi15 ? n44835 : n44840;
  assign n44842 = pi18 ? n32 : ~n23514;
  assign n44843 = pi17 ? n44842 : ~n2653;
  assign n44844 = pi16 ? n32 : n44843;
  assign n44845 = pi17 ? n2959 : ~n2653;
  assign n44846 = pi16 ? n32 : n44845;
  assign n44847 = pi15 ? n44844 : n44846;
  assign n44848 = pi14 ? n44841 : n44847;
  assign n44849 = pi13 ? n44832 : n44848;
  assign n44850 = pi12 ? n44830 : n44849;
  assign n44851 = pi18 ? n268 : n418;
  assign n44852 = pi17 ? n17463 : ~n44851;
  assign n44853 = pi16 ? n32 : n44852;
  assign n44854 = pi17 ? n32 : ~n2425;
  assign n44855 = pi16 ? n32 : n44854;
  assign n44856 = pi15 ? n44853 : n44855;
  assign n44857 = pi18 ? n237 : ~n33596;
  assign n44858 = pi17 ? n32 : n44857;
  assign n44859 = pi16 ? n32 : n44858;
  assign n44860 = pi15 ? n44859 : n31388;
  assign n44861 = pi14 ? n44856 : n44860;
  assign n44862 = pi18 ? n4428 : ~n2424;
  assign n44863 = pi17 ? n32 : n44862;
  assign n44864 = pi16 ? n32 : n44863;
  assign n44865 = pi15 ? n21755 : n44864;
  assign n44866 = pi14 ? n31394 : n44865;
  assign n44867 = pi13 ? n44861 : n44866;
  assign n44868 = pi18 ? n702 : ~n2424;
  assign n44869 = pi17 ? n32 : n44868;
  assign n44870 = pi16 ? n32 : n44869;
  assign n44871 = pi18 ? n1139 : n20848;
  assign n44872 = pi17 ? n32 : n44871;
  assign n44873 = pi16 ? n32 : n44872;
  assign n44874 = pi15 ? n44870 : n44873;
  assign n44875 = pi18 ? n863 : n4671;
  assign n44876 = pi17 ? n32 : n44875;
  assign n44877 = pi16 ? n32 : n44876;
  assign n44878 = pi15 ? n20982 : n44877;
  assign n44879 = pi14 ? n44874 : n44878;
  assign n44880 = pi18 ? n268 : n31409;
  assign n44881 = pi17 ? n32 : n44880;
  assign n44882 = pi16 ? n32 : n44881;
  assign n44883 = pi15 ? n44882 : n31415;
  assign n44884 = pi14 ? n44883 : n31417;
  assign n44885 = pi13 ? n44879 : n44884;
  assign n44886 = pi12 ? n44867 : n44885;
  assign n44887 = pi11 ? n44850 : n44886;
  assign n44888 = pi18 ? n16543 : n880;
  assign n44889 = pi18 ? n20717 : ~n32;
  assign n44890 = pi17 ? n44888 : n44889;
  assign n44891 = pi16 ? n1214 : ~n44890;
  assign n44892 = pi15 ? n31262 : n44891;
  assign n44893 = pi14 ? n32 : n44892;
  assign n44894 = pi13 ? n32 : n44893;
  assign n44895 = pi12 ? n32 : n44894;
  assign n44896 = pi18 ? n20725 : n32;
  assign n44897 = pi17 ? n2733 : ~n44896;
  assign n44898 = pi16 ? n1135 : ~n44897;
  assign n44899 = pi17 ? n20730 : ~n30107;
  assign n44900 = pi16 ? n1135 : ~n44899;
  assign n44901 = pi15 ? n44898 : n44900;
  assign n44902 = pi17 ? n20738 : n32;
  assign n44903 = pi16 ? n30460 : n44902;
  assign n44904 = pi15 ? n30109 : n44903;
  assign n44905 = pi14 ? n44901 : n44904;
  assign n44906 = pi15 ? n44903 : n29729;
  assign n44907 = pi15 ? n30941 : n29729;
  assign n44908 = pi14 ? n44906 : n44907;
  assign n44909 = pi13 ? n44905 : n44908;
  assign n44910 = pi17 ? n36949 : ~n1807;
  assign n44911 = pi16 ? n32 : n44910;
  assign n44912 = pi17 ? n44679 : ~n1807;
  assign n44913 = pi16 ? n32 : n44912;
  assign n44914 = pi15 ? n44911 : n44913;
  assign n44915 = pi19 ? n5694 : ~n9822;
  assign n44916 = pi18 ? n44915 : n350;
  assign n44917 = pi17 ? n3067 : ~n44916;
  assign n44918 = pi16 ? n32 : n44917;
  assign n44919 = pi18 ? n32 : ~n44687;
  assign n44920 = pi17 ? n32 : n44919;
  assign n44921 = pi17 ? n28644 : n2325;
  assign n44922 = pi16 ? n44920 : ~n44921;
  assign n44923 = pi15 ? n44918 : n44922;
  assign n44924 = pi14 ? n44914 : n44923;
  assign n44925 = pi18 ? n32 : ~n441;
  assign n44926 = pi17 ? n31659 : n44925;
  assign n44927 = pi16 ? n3438 : ~n44926;
  assign n44928 = pi17 ? n32 : n44925;
  assign n44929 = pi16 ? n1214 : ~n44928;
  assign n44930 = pi15 ? n44927 : n44929;
  assign n44931 = pi16 ? n19652 : ~n44928;
  assign n44932 = pi18 ? n566 : ~n31484;
  assign n44933 = pi17 ? n32 : n44932;
  assign n44934 = pi19 ? n11899 : n31488;
  assign n44935 = pi18 ? n44934 : ~n32;
  assign n44936 = pi17 ? n44935 : ~n2325;
  assign n44937 = pi16 ? n44933 : n44936;
  assign n44938 = pi15 ? n44931 : n44937;
  assign n44939 = pi14 ? n44930 : n44938;
  assign n44940 = pi13 ? n44924 : n44939;
  assign n44941 = pi12 ? n44909 : n44940;
  assign n44942 = pi11 ? n44895 : n44941;
  assign n44943 = pi10 ? n44887 : n44942;
  assign n44944 = pi09 ? n32 : n44943;
  assign n44945 = pi17 ? n32 : n36054;
  assign n44946 = pi16 ? n44945 : ~n2120;
  assign n44947 = pi15 ? n32 : n44946;
  assign n44948 = pi14 ? n32 : n44947;
  assign n44949 = pi20 ? n3523 : ~n18255;
  assign n44950 = pi19 ? n44949 : ~n32;
  assign n44951 = pi18 ? n44950 : ~n32;
  assign n44952 = pi17 ? n44951 : ~n2119;
  assign n44953 = pi16 ? n32 : n44952;
  assign n44954 = pi20 ? n428 : n6050;
  assign n44955 = pi19 ? n32 : n44954;
  assign n44956 = pi20 ? n29457 : ~n32;
  assign n44957 = pi19 ? n44956 : ~n32;
  assign n44958 = pi18 ? n44955 : n44957;
  assign n44959 = pi17 ? n44958 : ~n2653;
  assign n44960 = pi16 ? n32 : n44959;
  assign n44961 = pi15 ? n44953 : n44960;
  assign n44962 = pi14 ? n44961 : n44847;
  assign n44963 = pi13 ? n44948 : n44962;
  assign n44964 = pi12 ? n44830 : n44963;
  assign n44965 = pi18 ? n1139 : n21043;
  assign n44966 = pi17 ? n32 : n44965;
  assign n44967 = pi16 ? n32 : n44966;
  assign n44968 = pi15 ? n44870 : n44967;
  assign n44969 = pi14 ? n44968 : n44878;
  assign n44970 = pi18 ? n268 : n31505;
  assign n44971 = pi17 ? n32 : n44970;
  assign n44972 = pi16 ? n32 : n44971;
  assign n44973 = pi15 ? n44972 : n31511;
  assign n44974 = pi14 ? n44973 : n31516;
  assign n44975 = pi13 ? n44969 : n44974;
  assign n44976 = pi12 ? n44867 : n44975;
  assign n44977 = pi11 ? n44964 : n44976;
  assign n44978 = pi18 ? n20717 : ~n113;
  assign n44979 = pi17 ? n44888 : n44978;
  assign n44980 = pi16 ? n1214 : ~n44979;
  assign n44981 = pi15 ? n31533 : n44980;
  assign n44982 = pi14 ? n32 : n44981;
  assign n44983 = pi13 ? n32 : n44982;
  assign n44984 = pi12 ? n32 : n44983;
  assign n44985 = pi16 ? n270 : n44902;
  assign n44986 = pi15 ? n30109 : n44985;
  assign n44987 = pi14 ? n44901 : n44986;
  assign n44988 = pi15 ? n44985 : n29729;
  assign n44989 = pi14 ? n44988 : n44907;
  assign n44990 = pi13 ? n44987 : n44989;
  assign n44991 = pi17 ? n31659 : n2136;
  assign n44992 = pi16 ? n3438 : ~n44991;
  assign n44993 = pi16 ? n1214 : ~n2137;
  assign n44994 = pi15 ? n44992 : n44993;
  assign n44995 = pi18 ? n566 : ~n31549;
  assign n44996 = pi17 ? n32 : n44995;
  assign n44997 = pi20 ? n314 : ~n342;
  assign n44998 = pi19 ? n44997 : n31553;
  assign n44999 = pi18 ? n44998 : ~n32;
  assign n45000 = pi17 ? n44999 : ~n2325;
  assign n45001 = pi16 ? n44996 : n45000;
  assign n45002 = pi15 ? n44993 : n45001;
  assign n45003 = pi14 ? n44994 : n45002;
  assign n45004 = pi13 ? n44924 : n45003;
  assign n45005 = pi12 ? n44990 : n45004;
  assign n45006 = pi11 ? n44984 : n45005;
  assign n45007 = pi10 ? n44977 : n45006;
  assign n45008 = pi09 ? n32 : n45007;
  assign n45009 = pi08 ? n44944 : n45008;
  assign n45010 = pi07 ? n44827 : n45009;
  assign n45011 = pi06 ? n44554 : n45010;
  assign n45012 = pi14 ? n31717 : n31783;
  assign n45013 = pi13 ? n45012 : n20833;
  assign n45014 = pi18 ? n32 : n18710;
  assign n45015 = pi17 ? n32 : n45014;
  assign n45016 = pi16 ? n45015 : ~n2415;
  assign n45017 = pi17 ? n32 : n3447;
  assign n45018 = pi16 ? n45017 : ~n2120;
  assign n45019 = pi15 ? n45016 : n45018;
  assign n45020 = pi14 ? n20831 : n45019;
  assign n45021 = pi19 ? n208 : n236;
  assign n45022 = pi18 ? n45021 : ~n32;
  assign n45023 = pi17 ? n45022 : ~n2119;
  assign n45024 = pi16 ? n32 : n45023;
  assign n45025 = pi18 ? n4127 : ~n18532;
  assign n45026 = pi17 ? n45025 : ~n2653;
  assign n45027 = pi16 ? n32 : n45026;
  assign n45028 = pi15 ? n45024 : n45027;
  assign n45029 = pi19 ? n507 : n4406;
  assign n45030 = pi18 ? n32 : n45029;
  assign n45031 = pi17 ? n45030 : ~n2119;
  assign n45032 = pi16 ? n32 : n45031;
  assign n45033 = pi20 ? n8644 : n18834;
  assign n45034 = pi19 ? n45033 : n28076;
  assign n45035 = pi20 ? n820 : n1940;
  assign n45036 = pi19 ? n45035 : ~n32;
  assign n45037 = pi18 ? n45034 : ~n45036;
  assign n45038 = pi17 ? n32 : n45037;
  assign n45039 = pi16 ? n32 : n45038;
  assign n45040 = pi15 ? n45032 : n45039;
  assign n45041 = pi14 ? n45028 : n45040;
  assign n45042 = pi13 ? n45020 : n45041;
  assign n45043 = pi12 ? n45013 : n45042;
  assign n45044 = pi15 ? n31577 : n31583;
  assign n45045 = pi14 ? n31578 : n45044;
  assign n45046 = pi15 ? n31588 : n33101;
  assign n45047 = pi18 ? n508 : ~n605;
  assign n45048 = pi17 ? n32 : n45047;
  assign n45049 = pi16 ? n32 : n45048;
  assign n45050 = pi15 ? n45049 : n11426;
  assign n45051 = pi14 ? n45046 : n45050;
  assign n45052 = pi13 ? n45045 : n45051;
  assign n45053 = pi18 ? n496 : ~n5436;
  assign n45054 = pi17 ? n32 : n45053;
  assign n45055 = pi16 ? n32 : n45054;
  assign n45056 = pi15 ? n45055 : n20686;
  assign n45057 = pi14 ? n45056 : n31597;
  assign n45058 = pi18 ? n4722 : n13080;
  assign n45059 = pi17 ? n32 : n45058;
  assign n45060 = pi16 ? n32 : n45059;
  assign n45061 = pi15 ? n12098 : n45060;
  assign n45062 = pi14 ? n45061 : n32;
  assign n45063 = pi13 ? n45057 : n45062;
  assign n45064 = pi12 ? n45052 : n45063;
  assign n45065 = pi11 ? n45043 : n45064;
  assign n45066 = pi14 ? n32 : n146;
  assign n45067 = pi13 ? n45066 : n44299;
  assign n45068 = pi15 ? n32 : n31653;
  assign n45069 = pi17 ? n17463 : n1213;
  assign n45070 = pi16 ? n1135 : ~n45069;
  assign n45071 = pi18 ? n19202 : n209;
  assign n45072 = pi18 ? n14413 : n32;
  assign n45073 = pi17 ? n45071 : ~n45072;
  assign n45074 = pi16 ? n1471 : ~n45073;
  assign n45075 = pi15 ? n45070 : n45074;
  assign n45076 = pi14 ? n45068 : n45075;
  assign n45077 = pi13 ? n32 : n45076;
  assign n45078 = pi12 ? n45067 : n45077;
  assign n45079 = pi17 ? n2959 : ~n30877;
  assign n45080 = pi16 ? n1135 : ~n45079;
  assign n45081 = pi17 ? n20913 : ~n19529;
  assign n45082 = pi16 ? n1135 : ~n45081;
  assign n45083 = pi15 ? n45080 : n45082;
  assign n45084 = pi17 ? n269 : n32;
  assign n45085 = pi16 ? n18018 : n45084;
  assign n45086 = pi18 ? n341 : ~n20920;
  assign n45087 = pi17 ? n32 : n45086;
  assign n45088 = pi17 ? n20927 : ~n42923;
  assign n45089 = pi16 ? n45087 : ~n45088;
  assign n45090 = pi15 ? n45085 : n45089;
  assign n45091 = pi14 ? n45083 : n45090;
  assign n45092 = pi19 ? n33683 : n1385;
  assign n45093 = pi18 ? n341 : ~n45092;
  assign n45094 = pi17 ? n32 : n45093;
  assign n45095 = pi20 ? n18624 : ~n9641;
  assign n45096 = pi19 ? n30461 : ~n45095;
  assign n45097 = pi20 ? n17669 : n785;
  assign n45098 = pi19 ? n17641 : ~n45097;
  assign n45099 = pi18 ? n45096 : n45098;
  assign n45100 = pi20 ? n12884 : ~n20944;
  assign n45101 = pi19 ? n45100 : n7435;
  assign n45102 = pi18 ? n45101 : n350;
  assign n45103 = pi17 ? n45099 : n45102;
  assign n45104 = pi16 ? n45094 : ~n45103;
  assign n45105 = pi15 ? n45104 : n31684;
  assign n45106 = pi14 ? n45105 : n31688;
  assign n45107 = pi13 ? n45091 : n45106;
  assign n45108 = pi18 ? n5351 : n496;
  assign n45109 = pi19 ? n6887 : ~n32;
  assign n45110 = pi18 ? n32 : n45109;
  assign n45111 = pi17 ? n45108 : ~n45110;
  assign n45112 = pi16 ? n32 : n45111;
  assign n45113 = pi18 ? n32 : n28602;
  assign n45114 = pi17 ? n32 : n45113;
  assign n45115 = pi18 ? n19202 : n32;
  assign n45116 = pi17 ? n45115 : n1807;
  assign n45117 = pi16 ? n45114 : ~n45116;
  assign n45118 = pi15 ? n45112 : n45117;
  assign n45119 = pi14 ? n31696 : n45118;
  assign n45120 = pi18 ? n32 : n33017;
  assign n45121 = pi17 ? n32 : n45120;
  assign n45122 = pi19 ? n349 : ~n4982;
  assign n45123 = pi18 ? n45122 : ~n32;
  assign n45124 = pi17 ? n45123 : ~n2136;
  assign n45125 = pi16 ? n45121 : n45124;
  assign n45126 = pi15 ? n45125 : n20034;
  assign n45127 = pi17 ? n20165 : n2136;
  assign n45128 = pi16 ? n1135 : ~n45127;
  assign n45129 = pi18 ? n127 : ~n20172;
  assign n45130 = pi17 ? n32 : n45129;
  assign n45131 = pi16 ? n45130 : ~n2326;
  assign n45132 = pi15 ? n45128 : n45131;
  assign n45133 = pi14 ? n45126 : n45132;
  assign n45134 = pi13 ? n45119 : n45133;
  assign n45135 = pi12 ? n45107 : n45134;
  assign n45136 = pi11 ? n45078 : n45135;
  assign n45137 = pi10 ? n45065 : n45136;
  assign n45138 = pi09 ? n32 : n45137;
  assign n45139 = pi15 ? n20836 : n21232;
  assign n45140 = pi14 ? n45139 : n31783;
  assign n45141 = pi13 ? n45140 : n20968;
  assign n45142 = pi20 ? n175 : n820;
  assign n45143 = pi19 ? n32 : n45142;
  assign n45144 = pi18 ? n32 : n45143;
  assign n45145 = pi17 ? n32 : n45144;
  assign n45146 = pi16 ? n45145 : ~n2409;
  assign n45147 = pi15 ? n45146 : n45018;
  assign n45148 = pi14 ? n20836 : n45147;
  assign n45149 = pi17 ? n45025 : ~n2119;
  assign n45150 = pi16 ? n32 : n45149;
  assign n45151 = pi15 ? n45024 : n45150;
  assign n45152 = pi14 ? n45151 : n45040;
  assign n45153 = pi13 ? n45148 : n45152;
  assign n45154 = pi12 ? n45141 : n45153;
  assign n45155 = pi14 ? n31721 : n45044;
  assign n45156 = pi15 ? n31729 : n33101;
  assign n45157 = pi14 ? n45156 : n45050;
  assign n45158 = pi13 ? n45155 : n45157;
  assign n45159 = pi12 ? n45158 : n45063;
  assign n45160 = pi11 ? n45154 : n45159;
  assign n45161 = pi12 ? n32 : n45077;
  assign n45162 = pi16 ? n1233 : ~n45079;
  assign n45163 = pi16 ? n1233 : ~n45081;
  assign n45164 = pi15 ? n45162 : n45163;
  assign n45165 = pi14 ? n45164 : n45090;
  assign n45166 = pi14 ? n45105 : n31744;
  assign n45167 = pi13 ? n45165 : n45166;
  assign n45168 = pi21 ? n35 : n140;
  assign n45169 = pi20 ? n45168 : ~n32;
  assign n45170 = pi19 ? n45169 : ~n32;
  assign n45171 = pi18 ? n32 : n45170;
  assign n45172 = pi17 ? n45108 : ~n45171;
  assign n45173 = pi16 ? n32 : n45172;
  assign n45174 = pi15 ? n45173 : n45117;
  assign n45175 = pi14 ? n31696 : n45174;
  assign n45176 = pi16 ? n1233 : ~n45127;
  assign n45177 = pi15 ? n45176 : n45131;
  assign n45178 = pi14 ? n45126 : n45177;
  assign n45179 = pi13 ? n45175 : n45178;
  assign n45180 = pi12 ? n45167 : n45179;
  assign n45181 = pi11 ? n45161 : n45180;
  assign n45182 = pi10 ? n45160 : n45181;
  assign n45183 = pi09 ? n32 : n45182;
  assign n45184 = pi08 ? n45138 : n45183;
  assign n45185 = pi14 ? n23063 : n21553;
  assign n45186 = pi13 ? n45185 : n32;
  assign n45187 = pi16 ? n3165 : ~n2409;
  assign n45188 = pi17 ? n2177 : ~n2408;
  assign n45189 = pi16 ? n3438 : n45188;
  assign n45190 = pi15 ? n45187 : n45189;
  assign n45191 = pi14 ? n20836 : n45190;
  assign n45192 = pi18 ? n7038 : ~n18532;
  assign n45193 = pi17 ? n45192 : ~n2119;
  assign n45194 = pi16 ? n32 : n45193;
  assign n45195 = pi18 ? n32 : ~n21661;
  assign n45196 = pi17 ? n45195 : ~n2119;
  assign n45197 = pi16 ? n32 : n45196;
  assign n45198 = pi15 ? n45194 : n45197;
  assign n45199 = pi19 ? n44321 : ~n28076;
  assign n45200 = pi20 ? n18261 : n207;
  assign n45201 = pi19 ? n45200 : ~n32;
  assign n45202 = pi18 ? n45199 : n45201;
  assign n45203 = pi17 ? n17346 : ~n45202;
  assign n45204 = pi16 ? n32 : n45203;
  assign n45205 = pi15 ? n45204 : n13948;
  assign n45206 = pi14 ? n45198 : n45205;
  assign n45207 = pi13 ? n45191 : n45206;
  assign n45208 = pi12 ? n45186 : n45207;
  assign n45209 = pi18 ? n350 : ~n2413;
  assign n45210 = pi17 ? n18292 : n45209;
  assign n45211 = pi16 ? n32 : n45210;
  assign n45212 = pi15 ? n31767 : n45211;
  assign n45213 = pi14 ? n45212 : n31778;
  assign n45214 = pi18 ? n323 : ~n2413;
  assign n45215 = pi17 ? n32 : n45214;
  assign n45216 = pi16 ? n32 : n45215;
  assign n45217 = pi18 ? n4428 : ~n2413;
  assign n45218 = pi17 ? n32 : n45217;
  assign n45219 = pi16 ? n32 : n45218;
  assign n45220 = pi15 ? n45216 : n45219;
  assign n45221 = pi18 ? n508 : ~n2413;
  assign n45222 = pi17 ? n32 : n45221;
  assign n45223 = pi16 ? n32 : n45222;
  assign n45224 = pi15 ? n45223 : n22036;
  assign n45225 = pi14 ? n45220 : n45224;
  assign n45226 = pi13 ? n45213 : n45225;
  assign n45227 = pi18 ? n496 : ~n23217;
  assign n45228 = pi17 ? n32 : n45227;
  assign n45229 = pi16 ? n32 : n45228;
  assign n45230 = pi18 ? n863 : n21568;
  assign n45231 = pi17 ? n32 : n45230;
  assign n45232 = pi16 ? n32 : n45231;
  assign n45233 = pi15 ? n45229 : n45232;
  assign n45234 = pi14 ? n45233 : n31792;
  assign n45235 = pi20 ? n339 : ~n339;
  assign n45236 = pi19 ? n45235 : n32;
  assign n45237 = pi18 ? n4722 : n45236;
  assign n45238 = pi17 ? n32 : n45237;
  assign n45239 = pi16 ? n32 : n45238;
  assign n45240 = pi15 ? n12098 : n45239;
  assign n45241 = pi14 ? n45240 : n32;
  assign n45242 = pi13 ? n45234 : n45241;
  assign n45243 = pi12 ? n45226 : n45242;
  assign n45244 = pi11 ? n45208 : n45243;
  assign n45245 = pi15 ? n32 : n29519;
  assign n45246 = pi18 ? n21081 : ~n32;
  assign n45247 = pi17 ? n4261 : n45246;
  assign n45248 = pi16 ? n1135 : ~n45247;
  assign n45249 = pi18 ? n19350 : n863;
  assign n45250 = pi17 ? n45249 : ~n31659;
  assign n45251 = pi16 ? n1471 : ~n45250;
  assign n45252 = pi15 ? n45248 : n45251;
  assign n45253 = pi14 ? n45245 : n45252;
  assign n45254 = pi13 ? n32 : n45253;
  assign n45255 = pi12 ? n32 : n45254;
  assign n45256 = pi18 ? n15241 : n32;
  assign n45257 = pi17 ? n3164 : ~n45256;
  assign n45258 = pi16 ? n1135 : ~n45257;
  assign n45259 = pi17 ? n21095 : ~n19529;
  assign n45260 = pi16 ? n1135 : ~n45259;
  assign n45261 = pi15 ? n45258 : n45260;
  assign n45262 = pi17 ? n34856 : n32;
  assign n45263 = pi16 ? n18018 : n45262;
  assign n45264 = pi18 ? n341 : ~n21102;
  assign n45265 = pi17 ? n32 : n45264;
  assign n45266 = pi20 ? n9641 : n11107;
  assign n45267 = pi19 ? n21105 : n45266;
  assign n45268 = pi18 ? n45267 : n21109;
  assign n45269 = pi18 ? n21114 : ~n350;
  assign n45270 = pi17 ? n45268 : ~n45269;
  assign n45271 = pi16 ? n45265 : ~n45270;
  assign n45272 = pi15 ? n45263 : n45271;
  assign n45273 = pi14 ? n45261 : n45272;
  assign n45274 = pi19 ? n266 : n321;
  assign n45275 = pi18 ? n209 : ~n45274;
  assign n45276 = pi17 ? n32 : n45275;
  assign n45277 = pi16 ? n45276 : ~n31852;
  assign n45278 = pi15 ? n45277 : n31854;
  assign n45279 = pi14 ? n45278 : n31858;
  assign n45280 = pi13 ? n45273 : n45279;
  assign n45281 = pi18 ? n26660 : n496;
  assign n45282 = pi17 ? n45281 : ~n2537;
  assign n45283 = pi16 ? n32 : n45282;
  assign n45284 = pi19 ? n321 : ~n207;
  assign n45285 = pi18 ? n32 : n45284;
  assign n45286 = pi17 ? n32 : n45285;
  assign n45287 = pi18 ? n22885 : n32;
  assign n45288 = pi17 ? n45287 : n1807;
  assign n45289 = pi16 ? n45286 : ~n45288;
  assign n45290 = pi15 ? n45283 : n45289;
  assign n45291 = pi14 ? n31865 : n45290;
  assign n45292 = pi19 ? n236 : ~n16002;
  assign n45293 = pi18 ? n32 : n45292;
  assign n45294 = pi17 ? n32 : n45293;
  assign n45295 = pi19 ? n1757 : n4982;
  assign n45296 = pi18 ? n45295 : n32;
  assign n45297 = pi17 ? n45296 : n36008;
  assign n45298 = pi16 ? n45294 : ~n45297;
  assign n45299 = pi15 ? n45298 : n20034;
  assign n45300 = pi18 ? n366 : ~n20912;
  assign n45301 = pi17 ? n32 : n45300;
  assign n45302 = pi19 ? n31483 : ~n349;
  assign n45303 = pi18 ? n31879 : n45302;
  assign n45304 = pi17 ? n45303 : n2325;
  assign n45305 = pi16 ? n45301 : ~n45304;
  assign n45306 = pi18 ? n127 : ~n32;
  assign n45307 = pi17 ? n32 : n45306;
  assign n45308 = pi16 ? n45307 : ~n2137;
  assign n45309 = pi15 ? n45305 : n45308;
  assign n45310 = pi14 ? n45299 : n45309;
  assign n45311 = pi13 ? n45291 : n45310;
  assign n45312 = pi12 ? n45280 : n45311;
  assign n45313 = pi11 ? n45255 : n45312;
  assign n45314 = pi10 ? n45244 : n45313;
  assign n45315 = pi09 ? n32 : n45314;
  assign n45316 = pi14 ? n23063 : n21630;
  assign n45317 = pi13 ? n45316 : n32;
  assign n45318 = pi16 ? n3165 : ~n2293;
  assign n45319 = pi15 ? n45318 : n45189;
  assign n45320 = pi14 ? n14613 : n45319;
  assign n45321 = pi17 ? n45192 : ~n2408;
  assign n45322 = pi16 ? n32 : n45321;
  assign n45323 = pi15 ? n45322 : n45197;
  assign n45324 = pi14 ? n45323 : n45205;
  assign n45325 = pi13 ? n45320 : n45324;
  assign n45326 = pi12 ? n45317 : n45325;
  assign n45327 = pi18 ? n350 : ~n605;
  assign n45328 = pi17 ? n18292 : n45327;
  assign n45329 = pi16 ? n32 : n45328;
  assign n45330 = pi15 ? n31899 : n45329;
  assign n45331 = pi15 ? n31583 : n31588;
  assign n45332 = pi14 ? n45330 : n45331;
  assign n45333 = pi15 ? n33101 : n45219;
  assign n45334 = pi14 ? n45333 : n45224;
  assign n45335 = pi13 ? n45332 : n45334;
  assign n45336 = pi18 ? n863 : n27138;
  assign n45337 = pi17 ? n32 : n45336;
  assign n45338 = pi16 ? n32 : n45337;
  assign n45339 = pi15 ? n45229 : n45338;
  assign n45340 = pi14 ? n45339 : n31792;
  assign n45341 = pi20 ? n339 : ~n243;
  assign n45342 = pi19 ? n45341 : n32;
  assign n45343 = pi18 ? n4722 : n45342;
  assign n45344 = pi17 ? n32 : n45343;
  assign n45345 = pi16 ? n32 : n45344;
  assign n45346 = pi15 ? n12098 : n45345;
  assign n45347 = pi14 ? n45346 : n32;
  assign n45348 = pi13 ? n45340 : n45347;
  assign n45349 = pi12 ? n45335 : n45348;
  assign n45350 = pi11 ? n45326 : n45349;
  assign n45351 = pi15 ? n32 : n29676;
  assign n45352 = pi18 ? n21081 : ~n19966;
  assign n45353 = pi17 ? n4261 : n45352;
  assign n45354 = pi16 ? n1135 : ~n45353;
  assign n45355 = pi15 ? n45354 : n45251;
  assign n45356 = pi14 ? n45351 : n45355;
  assign n45357 = pi13 ? n32 : n45356;
  assign n45358 = pi12 ? n32 : n45357;
  assign n45359 = pi18 ? n366 : ~n21102;
  assign n45360 = pi17 ? n32 : n45359;
  assign n45361 = pi16 ? n45360 : ~n45270;
  assign n45362 = pi15 ? n45263 : n45361;
  assign n45363 = pi14 ? n45261 : n45362;
  assign n45364 = pi13 ? n45363 : n45279;
  assign n45365 = pi17 ? n45287 : n3337;
  assign n45366 = pi16 ? n45286 : ~n45365;
  assign n45367 = pi15 ? n45283 : n45366;
  assign n45368 = pi14 ? n31865 : n45367;
  assign n45369 = pi18 ? n366 : ~n31938;
  assign n45370 = pi17 ? n32 : n45369;
  assign n45371 = pi18 ? n31942 : n45302;
  assign n45372 = pi17 ? n45371 : n2325;
  assign n45373 = pi16 ? n45370 : ~n45372;
  assign n45374 = pi15 ? n45373 : n45308;
  assign n45375 = pi14 ? n45299 : n45374;
  assign n45376 = pi13 ? n45368 : n45375;
  assign n45377 = pi12 ? n45364 : n45376;
  assign n45378 = pi11 ? n45358 : n45377;
  assign n45379 = pi10 ? n45350 : n45378;
  assign n45380 = pi09 ? n32 : n45379;
  assign n45381 = pi08 ? n45315 : n45380;
  assign n45382 = pi07 ? n45184 : n45381;
  assign n45383 = pi15 ? n658 : n14613;
  assign n45384 = pi14 ? n45383 : n14613;
  assign n45385 = pi13 ? n45384 : n32;
  assign n45386 = pi19 ? n247 : n176;
  assign n45387 = pi18 ? n863 : ~n45386;
  assign n45388 = pi17 ? n32 : n45387;
  assign n45389 = pi16 ? n45388 : ~n2293;
  assign n45390 = pi15 ? n14613 : n45389;
  assign n45391 = pi19 ? n28477 : n31100;
  assign n45392 = pi18 ? n858 : n45391;
  assign n45393 = pi17 ? n32 : n45392;
  assign n45394 = pi16 ? n45393 : ~n2293;
  assign n45395 = pi20 ? n6621 : ~n246;
  assign n45396 = pi19 ? n19141 : n45395;
  assign n45397 = pi18 ? n45396 : ~n32;
  assign n45398 = pi17 ? n45397 : ~n2408;
  assign n45399 = pi16 ? n32 : n45398;
  assign n45400 = pi15 ? n45394 : n45399;
  assign n45401 = pi14 ? n45390 : n45400;
  assign n45402 = pi17 ? n36742 : ~n2408;
  assign n45403 = pi16 ? n32 : n45402;
  assign n45404 = pi20 ? n1331 : n2358;
  assign n45405 = pi19 ? n45404 : ~n32;
  assign n45406 = pi18 ? n45405 : ~n532;
  assign n45407 = pi17 ? n17346 : n45406;
  assign n45408 = pi16 ? n32 : n45407;
  assign n45409 = pi15 ? n45403 : n45408;
  assign n45410 = pi14 ? n45409 : n31963;
  assign n45411 = pi13 ? n45401 : n45410;
  assign n45412 = pi12 ? n45385 : n45411;
  assign n45413 = pi18 ? n28193 : ~n797;
  assign n45414 = pi17 ? n17705 : n45413;
  assign n45415 = pi16 ? n32 : n45414;
  assign n45416 = pi20 ? n1817 : n266;
  assign n45417 = pi19 ? n1817 : n45416;
  assign n45418 = pi20 ? n175 : ~n220;
  assign n45419 = pi19 ? n29444 : ~n45418;
  assign n45420 = pi18 ? n45417 : ~n45419;
  assign n45421 = pi18 ? n20605 : n797;
  assign n45422 = pi17 ? n45420 : ~n45421;
  assign n45423 = pi16 ? n21739 : n45422;
  assign n45424 = pi15 ? n45415 : n45423;
  assign n45425 = pi20 ? n17669 : n354;
  assign n45426 = pi19 ? n32 : n45425;
  assign n45427 = pi20 ? n3523 : n749;
  assign n45428 = pi19 ? n45427 : ~n32;
  assign n45429 = pi18 ? n45426 : ~n45428;
  assign n45430 = pi17 ? n32 : n45429;
  assign n45431 = pi16 ? n32 : n45430;
  assign n45432 = pi15 ? n45431 : n22167;
  assign n45433 = pi14 ? n45424 : n45432;
  assign n45434 = pi20 ? n428 : n518;
  assign n45435 = pi19 ? n45434 : ~n32;
  assign n45436 = pi18 ? n45435 : ~n797;
  assign n45437 = pi17 ? n32 : n45436;
  assign n45438 = pi16 ? n32 : n45437;
  assign n45439 = pi15 ? n45438 : n11856;
  assign n45440 = pi15 ? n22170 : n22162;
  assign n45441 = pi14 ? n45439 : n45440;
  assign n45442 = pi13 ? n45433 : n45441;
  assign n45443 = pi18 ? n8819 : ~n532;
  assign n45444 = pi17 ? n32 : n45443;
  assign n45445 = pi16 ? n32 : n45444;
  assign n45446 = pi15 ? n45445 : n13948;
  assign n45447 = pi14 ? n45446 : n31981;
  assign n45448 = pi18 ? n863 : n6059;
  assign n45449 = pi17 ? n32 : n45448;
  assign n45450 = pi16 ? n32 : n45449;
  assign n45451 = pi15 ? n45450 : n20477;
  assign n45452 = pi14 ? n45451 : n32;
  assign n45453 = pi13 ? n45447 : n45452;
  assign n45454 = pi12 ? n45442 : n45453;
  assign n45455 = pi11 ? n45412 : n45454;
  assign n45456 = pi16 ? n1233 : ~n32034;
  assign n45457 = pi15 ? n32 : n45456;
  assign n45458 = pi17 ? n18437 : n32041;
  assign n45459 = pi16 ? n1214 : ~n45458;
  assign n45460 = pi15 ? n32277 : n45459;
  assign n45461 = pi14 ? n45457 : n45460;
  assign n45462 = pi13 ? n32 : n45461;
  assign n45463 = pi12 ? n32 : n45462;
  assign n45464 = pi18 ? n21283 : n32;
  assign n45465 = pi17 ? n32 : ~n45464;
  assign n45466 = pi16 ? n1135 : ~n45465;
  assign n45467 = pi17 ? n21288 : ~n32;
  assign n45468 = pi16 ? n1135 : ~n45467;
  assign n45469 = pi15 ? n45466 : n45468;
  assign n45470 = pi18 ? n940 : ~n21292;
  assign n45471 = pi17 ? n32 : n45470;
  assign n45472 = pi18 ? n21299 : n6059;
  assign n45473 = pi17 ? n21298 : ~n45472;
  assign n45474 = pi16 ? n45471 : ~n45473;
  assign n45475 = pi15 ? n45474 : n31854;
  assign n45476 = pi14 ? n45469 : n45475;
  assign n45477 = pi15 ? n31854 : n30941;
  assign n45478 = pi16 ? n20208 : ~n2540;
  assign n45479 = pi20 ? n18261 : ~n32;
  assign n45480 = pi19 ? n45479 : ~n32;
  assign n45481 = pi18 ? n32 : n45480;
  assign n45482 = pi17 ? n32 : n45481;
  assign n45483 = pi18 ? n32 : n20345;
  assign n45484 = pi17 ? n32 : n45483;
  assign n45485 = pi16 ? n45482 : ~n45484;
  assign n45486 = pi15 ? n45478 : n45485;
  assign n45487 = pi14 ? n45477 : n45486;
  assign n45488 = pi13 ? n45476 : n45487;
  assign n45489 = pi19 ? n32082 : ~n9724;
  assign n45490 = pi18 ? n32081 : n45489;
  assign n45491 = pi17 ? n45490 : ~n2319;
  assign n45492 = pi16 ? n23483 : n45491;
  assign n45493 = pi19 ? n1464 : ~n208;
  assign n45494 = pi19 ? n5688 : ~n1757;
  assign n45495 = pi18 ? n45493 : n45494;
  assign n45496 = pi17 ? n45495 : ~n2319;
  assign n45497 = pi16 ? n23483 : n45496;
  assign n45498 = pi15 ? n45492 : n45497;
  assign n45499 = pi19 ? n32 : ~n4391;
  assign n45500 = pi18 ? n45499 : n684;
  assign n45501 = pi17 ? n45500 : ~n2319;
  assign n45502 = pi16 ? n32 : n45501;
  assign n45503 = pi19 ? n8622 : ~n18677;
  assign n45504 = pi18 ? n32 : n45503;
  assign n45505 = pi17 ? n32 : n45504;
  assign n45506 = pi19 ? n23895 : ~n5688;
  assign n45507 = pi19 ? n6988 : ~n349;
  assign n45508 = pi18 ? n45506 : ~n45507;
  assign n45509 = pi17 ? n45508 : ~n2537;
  assign n45510 = pi16 ? n45505 : n45509;
  assign n45511 = pi15 ? n45502 : n45510;
  assign n45512 = pi14 ? n45498 : n45511;
  assign n45513 = pi19 ? n221 : ~n8818;
  assign n45514 = pi18 ? n5667 : n45513;
  assign n45515 = pi17 ? n45514 : n2325;
  assign n45516 = pi16 ? n1135 : ~n45515;
  assign n45517 = pi15 ? n29135 : n45516;
  assign n45518 = pi18 ? n36293 : n31033;
  assign n45519 = pi17 ? n45518 : ~n2136;
  assign n45520 = pi16 ? n129 : n45519;
  assign n45521 = pi20 ? n1385 : ~n11107;
  assign n45522 = pi19 ? n349 : ~n45521;
  assign n45523 = pi18 ? n127 : n45522;
  assign n45524 = pi17 ? n32 : n45523;
  assign n45525 = pi17 ? n18017 : n2136;
  assign n45526 = pi16 ? n45524 : ~n45525;
  assign n45527 = pi15 ? n45520 : n45526;
  assign n45528 = pi14 ? n45517 : n45527;
  assign n45529 = pi13 ? n45512 : n45528;
  assign n45530 = pi12 ? n45488 : n45529;
  assign n45531 = pi11 ? n45463 : n45530;
  assign n45532 = pi10 ? n45455 : n45531;
  assign n45533 = pi09 ? n32 : n45532;
  assign n45534 = pi14 ? n21319 : n14613;
  assign n45535 = pi13 ? n45534 : n32;
  assign n45536 = pi16 ? n45388 : ~n3769;
  assign n45537 = pi15 ? n21319 : n45536;
  assign n45538 = pi20 ? n18415 : n18253;
  assign n45539 = pi19 ? n45538 : ~n31100;
  assign n45540 = pi18 ? n28770 : ~n45539;
  assign n45541 = pi17 ? n32 : n45540;
  assign n45542 = pi16 ? n45541 : ~n3769;
  assign n45543 = pi15 ? n45542 : n45399;
  assign n45544 = pi14 ? n45537 : n45543;
  assign n45545 = pi13 ? n45544 : n45410;
  assign n45546 = pi12 ? n45535 : n45545;
  assign n45547 = pi18 ? n28193 : ~n2291;
  assign n45548 = pi17 ? n17705 : n45547;
  assign n45549 = pi16 ? n32 : n45548;
  assign n45550 = pi15 ? n45549 : n45423;
  assign n45551 = pi19 ? n32 : n28893;
  assign n45552 = pi18 ? n45551 : ~n797;
  assign n45553 = pi17 ? n32 : n45552;
  assign n45554 = pi16 ? n32 : n45553;
  assign n45555 = pi15 ? n45554 : n22167;
  assign n45556 = pi14 ? n45550 : n45555;
  assign n45557 = pi13 ? n45556 : n45441;
  assign n45558 = pi14 ? n45446 : n12095;
  assign n45559 = pi15 ? n45450 : n13952;
  assign n45560 = pi14 ? n45559 : n32;
  assign n45561 = pi13 ? n45558 : n45560;
  assign n45562 = pi12 ? n45557 : n45561;
  assign n45563 = pi11 ? n45546 : n45562;
  assign n45564 = pi16 ? n1135 : ~n32034;
  assign n45565 = pi15 ? n32 : n45564;
  assign n45566 = pi15 ? n32039 : n45459;
  assign n45567 = pi14 ? n45565 : n45566;
  assign n45568 = pi13 ? n32 : n45567;
  assign n45569 = pi12 ? n32 : n45568;
  assign n45570 = pi15 ? n45474 : n32021;
  assign n45571 = pi14 ? n45469 : n45570;
  assign n45572 = pi16 ? n1233 : ~n1934;
  assign n45573 = pi16 ? n1233 : ~n45484;
  assign n45574 = pi15 ? n45572 : n45573;
  assign n45575 = pi16 ? n20208 : ~n2320;
  assign n45576 = pi15 ? n45575 : n45485;
  assign n45577 = pi14 ? n45574 : n45576;
  assign n45578 = pi13 ? n45571 : n45577;
  assign n45579 = pi17 ? n45508 : ~n3337;
  assign n45580 = pi16 ? n45505 : n45579;
  assign n45581 = pi15 ? n45502 : n45580;
  assign n45582 = pi14 ? n45498 : n45581;
  assign n45583 = pi16 ? n1233 : ~n45515;
  assign n45584 = pi15 ? n29135 : n45583;
  assign n45585 = pi16 ? n32 : n45519;
  assign n45586 = pi18 ? n32 : n45522;
  assign n45587 = pi17 ? n32 : n45586;
  assign n45588 = pi16 ? n45587 : ~n45525;
  assign n45589 = pi15 ? n45585 : n45588;
  assign n45590 = pi14 ? n45584 : n45589;
  assign n45591 = pi13 ? n45582 : n45590;
  assign n45592 = pi12 ? n45578 : n45591;
  assign n45593 = pi11 ? n45569 : n45592;
  assign n45594 = pi10 ? n45563 : n45593;
  assign n45595 = pi09 ? n32 : n45594;
  assign n45596 = pi08 ? n45533 : n45595;
  assign n45597 = pi14 ? n21389 : n21319;
  assign n45598 = pi13 ? n45597 : n32;
  assign n45599 = pi19 ? n32 : n32847;
  assign n45600 = pi18 ? n45599 : ~n9170;
  assign n45601 = pi17 ? n32 : n45600;
  assign n45602 = pi16 ? n45601 : ~n3769;
  assign n45603 = pi15 ? n21319 : n45602;
  assign n45604 = pi16 ? n32 : ~n3769;
  assign n45605 = pi18 ? n18668 : ~n248;
  assign n45606 = pi17 ? n45605 : ~n2408;
  assign n45607 = pi16 ? n32 : n45606;
  assign n45608 = pi15 ? n45604 : n45607;
  assign n45609 = pi14 ? n45603 : n45608;
  assign n45610 = pi19 ? n19116 : n32;
  assign n45611 = pi18 ? n45610 : n797;
  assign n45612 = pi17 ? n2512 : ~n45611;
  assign n45613 = pi16 ? n32 : n45612;
  assign n45614 = pi18 ? n508 : ~n22159;
  assign n45615 = pi17 ? n32 : n45614;
  assign n45616 = pi16 ? n32 : n45615;
  assign n45617 = pi15 ? n45613 : n45616;
  assign n45618 = pi14 ? n45617 : n32198;
  assign n45619 = pi13 ? n45609 : n45618;
  assign n45620 = pi12 ? n45598 : n45619;
  assign n45621 = pi19 ? n1844 : n3523;
  assign n45622 = pi18 ? n19082 : n45621;
  assign n45623 = pi17 ? n32 : n45622;
  assign n45624 = pi20 ? n339 : n354;
  assign n45625 = pi19 ? n339 : n45624;
  assign n45626 = pi20 ? n1331 : n357;
  assign n45627 = pi19 ? n45626 : n29002;
  assign n45628 = pi18 ? n45625 : ~n45627;
  assign n45629 = pi20 ? n310 : ~n32;
  assign n45630 = pi19 ? n45629 : ~n32;
  assign n45631 = pi18 ? n45630 : ~n2291;
  assign n45632 = pi17 ? n45628 : ~n45631;
  assign n45633 = pi16 ? n45623 : ~n45632;
  assign n45634 = pi15 ? n45633 : n32210;
  assign n45635 = pi18 ? n697 : ~n2291;
  assign n45636 = pi17 ? n32 : n45635;
  assign n45637 = pi16 ? n32 : n45636;
  assign n45638 = pi18 ? n702 : ~n2291;
  assign n45639 = pi17 ? n32 : n45638;
  assign n45640 = pi16 ? n32 : n45639;
  assign n45641 = pi15 ? n45637 : n45640;
  assign n45642 = pi14 ? n45634 : n45641;
  assign n45643 = pi18 ? n25110 : ~n2291;
  assign n45644 = pi17 ? n19803 : n45643;
  assign n45645 = pi16 ? n32 : n45644;
  assign n45646 = pi15 ? n45645 : n32210;
  assign n45647 = pi15 ? n45637 : n22313;
  assign n45648 = pi14 ? n45646 : n45647;
  assign n45649 = pi13 ? n45642 : n45648;
  assign n45650 = pi18 ? n8819 : ~n797;
  assign n45651 = pi17 ? n32 : n45650;
  assign n45652 = pi16 ? n32 : n45651;
  assign n45653 = pi15 ? n45652 : n13943;
  assign n45654 = pi14 ? n45653 : n32220;
  assign n45655 = pi15 ? n45450 : n32;
  assign n45656 = pi14 ? n45655 : n32;
  assign n45657 = pi13 ? n45654 : n45656;
  assign n45658 = pi12 ? n45649 : n45657;
  assign n45659 = pi11 ? n45620 : n45658;
  assign n45660 = pi20 ? n4279 : n1076;
  assign n45661 = pi20 ? n1076 : n4279;
  assign n45662 = pi19 ? n45660 : n45661;
  assign n45663 = pi18 ? n41883 : n45662;
  assign n45664 = pi17 ? n32 : n45663;
  assign n45665 = pi19 ? n4279 : n18133;
  assign n45666 = pi20 ? n287 : n310;
  assign n45667 = pi19 ? n6050 : n45666;
  assign n45668 = pi18 ? n45665 : ~n45667;
  assign n45669 = pi20 ? n785 : ~n2358;
  assign n45670 = pi19 ? n45669 : n29277;
  assign n45671 = pi18 ? n45670 : ~n618;
  assign n45672 = pi17 ? n45668 : n45671;
  assign n45673 = pi16 ? n45664 : n45672;
  assign n45674 = pi15 ? n45673 : n45456;
  assign n45675 = pi16 ? n1233 : ~n32038;
  assign n45676 = pi15 ? n45675 : n32279;
  assign n45677 = pi14 ? n45674 : n45676;
  assign n45678 = pi13 ? n32 : n45677;
  assign n45679 = pi12 ? n32 : n45678;
  assign n45680 = pi18 ? n21443 : ~n32;
  assign n45681 = pi17 ? n32 : n45680;
  assign n45682 = pi16 ? n1233 : ~n45681;
  assign n45683 = pi16 ? n1233 : ~n3436;
  assign n45684 = pi15 ? n45682 : n45683;
  assign n45685 = pi18 ? n18710 : ~n32025;
  assign n45686 = pi17 ? n32 : n45685;
  assign n45687 = pi16 ? n45686 : ~n2530;
  assign n45688 = pi15 ? n45687 : n32021;
  assign n45689 = pi14 ? n45684 : n45688;
  assign n45690 = pi19 ? n236 : ~n9007;
  assign n45691 = pi18 ? n341 : n45690;
  assign n45692 = pi17 ? n32 : n45691;
  assign n45693 = pi19 ? n207 : n9345;
  assign n45694 = pi18 ? n45693 : ~n20020;
  assign n45695 = pi17 ? n45694 : ~n1933;
  assign n45696 = pi16 ? n45692 : n45695;
  assign n45697 = pi15 ? n32021 : n45696;
  assign n45698 = pi18 ? n32 : ~n34006;
  assign n45699 = pi17 ? n32 : n45698;
  assign n45700 = pi17 ? n13946 : n1933;
  assign n45701 = pi16 ? n45699 : ~n45700;
  assign n45702 = pi19 ? n4982 : ~n22525;
  assign n45703 = pi18 ? n32 : n45702;
  assign n45704 = pi17 ? n32 : n45703;
  assign n45705 = pi18 ? n23073 : ~n32;
  assign n45706 = pi17 ? n45705 : ~n1933;
  assign n45707 = pi16 ? n45704 : n45706;
  assign n45708 = pi15 ? n45701 : n45707;
  assign n45709 = pi14 ? n45697 : n45708;
  assign n45710 = pi13 ? n45689 : n45709;
  assign n45711 = pi19 ? n32 : n20923;
  assign n45712 = pi18 ? n5657 : n45711;
  assign n45713 = pi17 ? n45712 : ~n1933;
  assign n45714 = pi16 ? n32 : n45713;
  assign n45715 = pi18 ? n618 : ~n344;
  assign n45716 = pi17 ? n32316 : n45715;
  assign n45717 = pi16 ? n32 : n45716;
  assign n45718 = pi15 ? n45714 : n45717;
  assign n45719 = pi18 ? n20164 : n880;
  assign n45720 = pi17 ? n45719 : ~n1933;
  assign n45721 = pi16 ? n32 : n45720;
  assign n45722 = pi20 ? n518 : ~n1685;
  assign n45723 = pi19 ? n9007 : ~n45722;
  assign n45724 = pi18 ? n863 : n45723;
  assign n45725 = pi17 ? n32 : n45724;
  assign n45726 = pi20 ? n1685 : ~n342;
  assign n45727 = pi19 ? n45726 : ~n322;
  assign n45728 = pi19 ? n18478 : ~n1757;
  assign n45729 = pi18 ? n45727 : n45728;
  assign n45730 = pi17 ? n45729 : ~n1807;
  assign n45731 = pi16 ? n45725 : n45730;
  assign n45732 = pi15 ? n45721 : n45731;
  assign n45733 = pi14 ? n45718 : n45732;
  assign n45734 = pi16 ? n20208 : ~n1808;
  assign n45735 = pi20 ? n1385 : ~n310;
  assign n45736 = pi20 ? n333 : ~n8644;
  assign n45737 = pi19 ? n45735 : ~n45736;
  assign n45738 = pi18 ? n936 : ~n45737;
  assign n45739 = pi17 ? n32 : n45738;
  assign n45740 = pi20 ? n8644 : n1076;
  assign n45741 = pi20 ? n7839 : n18245;
  assign n45742 = pi19 ? n45740 : ~n45741;
  assign n45743 = pi20 ? n321 : n18762;
  assign n45744 = pi19 ? n45743 : n8818;
  assign n45745 = pi18 ? n45742 : ~n45744;
  assign n45746 = pi20 ? n274 : ~n287;
  assign n45747 = pi19 ? n32 : n45746;
  assign n45748 = pi18 ? n45747 : ~n19654;
  assign n45749 = pi17 ? n45745 : n45748;
  assign n45750 = pi16 ? n45739 : ~n45749;
  assign n45751 = pi15 ? n45734 : n45750;
  assign n45752 = pi18 ? n14648 : n323;
  assign n45753 = pi17 ? n45752 : ~n2136;
  assign n45754 = pi16 ? n129 : n45753;
  assign n45755 = pi19 ? n349 : ~n5371;
  assign n45756 = pi18 ? n127 : n45755;
  assign n45757 = pi17 ? n32 : n45756;
  assign n45758 = pi16 ? n45757 : ~n45525;
  assign n45759 = pi15 ? n45754 : n45758;
  assign n45760 = pi14 ? n45751 : n45759;
  assign n45761 = pi13 ? n45733 : n45760;
  assign n45762 = pi12 ? n45710 : n45761;
  assign n45763 = pi11 ? n45679 : n45762;
  assign n45764 = pi10 ? n45659 : n45763;
  assign n45765 = pi09 ? n32 : n45764;
  assign n45766 = pi13 ? n45597 : n21466;
  assign n45767 = pi21 ? n8275 : ~n309;
  assign n45768 = pi20 ? n32 : n45767;
  assign n45769 = pi19 ? n32 : n45768;
  assign n45770 = pi18 ? n45769 : ~n9170;
  assign n45771 = pi17 ? n32 : n45770;
  assign n45772 = pi16 ? n45771 : ~n2756;
  assign n45773 = pi15 ? n21464 : n45772;
  assign n45774 = pi16 ? n32 : ~n2756;
  assign n45775 = pi17 ? n45605 : ~n2519;
  assign n45776 = pi16 ? n32 : n45775;
  assign n45777 = pi15 ? n45774 : n45776;
  assign n45778 = pi14 ? n45773 : n45777;
  assign n45779 = pi18 ? n45610 : n323;
  assign n45780 = pi17 ? n2512 : ~n45779;
  assign n45781 = pi16 ? n32 : n45780;
  assign n45782 = pi15 ? n45781 : n45616;
  assign n45783 = pi14 ? n45782 : n32198;
  assign n45784 = pi13 ? n45778 : n45783;
  assign n45785 = pi12 ? n45766 : n45784;
  assign n45786 = pi20 ? n820 : n339;
  assign n45787 = pi20 ? n339 : n18540;
  assign n45788 = pi19 ? n45786 : n45787;
  assign n45789 = pi20 ? n18415 : ~n6085;
  assign n45790 = pi19 ? n45789 : ~n28338;
  assign n45791 = pi18 ? n45788 : n45790;
  assign n45792 = pi18 ? n44957 : ~n323;
  assign n45793 = pi17 ? n45791 : ~n45792;
  assign n45794 = pi16 ? n45623 : ~n45793;
  assign n45795 = pi15 ? n45794 : n11856;
  assign n45796 = pi14 ? n45795 : n45641;
  assign n45797 = pi18 ? n25110 : ~n32919;
  assign n45798 = pi17 ? n19803 : n45797;
  assign n45799 = pi16 ? n32 : n45798;
  assign n45800 = pi15 ? n45799 : n32210;
  assign n45801 = pi14 ? n45800 : n45647;
  assign n45802 = pi13 ? n45796 : n45801;
  assign n45803 = pi18 ? n8819 : ~n2291;
  assign n45804 = pi17 ? n32 : n45803;
  assign n45805 = pi16 ? n32 : n45804;
  assign n45806 = pi15 ? n45805 : n13943;
  assign n45807 = pi14 ? n45806 : n32379;
  assign n45808 = pi20 ? n266 : n52;
  assign n45809 = pi19 ? n45808 : n32;
  assign n45810 = pi18 ? n863 : n45809;
  assign n45811 = pi17 ? n32 : n45810;
  assign n45812 = pi16 ? n32 : n45811;
  assign n45813 = pi15 ? n45812 : n32;
  assign n45814 = pi14 ? n45813 : n32;
  assign n45815 = pi13 ? n45807 : n45814;
  assign n45816 = pi12 ? n45802 : n45815;
  assign n45817 = pi11 ? n45785 : n45816;
  assign n45818 = pi20 ? n2019 : ~n501;
  assign n45819 = pi20 ? n501 : ~n2019;
  assign n45820 = pi19 ? n45818 : ~n45819;
  assign n45821 = pi18 ? n222 : ~n45820;
  assign n45822 = pi17 ? n32 : n45821;
  assign n45823 = pi21 ? n173 : n405;
  assign n45824 = pi20 ? n45823 : n17669;
  assign n45825 = pi19 ? n2019 : n45824;
  assign n45826 = pi20 ? n6050 : n29457;
  assign n45827 = pi20 ? n18624 : n1331;
  assign n45828 = pi19 ? n45826 : n45827;
  assign n45829 = pi18 ? n45825 : n45828;
  assign n45830 = pi20 ? n309 : n1377;
  assign n45831 = pi20 ? n6621 : ~n2385;
  assign n45832 = pi19 ? n45830 : ~n45831;
  assign n45833 = pi18 ? n45832 : n32390;
  assign n45834 = pi17 ? n45829 : n45833;
  assign n45835 = pi16 ? n45822 : ~n45834;
  assign n45836 = pi16 ? n1135 : ~n32415;
  assign n45837 = pi15 ? n45835 : n45836;
  assign n45838 = pi16 ? n1135 : ~n32419;
  assign n45839 = pi15 ? n45838 : n32423;
  assign n45840 = pi14 ? n45837 : n45839;
  assign n45841 = pi13 ? n32 : n45840;
  assign n45842 = pi12 ? n32 : n45841;
  assign n45843 = pi16 ? n1135 : ~n45681;
  assign n45844 = pi16 ? n1135 : ~n3436;
  assign n45845 = pi15 ? n45843 : n45844;
  assign n45846 = pi15 ? n45687 : n34377;
  assign n45847 = pi14 ? n45845 : n45846;
  assign n45848 = pi18 ? n127 : ~n34006;
  assign n45849 = pi17 ? n32 : n45848;
  assign n45850 = pi16 ? n45849 : ~n45700;
  assign n45851 = pi15 ? n45850 : n45707;
  assign n45852 = pi14 ? n45697 : n45851;
  assign n45853 = pi13 ? n45847 : n45852;
  assign n45854 = pi17 ? n32434 : n45715;
  assign n45855 = pi16 ? n32 : n45854;
  assign n45856 = pi15 ? n45714 : n45855;
  assign n45857 = pi14 ? n45856 : n45732;
  assign n45858 = pi20 ? n321 : ~n310;
  assign n45859 = pi20 ? n3523 : ~n785;
  assign n45860 = pi19 ? n45858 : ~n45859;
  assign n45861 = pi18 ? n32 : ~n45860;
  assign n45862 = pi17 ? n32 : n45861;
  assign n45863 = pi20 ? n785 : n501;
  assign n45864 = pi20 ? n7839 : n12884;
  assign n45865 = pi19 ? n45863 : ~n45864;
  assign n45866 = pi19 ? n22038 : n8818;
  assign n45867 = pi18 ? n45865 : ~n45866;
  assign n45868 = pi19 ? n8622 : n28957;
  assign n45869 = pi18 ? n45868 : ~n19654;
  assign n45870 = pi17 ? n45867 : n45869;
  assign n45871 = pi16 ? n45862 : ~n45870;
  assign n45872 = pi15 ? n45734 : n45871;
  assign n45873 = pi14 ? n45872 : n45759;
  assign n45874 = pi13 ? n45857 : n45873;
  assign n45875 = pi12 ? n45853 : n45874;
  assign n45876 = pi11 ? n45842 : n45875;
  assign n45877 = pi10 ? n45817 : n45876;
  assign n45878 = pi09 ? n32 : n45877;
  assign n45879 = pi08 ? n45765 : n45878;
  assign n45880 = pi07 ? n45596 : n45879;
  assign n45881 = pi06 ? n45382 : n45880;
  assign n45882 = pi05 ? n45011 : n45881;
  assign n45883 = pi04 ? n44020 : n45882;
  assign n45884 = pi03 ? n42476 : n45883;
  assign n45885 = pi14 ? n21543 : n21464;
  assign n45886 = pi18 ? n323 : n350;
  assign n45887 = pi17 ? n45886 : ~n2531;
  assign n45888 = pi16 ? n32 : n45887;
  assign n45889 = pi18 ? n32 : n39598;
  assign n45890 = pi17 ? n45886 : ~n45889;
  assign n45891 = pi16 ? n32 : n45890;
  assign n45892 = pi15 ? n45888 : n45891;
  assign n45893 = pi14 ? n32 : n45892;
  assign n45894 = pi13 ? n45885 : n45893;
  assign n45895 = pi20 ? n17669 : n17665;
  assign n45896 = pi19 ? n45895 : n30044;
  assign n45897 = pi18 ? n29681 : ~n45896;
  assign n45898 = pi17 ? n32 : n45897;
  assign n45899 = pi19 ? n18789 : n32;
  assign n45900 = pi18 ? n45899 : n32;
  assign n45901 = pi17 ? n45900 : n2755;
  assign n45902 = pi16 ? n45898 : ~n45901;
  assign n45903 = pi16 ? n1214 : ~n2756;
  assign n45904 = pi15 ? n45902 : n45903;
  assign n45905 = pi20 ? n206 : n220;
  assign n45906 = pi19 ? n45905 : n1248;
  assign n45907 = pi18 ? n863 : n45906;
  assign n45908 = pi17 ? n32 : n45907;
  assign n45909 = pi17 ? n18482 : n2755;
  assign n45910 = pi16 ? n45908 : ~n45909;
  assign n45911 = pi18 ? n32 : n25110;
  assign n45912 = pi18 ? n9012 : n323;
  assign n45913 = pi17 ? n45911 : ~n45912;
  assign n45914 = pi16 ? n18293 : n45913;
  assign n45915 = pi15 ? n45910 : n45914;
  assign n45916 = pi14 ? n45904 : n45915;
  assign n45917 = pi18 ? n1750 : ~n532;
  assign n45918 = pi17 ? n32 : n45917;
  assign n45919 = pi16 ? n32 : n45918;
  assign n45920 = pi15 ? n45919 : n20883;
  assign n45921 = pi14 ? n45920 : n32462;
  assign n45922 = pi13 ? n45916 : n45921;
  assign n45923 = pi12 ? n45894 : n45922;
  assign n45924 = pi19 ? n3692 : n321;
  assign n45925 = pi18 ? n222 : n45924;
  assign n45926 = pi17 ? n32 : n45925;
  assign n45927 = pi19 ? n1490 : n18390;
  assign n45928 = pi19 ? n1464 : n17766;
  assign n45929 = pi18 ? n45927 : n45928;
  assign n45930 = pi17 ? n45929 : n2519;
  assign n45931 = pi16 ? n45926 : ~n45930;
  assign n45932 = pi15 ? n45931 : n32468;
  assign n45933 = pi19 ? n322 : n4406;
  assign n45934 = pi18 ? n45933 : ~n323;
  assign n45935 = pi17 ? n32 : n45934;
  assign n45936 = pi16 ? n32 : n45935;
  assign n45937 = pi15 ? n45936 : n32468;
  assign n45938 = pi14 ? n45932 : n45937;
  assign n45939 = pi18 ? n496 : ~n323;
  assign n45940 = pi17 ? n32 : n45939;
  assign n45941 = pi16 ? n32 : n45940;
  assign n45942 = pi15 ? n32828 : n45941;
  assign n45943 = pi14 ? n45942 : n45941;
  assign n45944 = pi13 ? n45938 : n45943;
  assign n45945 = pi18 ? n32 : n32478;
  assign n45946 = pi17 ? n32 : n45945;
  assign n45947 = pi16 ? n32 : n45946;
  assign n45948 = pi15 ? n45947 : n20660;
  assign n45949 = pi14 ? n45948 : n32482;
  assign n45950 = pi13 ? n45949 : n32;
  assign n45951 = pi12 ? n45944 : n45950;
  assign n45952 = pi11 ? n45923 : n45951;
  assign n45953 = pi13 ? n20831 : n32;
  assign n45954 = pi18 ? n42797 : n6059;
  assign n45955 = pi17 ? n32 : n45954;
  assign n45956 = pi16 ? n32 : n45955;
  assign n45957 = pi15 ? n32 : n45956;
  assign n45958 = pi14 ? n32 : n45957;
  assign n45959 = pi17 ? n21582 : n1500;
  assign n45960 = pi16 ? n1135 : ~n45959;
  assign n45961 = pi15 ? n45960 : n32526;
  assign n45962 = pi18 ? n21595 : n237;
  assign n45963 = pi17 ? n32 : n45962;
  assign n45964 = pi16 ? n1135 : ~n45963;
  assign n45965 = pi15 ? n45964 : n32530;
  assign n45966 = pi14 ? n45961 : n45965;
  assign n45967 = pi13 ? n45958 : n45966;
  assign n45968 = pi12 ? n45953 : n45967;
  assign n45969 = pi16 ? n1214 : ~n2530;
  assign n45970 = pi15 ? n31056 : n45969;
  assign n45971 = pi14 ? n45970 : n32021;
  assign n45972 = pi16 ? n3625 : ~n2306;
  assign n45973 = pi15 ? n32021 : n45972;
  assign n45974 = pi14 ? n32154 : n45973;
  assign n45975 = pi13 ? n45971 : n45974;
  assign n45976 = pi18 ? n29802 : n496;
  assign n45977 = pi17 ? n45976 : ~n2305;
  assign n45978 = pi16 ? n32 : n45977;
  assign n45979 = pi18 ? n19232 : n2304;
  assign n45980 = pi17 ? n3164 : ~n45979;
  assign n45981 = pi16 ? n32 : n45980;
  assign n45982 = pi15 ? n45978 : n45981;
  assign n45983 = pi18 ? n16449 : n940;
  assign n45984 = pi17 ? n45983 : ~n1933;
  assign n45985 = pi16 ? n32 : n45984;
  assign n45986 = pi17 ? n18487 : n1807;
  assign n45987 = pi16 ? n1471 : ~n45986;
  assign n45988 = pi15 ? n45985 : n45987;
  assign n45989 = pi14 ? n45982 : n45988;
  assign n45990 = pi18 ? n1395 : ~n20164;
  assign n45991 = pi17 ? n32 : n45990;
  assign n45992 = pi19 ? n25120 : ~n4391;
  assign n45993 = pi18 ? n15241 : n45992;
  assign n45994 = pi17 ? n45993 : n1807;
  assign n45995 = pi16 ? n45991 : ~n45994;
  assign n45996 = pi19 ? n236 : ~n321;
  assign n45997 = pi18 ? n25760 : ~n45996;
  assign n45998 = pi17 ? n45997 : ~n1807;
  assign n45999 = pi16 ? n32 : n45998;
  assign n46000 = pi15 ? n45995 : n45999;
  assign n46001 = pi18 ? n463 : n30574;
  assign n46002 = pi17 ? n32 : n46001;
  assign n46003 = pi19 ? n32 : ~n5435;
  assign n46004 = pi19 ? n22652 : n207;
  assign n46005 = pi18 ? n46003 : n46004;
  assign n46006 = pi17 ? n46005 : ~n2314;
  assign n46007 = pi16 ? n46002 : n46006;
  assign n46008 = pi18 ? n463 : n15400;
  assign n46009 = pi17 ? n32 : n46008;
  assign n46010 = pi19 ? n9028 : ~n32;
  assign n46011 = pi18 ? n15570 : n46010;
  assign n46012 = pi17 ? n46011 : ~n1807;
  assign n46013 = pi16 ? n46009 : n46012;
  assign n46014 = pi15 ? n46007 : n46013;
  assign n46015 = pi14 ? n46000 : n46014;
  assign n46016 = pi13 ? n45989 : n46015;
  assign n46017 = pi12 ? n45975 : n46016;
  assign n46018 = pi11 ? n45968 : n46017;
  assign n46019 = pi10 ? n45952 : n46018;
  assign n46020 = pi09 ? n32 : n46019;
  assign n46021 = pi20 ? n32 : ~n382;
  assign n46022 = pi19 ? n46021 : ~n32;
  assign n46023 = pi18 ? n32 : n46022;
  assign n46024 = pi17 ? n45886 : ~n46023;
  assign n46025 = pi16 ? n32 : n46024;
  assign n46026 = pi15 ? n45888 : n46025;
  assign n46027 = pi14 ? n32 : n46026;
  assign n46028 = pi13 ? n45885 : n46027;
  assign n46029 = pi21 ? n1392 : n174;
  assign n46030 = pi20 ? n32 : n46029;
  assign n46031 = pi19 ? n32 : n46030;
  assign n46032 = pi18 ? n46031 : ~n45896;
  assign n46033 = pi17 ? n32 : n46032;
  assign n46034 = pi17 ? n45900 : n2517;
  assign n46035 = pi16 ? n46033 : ~n46034;
  assign n46036 = pi16 ? n1214 : ~n2518;
  assign n46037 = pi15 ? n46035 : n46036;
  assign n46038 = pi16 ? n45908 : ~n34661;
  assign n46039 = pi18 ? n9012 : n2754;
  assign n46040 = pi17 ? n45911 : ~n46039;
  assign n46041 = pi16 ? n18293 : n46040;
  assign n46042 = pi15 ? n46038 : n46041;
  assign n46043 = pi14 ? n46037 : n46042;
  assign n46044 = pi13 ? n46043 : n45921;
  assign n46045 = pi12 ? n46028 : n46044;
  assign n46046 = pi17 ? n45929 : n2755;
  assign n46047 = pi16 ? n45926 : ~n46046;
  assign n46048 = pi15 ? n46047 : n32468;
  assign n46049 = pi14 ? n46048 : n45937;
  assign n46050 = pi13 ? n46049 : n45943;
  assign n46051 = pi14 ? n45948 : n32614;
  assign n46052 = pi13 ? n46051 : n32;
  assign n46053 = pi12 ? n46050 : n46052;
  assign n46054 = pi11 ? n46045 : n46053;
  assign n46055 = pi15 ? n45960 : n32646;
  assign n46056 = pi14 ? n46055 : n45965;
  assign n46057 = pi13 ? n45958 : n46056;
  assign n46058 = pi12 ? n32 : n46057;
  assign n46059 = pi15 ? n31146 : n45969;
  assign n46060 = pi14 ? n46059 : n32021;
  assign n46061 = pi16 ? n3625 : ~n1934;
  assign n46062 = pi15 ? n32021 : n46061;
  assign n46063 = pi14 ? n32154 : n46062;
  assign n46064 = pi13 ? n46060 : n46063;
  assign n46065 = pi17 ? n45983 : ~n2305;
  assign n46066 = pi16 ? n32 : n46065;
  assign n46067 = pi15 ? n46066 : n45987;
  assign n46068 = pi14 ? n45982 : n46067;
  assign n46069 = pi16 ? n29305 : ~n45994;
  assign n46070 = pi15 ? n46069 : n45999;
  assign n46071 = pi18 ? n1012 : n30574;
  assign n46072 = pi17 ? n32 : n46071;
  assign n46073 = pi16 ? n46072 : n46006;
  assign n46074 = pi18 ? n1012 : n15400;
  assign n46075 = pi17 ? n32 : n46074;
  assign n46076 = pi16 ? n46075 : n46012;
  assign n46077 = pi15 ? n46073 : n46076;
  assign n46078 = pi14 ? n46070 : n46077;
  assign n46079 = pi13 ? n46068 : n46078;
  assign n46080 = pi12 ? n46064 : n46079;
  assign n46081 = pi11 ? n46058 : n46080;
  assign n46082 = pi10 ? n46054 : n46081;
  assign n46083 = pi09 ? n32 : n46082;
  assign n46084 = pi08 ? n46020 : n46083;
  assign n46085 = pi14 ? n21686 : n387;
  assign n46086 = pi18 ? n32 : n35545;
  assign n46087 = pi17 ? n45886 : ~n46086;
  assign n46088 = pi16 ? n32 : n46087;
  assign n46089 = pi15 ? n45888 : n46088;
  assign n46090 = pi14 ? n32 : n46089;
  assign n46091 = pi13 ? n46085 : n46090;
  assign n46092 = pi20 ? n10644 : ~n18762;
  assign n46093 = pi19 ? n19141 : n46092;
  assign n46094 = pi18 ? n46093 : ~n44474;
  assign n46095 = pi17 ? n46094 : ~n2517;
  assign n46096 = pi16 ? n32 : n46095;
  assign n46097 = pi19 ? n267 : n266;
  assign n46098 = pi18 ? n46097 : n605;
  assign n46099 = pi18 ? n21316 : n520;
  assign n46100 = pi17 ? n46098 : ~n46099;
  assign n46101 = pi16 ? n32 : n46100;
  assign n46102 = pi15 ? n46096 : n46101;
  assign n46103 = pi19 ? n32082 : n594;
  assign n46104 = pi18 ? n32 : n46103;
  assign n46105 = pi17 ? n32 : n46104;
  assign n46106 = pi19 ? n29145 : n5854;
  assign n46107 = pi19 ? n29294 : ~n358;
  assign n46108 = pi18 ? n46106 : n46107;
  assign n46109 = pi20 ? n333 : ~n2358;
  assign n46110 = pi19 ? n46109 : n1844;
  assign n46111 = pi18 ? n46110 : n520;
  assign n46112 = pi17 ? n46108 : ~n46111;
  assign n46113 = pi16 ? n46105 : n46112;
  assign n46114 = pi20 ? n220 : n10644;
  assign n46115 = pi19 ? n32 : n46114;
  assign n46116 = pi18 ? n32 : n46115;
  assign n46117 = pi18 ? n9008 : ~n323;
  assign n46118 = pi17 ? n46116 : n46117;
  assign n46119 = pi16 ? n32 : n46118;
  assign n46120 = pi15 ? n46113 : n46119;
  assign n46121 = pi14 ? n46102 : n46120;
  assign n46122 = pi18 ? n684 : ~n532;
  assign n46123 = pi17 ? n32 : n46122;
  assign n46124 = pi16 ? n32 : n46123;
  assign n46125 = pi15 ? n46124 : n20883;
  assign n46126 = pi14 ? n46125 : n32670;
  assign n46127 = pi13 ? n46121 : n46126;
  assign n46128 = pi12 ? n46091 : n46127;
  assign n46129 = pi20 ? n3523 : n1839;
  assign n46130 = pi19 ? n46129 : ~n32;
  assign n46131 = pi18 ? n356 : ~n46130;
  assign n46132 = pi17 ? n32 : n46131;
  assign n46133 = pi16 ? n32 : n46132;
  assign n46134 = pi15 ? n12083 : n46133;
  assign n46135 = pi14 ? n46134 : n12079;
  assign n46136 = pi18 ? n1741 : ~n2754;
  assign n46137 = pi17 ? n32 : n46136;
  assign n46138 = pi16 ? n32 : n46137;
  assign n46139 = pi15 ? n12083 : n46138;
  assign n46140 = pi18 ? n9038 : ~n2754;
  assign n46141 = pi17 ? n32 : n46140;
  assign n46142 = pi16 ? n32 : n46141;
  assign n46143 = pi18 ? n9029 : n33017;
  assign n46144 = pi17 ? n32 : n46143;
  assign n46145 = pi16 ? n32 : n46144;
  assign n46146 = pi15 ? n46142 : n46145;
  assign n46147 = pi14 ? n46139 : n46146;
  assign n46148 = pi13 ? n46135 : n46147;
  assign n46149 = pi15 ? n21346 : n32685;
  assign n46150 = pi14 ? n46149 : n32687;
  assign n46151 = pi13 ? n46150 : n32;
  assign n46152 = pi12 ? n46148 : n46151;
  assign n46153 = pi11 ? n46128 : n46152;
  assign n46154 = pi18 ? n15227 : n344;
  assign n46155 = pi17 ? n32 : n46154;
  assign n46156 = pi16 ? n1135 : ~n46155;
  assign n46157 = pi15 ? n32 : n46156;
  assign n46158 = pi14 ? n32 : n46157;
  assign n46159 = pi17 ? n17734 : n1500;
  assign n46160 = pi16 ? n1233 : ~n46159;
  assign n46161 = pi15 ? n46160 : n32741;
  assign n46162 = pi14 ? n46161 : n32748;
  assign n46163 = pi13 ? n46158 : n46162;
  assign n46164 = pi12 ? n32 : n46163;
  assign n46165 = pi18 ? n16389 : n350;
  assign n46166 = pi17 ? n32 : n46165;
  assign n46167 = pi16 ? n1135 : ~n46166;
  assign n46168 = pi15 ? n46167 : n32153;
  assign n46169 = pi16 ? n19652 : ~n2530;
  assign n46170 = pi14 ? n46168 : n46169;
  assign n46171 = pi15 ? n46169 : n45969;
  assign n46172 = pi16 ? n3625 : ~n2530;
  assign n46173 = pi15 ? n31828 : n46172;
  assign n46174 = pi14 ? n46171 : n46173;
  assign n46175 = pi13 ? n46170 : n46174;
  assign n46176 = pi19 ? n275 : n349;
  assign n46177 = pi18 ? n37120 : n46176;
  assign n46178 = pi17 ? n46177 : ~n2410;
  assign n46179 = pi16 ? n16983 : n46178;
  assign n46180 = pi18 ? n248 : n344;
  assign n46181 = pi17 ? n3164 : ~n46180;
  assign n46182 = pi16 ? n32 : n46181;
  assign n46183 = pi15 ? n46179 : n46182;
  assign n46184 = pi20 ? n428 : n266;
  assign n46185 = pi19 ? n32 : n46184;
  assign n46186 = pi18 ? n46185 : n12368;
  assign n46187 = pi17 ? n46186 : ~n1933;
  assign n46188 = pi16 ? n32 : n46187;
  assign n46189 = pi15 ? n46188 : n45987;
  assign n46190 = pi14 ? n46183 : n46189;
  assign n46191 = pi20 ? n5854 : n260;
  assign n46192 = pi19 ? n46191 : ~n5675;
  assign n46193 = pi18 ? n28748 : ~n46192;
  assign n46194 = pi17 ? n32 : n46193;
  assign n46195 = pi19 ? n1844 : n34188;
  assign n46196 = pi19 ? n22185 : ~n4391;
  assign n46197 = pi18 ? n46195 : ~n46196;
  assign n46198 = pi17 ? n46197 : ~n1807;
  assign n46199 = pi16 ? n46194 : n46198;
  assign n46200 = pi19 ? n22185 : ~n31490;
  assign n46201 = pi18 ? n39110 : ~n46200;
  assign n46202 = pi17 ? n46201 : ~n1807;
  assign n46203 = pi16 ? n17347 : n46202;
  assign n46204 = pi15 ? n46199 : n46203;
  assign n46205 = pi17 ? n32 : n34278;
  assign n46206 = pi20 ? n2385 : n18762;
  assign n46207 = pi19 ? n6057 : n46206;
  assign n46208 = pi20 ? n287 : ~n17665;
  assign n46209 = pi19 ? n23709 : n46208;
  assign n46210 = pi18 ? n46207 : n46209;
  assign n46211 = pi17 ? n46210 : ~n3337;
  assign n46212 = pi16 ? n46205 : n46211;
  assign n46213 = pi15 ? n46212 : n32;
  assign n46214 = pi14 ? n46204 : n46213;
  assign n46215 = pi13 ? n46190 : n46214;
  assign n46216 = pi12 ? n46175 : n46215;
  assign n46217 = pi11 ? n46164 : n46216;
  assign n46218 = pi10 ? n46153 : n46217;
  assign n46219 = pi09 ? n32 : n46218;
  assign n46220 = pi14 ? n21686 : n23466;
  assign n46221 = pi19 ? n41566 : ~n32;
  assign n46222 = pi18 ? n32 : n46221;
  assign n46223 = pi17 ? n45886 : ~n46222;
  assign n46224 = pi16 ? n32 : n46223;
  assign n46225 = pi15 ? n45888 : n46224;
  assign n46226 = pi14 ? n32 : n46225;
  assign n46227 = pi13 ? n46220 : n46226;
  assign n46228 = pi17 ? n46094 : ~n2748;
  assign n46229 = pi16 ? n32 : n46228;
  assign n46230 = pi18 ? n21316 : n2747;
  assign n46231 = pi17 ? n46098 : ~n46230;
  assign n46232 = pi16 ? n32 : n46231;
  assign n46233 = pi15 ? n46229 : n46232;
  assign n46234 = pi18 ? n46110 : n2747;
  assign n46235 = pi17 ? n46108 : ~n46234;
  assign n46236 = pi16 ? n46105 : n46235;
  assign n46237 = pi18 ? n9008 : ~n520;
  assign n46238 = pi17 ? n46116 : n46237;
  assign n46239 = pi16 ? n32 : n46238;
  assign n46240 = pi15 ? n46236 : n46239;
  assign n46241 = pi14 ? n46233 : n46240;
  assign n46242 = pi14 ? n46125 : n32822;
  assign n46243 = pi13 ? n46241 : n46242;
  assign n46244 = pi12 ? n46227 : n46243;
  assign n46245 = pi16 ? n32 : n529;
  assign n46246 = pi15 ? n32828 : n46245;
  assign n46247 = pi15 ? n32468 : n12079;
  assign n46248 = pi14 ? n46246 : n46247;
  assign n46249 = pi21 ? n2076 : n140;
  assign n46250 = pi20 ? n206 : ~n46249;
  assign n46251 = pi19 ? n46250 : n32;
  assign n46252 = pi18 ? n9029 : n46251;
  assign n46253 = pi17 ? n32 : n46252;
  assign n46254 = pi16 ? n32 : n46253;
  assign n46255 = pi15 ? n46142 : n46254;
  assign n46256 = pi14 ? n46139 : n46255;
  assign n46257 = pi13 ? n46248 : n46256;
  assign n46258 = pi20 ? n342 : ~n7013;
  assign n46259 = pi19 ? n46258 : n32;
  assign n46260 = pi18 ? n32 : n46259;
  assign n46261 = pi17 ? n32 : n46260;
  assign n46262 = pi16 ? n32 : n46261;
  assign n46263 = pi15 ? n46262 : n32685;
  assign n46264 = pi14 ? n46263 : n32687;
  assign n46265 = pi13 ? n46264 : n32;
  assign n46266 = pi12 ? n46257 : n46265;
  assign n46267 = pi11 ? n46244 : n46266;
  assign n46268 = pi19 ? n12947 : ~n32;
  assign n46269 = pi18 ? n15227 : n46268;
  assign n46270 = pi17 ? n32 : n46269;
  assign n46271 = pi16 ? n1135 : ~n46270;
  assign n46272 = pi15 ? n32 : n46271;
  assign n46273 = pi14 ? n32 : n46272;
  assign n46274 = pi16 ? n1135 : ~n46159;
  assign n46275 = pi15 ? n46274 : n32741;
  assign n46276 = pi14 ? n46275 : n32864;
  assign n46277 = pi13 ? n46273 : n46276;
  assign n46278 = pi12 ? n32 : n46277;
  assign n46279 = pi14 ? n46168 : n45969;
  assign n46280 = pi14 ? n45969 : n46173;
  assign n46281 = pi13 ? n46279 : n46280;
  assign n46282 = pi19 ? n29033 : n17641;
  assign n46283 = pi18 ? n1613 : n46282;
  assign n46284 = pi17 ? n32 : n46283;
  assign n46285 = pi18 ? n39110 : ~n46196;
  assign n46286 = pi17 ? n46285 : ~n32801;
  assign n46287 = pi16 ? n46284 : n46286;
  assign n46288 = pi15 ? n46287 : n46203;
  assign n46289 = pi18 ? n127 : n30574;
  assign n46290 = pi17 ? n32 : n46289;
  assign n46291 = pi17 ? n46210 : ~n1807;
  assign n46292 = pi16 ? n46290 : n46291;
  assign n46293 = pi15 ? n46292 : n130;
  assign n46294 = pi14 ? n46288 : n46293;
  assign n46295 = pi13 ? n46190 : n46294;
  assign n46296 = pi12 ? n46281 : n46295;
  assign n46297 = pi11 ? n46278 : n46296;
  assign n46298 = pi10 ? n46267 : n46297;
  assign n46299 = pi09 ? n32 : n46298;
  assign n46300 = pi08 ? n46219 : n46299;
  assign n46301 = pi07 ? n46084 : n46300;
  assign n46302 = pi14 ? n21853 : n21790;
  assign n46303 = pi15 ? n6215 : n34765;
  assign n46304 = pi14 ? n32 : n46303;
  assign n46305 = pi13 ? n46302 : n46304;
  assign n46306 = pi17 ? n2119 : ~n2748;
  assign n46307 = pi16 ? n32 : n46306;
  assign n46308 = pi18 ? n6163 : n2747;
  assign n46309 = pi17 ? n2750 : ~n46308;
  assign n46310 = pi16 ? n32 : n46309;
  assign n46311 = pi15 ? n46307 : n46310;
  assign n46312 = pi18 ? n684 : ~n2747;
  assign n46313 = pi17 ? n16390 : n46312;
  assign n46314 = pi16 ? n32 : n46313;
  assign n46315 = pi15 ? n46314 : n12289;
  assign n46316 = pi14 ? n46311 : n46315;
  assign n46317 = pi14 ? n32882 : n32885;
  assign n46318 = pi13 ? n46316 : n46317;
  assign n46319 = pi12 ? n46305 : n46318;
  assign n46320 = pi18 ? n209 : ~n520;
  assign n46321 = pi17 ? n32 : n46320;
  assign n46322 = pi16 ? n32 : n46321;
  assign n46323 = pi19 ? n38388 : n32;
  assign n46324 = pi18 ? n940 : n46323;
  assign n46325 = pi17 ? n32 : n46324;
  assign n46326 = pi16 ? n32 : n46325;
  assign n46327 = pi15 ? n46322 : n46326;
  assign n46328 = pi14 ? n12289 : n46327;
  assign n46329 = pi18 ? n32 : n46323;
  assign n46330 = pi17 ? n32 : n46329;
  assign n46331 = pi16 ? n32 : n46330;
  assign n46332 = pi15 ? n14152 : n21543;
  assign n46333 = pi14 ? n46331 : n46332;
  assign n46334 = pi13 ? n46328 : n46333;
  assign n46335 = pi13 ? n32900 : n32;
  assign n46336 = pi12 ? n46334 : n46335;
  assign n46337 = pi11 ? n46319 : n46336;
  assign n46338 = pi13 ? n21132 : n32;
  assign n46339 = pi18 ? n29802 : ~n32;
  assign n46340 = pi17 ? n32 : n46339;
  assign n46341 = pi16 ? n1471 : ~n46340;
  assign n46342 = pi18 ? n21888 : n532;
  assign n46343 = pi17 ? n32 : n46342;
  assign n46344 = pi16 ? n1233 : ~n46343;
  assign n46345 = pi15 ? n46341 : n46344;
  assign n46346 = pi14 ? n32 : n46345;
  assign n46347 = pi18 ? n21595 : ~n32;
  assign n46348 = pi17 ? n14392 : n46347;
  assign n46349 = pi16 ? n1135 : ~n46348;
  assign n46350 = pi15 ? n32937 : n46349;
  assign n46351 = pi14 ? n32935 : n46350;
  assign n46352 = pi13 ? n46346 : n46351;
  assign n46353 = pi12 ? n46338 : n46352;
  assign n46354 = pi16 ? n1233 : ~n2530;
  assign n46355 = pi20 ? n448 : n18253;
  assign n46356 = pi19 ? n46355 : n32;
  assign n46357 = pi18 ? n366 : ~n46356;
  assign n46358 = pi17 ? n32 : n46357;
  assign n46359 = pi20 ? n1091 : n406;
  assign n46360 = pi19 ? n1091 : n46359;
  assign n46361 = pi20 ? n14286 : n175;
  assign n46362 = pi19 ? n32633 : ~n46361;
  assign n46363 = pi18 ? n46360 : ~n46362;
  assign n46364 = pi17 ? n46363 : n2410;
  assign n46365 = pi16 ? n46358 : ~n46364;
  assign n46366 = pi15 ? n46354 : n46365;
  assign n46367 = pi14 ? n35162 : n46366;
  assign n46368 = pi18 ? n1395 : ~n6867;
  assign n46369 = pi17 ? n32 : n46368;
  assign n46370 = pi16 ? n46369 : ~n2530;
  assign n46371 = pi19 ? n15527 : n32;
  assign n46372 = pi18 ? n1395 : ~n46371;
  assign n46373 = pi17 ? n32 : n46372;
  assign n46374 = pi16 ? n46373 : ~n2530;
  assign n46375 = pi15 ? n46370 : n46374;
  assign n46376 = pi19 ? n4964 : ~n321;
  assign n46377 = pi18 ? n16847 : ~n46376;
  assign n46378 = pi17 ? n46377 : ~n2299;
  assign n46379 = pi16 ? n16849 : n46378;
  assign n46380 = pi15 ? n46379 : n44087;
  assign n46381 = pi14 ? n46375 : n46380;
  assign n46382 = pi13 ? n46367 : n46381;
  assign n46383 = pi18 ? n32 : n4519;
  assign n46384 = pi17 ? n32 : n46383;
  assign n46385 = pi17 ? n17119 : ~n32971;
  assign n46386 = pi16 ? n46384 : n46385;
  assign n46387 = pi15 ? n46386 : n32976;
  assign n46388 = pi19 ? n507 : ~n34031;
  assign n46389 = pi18 ? n940 : n46388;
  assign n46390 = pi17 ? n32 : n46389;
  assign n46391 = pi19 ? n321 : n18728;
  assign n46392 = pi19 ? n29186 : n16002;
  assign n46393 = pi18 ? n46391 : ~n46392;
  assign n46394 = pi17 ? n46393 : n1933;
  assign n46395 = pi16 ? n46390 : ~n46394;
  assign n46396 = pi15 ? n32980 : n46395;
  assign n46397 = pi14 ? n46387 : n46396;
  assign n46398 = pi18 ? n209 : ~n5747;
  assign n46399 = pi17 ? n32 : n46398;
  assign n46400 = pi19 ? n321 : n32;
  assign n46401 = pi18 ? n46400 : n32;
  assign n46402 = pi17 ? n46401 : n2537;
  assign n46403 = pi16 ? n46399 : ~n46402;
  assign n46404 = pi19 ? n5694 : n5707;
  assign n46405 = pi18 ? n880 : ~n46404;
  assign n46406 = pi18 ? n940 : n289;
  assign n46407 = pi17 ? n46405 : ~n46406;
  assign n46408 = pi16 ? n3165 : n46407;
  assign n46409 = pi15 ? n46403 : n46408;
  assign n46410 = pi14 ? n46409 : n130;
  assign n46411 = pi13 ? n46397 : n46410;
  assign n46412 = pi12 ? n46382 : n46411;
  assign n46413 = pi11 ? n46353 : n46412;
  assign n46414 = pi10 ? n46337 : n46413;
  assign n46415 = pi09 ? n32 : n46414;
  assign n46416 = pi15 ? n6215 : n34982;
  assign n46417 = pi14 ? n32 : n46416;
  assign n46418 = pi13 ? n46302 : n46417;
  assign n46419 = pi17 ? n2119 : ~n2512;
  assign n46420 = pi16 ? n32 : n46419;
  assign n46421 = pi18 ? n6163 : n508;
  assign n46422 = pi17 ? n2750 : ~n46421;
  assign n46423 = pi16 ? n32 : n46422;
  assign n46424 = pi15 ? n46420 : n46423;
  assign n46425 = pi18 ? n684 : ~n508;
  assign n46426 = pi17 ? n16390 : n46425;
  assign n46427 = pi16 ? n32 : n46426;
  assign n46428 = pi15 ? n46427 : n12289;
  assign n46429 = pi14 ? n46424 : n46428;
  assign n46430 = pi14 ? n33013 : n32885;
  assign n46431 = pi13 ? n46429 : n46430;
  assign n46432 = pi12 ? n46418 : n46431;
  assign n46433 = pi13 ? n33022 : n32;
  assign n46434 = pi12 ? n46334 : n46433;
  assign n46435 = pi11 ? n46432 : n46434;
  assign n46436 = pi16 ? n1135 : ~n46343;
  assign n46437 = pi15 ? n46341 : n46436;
  assign n46438 = pi14 ? n32 : n46437;
  assign n46439 = pi13 ? n46438 : n46351;
  assign n46440 = pi12 ? n32 : n46439;
  assign n46441 = pi16 ? n1135 : ~n2654;
  assign n46442 = pi15 ? n46441 : n35162;
  assign n46443 = pi20 ? n501 : n1331;
  assign n46444 = pi19 ? n46443 : ~n333;
  assign n46445 = pi18 ? n42338 : n46444;
  assign n46446 = pi17 ? n32 : n46445;
  assign n46447 = pi20 ? n2385 : n7839;
  assign n46448 = pi19 ? n2385 : n46447;
  assign n46449 = pi20 ? n1385 : n342;
  assign n46450 = pi19 ? n19191 : ~n46449;
  assign n46451 = pi18 ? n46448 : n46450;
  assign n46452 = pi20 ? n333 : ~n339;
  assign n46453 = pi19 ? n46452 : n32;
  assign n46454 = pi18 ? n46453 : n2298;
  assign n46455 = pi17 ? n46451 : ~n46454;
  assign n46456 = pi16 ? n46446 : n46455;
  assign n46457 = pi15 ? n31828 : n46456;
  assign n46458 = pi14 ? n46442 : n46457;
  assign n46459 = pi18 ? n209 : ~n6867;
  assign n46460 = pi17 ? n32 : n46459;
  assign n46461 = pi16 ? n46460 : ~n2300;
  assign n46462 = pi18 ? n209 : ~n46371;
  assign n46463 = pi17 ? n32 : n46462;
  assign n46464 = pi16 ? n46463 : ~n2300;
  assign n46465 = pi15 ? n46461 : n46464;
  assign n46466 = pi14 ? n46465 : n46380;
  assign n46467 = pi13 ? n46458 : n46466;
  assign n46468 = pi19 ? n29002 : n13939;
  assign n46469 = pi18 ? n858 : n46468;
  assign n46470 = pi17 ? n46469 : ~n32971;
  assign n46471 = pi16 ? n46384 : n46470;
  assign n46472 = pi15 ? n46471 : n33060;
  assign n46473 = pi15 ? n33064 : n46395;
  assign n46474 = pi14 ? n46472 : n46473;
  assign n46475 = pi17 ? n46401 : n1933;
  assign n46476 = pi16 ? n46399 : ~n46475;
  assign n46477 = pi18 ? n940 : n20267;
  assign n46478 = pi17 ? n46405 : ~n46477;
  assign n46479 = pi16 ? n3165 : n46478;
  assign n46480 = pi15 ? n46476 : n46479;
  assign n46481 = pi14 ? n46480 : n32;
  assign n46482 = pi13 ? n46474 : n46481;
  assign n46483 = pi12 ? n46467 : n46482;
  assign n46484 = pi11 ? n46440 : n46483;
  assign n46485 = pi10 ? n46435 : n46484;
  assign n46486 = pi09 ? n32 : n46485;
  assign n46487 = pi08 ? n46415 : n46486;
  assign n46488 = pi14 ? n14790 : n22133;
  assign n46489 = pi13 ? n46488 : n46417;
  assign n46490 = pi19 ? n32 : n6308;
  assign n46491 = pi18 ? n46490 : ~n13070;
  assign n46492 = pi17 ? n46491 : ~n2512;
  assign n46493 = pi16 ? n32 : n46492;
  assign n46494 = pi18 ? n23504 : n508;
  assign n46495 = pi17 ? n2750 : ~n46494;
  assign n46496 = pi16 ? n32 : n46495;
  assign n46497 = pi15 ? n46493 : n46496;
  assign n46498 = pi15 ? n46427 : n12283;
  assign n46499 = pi14 ? n46497 : n46498;
  assign n46500 = pi20 ? n207 : ~n17712;
  assign n46501 = pi19 ? n46500 : ~n32;
  assign n46502 = pi18 ? n32 : ~n46501;
  assign n46503 = pi17 ? n32 : n46502;
  assign n46504 = pi16 ? n32 : n46503;
  assign n46505 = pi15 ? n46504 : n12283;
  assign n46506 = pi14 ? n46505 : n12515;
  assign n46507 = pi13 ? n46499 : n46506;
  assign n46508 = pi12 ? n46489 : n46507;
  assign n46509 = pi20 ? n206 : ~n1319;
  assign n46510 = pi19 ? n46509 : n32;
  assign n46511 = pi18 ? n940 : n46510;
  assign n46512 = pi17 ? n32 : n46511;
  assign n46513 = pi16 ? n32 : n46512;
  assign n46514 = pi15 ? n12518 : n46513;
  assign n46515 = pi14 ? n12518 : n46514;
  assign n46516 = pi18 ? n32 : n46510;
  assign n46517 = pi17 ? n32 : n46516;
  assign n46518 = pi16 ? n32 : n46517;
  assign n46519 = pi15 ? n46518 : n35776;
  assign n46520 = pi15 ? n22469 : n22006;
  assign n46521 = pi14 ? n46519 : n46520;
  assign n46522 = pi13 ? n46515 : n46521;
  assign n46523 = pi13 ? n33089 : n32;
  assign n46524 = pi12 ? n46522 : n46523;
  assign n46525 = pi11 ? n46508 : n46524;
  assign n46526 = pi14 ? n20661 : n32;
  assign n46527 = pi13 ? n32 : n46526;
  assign n46528 = pi18 ? n29802 : ~n13945;
  assign n46529 = pi17 ? n32 : n46528;
  assign n46530 = pi16 ? n1471 : ~n46529;
  assign n46531 = pi18 ? n21888 : ~n13080;
  assign n46532 = pi17 ? n32 : n46531;
  assign n46533 = pi16 ? n1214 : ~n46532;
  assign n46534 = pi15 ? n46530 : n46533;
  assign n46535 = pi14 ? n32 : n46534;
  assign n46536 = pi20 ? n1324 : n342;
  assign n46537 = pi19 ? n32 : n46536;
  assign n46538 = pi18 ? n46537 : n418;
  assign n46539 = pi17 ? n22823 : n46538;
  assign n46540 = pi16 ? n1214 : ~n46539;
  assign n46541 = pi15 ? n33114 : n46540;
  assign n46542 = pi14 ? n33112 : n46541;
  assign n46543 = pi13 ? n46535 : n46542;
  assign n46544 = pi12 ? n46527 : n46543;
  assign n46545 = pi18 ? n4380 : n41276;
  assign n46546 = pi17 ? n32 : n46545;
  assign n46547 = pi19 ? n246 : n247;
  assign n46548 = pi19 ? n221 : n4670;
  assign n46549 = pi18 ? n46547 : n46548;
  assign n46550 = pi17 ? n46549 : n2531;
  assign n46551 = pi16 ? n46546 : ~n46550;
  assign n46552 = pi15 ? n35162 : n46551;
  assign n46553 = pi14 ? n46442 : n46552;
  assign n46554 = pi18 ? n341 : ~n4671;
  assign n46555 = pi17 ? n32 : n46554;
  assign n46556 = pi16 ? n46555 : ~n3625;
  assign n46557 = pi15 ? n35162 : n46556;
  assign n46558 = pi17 ? n46377 : ~n2531;
  assign n46559 = pi16 ? n16849 : n46558;
  assign n46560 = pi18 ? n350 : ~n532;
  assign n46561 = pi17 ? n32 : n46560;
  assign n46562 = pi16 ? n32 : n46561;
  assign n46563 = pi15 ? n46559 : n46562;
  assign n46564 = pi14 ? n46557 : n46563;
  assign n46565 = pi13 ? n46553 : n46564;
  assign n46566 = pi19 ? n5707 : n5371;
  assign n46567 = pi18 ? n341 : n46566;
  assign n46568 = pi17 ? n32 : n46567;
  assign n46569 = pi19 ? n342 : n4670;
  assign n46570 = pi18 ? n46569 : n29440;
  assign n46571 = pi17 ? n46570 : n1933;
  assign n46572 = pi16 ? n46568 : ~n46571;
  assign n46573 = pi15 ? n46572 : n33158;
  assign n46574 = pi19 ? n32 : n29790;
  assign n46575 = pi20 ? n357 : n2358;
  assign n46576 = pi19 ? n32 : n46575;
  assign n46577 = pi18 ? n46574 : n46576;
  assign n46578 = pi17 ? n32 : n46577;
  assign n46579 = pi19 ? n32336 : ~n11531;
  assign n46580 = pi20 ? n266 : ~n749;
  assign n46581 = pi19 ? n46580 : n17766;
  assign n46582 = pi18 ? n46579 : n46581;
  assign n46583 = pi17 ? n46582 : n1933;
  assign n46584 = pi16 ? n46578 : ~n46583;
  assign n46585 = pi15 ? n33158 : n46584;
  assign n46586 = pi14 ? n46573 : n46585;
  assign n46587 = pi18 ? n341 : ~n6669;
  assign n46588 = pi17 ? n32 : n46587;
  assign n46589 = pi16 ? n46588 : ~n46475;
  assign n46590 = pi19 ? n4982 : n4342;
  assign n46591 = pi18 ? n11884 : n46590;
  assign n46592 = pi18 ? n1592 : ~n19232;
  assign n46593 = pi17 ? n46591 : n46592;
  assign n46594 = pi16 ? n3165 : ~n46593;
  assign n46595 = pi15 ? n46589 : n46594;
  assign n46596 = pi14 ? n46595 : n130;
  assign n46597 = pi13 ? n46586 : n46596;
  assign n46598 = pi12 ? n46565 : n46597;
  assign n46599 = pi11 ? n46544 : n46598;
  assign n46600 = pi10 ? n46525 : n46599;
  assign n46601 = pi09 ? n32 : n46600;
  assign n46602 = pi14 ? n14790 : n476;
  assign n46603 = pi19 ? n27488 : ~n32;
  assign n46604 = pi18 ? n32 : n46603;
  assign n46605 = pi17 ? n1215 : ~n46604;
  assign n46606 = pi16 ? n32 : n46605;
  assign n46607 = pi17 ? n1215 : ~n2628;
  assign n46608 = pi16 ? n32 : n46607;
  assign n46609 = pi15 ? n46606 : n46608;
  assign n46610 = pi14 ? n32 : n46609;
  assign n46611 = pi13 ? n46602 : n46610;
  assign n46612 = pi17 ? n46491 : ~n2628;
  assign n46613 = pi16 ? n32 : n46612;
  assign n46614 = pi18 ? n23504 : n2627;
  assign n46615 = pi17 ? n2750 : ~n46614;
  assign n46616 = pi16 ? n32 : n46615;
  assign n46617 = pi15 ? n46613 : n46616;
  assign n46618 = pi18 ? n684 : ~n2627;
  assign n46619 = pi17 ? n16390 : n46618;
  assign n46620 = pi16 ? n32 : n46619;
  assign n46621 = pi18 ? n880 : ~n2627;
  assign n46622 = pi17 ? n32 : n46621;
  assign n46623 = pi16 ? n32 : n46622;
  assign n46624 = pi15 ? n46620 : n46623;
  assign n46625 = pi14 ? n46617 : n46624;
  assign n46626 = pi18 ? n32 : ~n37675;
  assign n46627 = pi17 ? n32 : n46626;
  assign n46628 = pi16 ? n32 : n46627;
  assign n46629 = pi15 ? n46628 : n12283;
  assign n46630 = pi14 ? n46629 : n12515;
  assign n46631 = pi13 ? n46625 : n46630;
  assign n46632 = pi12 ? n46611 : n46631;
  assign n46633 = pi15 ? n12518 : n46326;
  assign n46634 = pi14 ? n12518 : n46633;
  assign n46635 = pi13 ? n46634 : n46521;
  assign n46636 = pi12 ? n46635 : n46523;
  assign n46637 = pi11 ? n46632 : n46636;
  assign n46638 = pi18 ? n29802 : ~n21229;
  assign n46639 = pi17 ? n32 : n46638;
  assign n46640 = pi16 ? n1471 : ~n46639;
  assign n46641 = pi20 ? n207 : n52;
  assign n46642 = pi19 ? n46641 : n32;
  assign n46643 = pi18 ? n21888 : ~n46642;
  assign n46644 = pi17 ? n32 : n46643;
  assign n46645 = pi16 ? n1214 : ~n46644;
  assign n46646 = pi15 ? n46640 : n46645;
  assign n46647 = pi14 ? n32 : n46646;
  assign n46648 = pi18 ? n46537 : n2413;
  assign n46649 = pi17 ? n22823 : n46648;
  assign n46650 = pi16 ? n19652 : ~n46649;
  assign n46651 = pi15 ? n33207 : n46650;
  assign n46652 = pi14 ? n33205 : n46651;
  assign n46653 = pi13 ? n46647 : n46652;
  assign n46654 = pi12 ? n46527 : n46653;
  assign n46655 = pi16 ? n1233 : ~n2654;
  assign n46656 = pi14 ? n46655 : n46552;
  assign n46657 = pi13 ? n46656 : n46564;
  assign n46658 = pi18 ? n11884 : n46581;
  assign n46659 = pi19 ? n32 : n29002;
  assign n46660 = pi18 ? n46659 : n43756;
  assign n46661 = pi17 ? n46658 : n46660;
  assign n46662 = pi16 ? n33161 : ~n46661;
  assign n46663 = pi15 ? n33158 : n46662;
  assign n46664 = pi14 ? n46573 : n46663;
  assign n46665 = pi14 ? n46595 : n32;
  assign n46666 = pi13 ? n46664 : n46665;
  assign n46667 = pi12 ? n46657 : n46666;
  assign n46668 = pi11 ? n46654 : n46667;
  assign n46669 = pi10 ? n46637 : n46668;
  assign n46670 = pi09 ? n32 : n46669;
  assign n46671 = pi08 ? n46601 : n46670;
  assign n46672 = pi07 ? n46487 : n46671;
  assign n46673 = pi06 ? n46301 : n46672;
  assign n46674 = pi14 ? n15123 : n648;
  assign n46675 = pi16 ? n3061 : ~n2629;
  assign n46676 = pi17 ? n1219 : ~n2628;
  assign n46677 = pi16 ? n32 : n46676;
  assign n46678 = pi15 ? n46675 : n46677;
  assign n46679 = pi14 ? n32 : n46678;
  assign n46680 = pi13 ? n46674 : n46679;
  assign n46681 = pi18 ? n9012 : n2627;
  assign n46682 = pi17 ? n2512 : ~n46681;
  assign n46683 = pi16 ? n32 : n46682;
  assign n46684 = pi19 ? n5694 : n3692;
  assign n46685 = pi18 ? n46684 : n2627;
  assign n46686 = pi17 ? n2959 : ~n46685;
  assign n46687 = pi16 ? n32 : n46686;
  assign n46688 = pi15 ? n46683 : n46687;
  assign n46689 = pi19 ? n1844 : n322;
  assign n46690 = pi18 ? n46689 : ~n2627;
  assign n46691 = pi17 ? n17346 : n46690;
  assign n46692 = pi16 ? n32 : n46691;
  assign n46693 = pi19 ? n18464 : ~n32;
  assign n46694 = pi18 ? n940 : ~n46693;
  assign n46695 = pi17 ? n32 : n46694;
  assign n46696 = pi16 ? n32 : n46695;
  assign n46697 = pi15 ? n46692 : n46696;
  assign n46698 = pi14 ? n46688 : n46697;
  assign n46699 = pi15 ? n22650 : n12515;
  assign n46700 = pi15 ? n37814 : n33246;
  assign n46701 = pi14 ? n46699 : n46700;
  assign n46702 = pi13 ? n46698 : n46701;
  assign n46703 = pi12 ? n46680 : n46702;
  assign n46704 = pi19 ? n18678 : ~n32;
  assign n46705 = pi18 ? n940 : ~n46704;
  assign n46706 = pi17 ? n32 : n46705;
  assign n46707 = pi16 ? n32 : n46706;
  assign n46708 = pi15 ? n33253 : n46707;
  assign n46709 = pi19 ? n45905 : n32;
  assign n46710 = pi18 ? n32 : n46709;
  assign n46711 = pi17 ? n32 : n46710;
  assign n46712 = pi16 ? n32 : n46711;
  assign n46713 = pi18 ? n863 : n5357;
  assign n46714 = pi17 ? n32 : n46713;
  assign n46715 = pi16 ? n32 : n46714;
  assign n46716 = pi15 ? n46712 : n46715;
  assign n46717 = pi14 ? n46708 : n46716;
  assign n46718 = pi18 ? n940 : n33508;
  assign n46719 = pi17 ? n32 : n46718;
  assign n46720 = pi16 ? n32 : n46719;
  assign n46721 = pi18 ? n209 : n24195;
  assign n46722 = pi17 ? n32 : n46721;
  assign n46723 = pi16 ? n32 : n46722;
  assign n46724 = pi15 ? n46720 : n46723;
  assign n46725 = pi19 ? n37871 : n32;
  assign n46726 = pi18 ? n32 : n46725;
  assign n46727 = pi17 ? n32 : n46726;
  assign n46728 = pi16 ? n32 : n46727;
  assign n46729 = pi15 ? n14147 : n46728;
  assign n46730 = pi14 ? n46724 : n46729;
  assign n46731 = pi13 ? n46717 : n46730;
  assign n46732 = pi15 ? n14394 : n21543;
  assign n46733 = pi14 ? n46732 : n32;
  assign n46734 = pi13 ? n46733 : n32;
  assign n46735 = pi12 ? n46731 : n46734;
  assign n46736 = pi11 ? n46703 : n46735;
  assign n46737 = pi14 ? n21467 : n32;
  assign n46738 = pi13 ? n46737 : n32;
  assign n46739 = pi19 ? n322 : n5694;
  assign n46740 = pi18 ? n32 : n46739;
  assign n46741 = pi17 ? n46740 : n1480;
  assign n46742 = pi16 ? n1471 : ~n46741;
  assign n46743 = pi18 ? n15844 : n33304;
  assign n46744 = pi17 ? n32 : n46743;
  assign n46745 = pi16 ? n1233 : ~n46744;
  assign n46746 = pi18 ? n496 : ~n13945;
  assign n46747 = pi17 ? n32 : n46746;
  assign n46748 = pi16 ? n1471 : ~n46747;
  assign n46749 = pi15 ? n46745 : n46748;
  assign n46750 = pi14 ? n46742 : n46749;
  assign n46751 = pi17 ? n23931 : n2414;
  assign n46752 = pi16 ? n1214 : ~n46751;
  assign n46753 = pi15 ? n33320 : n46752;
  assign n46754 = pi14 ? n33317 : n46753;
  assign n46755 = pi13 ? n46750 : n46754;
  assign n46756 = pi12 ? n46738 : n46755;
  assign n46757 = pi19 ? n594 : ~n45479;
  assign n46758 = pi18 ? n341 : ~n46757;
  assign n46759 = pi17 ? n32 : n46758;
  assign n46760 = pi20 ? n428 : ~n18245;
  assign n46761 = pi19 ? n46760 : ~n18245;
  assign n46762 = pi20 ? n18540 : ~n175;
  assign n46763 = pi20 ? n207 : ~n9863;
  assign n46764 = pi19 ? n46762 : n46763;
  assign n46765 = pi18 ? n46761 : ~n46764;
  assign n46766 = pi18 ? n19232 : n532;
  assign n46767 = pi17 ? n46765 : n46766;
  assign n46768 = pi16 ? n46759 : ~n46767;
  assign n46769 = pi18 ? n341 : ~n13975;
  assign n46770 = pi17 ? n32 : n46769;
  assign n46771 = pi16 ? n46770 : ~n3625;
  assign n46772 = pi15 ? n46768 : n46771;
  assign n46773 = pi14 ? n35162 : n46772;
  assign n46774 = pi16 ? n1135 : ~n3788;
  assign n46775 = pi18 ? n8966 : ~n3786;
  assign n46776 = pi17 ? n14154 : n46775;
  assign n46777 = pi16 ? n32 : n46776;
  assign n46778 = pi18 ? n248 : n14153;
  assign n46779 = pi18 ? n13080 : n532;
  assign n46780 = pi17 ? n46778 : ~n46779;
  assign n46781 = pi16 ? n32 : n46780;
  assign n46782 = pi15 ? n46777 : n46781;
  assign n46783 = pi14 ? n46774 : n46782;
  assign n46784 = pi13 ? n46773 : n46783;
  assign n46785 = pi16 ? n33623 : ~n3625;
  assign n46786 = pi15 ? n46785 : n33358;
  assign n46787 = pi14 ? n46786 : n33365;
  assign n46788 = pi19 ? n321 : ~n208;
  assign n46789 = pi18 ? n222 : ~n46788;
  assign n46790 = pi17 ? n32 : n46789;
  assign n46791 = pi16 ? n46790 : n33371;
  assign n46792 = pi17 ? n32 : n17951;
  assign n46793 = pi16 ? n1014 : n46792;
  assign n46794 = pi15 ? n46791 : n46793;
  assign n46795 = pi14 ? n46794 : n130;
  assign n46796 = pi13 ? n46787 : n46795;
  assign n46797 = pi12 ? n46784 : n46796;
  assign n46798 = pi11 ? n46756 : n46797;
  assign n46799 = pi10 ? n46736 : n46798;
  assign n46800 = pi09 ? n32 : n46799;
  assign n46801 = pi14 ? n15123 : n22257;
  assign n46802 = pi16 ? n3061 : ~n3946;
  assign n46803 = pi17 ? n1219 : ~n2618;
  assign n46804 = pi16 ? n32 : n46803;
  assign n46805 = pi15 ? n46802 : n46804;
  assign n46806 = pi14 ? n32 : n46805;
  assign n46807 = pi13 ? n46801 : n46806;
  assign n46808 = pi18 ? n9012 : n595;
  assign n46809 = pi17 ? n2512 : ~n46808;
  assign n46810 = pi16 ? n32 : n46809;
  assign n46811 = pi18 ? n46684 : n595;
  assign n46812 = pi17 ? n2959 : ~n46811;
  assign n46813 = pi16 ? n32 : n46812;
  assign n46814 = pi15 ? n46810 : n46813;
  assign n46815 = pi18 ? n46689 : ~n595;
  assign n46816 = pi17 ? n17346 : n46815;
  assign n46817 = pi16 ? n32 : n46816;
  assign n46818 = pi15 ? n46817 : n46696;
  assign n46819 = pi14 ? n46814 : n46818;
  assign n46820 = pi15 ? n22749 : n12515;
  assign n46821 = pi18 ? n4127 : ~n2627;
  assign n46822 = pi17 ? n32 : n46821;
  assign n46823 = pi16 ? n32 : n46822;
  assign n46824 = pi15 ? n46823 : n33399;
  assign n46825 = pi14 ? n46820 : n46824;
  assign n46826 = pi13 ? n46819 : n46825;
  assign n46827 = pi12 ? n46807 : n46826;
  assign n46828 = pi15 ? n33246 : n46707;
  assign n46829 = pi14 ? n46828 : n46716;
  assign n46830 = pi21 ? n259 : n242;
  assign n46831 = pi20 ? n32 : ~n46830;
  assign n46832 = pi19 ? n46831 : n32;
  assign n46833 = pi18 ? n32 : n46832;
  assign n46834 = pi17 ? n32 : n46833;
  assign n46835 = pi16 ? n32 : n46834;
  assign n46836 = pi15 ? n14147 : n46835;
  assign n46837 = pi14 ? n46724 : n46836;
  assign n46838 = pi13 ? n46829 : n46837;
  assign n46839 = pi15 ? n14394 : n21686;
  assign n46840 = pi14 ? n46839 : n32;
  assign n46841 = pi13 ? n46840 : n32;
  assign n46842 = pi12 ? n46838 : n46841;
  assign n46843 = pi11 ? n46827 : n46842;
  assign n46844 = pi16 ? n1135 : ~n46744;
  assign n46845 = pi15 ? n46844 : n46748;
  assign n46846 = pi14 ? n46742 : n46845;
  assign n46847 = pi17 ? n23931 : n2119;
  assign n46848 = pi16 ? n1214 : ~n46847;
  assign n46849 = pi15 ? n33320 : n46848;
  assign n46850 = pi14 ? n33317 : n46849;
  assign n46851 = pi13 ? n46846 : n46850;
  assign n46852 = pi12 ? n32 : n46851;
  assign n46853 = pi20 ? n6085 : n1611;
  assign n46854 = pi20 ? n1611 : n314;
  assign n46855 = pi19 ? n46853 : ~n46854;
  assign n46856 = pi18 ? n356 : ~n46855;
  assign n46857 = pi17 ? n32 : n46856;
  assign n46858 = pi20 ? n13171 : n12884;
  assign n46859 = pi19 ? n46858 : n12884;
  assign n46860 = pi20 ? n12882 : ~n342;
  assign n46861 = pi20 ? n207 : ~n1685;
  assign n46862 = pi19 ? n46860 : n46861;
  assign n46863 = pi18 ? n46859 : n46862;
  assign n46864 = pi20 ? n246 : ~n18415;
  assign n46865 = pi19 ? n46864 : n5614;
  assign n46866 = pi18 ? n46865 : n532;
  assign n46867 = pi17 ? n46863 : ~n46866;
  assign n46868 = pi16 ? n46857 : n46867;
  assign n46869 = pi20 ? n357 : ~n32;
  assign n46870 = pi19 ? n46869 : ~n32;
  assign n46871 = pi18 ? n32 : n46870;
  assign n46872 = pi17 ? n32 : n46871;
  assign n46873 = pi16 ? n46770 : ~n46872;
  assign n46874 = pi15 ? n46868 : n46873;
  assign n46875 = pi14 ? n35359 : n46874;
  assign n46876 = pi18 ? n13080 : n3786;
  assign n46877 = pi17 ? n46778 : ~n46876;
  assign n46878 = pi16 ? n32 : n46877;
  assign n46879 = pi15 ? n46777 : n46878;
  assign n46880 = pi14 ? n35162 : n46879;
  assign n46881 = pi13 ? n46875 : n46880;
  assign n46882 = pi16 ? n33354 : ~n3788;
  assign n46883 = pi15 ? n46882 : n33459;
  assign n46884 = pi14 ? n46883 : n33365;
  assign n46885 = pi15 ? n46791 : n1015;
  assign n46886 = pi14 ? n46885 : n131;
  assign n46887 = pi13 ? n46884 : n46886;
  assign n46888 = pi12 ? n46881 : n46887;
  assign n46889 = pi11 ? n46852 : n46888;
  assign n46890 = pi10 ? n46843 : n46889;
  assign n46891 = pi09 ? n32 : n46890;
  assign n46892 = pi08 ? n46800 : n46891;
  assign n46893 = pi14 ? n22347 : n23604;
  assign n46894 = pi16 ? n2958 : ~n3946;
  assign n46895 = pi17 ? n38528 : ~n2618;
  assign n46896 = pi16 ? n32 : n46895;
  assign n46897 = pi15 ? n46894 : n46896;
  assign n46898 = pi14 ? n32 : n46897;
  assign n46899 = pi13 ? n46893 : n46898;
  assign n46900 = pi20 ? n206 : ~n357;
  assign n46901 = pi19 ? n507 : n46900;
  assign n46902 = pi18 ? n32 : n46901;
  assign n46903 = pi19 ? n267 : n16294;
  assign n46904 = pi18 ? n46903 : n595;
  assign n46905 = pi17 ? n46902 : ~n46904;
  assign n46906 = pi16 ? n32 : n46905;
  assign n46907 = pi19 ? n4982 : n3692;
  assign n46908 = pi18 ? n46907 : n595;
  assign n46909 = pi17 ? n4302 : ~n46908;
  assign n46910 = pi16 ? n32 : n46909;
  assign n46911 = pi15 ? n46906 : n46910;
  assign n46912 = pi18 ? n940 : ~n595;
  assign n46913 = pi17 ? n17346 : n46912;
  assign n46914 = pi16 ? n32 : n46913;
  assign n46915 = pi19 ? n18489 : ~n32;
  assign n46916 = pi18 ? n940 : ~n46915;
  assign n46917 = pi17 ? n32 : n46916;
  assign n46918 = pi16 ? n32 : n46917;
  assign n46919 = pi15 ? n46914 : n46918;
  assign n46920 = pi14 ? n46911 : n46919;
  assign n46921 = pi15 ? n22650 : n12764;
  assign n46922 = pi20 ? n785 : n22331;
  assign n46923 = pi19 ? n46922 : n32;
  assign n46924 = pi18 ? n32 : n46923;
  assign n46925 = pi17 ? n32 : n46924;
  assign n46926 = pi16 ? n32 : n46925;
  assign n46927 = pi15 ? n33479 : n46926;
  assign n46928 = pi14 ? n46921 : n46927;
  assign n46929 = pi13 ? n46920 : n46928;
  assign n46930 = pi12 ? n46899 : n46929;
  assign n46931 = pi22 ? n84 : ~n50;
  assign n46932 = pi21 ? n32 : ~n46931;
  assign n46933 = pi20 ? n246 : n46932;
  assign n46934 = pi19 ? n46933 : ~n32;
  assign n46935 = pi18 ? n940 : ~n46934;
  assign n46936 = pi17 ? n32 : n46935;
  assign n46937 = pi16 ? n32 : n46936;
  assign n46938 = pi15 ? n20608 : n46937;
  assign n46939 = pi21 ? n32 : n46931;
  assign n46940 = pi20 ? n321 : ~n46939;
  assign n46941 = pi19 ? n46940 : ~n32;
  assign n46942 = pi18 ? n32 : ~n46941;
  assign n46943 = pi17 ? n32 : n46942;
  assign n46944 = pi16 ? n32 : n46943;
  assign n46945 = pi18 ? n863 : n39697;
  assign n46946 = pi17 ? n32 : n46945;
  assign n46947 = pi16 ? n32 : n46946;
  assign n46948 = pi15 ? n46944 : n46947;
  assign n46949 = pi14 ? n46938 : n46948;
  assign n46950 = pi20 ? n974 : ~n2140;
  assign n46951 = pi19 ? n46950 : n32;
  assign n46952 = pi18 ? n940 : n46951;
  assign n46953 = pi17 ? n32 : n46952;
  assign n46954 = pi16 ? n32 : n46953;
  assign n46955 = pi20 ? n5854 : n2140;
  assign n46956 = pi19 ? n46955 : ~n32;
  assign n46957 = pi18 ? n209 : ~n46956;
  assign n46958 = pi17 ? n32 : n46957;
  assign n46959 = pi16 ? n32 : n46958;
  assign n46960 = pi15 ? n46954 : n46959;
  assign n46961 = pi20 ? n339 : n2140;
  assign n46962 = pi19 ? n46961 : ~n32;
  assign n46963 = pi18 ? n4127 : ~n46962;
  assign n46964 = pi17 ? n32 : n46963;
  assign n46965 = pi16 ? n32 : n46964;
  assign n46966 = pi15 ? n46965 : n33511;
  assign n46967 = pi14 ? n46960 : n46966;
  assign n46968 = pi13 ? n46949 : n46967;
  assign n46969 = pi15 ? n14147 : n32;
  assign n46970 = pi14 ? n46969 : n21319;
  assign n46971 = pi13 ? n46970 : n32;
  assign n46972 = pi12 ? n46968 : n46971;
  assign n46973 = pi11 ? n46930 : n46972;
  assign n46974 = pi18 ? n702 : ~n13940;
  assign n46975 = pi17 ? n46740 : n46974;
  assign n46976 = pi16 ? n1471 : ~n46975;
  assign n46977 = pi15 ? n46742 : n46976;
  assign n46978 = pi18 ? n15844 : n33579;
  assign n46979 = pi17 ? n32 : n46978;
  assign n46980 = pi16 ? n1135 : ~n46979;
  assign n46981 = pi18 ? n496 : ~n13940;
  assign n46982 = pi17 ? n32 : n46981;
  assign n46983 = pi16 ? n1471 : ~n46982;
  assign n46984 = pi15 ? n46980 : n46983;
  assign n46985 = pi14 ? n46977 : n46984;
  assign n46986 = pi17 ? n24698 : n2119;
  assign n46987 = pi16 ? n1135 : ~n46986;
  assign n46988 = pi14 ? n33586 : n46987;
  assign n46989 = pi13 ? n46985 : n46988;
  assign n46990 = pi12 ? n32 : n46989;
  assign n46991 = pi16 ? n1135 : ~n2426;
  assign n46992 = pi15 ? n46991 : n46441;
  assign n46993 = pi19 ? n266 : n1464;
  assign n46994 = pi18 ? n209 : n46993;
  assign n46995 = pi17 ? n32 : n46994;
  assign n46996 = pi19 ? n5371 : ~n266;
  assign n46997 = pi18 ? n46996 : ~n33637;
  assign n46998 = pi17 ? n46997 : ~n2653;
  assign n46999 = pi16 ? n46995 : n46998;
  assign n47000 = pi18 ? n209 : ~n13975;
  assign n47001 = pi17 ? n32 : n47000;
  assign n47002 = pi16 ? n47001 : ~n2654;
  assign n47003 = pi15 ? n46999 : n47002;
  assign n47004 = pi14 ? n46992 : n47003;
  assign n47005 = pi18 ? n8966 : ~n532;
  assign n47006 = pi17 ? n14154 : n47005;
  assign n47007 = pi16 ? n32 : n47006;
  assign n47008 = pi18 ? n4380 : n46993;
  assign n47009 = pi17 ? n32 : n47008;
  assign n47010 = pi19 ? n9822 : n342;
  assign n47011 = pi20 ? n246 : ~n1324;
  assign n47012 = pi19 ? n47011 : n5748;
  assign n47013 = pi18 ? n47010 : n47012;
  assign n47014 = pi18 ? n20611 : n532;
  assign n47015 = pi17 ? n47013 : ~n47014;
  assign n47016 = pi16 ? n47009 : n47015;
  assign n47017 = pi15 ? n47007 : n47016;
  assign n47018 = pi14 ? n46441 : n47017;
  assign n47019 = pi13 ? n47004 : n47018;
  assign n47020 = pi15 ? n46785 : n33627;
  assign n47021 = pi14 ? n47020 : n33634;
  assign n47022 = pi19 ? n266 : n322;
  assign n47023 = pi18 ? n312 : n47022;
  assign n47024 = pi17 ? n32 : n47023;
  assign n47025 = pi20 ? n1817 : n274;
  assign n47026 = pi19 ? n47025 : ~n22525;
  assign n47027 = pi18 ? n46376 : ~n47026;
  assign n47028 = pi20 ? n339 : n207;
  assign n47029 = pi19 ? n47028 : ~n32;
  assign n47030 = pi18 ? n47029 : ~n344;
  assign n47031 = pi17 ? n47027 : n47030;
  assign n47032 = pi16 ? n47024 : n47031;
  assign n47033 = pi15 ? n47032 : n130;
  assign n47034 = pi14 ? n47033 : n130;
  assign n47035 = pi13 ? n47021 : n47034;
  assign n47036 = pi12 ? n47019 : n47035;
  assign n47037 = pi11 ? n46990 : n47036;
  assign n47038 = pi10 ? n46973 : n47037;
  assign n47039 = pi09 ? n32 : n47038;
  assign n47040 = pi14 ? n22347 : n15123;
  assign n47041 = pi16 ? n2958 : ~n4100;
  assign n47042 = pi17 ? n38528 : ~n4099;
  assign n47043 = pi16 ? n32 : n47042;
  assign n47044 = pi15 ? n47041 : n47043;
  assign n47045 = pi14 ? n32 : n47044;
  assign n47046 = pi13 ? n47040 : n47045;
  assign n47047 = pi18 ? n46903 : n4098;
  assign n47048 = pi17 ? n46902 : ~n47047;
  assign n47049 = pi16 ? n32 : n47048;
  assign n47050 = pi18 ? n46907 : n4098;
  assign n47051 = pi17 ? n4302 : ~n47050;
  assign n47052 = pi16 ? n32 : n47051;
  assign n47053 = pi15 ? n47049 : n47052;
  assign n47054 = pi17 ? n17346 : n12754;
  assign n47055 = pi16 ? n32 : n47054;
  assign n47056 = pi15 ? n47055 : n46918;
  assign n47057 = pi14 ? n47053 : n47056;
  assign n47058 = pi20 ? n785 : n21111;
  assign n47059 = pi19 ? n47058 : n32;
  assign n47060 = pi18 ? n32 : n47059;
  assign n47061 = pi17 ? n32 : n47060;
  assign n47062 = pi16 ? n32 : n47061;
  assign n47063 = pi15 ? n33479 : n47062;
  assign n47064 = pi14 ? n46921 : n47063;
  assign n47065 = pi13 ? n47057 : n47064;
  assign n47066 = pi12 ? n47046 : n47065;
  assign n47067 = pi20 ? n246 : n1076;
  assign n47068 = pi19 ? n47067 : ~n32;
  assign n47069 = pi18 ? n940 : ~n47068;
  assign n47070 = pi17 ? n32 : n47069;
  assign n47071 = pi16 ? n32 : n47070;
  assign n47072 = pi15 ? n20608 : n47071;
  assign n47073 = pi20 ? n321 : ~n3523;
  assign n47074 = pi19 ? n47073 : ~n32;
  assign n47075 = pi18 ? n32 : ~n47074;
  assign n47076 = pi17 ? n32 : n47075;
  assign n47077 = pi16 ? n32 : n47076;
  assign n47078 = pi18 ? n863 : n23871;
  assign n47079 = pi17 ? n32 : n47078;
  assign n47080 = pi16 ? n32 : n47079;
  assign n47081 = pi15 ? n47077 : n47080;
  assign n47082 = pi14 ? n47072 : n47081;
  assign n47083 = pi15 ? n46965 : n33678;
  assign n47084 = pi14 ? n46960 : n47083;
  assign n47085 = pi13 ? n47082 : n47084;
  assign n47086 = pi14 ? n46969 : n32;
  assign n47087 = pi13 ? n47086 : n32;
  assign n47088 = pi12 ? n47085 : n47087;
  assign n47089 = pi11 ? n47066 : n47088;
  assign n47090 = pi18 ? n15844 : n33702;
  assign n47091 = pi17 ? n32 : n47090;
  assign n47092 = pi16 ? n1233 : ~n47091;
  assign n47093 = pi15 ? n47092 : n46983;
  assign n47094 = pi14 ? n46977 : n47093;
  assign n47095 = pi17 ? n24698 : n2408;
  assign n47096 = pi16 ? n1135 : ~n47095;
  assign n47097 = pi15 ? n47096 : n46987;
  assign n47098 = pi14 ? n33709 : n47097;
  assign n47099 = pi13 ? n47094 : n47098;
  assign n47100 = pi12 ? n32 : n47099;
  assign n47101 = pi15 ? n36601 : n46655;
  assign n47102 = pi18 ? n1395 : n46993;
  assign n47103 = pi17 ? n32 : n47102;
  assign n47104 = pi16 ? n47103 : n46998;
  assign n47105 = pi18 ? n1395 : ~n13975;
  assign n47106 = pi17 ? n32 : n47105;
  assign n47107 = pi16 ? n47106 : ~n2654;
  assign n47108 = pi15 ? n47104 : n47107;
  assign n47109 = pi14 ? n47101 : n47108;
  assign n47110 = pi15 ? n46655 : n46441;
  assign n47111 = pi14 ? n47110 : n47017;
  assign n47112 = pi13 ? n47109 : n47111;
  assign n47113 = pi16 ? n33354 : ~n3625;
  assign n47114 = pi15 ? n47113 : n33627;
  assign n47115 = pi14 ? n47114 : n33634;
  assign n47116 = pi14 ? n47033 : n131;
  assign n47117 = pi13 ? n47115 : n47116;
  assign n47118 = pi12 ? n47112 : n47117;
  assign n47119 = pi11 ? n47100 : n47118;
  assign n47120 = pi10 ? n47089 : n47119;
  assign n47121 = pi09 ? n32 : n47120;
  assign n47122 = pi08 ? n47039 : n47121;
  assign n47123 = pi07 ? n46892 : n47122;
  assign n47124 = pi15 ? n23443 : n22540;
  assign n47125 = pi14 ? n47124 : n22424;
  assign n47126 = pi18 ? n32 : ~n41055;
  assign n47127 = pi17 ? n35241 : n47126;
  assign n47128 = pi16 ? n32 : n47127;
  assign n47129 = pi15 ? n32 : n47128;
  assign n47130 = pi18 ? n9461 : ~n4343;
  assign n47131 = pi17 ? n47130 : ~n2618;
  assign n47132 = pi16 ? n32 : n47131;
  assign n47133 = pi18 ? n496 : ~n4343;
  assign n47134 = pi17 ? n47133 : ~n2512;
  assign n47135 = pi16 ? n32 : n47134;
  assign n47136 = pi15 ? n47132 : n47135;
  assign n47137 = pi14 ? n47129 : n47136;
  assign n47138 = pi13 ? n47125 : n47137;
  assign n47139 = pi19 ? n32 : n17757;
  assign n47140 = pi18 ? n32 : n47139;
  assign n47141 = pi20 ? n5854 : ~n342;
  assign n47142 = pi20 ? n357 : n321;
  assign n47143 = pi19 ? n47141 : ~n47142;
  assign n47144 = pi19 ? n18982 : ~n32;
  assign n47145 = pi18 ? n47143 : n47144;
  assign n47146 = pi17 ? n47140 : ~n47145;
  assign n47147 = pi16 ? n32 : n47146;
  assign n47148 = pi18 ? n28382 : ~n47144;
  assign n47149 = pi17 ? n3164 : n47148;
  assign n47150 = pi16 ? n32 : n47149;
  assign n47151 = pi15 ? n47147 : n47150;
  assign n47152 = pi17 ? n23052 : n12759;
  assign n47153 = pi16 ? n32 : n47152;
  assign n47154 = pi19 ? n507 : n18396;
  assign n47155 = pi18 ? n32 : n47154;
  assign n47156 = pi19 ? n246 : n4126;
  assign n47157 = pi18 ? n47156 : ~n595;
  assign n47158 = pi17 ? n47155 : n47157;
  assign n47159 = pi16 ? n32 : n47158;
  assign n47160 = pi15 ? n47153 : n47159;
  assign n47161 = pi14 ? n47151 : n47160;
  assign n47162 = pi17 ? n26267 : n46912;
  assign n47163 = pi16 ? n32 : n47162;
  assign n47164 = pi18 ? n880 : ~n595;
  assign n47165 = pi17 ? n17346 : n47164;
  assign n47166 = pi16 ? n32 : n47165;
  assign n47167 = pi15 ? n47163 : n47166;
  assign n47168 = pi18 ? n863 : ~n595;
  assign n47169 = pi17 ? n32 : n47168;
  assign n47170 = pi16 ? n32 : n47169;
  assign n47171 = pi20 ? n220 : ~n3695;
  assign n47172 = pi19 ? n47171 : ~n32;
  assign n47173 = pi18 ? n936 : ~n47172;
  assign n47174 = pi17 ? n32 : n47173;
  assign n47175 = pi16 ? n32 : n47174;
  assign n47176 = pi15 ? n47170 : n47175;
  assign n47177 = pi14 ? n47167 : n47176;
  assign n47178 = pi13 ? n47161 : n47177;
  assign n47179 = pi12 ? n47138 : n47178;
  assign n47180 = pi20 ? n342 : n12884;
  assign n47181 = pi19 ? n47180 : n32;
  assign n47182 = pi18 ? n32 : n47181;
  assign n47183 = pi17 ? n32 : n47182;
  assign n47184 = pi16 ? n32 : n47183;
  assign n47185 = pi15 ? n47184 : n23037;
  assign n47186 = pi17 ? n32 : n46912;
  assign n47187 = pi16 ? n32 : n47186;
  assign n47188 = pi18 ? n32 : n17767;
  assign n47189 = pi18 ? n4392 : ~n34621;
  assign n47190 = pi17 ? n47188 : n47189;
  assign n47191 = pi16 ? n32 : n47190;
  assign n47192 = pi15 ? n47187 : n47191;
  assign n47193 = pi14 ? n47185 : n47192;
  assign n47194 = pi20 ? n3523 : n206;
  assign n47195 = pi19 ? n32 : ~n47194;
  assign n47196 = pi18 ? n20164 : n47195;
  assign n47197 = pi19 ? n5435 : n236;
  assign n47198 = pi18 ? n47197 : ~n595;
  assign n47199 = pi17 ? n47196 : n47198;
  assign n47200 = pi16 ? n32 : n47199;
  assign n47201 = pi19 ? n23489 : ~n32;
  assign n47202 = pi18 ? n880 : ~n47201;
  assign n47203 = pi17 ? n32 : n47202;
  assign n47204 = pi16 ? n32 : n47203;
  assign n47205 = pi15 ? n47200 : n47204;
  assign n47206 = pi20 ? n339 : ~n11107;
  assign n47207 = pi19 ? n47206 : n32;
  assign n47208 = pi18 ? n18710 : n47207;
  assign n47209 = pi17 ? n32 : n47208;
  assign n47210 = pi16 ? n32 : n47209;
  assign n47211 = pi20 ? n518 : ~n206;
  assign n47212 = pi19 ? n47211 : n32;
  assign n47213 = pi18 ? n32 : n47212;
  assign n47214 = pi17 ? n32 : n47213;
  assign n47215 = pi16 ? n32 : n47214;
  assign n47216 = pi15 ? n47210 : n47215;
  assign n47217 = pi14 ? n47205 : n47216;
  assign n47218 = pi13 ? n47193 : n47217;
  assign n47219 = pi14 ? n32 : n21790;
  assign n47220 = pi13 ? n32 : n47219;
  assign n47221 = pi12 ? n47218 : n47220;
  assign n47222 = pi11 ? n47179 : n47221;
  assign n47223 = pi15 ? n21786 : n21543;
  assign n47224 = pi14 ? n47223 : n32;
  assign n47225 = pi13 ? n47224 : n32;
  assign n47226 = pi17 ? n46740 : n1978;
  assign n47227 = pi16 ? n1471 : ~n47226;
  assign n47228 = pi18 ? n880 : ~n13058;
  assign n47229 = pi17 ? n32 : n47228;
  assign n47230 = pi16 ? n1135 : ~n47229;
  assign n47231 = pi15 ? n47227 : n47230;
  assign n47232 = pi18 ? n684 : ~n5164;
  assign n47233 = pi17 ? n32 : n47232;
  assign n47234 = pi16 ? n1135 : ~n47233;
  assign n47235 = pi18 ? n940 : ~n20164;
  assign n47236 = pi17 ? n32 : n47235;
  assign n47237 = pi19 ? n4126 : n4721;
  assign n47238 = pi18 ? n9012 : n47237;
  assign n47239 = pi19 ? n4342 : n1757;
  assign n47240 = pi19 ? n46580 : n32;
  assign n47241 = pi18 ? n47239 : n47240;
  assign n47242 = pi17 ? n47238 : n47241;
  assign n47243 = pi16 ? n47236 : n47242;
  assign n47244 = pi15 ? n47234 : n47243;
  assign n47245 = pi14 ? n47231 : n47244;
  assign n47246 = pi18 ? n1379 : n33824;
  assign n47247 = pi17 ? n32 : n47246;
  assign n47248 = pi16 ? n1233 : ~n47247;
  assign n47249 = pi15 ? n33822 : n47248;
  assign n47250 = pi17 ? n25761 : n2119;
  assign n47251 = pi16 ? n1214 : ~n47250;
  assign n47252 = pi15 ? n33830 : n47251;
  assign n47253 = pi14 ? n47249 : n47252;
  assign n47254 = pi13 ? n47245 : n47253;
  assign n47255 = pi12 ? n47225 : n47254;
  assign n47256 = pi16 ? n1135 : ~n2120;
  assign n47257 = pi18 ? n209 : ~n15849;
  assign n47258 = pi17 ? n32 : n47257;
  assign n47259 = pi16 ? n47258 : ~n2654;
  assign n47260 = pi15 ? n47256 : n47259;
  assign n47261 = pi16 ? n1214 : ~n3625;
  assign n47262 = pi15 ? n47261 : n35162;
  assign n47263 = pi14 ? n47260 : n47262;
  assign n47264 = pi16 ? n1214 : ~n2654;
  assign n47265 = pi15 ? n47264 : n46441;
  assign n47266 = pi14 ? n46441 : n47265;
  assign n47267 = pi13 ? n47263 : n47266;
  assign n47268 = pi15 ? n47261 : n33870;
  assign n47269 = pi19 ? n35996 : ~n32;
  assign n47270 = pi18 ? n222 : ~n47269;
  assign n47271 = pi17 ? n32 : n47270;
  assign n47272 = pi16 ? n47271 : ~n33880;
  assign n47273 = pi15 ? n33135 : n47272;
  assign n47274 = pi14 ? n47268 : n47273;
  assign n47275 = pi15 ? n32 : n130;
  assign n47276 = pi14 ? n47275 : n130;
  assign n47277 = pi13 ? n47274 : n47276;
  assign n47278 = pi12 ? n47267 : n47277;
  assign n47279 = pi11 ? n47255 : n47278;
  assign n47280 = pi10 ? n47222 : n47279;
  assign n47281 = pi09 ? n32 : n47280;
  assign n47282 = pi17 ? n47130 : ~n2750;
  assign n47283 = pi16 ? n32 : n47282;
  assign n47284 = pi17 ? n47133 : ~n2861;
  assign n47285 = pi16 ? n32 : n47284;
  assign n47286 = pi15 ? n47283 : n47285;
  assign n47287 = pi14 ? n47129 : n47286;
  assign n47288 = pi13 ? n47125 : n47287;
  assign n47289 = pi18 ? n47143 : n2684;
  assign n47290 = pi17 ? n47140 : ~n47289;
  assign n47291 = pi16 ? n32 : n47290;
  assign n47292 = pi18 ? n28382 : ~n2684;
  assign n47293 = pi17 ? n3164 : n47292;
  assign n47294 = pi16 ? n32 : n47293;
  assign n47295 = pi15 ? n47291 : n47294;
  assign n47296 = pi18 ? n863 : ~n702;
  assign n47297 = pi17 ? n23052 : n47296;
  assign n47298 = pi16 ? n32 : n47297;
  assign n47299 = pi15 ? n47298 : n47159;
  assign n47300 = pi14 ? n47295 : n47299;
  assign n47301 = pi21 ? n309 : ~n100;
  assign n47302 = pi20 ? n220 : ~n47301;
  assign n47303 = pi19 ? n47302 : ~n32;
  assign n47304 = pi18 ? n936 : ~n47303;
  assign n47305 = pi17 ? n32 : n47304;
  assign n47306 = pi16 ? n32 : n47305;
  assign n47307 = pi15 ? n47170 : n47306;
  assign n47308 = pi14 ? n47167 : n47307;
  assign n47309 = pi13 ? n47300 : n47308;
  assign n47310 = pi12 ? n47288 : n47309;
  assign n47311 = pi20 ? n20944 : ~n11107;
  assign n47312 = pi19 ? n47311 : n32;
  assign n47313 = pi18 ? n1379 : n47312;
  assign n47314 = pi17 ? n32 : n47313;
  assign n47315 = pi16 ? n32 : n47314;
  assign n47316 = pi15 ? n47315 : n47215;
  assign n47317 = pi14 ? n47205 : n47316;
  assign n47318 = pi13 ? n47193 : n47317;
  assign n47319 = pi12 ? n47318 : n32;
  assign n47320 = pi11 ? n47310 : n47319;
  assign n47321 = pi14 ? n21681 : n32;
  assign n47322 = pi13 ? n47321 : n32;
  assign n47323 = pi18 ? n880 : ~n23548;
  assign n47324 = pi17 ? n32 : n47323;
  assign n47325 = pi16 ? n1233 : ~n47324;
  assign n47326 = pi15 ? n47227 : n47325;
  assign n47327 = pi16 ? n1233 : ~n47233;
  assign n47328 = pi15 ? n47327 : n47243;
  assign n47329 = pi14 ? n47326 : n47328;
  assign n47330 = pi20 ? n3523 : ~n274;
  assign n47331 = pi19 ? n47330 : ~n32;
  assign n47332 = pi18 ? n863 : n47331;
  assign n47333 = pi17 ? n32 : n47332;
  assign n47334 = pi16 ? n1135 : ~n47333;
  assign n47335 = pi15 ? n33822 : n47334;
  assign n47336 = pi14 ? n47335 : n47252;
  assign n47337 = pi13 ? n47329 : n47336;
  assign n47338 = pi12 ? n47322 : n47337;
  assign n47339 = pi15 ? n47261 : n35359;
  assign n47340 = pi14 ? n47260 : n47339;
  assign n47341 = pi16 ? n1214 : ~n2426;
  assign n47342 = pi15 ? n47341 : n46441;
  assign n47343 = pi14 ? n46991 : n47342;
  assign n47344 = pi13 ? n47340 : n47343;
  assign n47345 = pi12 ? n47344 : n47277;
  assign n47346 = pi11 ? n47338 : n47345;
  assign n47347 = pi10 ? n47320 : n47346;
  assign n47348 = pi09 ? n32 : n47347;
  assign n47349 = pi08 ? n47281 : n47348;
  assign n47350 = pi15 ? n25001 : n23011;
  assign n47351 = pi14 ? n47350 : n22540;
  assign n47352 = pi20 ? n18129 : ~n9491;
  assign n47353 = pi19 ? n47352 : ~n36874;
  assign n47354 = pi18 ? n32 : n47353;
  assign n47355 = pi17 ? n32 : n47354;
  assign n47356 = pi19 ? n23644 : n247;
  assign n47357 = pi18 ? n47356 : n20020;
  assign n47358 = pi17 ? n47357 : n2618;
  assign n47359 = pi16 ? n47355 : ~n47358;
  assign n47360 = pi15 ? n32 : n47359;
  assign n47361 = pi18 ? n9461 : ~n30986;
  assign n47362 = pi19 ? n267 : n8622;
  assign n47363 = pi18 ? n47362 : n702;
  assign n47364 = pi17 ? n47361 : ~n47363;
  assign n47365 = pi16 ? n32 : n47364;
  assign n47366 = pi18 ? n1758 : ~n4343;
  assign n47367 = pi17 ? n47366 : ~n2750;
  assign n47368 = pi16 ? n32 : n47367;
  assign n47369 = pi15 ? n47365 : n47368;
  assign n47370 = pi14 ? n47360 : n47369;
  assign n47371 = pi13 ? n47351 : n47370;
  assign n47372 = pi19 ? n507 : n207;
  assign n47373 = pi18 ? n47372 : n18891;
  assign n47374 = pi19 ? n221 : n34188;
  assign n47375 = pi18 ? n47374 : n702;
  assign n47376 = pi17 ? n47373 : ~n47375;
  assign n47377 = pi16 ? n32 : n47376;
  assign n47378 = pi19 ? n32082 : n507;
  assign n47379 = pi18 ? n47378 : ~n702;
  assign n47380 = pi17 ? n3164 : n47379;
  assign n47381 = pi16 ? n32 : n47380;
  assign n47382 = pi15 ? n47377 : n47381;
  assign n47383 = pi20 ? n266 : n5854;
  assign n47384 = pi20 ? n246 : ~n220;
  assign n47385 = pi19 ? n47383 : n47384;
  assign n47386 = pi18 ? n47385 : ~n702;
  assign n47387 = pi17 ? n34459 : n47386;
  assign n47388 = pi16 ? n32 : n47387;
  assign n47389 = pi19 ? n6327 : n207;
  assign n47390 = pi18 ? n222 : n47389;
  assign n47391 = pi18 ? n16449 : n595;
  assign n47392 = pi17 ? n47390 : ~n47391;
  assign n47393 = pi16 ? n16605 : n47392;
  assign n47394 = pi15 ? n47388 : n47393;
  assign n47395 = pi14 ? n47382 : n47394;
  assign n47396 = pi19 ? n22185 : ~n804;
  assign n47397 = pi18 ? n47396 : n595;
  assign n47398 = pi17 ? n2959 : ~n47397;
  assign n47399 = pi16 ? n32 : n47398;
  assign n47400 = pi19 ? n462 : n1325;
  assign n47401 = pi18 ? n47400 : ~n595;
  assign n47402 = pi17 ? n32 : n47401;
  assign n47403 = pi16 ? n32 : n47402;
  assign n47404 = pi15 ? n47399 : n47403;
  assign n47405 = pi18 ? n32 : n24751;
  assign n47406 = pi17 ? n32 : n47405;
  assign n47407 = pi16 ? n32 : n47406;
  assign n47408 = pi15 ? n47170 : n47407;
  assign n47409 = pi14 ? n47404 : n47408;
  assign n47410 = pi13 ? n47395 : n47409;
  assign n47411 = pi12 ? n47371 : n47410;
  assign n47412 = pi18 ? n32 : ~n47144;
  assign n47413 = pi17 ? n32 : n47412;
  assign n47414 = pi16 ? n32 : n47413;
  assign n47415 = pi15 ? n35668 : n47414;
  assign n47416 = pi18 ? n940 : ~n47144;
  assign n47417 = pi17 ? n32 : n47416;
  assign n47418 = pi16 ? n32 : n47417;
  assign n47419 = pi19 ? n32 : n32340;
  assign n47420 = pi20 ? n32 : ~n13387;
  assign n47421 = pi19 ? n47420 : ~n32;
  assign n47422 = pi18 ? n47419 : ~n47421;
  assign n47423 = pi17 ? n16450 : n47422;
  assign n47424 = pi16 ? n32 : n47423;
  assign n47425 = pi15 ? n47418 : n47424;
  assign n47426 = pi14 ? n47415 : n47425;
  assign n47427 = pi19 ? n175 : ~n32;
  assign n47428 = pi18 ? n34445 : n47427;
  assign n47429 = pi19 ? n4391 : n236;
  assign n47430 = pi18 ? n47429 : ~n4098;
  assign n47431 = pi17 ? n47428 : n47430;
  assign n47432 = pi16 ? n16391 : n47431;
  assign n47433 = pi17 ? n34426 : n12068;
  assign n47434 = pi16 ? n32 : n47433;
  assign n47435 = pi15 ? n47432 : n47434;
  assign n47436 = pi15 ? n35650 : n24539;
  assign n47437 = pi14 ? n47435 : n47436;
  assign n47438 = pi13 ? n47426 : n47437;
  assign n47439 = pi12 ? n47438 : n32;
  assign n47440 = pi11 ? n47411 : n47439;
  assign n47441 = pi17 ? n17119 : n47323;
  assign n47442 = pi16 ? n1135 : ~n47441;
  assign n47443 = pi15 ? n47227 : n47442;
  assign n47444 = pi18 ? n209 : ~n5005;
  assign n47445 = pi17 ? n17433 : n47444;
  assign n47446 = pi16 ? n1135 : ~n47445;
  assign n47447 = pi19 ? n3692 : ~n33526;
  assign n47448 = pi18 ? n34030 : ~n47447;
  assign n47449 = pi19 ? n18489 : n208;
  assign n47450 = pi18 ? n47449 : ~n13945;
  assign n47451 = pi17 ? n47448 : ~n47450;
  assign n47452 = pi16 ? n1471 : n47451;
  assign n47453 = pi15 ? n47446 : n47452;
  assign n47454 = pi14 ? n47443 : n47453;
  assign n47455 = pi20 ? n357 : ~n274;
  assign n47456 = pi19 ? n47455 : ~n32;
  assign n47457 = pi18 ? n17848 : n47456;
  assign n47458 = pi17 ? n32 : n47457;
  assign n47459 = pi16 ? n1135 : ~n47458;
  assign n47460 = pi15 ? n47459 : n34044;
  assign n47461 = pi17 ? n16802 : n2408;
  assign n47462 = pi16 ? n1135 : ~n47461;
  assign n47463 = pi15 ? n34047 : n47462;
  assign n47464 = pi14 ? n47460 : n47463;
  assign n47465 = pi13 ? n47454 : n47464;
  assign n47466 = pi12 ? n32 : n47465;
  assign n47467 = pi18 ? n341 : ~n15849;
  assign n47468 = pi17 ? n32 : n47467;
  assign n47469 = pi16 ? n47468 : ~n2120;
  assign n47470 = pi15 ? n47256 : n47469;
  assign n47471 = pi16 ? n1214 : ~n2120;
  assign n47472 = pi15 ? n47256 : n47471;
  assign n47473 = pi14 ? n47470 : n47472;
  assign n47474 = pi17 ? n14395 : n2653;
  assign n47475 = pi16 ? n1214 : ~n47474;
  assign n47476 = pi17 ? n17119 : n2653;
  assign n47477 = pi16 ? n1214 : ~n47476;
  assign n47478 = pi15 ? n47475 : n47477;
  assign n47479 = pi14 ? n47264 : n47478;
  assign n47480 = pi13 ? n47473 : n47479;
  assign n47481 = pi19 ? n45626 : n32;
  assign n47482 = pi18 ? n28770 : n47481;
  assign n47483 = pi17 ? n32 : n47482;
  assign n47484 = pi16 ? n47483 : n34089;
  assign n47485 = pi15 ? n46441 : n47484;
  assign n47486 = pi19 ? n18111 : n34100;
  assign n47487 = pi18 ? n34098 : n47486;
  assign n47488 = pi17 ? n47487 : n34104;
  assign n47489 = pi16 ? n23249 : n47488;
  assign n47490 = pi15 ? n33135 : n47489;
  assign n47491 = pi14 ? n47485 : n47490;
  assign n47492 = pi15 ? n32 : n466;
  assign n47493 = pi14 ? n47492 : n1015;
  assign n47494 = pi13 ? n47491 : n47493;
  assign n47495 = pi12 ? n47480 : n47494;
  assign n47496 = pi11 ? n47466 : n47495;
  assign n47497 = pi10 ? n47440 : n47496;
  assign n47498 = pi09 ? n32 : n47497;
  assign n47499 = pi18 ? n47362 : n2622;
  assign n47500 = pi17 ? n47361 : ~n47499;
  assign n47501 = pi16 ? n32 : n47500;
  assign n47502 = pi17 ? n47366 : ~n2623;
  assign n47503 = pi16 ? n32 : n47502;
  assign n47504 = pi15 ? n47501 : n47503;
  assign n47505 = pi14 ? n47360 : n47504;
  assign n47506 = pi13 ? n47351 : n47505;
  assign n47507 = pi18 ? n47374 : n2622;
  assign n47508 = pi17 ? n47373 : ~n47507;
  assign n47509 = pi16 ? n32 : n47508;
  assign n47510 = pi18 ? n47378 : ~n2622;
  assign n47511 = pi17 ? n3164 : n47510;
  assign n47512 = pi16 ? n32 : n47511;
  assign n47513 = pi15 ? n47509 : n47512;
  assign n47514 = pi18 ? n47385 : ~n2622;
  assign n47515 = pi17 ? n34459 : n47514;
  assign n47516 = pi16 ? n32 : n47515;
  assign n47517 = pi18 ? n16449 : n702;
  assign n47518 = pi17 ? n47390 : ~n47517;
  assign n47519 = pi16 ? n16605 : n47518;
  assign n47520 = pi15 ? n47516 : n47519;
  assign n47521 = pi14 ? n47513 : n47520;
  assign n47522 = pi19 ? n462 : n1464;
  assign n47523 = pi20 ? n1331 : n1817;
  assign n47524 = pi19 ? n47523 : ~n32;
  assign n47525 = pi18 ? n47522 : ~n47524;
  assign n47526 = pi17 ? n32 : n47525;
  assign n47527 = pi16 ? n32 : n47526;
  assign n47528 = pi15 ? n47399 : n47527;
  assign n47529 = pi15 ? n47170 : n13904;
  assign n47530 = pi14 ? n47528 : n47529;
  assign n47531 = pi13 ? n47521 : n47530;
  assign n47532 = pi12 ? n47506 : n47531;
  assign n47533 = pi11 ? n47532 : n47439;
  assign n47534 = pi18 ? n880 : ~n23700;
  assign n47535 = pi17 ? n17119 : n47534;
  assign n47536 = pi16 ? n1233 : ~n47535;
  assign n47537 = pi15 ? n47227 : n47536;
  assign n47538 = pi18 ? n209 : ~n39705;
  assign n47539 = pi17 ? n17433 : n47538;
  assign n47540 = pi16 ? n1233 : ~n47539;
  assign n47541 = pi15 ? n47540 : n47452;
  assign n47542 = pi14 ? n47537 : n47541;
  assign n47543 = pi18 ? n17848 : n28193;
  assign n47544 = pi17 ? n32 : n47543;
  assign n47545 = pi16 ? n1135 : ~n47544;
  assign n47546 = pi15 ? n47545 : n34146;
  assign n47547 = pi14 ? n47546 : n47463;
  assign n47548 = pi13 ? n47542 : n47547;
  assign n47549 = pi12 ? n32 : n47548;
  assign n47550 = pi19 ? n6120 : n32;
  assign n47551 = pi18 ? n32 : ~n47550;
  assign n47552 = pi17 ? n32 : n47551;
  assign n47553 = pi16 ? n47468 : ~n47552;
  assign n47554 = pi15 ? n47256 : n47553;
  assign n47555 = pi16 ? n19652 : ~n2120;
  assign n47556 = pi15 ? n47256 : n47555;
  assign n47557 = pi14 ? n47554 : n47556;
  assign n47558 = pi13 ? n47557 : n47479;
  assign n47559 = pi18 ? n858 : n7221;
  assign n47560 = pi17 ? n32 : n47559;
  assign n47561 = pi16 ? n47560 : n34089;
  assign n47562 = pi15 ? n46441 : n47561;
  assign n47563 = pi18 ? n34098 : n4671;
  assign n47564 = pi20 ? n5854 : ~n206;
  assign n47565 = pi19 ? n32 : ~n47564;
  assign n47566 = pi18 ? n47565 : n6059;
  assign n47567 = pi17 ? n47563 : n47566;
  assign n47568 = pi16 ? n23249 : n47567;
  assign n47569 = pi15 ? n33135 : n47568;
  assign n47570 = pi14 ? n47562 : n47569;
  assign n47571 = pi14 ? n47492 : n466;
  assign n47572 = pi13 ? n47570 : n47571;
  assign n47573 = pi12 ? n47558 : n47572;
  assign n47574 = pi11 ? n47549 : n47573;
  assign n47575 = pi10 ? n47533 : n47574;
  assign n47576 = pi09 ? n32 : n47575;
  assign n47577 = pi08 ? n47498 : n47576;
  assign n47578 = pi07 ? n47349 : n47577;
  assign n47579 = pi06 ? n47123 : n47578;
  assign n47580 = pi05 ? n46673 : n47579;
  assign n47581 = pi13 ? n32 : n24328;
  assign n47582 = pi12 ? n32 : n47581;
  assign n47583 = pi11 ? n32 : n47582;
  assign n47584 = pi10 ? n32 : n47583;
  assign n47585 = pi14 ? n22923 : n1110;
  assign n47586 = pi19 ? n349 : ~n17757;
  assign n47587 = pi18 ? n17118 : ~n47586;
  assign n47588 = pi20 ? n5854 : n207;
  assign n47589 = pi20 ? n6621 : ~n2358;
  assign n47590 = pi19 ? n47588 : n47589;
  assign n47591 = pi20 ? n207 : ~n12019;
  assign n47592 = pi19 ? n47591 : n32;
  assign n47593 = pi18 ? n47590 : ~n47592;
  assign n47594 = pi17 ? n47587 : ~n47593;
  assign n47595 = pi16 ? n32 : n47594;
  assign n47596 = pi15 ? n32 : n47595;
  assign n47597 = pi20 ? n3843 : ~n18408;
  assign n47598 = pi19 ? n47597 : n36181;
  assign n47599 = pi18 ? n32 : n47598;
  assign n47600 = pi17 ? n32 : n47599;
  assign n47601 = pi19 ? n36182 : n4670;
  assign n47602 = pi19 ? n18678 : n4670;
  assign n47603 = pi18 ? n47601 : n47602;
  assign n47604 = pi18 ? n22554 : n2622;
  assign n47605 = pi17 ? n47603 : n47604;
  assign n47606 = pi16 ? n47600 : ~n47605;
  assign n47607 = pi19 ? n594 : n207;
  assign n47608 = pi18 ? n47607 : n18891;
  assign n47609 = pi19 ? n1464 : n35996;
  assign n47610 = pi18 ? n47609 : n2622;
  assign n47611 = pi17 ? n47608 : ~n47610;
  assign n47612 = pi16 ? n32 : n47611;
  assign n47613 = pi15 ? n47606 : n47612;
  assign n47614 = pi14 ? n47596 : n47613;
  assign n47615 = pi13 ? n47585 : n47614;
  assign n47616 = pi17 ? n23052 : n47510;
  assign n47617 = pi16 ? n32 : n47616;
  assign n47618 = pi20 ? n32 : ~n9488;
  assign n47619 = pi19 ? n32 : n47618;
  assign n47620 = pi18 ? n32 : n47619;
  assign n47621 = pi17 ? n32 : n47620;
  assign n47622 = pi19 ? n31202 : ~n35706;
  assign n47623 = pi20 ? n9491 : n2358;
  assign n47624 = pi19 ? n47623 : ~n266;
  assign n47625 = pi18 ? n47622 : n47624;
  assign n47626 = pi20 ? n220 : ~n1611;
  assign n47627 = pi20 ? n1076 : ~n342;
  assign n47628 = pi19 ? n47626 : ~n47627;
  assign n47629 = pi18 ? n47628 : n13318;
  assign n47630 = pi17 ? n47625 : n47629;
  assign n47631 = pi16 ? n47621 : n47630;
  assign n47632 = pi15 ? n47617 : n47631;
  assign n47633 = pi19 ? n32 : ~n24055;
  assign n47634 = pi18 ? n863 : n47633;
  assign n47635 = pi19 ? n17641 : n1138;
  assign n47636 = pi18 ? n47635 : ~n2622;
  assign n47637 = pi17 ? n47634 : n47636;
  assign n47638 = pi16 ? n32 : n47637;
  assign n47639 = pi17 ? n2954 : n47296;
  assign n47640 = pi16 ? n32 : n47639;
  assign n47641 = pi15 ? n47638 : n47640;
  assign n47642 = pi14 ? n47632 : n47641;
  assign n47643 = pi19 ? n9007 : n1508;
  assign n47644 = pi18 ? n47643 : ~n702;
  assign n47645 = pi17 ? n23052 : n47644;
  assign n47646 = pi16 ? n16836 : n47645;
  assign n47647 = pi19 ? n358 : ~n32;
  assign n47648 = pi18 ? n863 : ~n47647;
  assign n47649 = pi17 ? n32 : n47648;
  assign n47650 = pi16 ? n32 : n47649;
  assign n47651 = pi15 ? n47646 : n47650;
  assign n47652 = pi15 ? n13620 : n25846;
  assign n47653 = pi14 ? n47651 : n47652;
  assign n47654 = pi13 ? n47642 : n47653;
  assign n47655 = pi12 ? n47615 : n47654;
  assign n47656 = pi20 ? n3523 : ~n18415;
  assign n47657 = pi19 ? n32 : n47656;
  assign n47658 = pi18 ? n32 : n47657;
  assign n47659 = pi19 ? n33526 : ~n29761;
  assign n47660 = pi18 ? n47659 : n37093;
  assign n47661 = pi17 ? n47658 : ~n47660;
  assign n47662 = pi16 ? n32 : n47661;
  assign n47663 = pi15 ? n22817 : n47662;
  assign n47664 = pi20 ? n321 : ~n1611;
  assign n47665 = pi19 ? n32 : n47664;
  assign n47666 = pi18 ? n32 : n47665;
  assign n47667 = pi19 ? n5741 : ~n32;
  assign n47668 = pi18 ? n37537 : n47667;
  assign n47669 = pi17 ? n47666 : ~n47668;
  assign n47670 = pi16 ? n32 : n47669;
  assign n47671 = pi18 ? n32 : n18183;
  assign n47672 = pi19 ? n18502 : ~n1740;
  assign n47673 = pi19 ? n36903 : ~n32;
  assign n47674 = pi18 ? n47672 : n47673;
  assign n47675 = pi17 ? n47671 : ~n47674;
  assign n47676 = pi16 ? n32 : n47675;
  assign n47677 = pi15 ? n47670 : n47676;
  assign n47678 = pi14 ? n47663 : n47677;
  assign n47679 = pi18 ? n4380 : ~n6500;
  assign n47680 = pi17 ? n17346 : n47679;
  assign n47681 = pi16 ? n32 : n47680;
  assign n47682 = pi20 ? n274 : n342;
  assign n47683 = pi19 ? n47682 : ~n32;
  assign n47684 = pi18 ? n936 : ~n47683;
  assign n47685 = pi17 ? n32 : n47684;
  assign n47686 = pi16 ? n32 : n47685;
  assign n47687 = pi15 ? n47681 : n47686;
  assign n47688 = pi15 ? n14156 : n32;
  assign n47689 = pi14 ? n47687 : n47688;
  assign n47690 = pi13 ? n47678 : n47689;
  assign n47691 = pi14 ? n32 : n648;
  assign n47692 = pi13 ? n32 : n47691;
  assign n47693 = pi12 ? n47690 : n47692;
  assign n47694 = pi11 ? n47655 : n47693;
  assign n47695 = pi17 ? n16848 : n1697;
  assign n47696 = pi16 ? n3068 : ~n47695;
  assign n47697 = pi14 ? n32 : n47696;
  assign n47698 = pi13 ? n32 : n47697;
  assign n47699 = pi15 ? n29676 : n42583;
  assign n47700 = pi17 ? n17346 : n1706;
  assign n47701 = pi16 ? n1214 : ~n47700;
  assign n47702 = pi19 ? n22501 : n4342;
  assign n47703 = pi18 ? n341 : n47702;
  assign n47704 = pi17 ? n32 : n47703;
  assign n47705 = pi17 ? n26426 : n47444;
  assign n47706 = pi16 ? n47704 : ~n47705;
  assign n47707 = pi15 ? n47701 : n47706;
  assign n47708 = pi14 ? n47699 : n47707;
  assign n47709 = pi16 ? n28804 : ~n3769;
  assign n47710 = pi16 ? n1135 : ~n3769;
  assign n47711 = pi15 ? n47709 : n47710;
  assign n47712 = pi19 ? n18496 : ~n9345;
  assign n47713 = pi18 ? n268 : ~n47712;
  assign n47714 = pi17 ? n32 : n47713;
  assign n47715 = pi17 ? n23052 : n2519;
  assign n47716 = pi16 ? n47714 : ~n47715;
  assign n47717 = pi18 ? n209 : ~n6059;
  assign n47718 = pi17 ? n32 : n47717;
  assign n47719 = pi17 ? n46383 : n2119;
  assign n47720 = pi16 ? n47718 : ~n47719;
  assign n47721 = pi15 ? n47716 : n47720;
  assign n47722 = pi14 ? n47711 : n47721;
  assign n47723 = pi13 ? n47708 : n47722;
  assign n47724 = pi12 ? n47698 : n47723;
  assign n47725 = pi20 ? n18832 : n9491;
  assign n47726 = pi20 ? n17652 : n18253;
  assign n47727 = pi19 ? n47725 : n47726;
  assign n47728 = pi18 ? n41321 : ~n47727;
  assign n47729 = pi17 ? n32 : n47728;
  assign n47730 = pi19 ? n9863 : n1076;
  assign n47731 = pi20 ? n1076 : n1817;
  assign n47732 = pi19 ? n47731 : n5614;
  assign n47733 = pi18 ? n47730 : n47732;
  assign n47734 = pi20 ? n14286 : ~n339;
  assign n47735 = pi19 ? n47734 : n32;
  assign n47736 = pi18 ? n47735 : n605;
  assign n47737 = pi17 ? n47733 : n47736;
  assign n47738 = pi16 ? n47729 : ~n47737;
  assign n47739 = pi19 ? n18722 : n32;
  assign n47740 = pi18 ? n209 : ~n47739;
  assign n47741 = pi17 ? n32 : n47740;
  assign n47742 = pi16 ? n47741 : ~n2120;
  assign n47743 = pi15 ? n47738 : n47742;
  assign n47744 = pi19 ? n4391 : ~n322;
  assign n47745 = pi18 ? n209 : n47744;
  assign n47746 = pi17 ? n32 : n47745;
  assign n47747 = pi18 ? n8192 : n4343;
  assign n47748 = pi17 ? n47747 : n2119;
  assign n47749 = pi16 ? n47746 : ~n47748;
  assign n47750 = pi19 ? n1757 : n322;
  assign n47751 = pi18 ? n940 : ~n47750;
  assign n47752 = pi17 ? n32 : n47751;
  assign n47753 = pi19 ? n9007 : n18478;
  assign n47754 = pi19 ? n4342 : ~n18502;
  assign n47755 = pi18 ? n47753 : n47754;
  assign n47756 = pi19 ? n247 : ~n236;
  assign n47757 = pi18 ? n47756 : n605;
  assign n47758 = pi17 ? n47755 : n47757;
  assign n47759 = pi16 ? n47752 : ~n47758;
  assign n47760 = pi15 ? n47749 : n47759;
  assign n47761 = pi14 ? n47743 : n47760;
  assign n47762 = pi19 ? n32 : ~n24349;
  assign n47763 = pi18 ? n18710 : ~n47762;
  assign n47764 = pi17 ? n32 : n47763;
  assign n47765 = pi18 ? n18891 : ~n32;
  assign n47766 = pi17 ? n47765 : ~n2119;
  assign n47767 = pi16 ? n47764 : n47766;
  assign n47768 = pi19 ? n322 : n18390;
  assign n47769 = pi18 ? n32 : n47768;
  assign n47770 = pi17 ? n32 : n47769;
  assign n47771 = pi19 ? n23895 : ~n22525;
  assign n47772 = pi19 ? n247 : n221;
  assign n47773 = pi18 ? n47771 : n47772;
  assign n47774 = pi19 ? n32733 : n32;
  assign n47775 = pi18 ? n47774 : n605;
  assign n47776 = pi17 ? n47773 : n47775;
  assign n47777 = pi16 ? n47770 : ~n47776;
  assign n47778 = pi15 ? n47767 : n47777;
  assign n47779 = pi19 ? n9007 : n24055;
  assign n47780 = pi19 ? n9037 : n6339;
  assign n47781 = pi18 ? n47779 : n47780;
  assign n47782 = pi19 ? n3692 : ~n349;
  assign n47783 = pi18 ? n47782 : n605;
  assign n47784 = pi17 ? n47781 : n47783;
  assign n47785 = pi16 ? n34526 : ~n47784;
  assign n47786 = pi19 ? n246 : n22652;
  assign n47787 = pi18 ? n18199 : ~n47786;
  assign n47788 = pi17 ? n32 : n47787;
  assign n47789 = pi20 ? n3843 : ~n501;
  assign n47790 = pi19 ? n2358 : ~n47789;
  assign n47791 = pi19 ? n19583 : ~n17649;
  assign n47792 = pi18 ? n47790 : n47791;
  assign n47793 = pi18 ? n248 : n430;
  assign n47794 = pi17 ? n47792 : ~n47793;
  assign n47795 = pi16 ? n47788 : n47794;
  assign n47796 = pi15 ? n47785 : n47795;
  assign n47797 = pi14 ? n47778 : n47796;
  assign n47798 = pi13 ? n47761 : n47797;
  assign n47799 = pi20 ? n354 : ~n266;
  assign n47800 = pi20 ? n266 : n287;
  assign n47801 = pi19 ? n47799 : n47800;
  assign n47802 = pi18 ? n268 : ~n47801;
  assign n47803 = pi17 ? n32 : n47802;
  assign n47804 = pi20 ? n3523 : ~n9491;
  assign n47805 = pi19 ? n266 : n47804;
  assign n47806 = pi19 ? n6314 : n1165;
  assign n47807 = pi18 ? n47805 : n47806;
  assign n47808 = pi18 ? n4492 : n532;
  assign n47809 = pi17 ? n47807 : n47808;
  assign n47810 = pi16 ? n47803 : ~n47809;
  assign n47811 = pi15 ? n47810 : n34308;
  assign n47812 = pi15 ? n34312 : n32;
  assign n47813 = pi14 ? n47811 : n47812;
  assign n47814 = pi16 ? n129 : n179;
  assign n47815 = pi15 ? n32 : n47814;
  assign n47816 = pi14 ? n47815 : n47814;
  assign n47817 = pi13 ? n47813 : n47816;
  assign n47818 = pi12 ? n47798 : n47817;
  assign n47819 = pi11 ? n47724 : n47818;
  assign n47820 = pi10 ? n47694 : n47819;
  assign n47821 = pi09 ? n47584 : n47820;
  assign n47822 = pi18 ? n47590 : ~n13335;
  assign n47823 = pi17 ? n47587 : ~n47822;
  assign n47824 = pi16 ? n32 : n47823;
  assign n47825 = pi15 ? n32 : n47824;
  assign n47826 = pi20 ? n1331 : ~n18408;
  assign n47827 = pi19 ? n47826 : n36181;
  assign n47828 = pi18 ? n32 : n47827;
  assign n47829 = pi17 ? n32 : n47828;
  assign n47830 = pi18 ? n22554 : n1750;
  assign n47831 = pi17 ? n47603 : n47830;
  assign n47832 = pi16 ? n47829 : ~n47831;
  assign n47833 = pi18 ? n47609 : n1750;
  assign n47834 = pi17 ? n47608 : ~n47833;
  assign n47835 = pi16 ? n32 : n47834;
  assign n47836 = pi15 ? n47832 : n47835;
  assign n47837 = pi14 ? n47825 : n47836;
  assign n47838 = pi13 ? n23089 : n47837;
  assign n47839 = pi18 ? n47378 : ~n1750;
  assign n47840 = pi17 ? n23052 : n47839;
  assign n47841 = pi16 ? n32 : n47840;
  assign n47842 = pi19 ? n236 : ~n617;
  assign n47843 = pi18 ? n47628 : n47842;
  assign n47844 = pi17 ? n47625 : n47843;
  assign n47845 = pi16 ? n47621 : n47844;
  assign n47846 = pi15 ? n47841 : n47845;
  assign n47847 = pi18 ? n47635 : ~n702;
  assign n47848 = pi17 ? n47634 : n47847;
  assign n47849 = pi16 ? n32 : n47848;
  assign n47850 = pi15 ? n47849 : n47640;
  assign n47851 = pi14 ? n47846 : n47850;
  assign n47852 = pi19 ? n1248 : ~n1105;
  assign n47853 = pi18 ? n32 : n47852;
  assign n47854 = pi17 ? n32 : n47853;
  assign n47855 = pi16 ? n32 : n47854;
  assign n47856 = pi15 ? n35947 : n47855;
  assign n47857 = pi14 ? n47651 : n47856;
  assign n47858 = pi13 ? n47851 : n47857;
  assign n47859 = pi12 ? n47838 : n47858;
  assign n47860 = pi18 ? n4380 : ~n702;
  assign n47861 = pi17 ? n17346 : n47860;
  assign n47862 = pi16 ? n32 : n47861;
  assign n47863 = pi18 ? n32 : ~n46915;
  assign n47864 = pi17 ? n32 : n47863;
  assign n47865 = pi16 ? n32 : n47864;
  assign n47866 = pi15 ? n47862 : n47865;
  assign n47867 = pi14 ? n47866 : n47688;
  assign n47868 = pi13 ? n47678 : n47867;
  assign n47869 = pi14 ? n22424 : n32;
  assign n47870 = pi13 ? n47869 : n32;
  assign n47871 = pi12 ? n47868 : n47870;
  assign n47872 = pi11 ? n47859 : n47871;
  assign n47873 = pi16 ? n1233 : ~n42582;
  assign n47874 = pi15 ? n29519 : n47873;
  assign n47875 = pi16 ? n19652 : ~n47700;
  assign n47876 = pi15 ? n47875 : n47706;
  assign n47877 = pi14 ? n47874 : n47876;
  assign n47878 = pi13 ? n47877 : n47722;
  assign n47879 = pi12 ? n47698 : n47878;
  assign n47880 = pi20 ? n18173 : n314;
  assign n47881 = pi20 ? n17652 : ~n1331;
  assign n47882 = pi19 ? n47880 : n47881;
  assign n47883 = pi18 ? n312 : ~n47882;
  assign n47884 = pi17 ? n32 : n47883;
  assign n47885 = pi19 ? n1685 : n321;
  assign n47886 = pi20 ? n6621 : n6085;
  assign n47887 = pi19 ? n18390 : n47886;
  assign n47888 = pi18 ? n47885 : n47887;
  assign n47889 = pi20 ? n3695 : ~n18624;
  assign n47890 = pi19 ? n47889 : n32;
  assign n47891 = pi18 ? n47890 : n605;
  assign n47892 = pi17 ? n47888 : n47891;
  assign n47893 = pi16 ? n47884 : ~n47892;
  assign n47894 = pi15 ? n47893 : n47742;
  assign n47895 = pi14 ? n47894 : n47760;
  assign n47896 = pi18 ? n47774 : n2413;
  assign n47897 = pi17 ? n47773 : n47896;
  assign n47898 = pi16 ? n47770 : ~n47897;
  assign n47899 = pi15 ? n47767 : n47898;
  assign n47900 = pi18 ? n4127 : ~n47786;
  assign n47901 = pi17 ? n32 : n47900;
  assign n47902 = pi16 ? n47901 : n47794;
  assign n47903 = pi15 ? n47785 : n47902;
  assign n47904 = pi14 ? n47899 : n47903;
  assign n47905 = pi13 ? n47895 : n47904;
  assign n47906 = pi13 ? n47813 : n47276;
  assign n47907 = pi12 ? n47905 : n47906;
  assign n47908 = pi11 ? n47879 : n47907;
  assign n47909 = pi10 ? n47872 : n47908;
  assign n47910 = pi09 ? n47584 : n47909;
  assign n47911 = pi08 ? n47821 : n47910;
  assign n47912 = pi13 ? n32 : n24608;
  assign n47913 = pi12 ? n32 : n47912;
  assign n47914 = pi11 ? n32 : n47913;
  assign n47915 = pi10 ? n32 : n47914;
  assign n47916 = pi15 ? n15518 : n15665;
  assign n47917 = pi14 ? n47916 : n32;
  assign n47918 = pi18 ? n237 : ~n23514;
  assign n47919 = pi17 ? n32 : ~n47918;
  assign n47920 = pi16 ? n32 : n47919;
  assign n47921 = pi15 ? n32 : n47920;
  assign n47922 = pi18 ? n18891 : n1750;
  assign n47923 = pi17 ? n32 : ~n47922;
  assign n47924 = pi16 ? n32 : n47923;
  assign n47925 = pi15 ? n25790 : n47924;
  assign n47926 = pi14 ? n47921 : n47925;
  assign n47927 = pi13 ? n47917 : n47926;
  assign n47928 = pi18 ? n32 : ~n1750;
  assign n47929 = pi17 ? n32 : n47928;
  assign n47930 = pi16 ? n32 : n47929;
  assign n47931 = pi18 ? n248 : n25787;
  assign n47932 = pi17 ? n2954 : n47931;
  assign n47933 = pi16 ? n32 : n47932;
  assign n47934 = pi15 ? n47930 : n47933;
  assign n47935 = pi19 ? n29286 : n6327;
  assign n47936 = pi18 ? n47935 : ~n702;
  assign n47937 = pi17 ? n36403 : n47936;
  assign n47938 = pi16 ? n32 : n47937;
  assign n47939 = pi15 ? n47938 : n47640;
  assign n47940 = pi14 ? n47934 : n47939;
  assign n47941 = pi19 ? n4558 : n32;
  assign n47942 = pi18 ? n32 : n47941;
  assign n47943 = pi17 ? n32 : n47942;
  assign n47944 = pi16 ? n32 : n47943;
  assign n47945 = pi15 ? n47944 : n35650;
  assign n47946 = pi19 ? n5741 : ~n1105;
  assign n47947 = pi18 ? n32 : n47946;
  assign n47948 = pi17 ? n32 : n47947;
  assign n47949 = pi16 ? n32 : n47948;
  assign n47950 = pi15 ? n47949 : n15119;
  assign n47951 = pi14 ? n47945 : n47950;
  assign n47952 = pi13 ? n47940 : n47951;
  assign n47953 = pi12 ? n47927 : n47952;
  assign n47954 = pi19 ? n5741 : n1105;
  assign n47955 = pi18 ? n32 : ~n47954;
  assign n47956 = pi17 ? n32 : n47955;
  assign n47957 = pi16 ? n32 : n47956;
  assign n47958 = pi15 ? n23011 : n47957;
  assign n47959 = pi18 ? n1613 : ~n47954;
  assign n47960 = pi17 ? n32 : n47959;
  assign n47961 = pi16 ? n32 : n47960;
  assign n47962 = pi19 ? n4964 : n1105;
  assign n47963 = pi18 ? n32 : ~n47962;
  assign n47964 = pi17 ? n32 : n47963;
  assign n47965 = pi16 ? n32 : n47964;
  assign n47966 = pi15 ? n47961 : n47965;
  assign n47967 = pi14 ? n47958 : n47966;
  assign n47968 = pi15 ? n13032 : n13629;
  assign n47969 = pi14 ? n47968 : n32;
  assign n47970 = pi13 ? n47967 : n47969;
  assign n47971 = pi13 ? n21930 : n32;
  assign n47972 = pi12 ? n47970 : n47971;
  assign n47973 = pi11 ? n47953 : n47972;
  assign n47974 = pi14 ? n21320 : n47696;
  assign n47975 = pi13 ? n32 : n47974;
  assign n47976 = pi19 ? n32 : n19582;
  assign n47977 = pi18 ? n47976 : ~n32;
  assign n47978 = pi17 ? n32 : n47977;
  assign n47979 = pi17 ? n23052 : n1470;
  assign n47980 = pi16 ? n47978 : ~n47979;
  assign n47981 = pi20 ? n32 : n6050;
  assign n47982 = pi19 ? n32 : n47981;
  assign n47983 = pi18 ? n47982 : ~n32;
  assign n47984 = pi17 ? n32 : n47983;
  assign n47985 = pi16 ? n47984 : ~n47979;
  assign n47986 = pi15 ? n47980 : n47985;
  assign n47987 = pi19 ? n21740 : ~n1757;
  assign n47988 = pi18 ? n32 : n47987;
  assign n47989 = pi17 ? n32 : n47988;
  assign n47990 = pi17 ? n17346 : n1470;
  assign n47991 = pi16 ? n47989 : ~n47990;
  assign n47992 = pi20 ? n32 : n18073;
  assign n47993 = pi19 ? n32 : n47992;
  assign n47994 = pi20 ? n9491 : n2180;
  assign n47995 = pi19 ? n47994 : n20884;
  assign n47996 = pi18 ? n47993 : n47995;
  assign n47997 = pi17 ? n32 : n47996;
  assign n47998 = pi17 ? n32 : ~n10245;
  assign n47999 = pi16 ? n47997 : ~n47998;
  assign n48000 = pi15 ? n47991 : n47999;
  assign n48001 = pi14 ? n47986 : n48000;
  assign n48002 = pi18 ? n833 : ~n5657;
  assign n48003 = pi17 ? n32 : n48002;
  assign n48004 = pi16 ? n48003 : ~n2756;
  assign n48005 = pi19 ? n21655 : n1077;
  assign n48006 = pi18 ? n858 : n48005;
  assign n48007 = pi17 ? n32 : n48006;
  assign n48008 = pi16 ? n48007 : ~n2756;
  assign n48009 = pi15 ? n48004 : n48008;
  assign n48010 = pi20 ? n266 : ~n29457;
  assign n48011 = pi19 ? n29476 : n48010;
  assign n48012 = pi18 ? n312 : n48011;
  assign n48013 = pi17 ? n32 : n48012;
  assign n48014 = pi18 ? n237 : ~n2754;
  assign n48015 = pi17 ? n32 : ~n48014;
  assign n48016 = pi16 ? n48013 : ~n48015;
  assign n48017 = pi17 ? n3164 : n2519;
  assign n48018 = pi16 ? n42252 : ~n48017;
  assign n48019 = pi15 ? n48016 : n48018;
  assign n48020 = pi14 ? n48009 : n48019;
  assign n48021 = pi13 ? n48001 : n48020;
  assign n48022 = pi12 ? n47975 : n48021;
  assign n48023 = pi19 ? n9007 : ~n7168;
  assign n48024 = pi19 ? n1331 : ~n18496;
  assign n48025 = pi18 ? n48023 : n48024;
  assign n48026 = pi19 ? n18497 : ~n1757;
  assign n48027 = pi18 ? n48026 : ~n797;
  assign n48028 = pi17 ? n48025 : n48027;
  assign n48029 = pi16 ? n32 : n48028;
  assign n48030 = pi20 ? n321 : n6050;
  assign n48031 = pi19 ? n48030 : ~n21329;
  assign n48032 = pi18 ? n940 : n48031;
  assign n48033 = pi17 ? n32 : n48032;
  assign n48034 = pi17 ? n1028 : ~n2408;
  assign n48035 = pi16 ? n48033 : n48034;
  assign n48036 = pi15 ? n48029 : n48035;
  assign n48037 = pi18 ? n940 : n47744;
  assign n48038 = pi17 ? n32 : n48037;
  assign n48039 = pi17 ? n47747 : n5945;
  assign n48040 = pi16 ? n48038 : ~n48039;
  assign n48041 = pi18 ? n940 : ~n28382;
  assign n48042 = pi17 ? n32 : n48041;
  assign n48043 = pi20 ? n3523 : ~n1076;
  assign n48044 = pi19 ? n9007 : ~n48043;
  assign n48045 = pi19 ? n47731 : ~n24343;
  assign n48046 = pi18 ? n48044 : n48045;
  assign n48047 = pi19 ? n18497 : ~n4391;
  assign n48048 = pi18 ? n48047 : n605;
  assign n48049 = pi17 ? n48046 : n48048;
  assign n48050 = pi16 ? n48042 : ~n48049;
  assign n48051 = pi15 ? n48040 : n48050;
  assign n48052 = pi14 ? n48036 : n48051;
  assign n48053 = pi20 ? n7939 : n501;
  assign n48054 = pi19 ? n6339 : ~n48053;
  assign n48055 = pi18 ? n1613 : ~n48054;
  assign n48056 = pi17 ? n32 : n48055;
  assign n48057 = pi19 ? n321 : ~n342;
  assign n48058 = pi19 ? n4670 : n18084;
  assign n48059 = pi18 ? n48057 : ~n48058;
  assign n48060 = pi18 ? n13945 : n2413;
  assign n48061 = pi17 ? n48059 : ~n48060;
  assign n48062 = pi16 ? n48056 : n48061;
  assign n48063 = pi19 ? n11879 : ~n23895;
  assign n48064 = pi19 ? n4670 : n1464;
  assign n48065 = pi18 ? n48063 : n48064;
  assign n48066 = pi18 ? n28162 : n2413;
  assign n48067 = pi17 ? n48065 : n48066;
  assign n48068 = pi16 ? n47770 : ~n48067;
  assign n48069 = pi15 ? n48062 : n48068;
  assign n48070 = pi18 ? n127 : ~n248;
  assign n48071 = pi17 ? n32 : n48070;
  assign n48072 = pi19 ? n267 : n342;
  assign n48073 = pi18 ? n48072 : n4380;
  assign n48074 = pi17 ? n48073 : n2119;
  assign n48075 = pi16 ? n48071 : ~n48074;
  assign n48076 = pi19 ? n18390 : n45905;
  assign n48077 = pi18 ? n32 : ~n48076;
  assign n48078 = pi17 ? n32 : n48077;
  assign n48079 = pi19 ? n342 : ~n20555;
  assign n48080 = pi19 ? n5435 : ~n321;
  assign n48081 = pi18 ? n48079 : n48080;
  assign n48082 = pi20 ? n4279 : n274;
  assign n48083 = pi19 ? n48082 : n32;
  assign n48084 = pi18 ? n48083 : n605;
  assign n48085 = pi17 ? n48081 : ~n48084;
  assign n48086 = pi16 ? n48078 : n48085;
  assign n48087 = pi15 ? n48075 : n48086;
  assign n48088 = pi14 ? n48069 : n48087;
  assign n48089 = pi13 ? n48052 : n48088;
  assign n48090 = pi14 ? n34515 : n32;
  assign n48091 = pi13 ? n48090 : n47276;
  assign n48092 = pi12 ? n48089 : n48091;
  assign n48093 = pi11 ? n48022 : n48092;
  assign n48094 = pi10 ? n47973 : n48093;
  assign n48095 = pi09 ? n47915 : n48094;
  assign n48096 = pi14 ? n15518 : n32;
  assign n48097 = pi19 ? n236 : n5626;
  assign n48098 = pi18 ? n237 : ~n48097;
  assign n48099 = pi17 ? n32 : ~n48098;
  assign n48100 = pi16 ? n32 : n48099;
  assign n48101 = pi15 ? n32 : n48100;
  assign n48102 = pi18 ? n18891 : n2615;
  assign n48103 = pi17 ? n32 : ~n48102;
  assign n48104 = pi16 ? n32 : n48103;
  assign n48105 = pi15 ? n25840 : n48104;
  assign n48106 = pi14 ? n48101 : n48105;
  assign n48107 = pi13 ? n48096 : n48106;
  assign n48108 = pi18 ? n32 : ~n2615;
  assign n48109 = pi17 ? n32 : n48108;
  assign n48110 = pi16 ? n32 : n48109;
  assign n48111 = pi18 ? n248 : n25837;
  assign n48112 = pi17 ? n2954 : n48111;
  assign n48113 = pi16 ? n32 : n48112;
  assign n48114 = pi15 ? n48110 : n48113;
  assign n48115 = pi14 ? n48114 : n47939;
  assign n48116 = pi15 ? n13904 : n35650;
  assign n48117 = pi19 ? n5741 : ~n617;
  assign n48118 = pi18 ? n32 : n48117;
  assign n48119 = pi17 ? n32 : n48118;
  assign n48120 = pi16 ? n32 : n48119;
  assign n48121 = pi15 ? n48120 : n15119;
  assign n48122 = pi14 ? n48116 : n48121;
  assign n48123 = pi13 ? n48115 : n48122;
  assign n48124 = pi12 ? n48107 : n48123;
  assign n48125 = pi18 ? n32 : ~n47667;
  assign n48126 = pi17 ? n32 : n48125;
  assign n48127 = pi16 ? n32 : n48126;
  assign n48128 = pi15 ? n22817 : n48127;
  assign n48129 = pi14 ? n48128 : n47966;
  assign n48130 = pi13 ? n48129 : n47969;
  assign n48131 = pi12 ? n48130 : n47971;
  assign n48132 = pi11 ? n48124 : n48131;
  assign n48133 = pi14 ? n659 : n47696;
  assign n48134 = pi13 ? n32 : n48133;
  assign n48135 = pi18 ? n940 : ~n2093;
  assign n48136 = pi17 ? n23052 : n48135;
  assign n48137 = pi16 ? n47978 : ~n48136;
  assign n48138 = pi16 ? n47984 : ~n48136;
  assign n48139 = pi15 ? n48137 : n48138;
  assign n48140 = pi17 ? n17346 : n48135;
  assign n48141 = pi16 ? n47989 : ~n48140;
  assign n48142 = pi20 ? n9491 : n1076;
  assign n48143 = pi19 ? n48142 : n20884;
  assign n48144 = pi18 ? n38852 : n48143;
  assign n48145 = pi17 ? n32 : n48144;
  assign n48146 = pi16 ? n48145 : ~n47998;
  assign n48147 = pi15 ? n48141 : n48146;
  assign n48148 = pi14 ? n48139 : n48147;
  assign n48149 = pi16 ? n48003 : ~n2518;
  assign n48150 = pi16 ? n48007 : ~n2518;
  assign n48151 = pi15 ? n48149 : n48150;
  assign n48152 = pi18 ? n237 : ~n520;
  assign n48153 = pi17 ? n32 : ~n48152;
  assign n48154 = pi16 ? n48013 : ~n48153;
  assign n48155 = pi15 ? n48154 : n48018;
  assign n48156 = pi14 ? n48151 : n48155;
  assign n48157 = pi13 ? n48148 : n48156;
  assign n48158 = pi12 ? n48134 : n48157;
  assign n48159 = pi18 ? n13945 : n797;
  assign n48160 = pi17 ? n48059 : ~n48159;
  assign n48161 = pi16 ? n48056 : n48160;
  assign n48162 = pi18 ? n28162 : n605;
  assign n48163 = pi17 ? n48065 : n48162;
  assign n48164 = pi16 ? n47770 : ~n48163;
  assign n48165 = pi15 ? n48161 : n48164;
  assign n48166 = pi18 ? n32 : ~n248;
  assign n48167 = pi17 ? n32 : n48166;
  assign n48168 = pi16 ? n48167 : ~n48074;
  assign n48169 = pi15 ? n48168 : n48086;
  assign n48170 = pi14 ? n48165 : n48169;
  assign n48171 = pi13 ? n48052 : n48170;
  assign n48172 = pi14 ? n34580 : n32;
  assign n48173 = pi14 ? n47275 : n32;
  assign n48174 = pi13 ? n48172 : n48173;
  assign n48175 = pi12 ? n48171 : n48174;
  assign n48176 = pi11 ? n48158 : n48175;
  assign n48177 = pi10 ? n48132 : n48176;
  assign n48178 = pi09 ? n47915 : n48177;
  assign n48179 = pi08 ? n48095 : n48178;
  assign n48180 = pi07 ? n47911 : n48179;
  assign n48181 = pi15 ? n32 : n23250;
  assign n48182 = pi14 ? n32 : n48181;
  assign n48183 = pi13 ? n32 : n48182;
  assign n48184 = pi12 ? n32 : n48183;
  assign n48185 = pi11 ? n32 : n48184;
  assign n48186 = pi10 ? n32 : n48185;
  assign n48187 = pi15 ? n22817 : n32;
  assign n48188 = pi14 ? n48187 : n25840;
  assign n48189 = pi13 ? n23426 : n48188;
  assign n48190 = pi19 ? n236 : ~n2614;
  assign n48191 = pi18 ? n32 : n48190;
  assign n48192 = pi17 ? n32 : n48191;
  assign n48193 = pi16 ? n32 : n48192;
  assign n48194 = pi15 ? n25840 : n48193;
  assign n48195 = pi15 ? n47930 : n25790;
  assign n48196 = pi14 ? n48194 : n48195;
  assign n48197 = pi15 ? n13620 : n13904;
  assign n48198 = pi15 ? n24528 : n15382;
  assign n48199 = pi14 ? n48197 : n48198;
  assign n48200 = pi13 ? n48196 : n48199;
  assign n48201 = pi12 ? n48189 : n48200;
  assign n48202 = pi20 ? n220 : n2358;
  assign n48203 = pi19 ? n48202 : ~n617;
  assign n48204 = pi18 ? n6118 : n48203;
  assign n48205 = pi17 ? n2954 : n48204;
  assign n48206 = pi16 ? n32 : n48205;
  assign n48207 = pi15 ? n24528 : n48206;
  assign n48208 = pi18 ? n863 : n34613;
  assign n48209 = pi17 ? n32 : n48208;
  assign n48210 = pi16 ? n32 : n48209;
  assign n48211 = pi17 ? n2954 : n25788;
  assign n48212 = pi16 ? n32 : n48211;
  assign n48213 = pi15 ? n48210 : n48212;
  assign n48214 = pi14 ? n48207 : n48213;
  assign n48215 = pi19 ? n4558 : ~n617;
  assign n48216 = pi18 ? n32 : n48215;
  assign n48217 = pi17 ? n32 : n48216;
  assign n48218 = pi16 ? n32 : n48217;
  assign n48219 = pi15 ? n48218 : n32;
  assign n48220 = pi14 ? n48219 : n32;
  assign n48221 = pi13 ? n48214 : n48220;
  assign n48222 = pi14 ? n22541 : n32;
  assign n48223 = pi13 ? n48222 : n32;
  assign n48224 = pi12 ? n48221 : n48223;
  assign n48225 = pi11 ? n48201 : n48224;
  assign n48226 = pi16 ? n3068 : ~n4729;
  assign n48227 = pi16 ? n3068 : ~n1683;
  assign n48228 = pi15 ? n48226 : n48227;
  assign n48229 = pi14 ? n32 : n48228;
  assign n48230 = pi13 ? n33386 : n48229;
  assign n48231 = pi18 ? n32 : n20007;
  assign n48232 = pi17 ? n32 : n48231;
  assign n48233 = pi16 ? n48232 : ~n1683;
  assign n48234 = pi20 ? n1817 : n321;
  assign n48235 = pi19 ? n32 : n48234;
  assign n48236 = pi18 ? n350 : ~n48235;
  assign n48237 = pi19 ? n4342 : n261;
  assign n48238 = pi18 ? n48237 : ~n32;
  assign n48239 = pi17 ? n48236 : ~n48238;
  assign n48240 = pi16 ? n32 : n48239;
  assign n48241 = pi15 ? n48233 : n48240;
  assign n48242 = pi19 ? n247 : n462;
  assign n48243 = pi18 ? n48242 : ~n8908;
  assign n48244 = pi17 ? n1215 : ~n48243;
  assign n48245 = pi16 ? n32 : n48244;
  assign n48246 = pi15 ? n48245 : n34658;
  assign n48247 = pi14 ? n48241 : n48246;
  assign n48248 = pi18 ? n32 : n41687;
  assign n48249 = pi17 ? n32 : n48248;
  assign n48250 = pi16 ? n48249 : ~n34661;
  assign n48251 = pi17 ? n1500 : ~n2517;
  assign n48252 = pi16 ? n32 : n48251;
  assign n48253 = pi15 ? n48250 : n48252;
  assign n48254 = pi18 ? n8975 : ~n32;
  assign n48255 = pi18 ? n19811 : n520;
  assign n48256 = pi17 ? n48254 : ~n48255;
  assign n48257 = pi16 ? n32 : n48256;
  assign n48258 = pi17 ? n32 : n36403;
  assign n48259 = pi19 ? n6173 : n236;
  assign n48260 = pi18 ? n48259 : ~n32;
  assign n48261 = pi18 ? n6059 : n323;
  assign n48262 = pi17 ? n48260 : ~n48261;
  assign n48263 = pi16 ? n48258 : n48262;
  assign n48264 = pi15 ? n48257 : n48263;
  assign n48265 = pi14 ? n48253 : n48264;
  assign n48266 = pi13 ? n48247 : n48265;
  assign n48267 = pi12 ? n48230 : n48266;
  assign n48268 = pi17 ? n16450 : n32208;
  assign n48269 = pi16 ? n32 : n48268;
  assign n48270 = pi19 ? n5694 : ~n32;
  assign n48271 = pi18 ? n48270 : ~n32;
  assign n48272 = pi17 ? n48271 : ~n2292;
  assign n48273 = pi16 ? n32 : n48272;
  assign n48274 = pi15 ? n48269 : n48273;
  assign n48275 = pi18 ? n32 : n20166;
  assign n48276 = pi17 ? n32 : n48275;
  assign n48277 = pi17 ? n1219 : ~n32217;
  assign n48278 = pi16 ? n48276 : ~n48277;
  assign n48279 = pi17 ? n1500 : ~n12775;
  assign n48280 = pi16 ? n16849 : ~n48279;
  assign n48281 = pi15 ? n48278 : n48280;
  assign n48282 = pi14 ? n48274 : n48281;
  assign n48283 = pi17 ? n1682 : ~n12775;
  assign n48284 = pi16 ? n32 : ~n48283;
  assign n48285 = pi17 ? n20200 : n34692;
  assign n48286 = pi16 ? n32 : ~n48285;
  assign n48287 = pi15 ? n48284 : n48286;
  assign n48288 = pi18 ? n13945 : n605;
  assign n48289 = pi17 ? n48271 : ~n48288;
  assign n48290 = pi16 ? n32 : n48289;
  assign n48291 = pi19 ? n17766 : ~n1757;
  assign n48292 = pi18 ? n48291 : ~n32;
  assign n48293 = pi17 ? n48292 : n34700;
  assign n48294 = pi16 ? n32 : n48293;
  assign n48295 = pi15 ? n48290 : n48294;
  assign n48296 = pi14 ? n48287 : n48295;
  assign n48297 = pi13 ? n48282 : n48296;
  assign n48298 = pi14 ? n34709 : n32;
  assign n48299 = pi19 ? n25120 : n32;
  assign n48300 = pi18 ? n4127 : n48299;
  assign n48301 = pi17 ? n32 : n48300;
  assign n48302 = pi16 ? n48301 : n32;
  assign n48303 = pi15 ? n48302 : n1015;
  assign n48304 = pi16 ? n1014 : n18083;
  assign n48305 = pi14 ? n48303 : n48304;
  assign n48306 = pi13 ? n48298 : n48305;
  assign n48307 = pi12 ? n48297 : n48306;
  assign n48308 = pi11 ? n48267 : n48307;
  assign n48309 = pi10 ? n48225 : n48308;
  assign n48310 = pi09 ? n48186 : n48309;
  assign n48311 = pi15 ? n22817 : n15655;
  assign n48312 = pi14 ? n48311 : n35393;
  assign n48313 = pi13 ? n23426 : n48312;
  assign n48314 = pi19 ? n236 : ~n236;
  assign n48315 = pi18 ? n32 : n48314;
  assign n48316 = pi17 ? n32 : n48315;
  assign n48317 = pi16 ? n32 : n48316;
  assign n48318 = pi15 ? n35393 : n48317;
  assign n48319 = pi14 ? n48318 : n48195;
  assign n48320 = pi14 ? n48197 : n15518;
  assign n48321 = pi13 ? n48319 : n48320;
  assign n48322 = pi12 ? n48313 : n48321;
  assign n48323 = pi15 ? n22923 : n48206;
  assign n48324 = pi14 ? n48323 : n48213;
  assign n48325 = pi15 ? n34616 : n32;
  assign n48326 = pi14 ? n48325 : n32;
  assign n48327 = pi13 ? n48324 : n48326;
  assign n48328 = pi15 ? n1109 : n22728;
  assign n48329 = pi14 ? n48328 : n32;
  assign n48330 = pi13 ? n48329 : n32;
  assign n48331 = pi12 ? n48327 : n48330;
  assign n48332 = pi11 ? n48322 : n48331;
  assign n48333 = pi18 ? n48242 : ~n13341;
  assign n48334 = pi17 ? n1215 : ~n48333;
  assign n48335 = pi16 ? n32 : n48334;
  assign n48336 = pi15 ? n48335 : n34759;
  assign n48337 = pi14 ? n48241 : n48336;
  assign n48338 = pi16 ? n48249 : ~n34762;
  assign n48339 = pi17 ? n1500 : ~n2748;
  assign n48340 = pi16 ? n32 : n48339;
  assign n48341 = pi15 ? n48338 : n48340;
  assign n48342 = pi18 ? n19811 : n2747;
  assign n48343 = pi17 ? n48254 : ~n48342;
  assign n48344 = pi16 ? n32 : n48343;
  assign n48345 = pi18 ? n6059 : n520;
  assign n48346 = pi17 ? n48260 : ~n48345;
  assign n48347 = pi16 ? n48258 : n48346;
  assign n48348 = pi15 ? n48344 : n48347;
  assign n48349 = pi14 ? n48341 : n48348;
  assign n48350 = pi13 ? n48337 : n48349;
  assign n48351 = pi12 ? n48230 : n48350;
  assign n48352 = pi17 ? n16450 : n11854;
  assign n48353 = pi16 ? n32 : n48352;
  assign n48354 = pi17 ? n48271 : ~n2408;
  assign n48355 = pi16 ? n32 : n48354;
  assign n48356 = pi15 ? n48353 : n48355;
  assign n48357 = pi17 ? n1500 : ~n34778;
  assign n48358 = pi16 ? n16849 : ~n48357;
  assign n48359 = pi15 ? n48278 : n48358;
  assign n48360 = pi14 ? n48356 : n48359;
  assign n48361 = pi17 ? n1682 : ~n34778;
  assign n48362 = pi16 ? n32 : ~n48361;
  assign n48363 = pi17 ? n20200 : n34783;
  assign n48364 = pi16 ? n32 : ~n48363;
  assign n48365 = pi15 ? n48362 : n48364;
  assign n48366 = pi14 ? n48365 : n48295;
  assign n48367 = pi13 ? n48360 : n48366;
  assign n48368 = pi14 ? n34789 : n32;
  assign n48369 = pi13 ? n48368 : n48305;
  assign n48370 = pi12 ? n48367 : n48369;
  assign n48371 = pi11 ? n48351 : n48370;
  assign n48372 = pi10 ? n48332 : n48371;
  assign n48373 = pi09 ? n48186 : n48372;
  assign n48374 = pi08 ? n48310 : n48373;
  assign n48375 = pi14 ? n32 : n16108;
  assign n48376 = pi13 ? n32 : n48375;
  assign n48377 = pi12 ? n32 : n48376;
  assign n48378 = pi11 ? n32 : n48377;
  assign n48379 = pi10 ? n32 : n48378;
  assign n48380 = pi18 ? n3496 : n6140;
  assign n48381 = pi17 ? n32 : n48380;
  assign n48382 = pi16 ? n32 : n48381;
  assign n48383 = pi15 ? n32 : n48382;
  assign n48384 = pi14 ? n23631 : n48383;
  assign n48385 = pi15 ? n32 : n23484;
  assign n48386 = pi19 ? n349 : n358;
  assign n48387 = pi18 ? n32 : n48386;
  assign n48388 = pi17 ? n32 : n48387;
  assign n48389 = pi16 ? n32 : n48388;
  assign n48390 = pi14 ? n48385 : n48389;
  assign n48391 = pi13 ? n48384 : n48390;
  assign n48392 = pi18 ? n23440 : n6132;
  assign n48393 = pi17 ? n32 : n48392;
  assign n48394 = pi16 ? n32 : n48393;
  assign n48395 = pi18 ? n359 : n48190;
  assign n48396 = pi17 ? n32 : n48395;
  assign n48397 = pi16 ? n32 : n48396;
  assign n48398 = pi15 ? n48394 : n48397;
  assign n48399 = pi19 ? n32 : n1331;
  assign n48400 = pi18 ? n32 : n48399;
  assign n48401 = pi20 ? n1611 : n246;
  assign n48402 = pi20 ? n333 : n342;
  assign n48403 = pi19 ? n48401 : n48402;
  assign n48404 = pi18 ? n48403 : ~n2615;
  assign n48405 = pi17 ? n48400 : n48404;
  assign n48406 = pi16 ? n32 : n48405;
  assign n48407 = pi19 ? n589 : ~n2614;
  assign n48408 = pi18 ? n32 : n48407;
  assign n48409 = pi17 ? n32 : n48408;
  assign n48410 = pi16 ? n32 : n48409;
  assign n48411 = pi15 ? n48406 : n48410;
  assign n48412 = pi14 ? n48398 : n48411;
  assign n48413 = pi15 ? n25790 : n13904;
  assign n48414 = pi15 ? n23160 : n23250;
  assign n48415 = pi14 ? n48413 : n48414;
  assign n48416 = pi13 ? n48412 : n48415;
  assign n48417 = pi12 ? n48391 : n48416;
  assign n48418 = pi19 ? n6018 : ~n2614;
  assign n48419 = pi18 ? n32 : n48418;
  assign n48420 = pi17 ? n32 : n48419;
  assign n48421 = pi16 ? n32 : n48420;
  assign n48422 = pi15 ? n34806 : n48421;
  assign n48423 = pi15 ? n23836 : n25840;
  assign n48424 = pi14 ? n48422 : n48423;
  assign n48425 = pi13 ? n48424 : n48326;
  assign n48426 = pi12 ? n48425 : n32;
  assign n48427 = pi11 ? n48417 : n48426;
  assign n48428 = pi18 ? n32 : n9461;
  assign n48429 = pi17 ? n32 : n48428;
  assign n48430 = pi18 ? n19082 : ~n32;
  assign n48431 = pi17 ? n32 : n48430;
  assign n48432 = pi16 ? n48429 : ~n48431;
  assign n48433 = pi15 ? n48226 : n48432;
  assign n48434 = pi14 ? n32 : n48433;
  assign n48435 = pi13 ? n22425 : n48434;
  assign n48436 = pi18 ? n237 : ~n4281;
  assign n48437 = pi18 ? n23363 : ~n32;
  assign n48438 = pi17 ? n48436 : ~n48437;
  assign n48439 = pi16 ? n32 : n48438;
  assign n48440 = pi20 ? n321 : n1324;
  assign n48441 = pi19 ? n32 : n48440;
  assign n48442 = pi18 ? n350 : ~n48441;
  assign n48443 = pi19 ? n16542 : n20006;
  assign n48444 = pi18 ? n48443 : ~n32;
  assign n48445 = pi17 ? n48442 : ~n48444;
  assign n48446 = pi16 ? n32 : n48445;
  assign n48447 = pi15 ? n48439 : n48446;
  assign n48448 = pi18 ? n13668 : n520;
  assign n48449 = pi17 ? n1215 : ~n48448;
  assign n48450 = pi16 ? n32 : n48449;
  assign n48451 = pi15 ? n48450 : n34865;
  assign n48452 = pi14 ? n48447 : n48451;
  assign n48453 = pi15 ? n48250 : n48340;
  assign n48454 = pi18 ? n13080 : n2747;
  assign n48455 = pi17 ? n1978 : ~n48454;
  assign n48456 = pi16 ? n32 : n48455;
  assign n48457 = pi18 ? n13080 : n24036;
  assign n48458 = pi17 ? n1978 : ~n48457;
  assign n48459 = pi16 ? n32 : n48458;
  assign n48460 = pi15 ? n48456 : n48459;
  assign n48461 = pi14 ? n48453 : n48460;
  assign n48462 = pi13 ? n48452 : n48461;
  assign n48463 = pi12 ? n48435 : n48462;
  assign n48464 = pi17 ? n16802 : n45939;
  assign n48465 = pi16 ? n32 : n48464;
  assign n48466 = pi15 ? n48465 : n48273;
  assign n48467 = pi17 ? n1219 : ~n34677;
  assign n48468 = pi16 ? n16396 : ~n48467;
  assign n48469 = pi15 ? n48468 : n48358;
  assign n48470 = pi14 ? n48466 : n48469;
  assign n48471 = pi16 ? n16836 : ~n48361;
  assign n48472 = pi19 ? n322 : n4342;
  assign n48473 = pi18 ? n48472 : n32;
  assign n48474 = pi17 ? n48473 : n34887;
  assign n48475 = pi16 ? n32 : ~n48474;
  assign n48476 = pi15 ? n48471 : n48475;
  assign n48477 = pi20 ? n339 : n342;
  assign n48478 = pi19 ? n48477 : n32;
  assign n48479 = pi18 ? n48478 : n32;
  assign n48480 = pi17 ? n48479 : n2292;
  assign n48481 = pi16 ? n16605 : ~n48480;
  assign n48482 = pi19 ? n1818 : n11546;
  assign n48483 = pi18 ? n48482 : ~n32;
  assign n48484 = pi17 ? n48483 : n34894;
  assign n48485 = pi16 ? n32 : n48484;
  assign n48486 = pi15 ? n48481 : n48485;
  assign n48487 = pi14 ? n48476 : n48486;
  assign n48488 = pi13 ? n48470 : n48487;
  assign n48489 = pi14 ? n34903 : n32;
  assign n48490 = pi20 ? n20396 : ~n765;
  assign n48491 = pi19 ? n32 : ~n48490;
  assign n48492 = pi18 ? n341 : ~n48491;
  assign n48493 = pi17 ? n32 : n48492;
  assign n48494 = pi20 ? n310 : ~n357;
  assign n48495 = pi20 ? n339 : ~n3523;
  assign n48496 = pi19 ? n48494 : n48495;
  assign n48497 = pi20 ? n785 : ~n1331;
  assign n48498 = pi19 ? n18256 : n48497;
  assign n48499 = pi18 ? n48496 : n48498;
  assign n48500 = pi20 ? n287 : ~n428;
  assign n48501 = pi19 ? n48500 : ~n358;
  assign n48502 = pi18 ? n48501 : ~n32;
  assign n48503 = pi17 ? n48499 : n48502;
  assign n48504 = pi16 ? n48493 : ~n48503;
  assign n48505 = pi15 ? n48504 : n130;
  assign n48506 = pi14 ? n48505 : n130;
  assign n48507 = pi13 ? n48489 : n48506;
  assign n48508 = pi12 ? n48488 : n48507;
  assign n48509 = pi11 ? n48463 : n48508;
  assign n48510 = pi10 ? n48427 : n48509;
  assign n48511 = pi09 ? n48379 : n48510;
  assign n48512 = pi14 ? n23741 : n48383;
  assign n48513 = pi19 ? n349 : n7502;
  assign n48514 = pi18 ? n32 : n48513;
  assign n48515 = pi17 ? n32 : n48514;
  assign n48516 = pi16 ? n32 : n48515;
  assign n48517 = pi14 ? n23750 : n48516;
  assign n48518 = pi13 ? n48512 : n48517;
  assign n48519 = pi18 ? n23440 : n37589;
  assign n48520 = pi17 ? n32 : n48519;
  assign n48521 = pi16 ? n32 : n48520;
  assign n48522 = pi15 ? n48521 : n48317;
  assign n48523 = pi18 ? n48403 : ~n697;
  assign n48524 = pi17 ? n32 : n48523;
  assign n48525 = pi16 ? n32 : n48524;
  assign n48526 = pi19 ? n32340 : ~n236;
  assign n48527 = pi18 ? n32 : n48526;
  assign n48528 = pi17 ? n32 : n48527;
  assign n48529 = pi16 ? n32 : n48528;
  assign n48530 = pi15 ? n48525 : n48529;
  assign n48531 = pi14 ? n48522 : n48530;
  assign n48532 = pi19 ? n343 : n358;
  assign n48533 = pi18 ? n32 : n48532;
  assign n48534 = pi17 ? n32 : n48533;
  assign n48535 = pi16 ? n32 : n48534;
  assign n48536 = pi15 ? n35393 : n48535;
  assign n48537 = pi14 ? n48536 : n15655;
  assign n48538 = pi13 ? n48531 : n48537;
  assign n48539 = pi12 ? n48518 : n48538;
  assign n48540 = pi19 ? n6018 : ~n617;
  assign n48541 = pi18 ? n32 : n48540;
  assign n48542 = pi17 ? n32 : n48541;
  assign n48543 = pi16 ? n32 : n48542;
  assign n48544 = pi15 ? n34950 : n48543;
  assign n48545 = pi19 ? n349 : n5626;
  assign n48546 = pi18 ? n32 : n48545;
  assign n48547 = pi17 ? n32 : n48546;
  assign n48548 = pi16 ? n32 : n48547;
  assign n48549 = pi15 ? n23836 : n48548;
  assign n48550 = pi14 ? n48544 : n48549;
  assign n48551 = pi13 ? n48550 : n48326;
  assign n48552 = pi12 ? n48551 : n32;
  assign n48553 = pi11 ? n48539 : n48552;
  assign n48554 = pi13 ? n32 : n48434;
  assign n48555 = pi18 ? n23363 : ~n645;
  assign n48556 = pi17 ? n48436 : ~n48555;
  assign n48557 = pi16 ? n32 : n48556;
  assign n48558 = pi18 ? n48443 : ~n645;
  assign n48559 = pi17 ? n48442 : ~n48558;
  assign n48560 = pi16 ? n32 : n48559;
  assign n48561 = pi15 ? n48557 : n48560;
  assign n48562 = pi18 ? n13668 : n508;
  assign n48563 = pi17 ? n1215 : ~n48562;
  assign n48564 = pi16 ? n32 : n48563;
  assign n48565 = pi15 ? n48564 : n5843;
  assign n48566 = pi14 ? n48561 : n48565;
  assign n48567 = pi17 ? n18482 : n2512;
  assign n48568 = pi16 ? n48249 : ~n48567;
  assign n48569 = pi17 ? n1500 : ~n2512;
  assign n48570 = pi16 ? n32 : n48569;
  assign n48571 = pi15 ? n48568 : n48570;
  assign n48572 = pi18 ? n13080 : n520;
  assign n48573 = pi17 ? n1978 : ~n48572;
  assign n48574 = pi16 ? n32 : n48573;
  assign n48575 = pi18 ? n13080 : n323;
  assign n48576 = pi17 ? n1978 : ~n48575;
  assign n48577 = pi16 ? n32 : n48576;
  assign n48578 = pi15 ? n48574 : n48577;
  assign n48579 = pi14 ? n48571 : n48578;
  assign n48580 = pi13 ? n48566 : n48579;
  assign n48581 = pi12 ? n48554 : n48580;
  assign n48582 = pi17 ? n48271 : ~n2519;
  assign n48583 = pi16 ? n32 : n48582;
  assign n48584 = pi15 ? n48465 : n48583;
  assign n48585 = pi17 ? n1219 : ~n32826;
  assign n48586 = pi16 ? n16396 : ~n48585;
  assign n48587 = pi17 ? n1500 : ~n12771;
  assign n48588 = pi16 ? n16849 : ~n48587;
  assign n48589 = pi15 ? n48586 : n48588;
  assign n48590 = pi14 ? n48584 : n48589;
  assign n48591 = pi16 ? n16836 : ~n48283;
  assign n48592 = pi17 ? n48473 : n34997;
  assign n48593 = pi16 ? n32 : ~n48592;
  assign n48594 = pi15 ? n48591 : n48593;
  assign n48595 = pi19 ? n1818 : n429;
  assign n48596 = pi18 ? n48595 : ~n32;
  assign n48597 = pi17 ? n48596 : n35001;
  assign n48598 = pi16 ? n32 : n48597;
  assign n48599 = pi15 ? n48481 : n48598;
  assign n48600 = pi14 ? n48594 : n48599;
  assign n48601 = pi13 ? n48590 : n48600;
  assign n48602 = pi18 ? n341 : ~n28927;
  assign n48603 = pi17 ? n32 : n48602;
  assign n48604 = pi19 ? n34921 : n236;
  assign n48605 = pi18 ? n48604 : ~n32;
  assign n48606 = pi17 ? n34920 : n48605;
  assign n48607 = pi16 ? n48603 : ~n48606;
  assign n48608 = pi15 ? n48607 : n130;
  assign n48609 = pi14 ? n48608 : n32;
  assign n48610 = pi13 ? n48489 : n48609;
  assign n48611 = pi12 ? n48601 : n48610;
  assign n48612 = pi11 ? n48581 : n48611;
  assign n48613 = pi10 ? n48553 : n48612;
  assign n48614 = pi09 ? n48379 : n48613;
  assign n48615 = pi08 ? n48511 : n48614;
  assign n48616 = pi07 ? n48374 : n48615;
  assign n48617 = pi06 ? n48180 : n48616;
  assign n48618 = pi14 ? n32 : n23574;
  assign n48619 = pi13 ? n32 : n48618;
  assign n48620 = pi12 ? n32 : n48619;
  assign n48621 = pi11 ? n32 : n48620;
  assign n48622 = pi10 ? n32 : n48621;
  assign n48623 = pi19 ? n29103 : n358;
  assign n48624 = pi18 ? n16449 : n48623;
  assign n48625 = pi17 ? n32 : n48624;
  assign n48626 = pi16 ? n32 : n48625;
  assign n48627 = pi15 ? n32 : n48626;
  assign n48628 = pi14 ? n23576 : n48627;
  assign n48629 = pi15 ? n23250 : n25466;
  assign n48630 = pi19 ? n246 : ~n343;
  assign n48631 = pi18 ? n48630 : n37589;
  assign n48632 = pi17 ? n32 : n48631;
  assign n48633 = pi16 ? n32 : n48632;
  assign n48634 = pi19 ? n236 : ~n1941;
  assign n48635 = pi18 ? n31093 : n48634;
  assign n48636 = pi17 ? n36573 : n48635;
  assign n48637 = pi16 ? n32 : n48636;
  assign n48638 = pi15 ? n48633 : n48637;
  assign n48639 = pi14 ? n48629 : n48638;
  assign n48640 = pi13 ? n48628 : n48639;
  assign n48641 = pi19 ? n322 : ~n288;
  assign n48642 = pi18 ? n48641 : n37589;
  assign n48643 = pi17 ? n32 : n48642;
  assign n48644 = pi16 ? n32 : n48643;
  assign n48645 = pi18 ? n20172 : n6132;
  assign n48646 = pi17 ? n32 : n48645;
  assign n48647 = pi16 ? n32 : n48646;
  assign n48648 = pi15 ? n48644 : n48647;
  assign n48649 = pi19 ? n813 : ~n236;
  assign n48650 = pi18 ? n20172 : n48649;
  assign n48651 = pi17 ? n32 : n48650;
  assign n48652 = pi16 ? n32 : n48651;
  assign n48653 = pi15 ? n48652 : n35452;
  assign n48654 = pi14 ? n48648 : n48653;
  assign n48655 = pi15 ? n13904 : n14156;
  assign n48656 = pi15 ? n23484 : n35023;
  assign n48657 = pi14 ? n48655 : n48656;
  assign n48658 = pi13 ? n48654 : n48657;
  assign n48659 = pi12 ? n48640 : n48658;
  assign n48660 = pi19 ? n18665 : n5614;
  assign n48661 = pi19 ? n6173 : ~n236;
  assign n48662 = pi18 ? n48660 : n48661;
  assign n48663 = pi17 ? n48400 : n48662;
  assign n48664 = pi16 ? n32 : n48663;
  assign n48665 = pi15 ? n35393 : n48664;
  assign n48666 = pi19 ? n207 : ~n236;
  assign n48667 = pi18 ? n32 : n48666;
  assign n48668 = pi17 ? n32 : n48667;
  assign n48669 = pi16 ? n32 : n48668;
  assign n48670 = pi19 ? n16542 : ~n236;
  assign n48671 = pi18 ? n32 : n48670;
  assign n48672 = pi17 ? n32 : n48671;
  assign n48673 = pi16 ? n32 : n48672;
  assign n48674 = pi15 ? n48669 : n48673;
  assign n48675 = pi14 ? n48665 : n48674;
  assign n48676 = pi14 ? n21558 : n32;
  assign n48677 = pi13 ? n48675 : n48676;
  assign n48678 = pi14 ? n24327 : n32;
  assign n48679 = pi14 ? n1110 : n32;
  assign n48680 = pi13 ? n48678 : n48679;
  assign n48681 = pi12 ? n48677 : n48680;
  assign n48682 = pi11 ? n48659 : n48681;
  assign n48683 = pi15 ? n15123 : n39582;
  assign n48684 = pi17 ? n18482 : n1580;
  assign n48685 = pi16 ? n32 : ~n48684;
  assign n48686 = pi17 ? n1227 : ~n28029;
  assign n48687 = pi16 ? n17486 : n48686;
  assign n48688 = pi15 ? n48685 : n48687;
  assign n48689 = pi14 ? n48683 : n48688;
  assign n48690 = pi13 ? n32 : n48689;
  assign n48691 = pi18 ? n4380 : n24344;
  assign n48692 = pi17 ? n4429 : ~n48691;
  assign n48693 = pi16 ? n32 : n48692;
  assign n48694 = pi18 ? n880 : ~n19202;
  assign n48695 = pi19 ? n23895 : ~n349;
  assign n48696 = pi18 ? n48695 : n2627;
  assign n48697 = pi17 ? n48694 : ~n48696;
  assign n48698 = pi16 ? n32 : n48697;
  assign n48699 = pi15 ? n48693 : n48698;
  assign n48700 = pi18 ? n35082 : ~n18882;
  assign n48701 = pi17 ? n48700 : ~n2628;
  assign n48702 = pi16 ? n32 : n48701;
  assign n48703 = pi15 ? n48702 : n35090;
  assign n48704 = pi14 ? n48699 : n48703;
  assign n48705 = pi19 ? n32 : n5675;
  assign n48706 = pi18 ? n32 : n48705;
  assign n48707 = pi17 ? n32 : n48706;
  assign n48708 = pi17 ? n18482 : n2628;
  assign n48709 = pi16 ? n48707 : ~n48708;
  assign n48710 = pi15 ? n48709 : n35095;
  assign n48711 = pi19 ? n9037 : n349;
  assign n48712 = pi18 ? n32 : n48711;
  assign n48713 = pi18 ? n13940 : n520;
  assign n48714 = pi17 ? n48712 : ~n48713;
  assign n48715 = pi16 ? n32 : n48714;
  assign n48716 = pi19 ? n13939 : n247;
  assign n48717 = pi18 ? n48716 : n520;
  assign n48718 = pi17 ? n48712 : ~n48717;
  assign n48719 = pi16 ? n32 : n48718;
  assign n48720 = pi15 ? n48715 : n48719;
  assign n48721 = pi14 ? n48710 : n48720;
  assign n48722 = pi13 ? n48704 : n48721;
  assign n48723 = pi12 ? n48690 : n48722;
  assign n48724 = pi17 ? n17346 : n32826;
  assign n48725 = pi16 ? n32 : n48724;
  assign n48726 = pi18 ? n32 : n34283;
  assign n48727 = pi18 ? n20164 : n323;
  assign n48728 = pi17 ? n48726 : ~n48727;
  assign n48729 = pi16 ? n32 : n48728;
  assign n48730 = pi15 ? n48725 : n48729;
  assign n48731 = pi18 ? n20164 : n532;
  assign n48732 = pi19 ? n321 : ~n349;
  assign n48733 = pi18 ? n48732 : n35111;
  assign n48734 = pi17 ? n48731 : ~n48733;
  assign n48735 = pi16 ? n3165 : ~n48734;
  assign n48736 = pi19 ? n4982 : ~n32;
  assign n48737 = pi18 ? n5657 : n48736;
  assign n48738 = pi19 ? n5004 : ~n6158;
  assign n48739 = pi18 ? n48738 : ~n323;
  assign n48740 = pi17 ? n48737 : ~n48739;
  assign n48741 = pi16 ? n3165 : ~n48740;
  assign n48742 = pi15 ? n48735 : n48741;
  assign n48743 = pi14 ? n48730 : n48742;
  assign n48744 = pi18 ? n46739 : n323;
  assign n48745 = pi17 ? n32 : n48744;
  assign n48746 = pi16 ? n1471 : ~n48745;
  assign n48747 = pi16 ? n1214 : ~n3769;
  assign n48748 = pi15 ? n48746 : n48747;
  assign n48749 = pi20 ? n287 : ~n220;
  assign n48750 = pi19 ? n246 : ~n48749;
  assign n48751 = pi18 ? n48750 : ~n5749;
  assign n48752 = pi17 ? n48751 : ~n2519;
  assign n48753 = pi16 ? n17434 : n48752;
  assign n48754 = pi15 ? n48753 : n35138;
  assign n48755 = pi14 ? n48748 : n48754;
  assign n48756 = pi13 ? n48743 : n48755;
  assign n48757 = pi15 ? n369 : n130;
  assign n48758 = pi14 ? n48757 : n130;
  assign n48759 = pi13 ? n32 : n48758;
  assign n48760 = pi12 ? n48756 : n48759;
  assign n48761 = pi11 ? n48723 : n48760;
  assign n48762 = pi10 ? n48682 : n48761;
  assign n48763 = pi09 ? n48622 : n48762;
  assign n48764 = pi15 ? n23250 : n25598;
  assign n48765 = pi18 ? n48630 : n24310;
  assign n48766 = pi17 ? n32 : n48765;
  assign n48767 = pi16 ? n32 : n48766;
  assign n48768 = pi19 ? n236 : ~n813;
  assign n48769 = pi18 ? n31093 : n48768;
  assign n48770 = pi17 ? n36573 : n48769;
  assign n48771 = pi16 ? n32 : n48770;
  assign n48772 = pi15 ? n48767 : n48771;
  assign n48773 = pi14 ? n48764 : n48772;
  assign n48774 = pi13 ? n48628 : n48773;
  assign n48775 = pi18 ? n48641 : n24310;
  assign n48776 = pi17 ? n32 : n48775;
  assign n48777 = pi16 ? n32 : n48776;
  assign n48778 = pi18 ? n20172 : n37589;
  assign n48779 = pi17 ? n32 : n48778;
  assign n48780 = pi16 ? n32 : n48779;
  assign n48781 = pi15 ? n48777 : n48780;
  assign n48782 = pi14 ? n48781 : n48653;
  assign n48783 = pi14 ? n48655 : n35177;
  assign n48784 = pi13 ? n48782 : n48783;
  assign n48785 = pi12 ? n48774 : n48784;
  assign n48786 = pi17 ? n32 : n48662;
  assign n48787 = pi16 ? n32 : n48786;
  assign n48788 = pi15 ? n35393 : n48787;
  assign n48789 = pi18 ? n32 : n31850;
  assign n48790 = pi17 ? n32 : n48789;
  assign n48791 = pi16 ? n32 : n48790;
  assign n48792 = pi15 ? n48669 : n48791;
  assign n48793 = pi14 ? n48788 : n48792;
  assign n48794 = pi13 ? n48793 : n48676;
  assign n48795 = pi15 ? n23160 : n22923;
  assign n48796 = pi14 ? n48795 : n32;
  assign n48797 = pi13 ? n48796 : n32;
  assign n48798 = pi12 ? n48794 : n48797;
  assign n48799 = pi11 ? n48785 : n48798;
  assign n48800 = pi15 ? n32 : n21853;
  assign n48801 = pi14 ? n48800 : n48688;
  assign n48802 = pi13 ? n1111 : n48801;
  assign n48803 = pi17 ? n48700 : ~n2512;
  assign n48804 = pi16 ? n32 : n48803;
  assign n48805 = pi15 ? n48804 : n35090;
  assign n48806 = pi14 ? n48699 : n48805;
  assign n48807 = pi16 ? n48707 : ~n48567;
  assign n48808 = pi15 ? n48807 : n35095;
  assign n48809 = pi14 ? n48808 : n48720;
  assign n48810 = pi13 ? n48806 : n48809;
  assign n48811 = pi12 ? n48802 : n48810;
  assign n48812 = pi18 ? n48738 : ~n2754;
  assign n48813 = pi17 ? n48737 : ~n48812;
  assign n48814 = pi16 ? n3165 : ~n48813;
  assign n48815 = pi15 ? n48735 : n48814;
  assign n48816 = pi14 ? n48730 : n48815;
  assign n48817 = pi13 ? n48816 : n48755;
  assign n48818 = pi12 ? n48817 : n48759;
  assign n48819 = pi11 ? n48811 : n48818;
  assign n48820 = pi10 ? n48799 : n48819;
  assign n48821 = pi09 ? n48622 : n48820;
  assign n48822 = pi08 ? n48763 : n48821;
  assign n48823 = pi14 ? n32 : n23725;
  assign n48824 = pi13 ? n32 : n48823;
  assign n48825 = pi12 ? n32 : n48824;
  assign n48826 = pi11 ? n32 : n48825;
  assign n48827 = pi10 ? n32 : n48826;
  assign n48828 = pi15 ? n24905 : n23569;
  assign n48829 = pi14 ? n48828 : n32;
  assign n48830 = pi15 ? n32 : n25598;
  assign n48831 = pi18 ? n32 : ~n24310;
  assign n48832 = pi17 ? n2736 : ~n48831;
  assign n48833 = pi16 ? n32 : n48832;
  assign n48834 = pi18 ? n32 : n22526;
  assign n48835 = pi18 ? n32 : ~n48768;
  assign n48836 = pi17 ? n48834 : ~n48835;
  assign n48837 = pi16 ? n32 : n48836;
  assign n48838 = pi15 ? n48833 : n48837;
  assign n48839 = pi14 ? n48830 : n48838;
  assign n48840 = pi13 ? n48829 : n48839;
  assign n48841 = pi19 ? n208 : ~n4721;
  assign n48842 = pi18 ? n48841 : n24310;
  assign n48843 = pi17 ? n32 : n48842;
  assign n48844 = pi16 ? n32 : n48843;
  assign n48845 = pi19 ? n24055 : n11027;
  assign n48846 = pi19 ? n617 : ~n236;
  assign n48847 = pi18 ? n48845 : ~n48846;
  assign n48848 = pi17 ? n32 : ~n48847;
  assign n48849 = pi16 ? n32 : n48848;
  assign n48850 = pi15 ? n48844 : n48849;
  assign n48851 = pi18 ? n24697 : n48314;
  assign n48852 = pi17 ? n32 : n48851;
  assign n48853 = pi16 ? n32 : n48852;
  assign n48854 = pi15 ? n48853 : n35452;
  assign n48855 = pi14 ? n48850 : n48854;
  assign n48856 = pi15 ? n13904 : n14397;
  assign n48857 = pi14 ? n48856 : n35226;
  assign n48858 = pi13 ? n48855 : n48857;
  assign n48859 = pi12 ? n48840 : n48858;
  assign n48860 = pi18 ? n936 : n37589;
  assign n48861 = pi17 ? n32 : n48860;
  assign n48862 = pi16 ? n32 : n48861;
  assign n48863 = pi19 ? n1464 : n594;
  assign n48864 = pi19 ? n6173 : ~n1941;
  assign n48865 = pi18 ? n48863 : n48864;
  assign n48866 = pi17 ? n32 : n48865;
  assign n48867 = pi16 ? n32 : n48866;
  assign n48868 = pi15 ? n48862 : n48867;
  assign n48869 = pi18 ? n6145 : n37589;
  assign n48870 = pi17 ? n32 : n48869;
  assign n48871 = pi16 ? n32 : n48870;
  assign n48872 = pi15 ? n48871 : n23250;
  assign n48873 = pi14 ? n48868 : n48872;
  assign n48874 = pi13 ? n48873 : n32;
  assign n48875 = pi14 ? n32 : n22540;
  assign n48876 = pi13 ? n48875 : n32;
  assign n48877 = pi12 ? n48874 : n48876;
  assign n48878 = pi11 ? n48859 : n48877;
  assign n48879 = pi18 ? n23660 : ~n618;
  assign n48880 = pi17 ? n1219 : n48879;
  assign n48881 = pi16 ? n32 : n48880;
  assign n48882 = pi15 ? n48685 : n48881;
  assign n48883 = pi14 ? n32 : n48882;
  assign n48884 = pi13 ? n32 : n48883;
  assign n48885 = pi18 ? n9346 : ~n32;
  assign n48886 = pi20 ? n749 : ~n274;
  assign n48887 = pi19 ? n48886 : ~n32;
  assign n48888 = pi18 ? n32 : n48887;
  assign n48889 = pi17 ? n48885 : ~n48888;
  assign n48890 = pi16 ? n32 : n48889;
  assign n48891 = pi18 ? n880 : ~n22885;
  assign n48892 = pi19 ? n11879 : ~n236;
  assign n48893 = pi18 ? n48892 : n595;
  assign n48894 = pi17 ? n48891 : ~n48893;
  assign n48895 = pi16 ? n32 : n48894;
  assign n48896 = pi15 ? n48890 : n48895;
  assign n48897 = pi18 ? n4380 : ~n4343;
  assign n48898 = pi18 ? n20912 : n595;
  assign n48899 = pi17 ? n48897 : ~n48898;
  assign n48900 = pi16 ? n32 : n48899;
  assign n48901 = pi15 ? n48900 : n35294;
  assign n48902 = pi14 ? n48896 : n48901;
  assign n48903 = pi18 ? n36192 : n289;
  assign n48904 = pi17 ? n48903 : ~n2618;
  assign n48905 = pi16 ? n3283 : n48904;
  assign n48906 = pi17 ? n1978 : ~n2512;
  assign n48907 = pi16 ? n32 : n48906;
  assign n48908 = pi15 ? n48905 : n48907;
  assign n48909 = pi18 ? n4983 : n508;
  assign n48910 = pi17 ? n35304 : ~n48909;
  assign n48911 = pi16 ? n32 : n48910;
  assign n48912 = pi19 ? n4982 : n247;
  assign n48913 = pi18 ? n48912 : n520;
  assign n48914 = pi17 ? n8859 : ~n48913;
  assign n48915 = pi16 ? n32 : n48914;
  assign n48916 = pi15 ? n48911 : n48915;
  assign n48917 = pi14 ? n48908 : n48916;
  assign n48918 = pi13 ? n48902 : n48917;
  assign n48919 = pi12 ? n48884 : n48918;
  assign n48920 = pi17 ? n23052 : n32826;
  assign n48921 = pi16 ? n32 : n48920;
  assign n48922 = pi15 ? n48921 : n48729;
  assign n48923 = pi18 ? n48732 : ~n34229;
  assign n48924 = pi17 ? n48731 : ~n48923;
  assign n48925 = pi16 ? n3165 : ~n48924;
  assign n48926 = pi19 ? n9007 : ~n1757;
  assign n48927 = pi18 ? n32 : n48926;
  assign n48928 = pi19 ? n47800 : n343;
  assign n48929 = pi18 ? n48928 : n2754;
  assign n48930 = pi17 ? n48927 : n48929;
  assign n48931 = pi16 ? n3165 : ~n48930;
  assign n48932 = pi15 ? n48925 : n48931;
  assign n48933 = pi14 ? n48922 : n48932;
  assign n48934 = pi18 ? n46739 : n2754;
  assign n48935 = pi17 ? n32 : n48934;
  assign n48936 = pi16 ? n1471 : ~n48935;
  assign n48937 = pi18 ? n20020 : n2754;
  assign n48938 = pi17 ? n19886 : n48937;
  assign n48939 = pi16 ? n1214 : ~n48938;
  assign n48940 = pi15 ? n48936 : n48939;
  assign n48941 = pi20 ? n246 : n12884;
  assign n48942 = pi20 ? n17669 : n1324;
  assign n48943 = pi19 ? n48941 : n48942;
  assign n48944 = pi20 ? n310 : ~n1091;
  assign n48945 = pi19 ? n48944 : ~n32;
  assign n48946 = pi18 ? n48943 : n48945;
  assign n48947 = pi18 ? n22554 : n2754;
  assign n48948 = pi17 ? n48946 : ~n48947;
  assign n48949 = pi16 ? n32 : n48948;
  assign n48950 = pi18 ? n24540 : n323;
  assign n48951 = pi17 ? n2512 : ~n48950;
  assign n48952 = pi16 ? n465 : n48951;
  assign n48953 = pi15 ? n48949 : n48952;
  assign n48954 = pi14 ? n48940 : n48953;
  assign n48955 = pi13 ? n48933 : n48954;
  assign n48956 = pi21 ? n124 : ~n259;
  assign n48957 = pi20 ? n32 : n48956;
  assign n48958 = pi19 ? n32 : n48957;
  assign n48959 = pi18 ? n48958 : n32;
  assign n48960 = pi17 ? n32 : n48959;
  assign n48961 = pi16 ? n48960 : n32;
  assign n48962 = pi15 ? n48961 : n13952;
  assign n48963 = pi14 ? n370 : n48962;
  assign n48964 = pi13 ? n924 : n48963;
  assign n48965 = pi12 ? n48955 : n48964;
  assign n48966 = pi11 ? n48919 : n48965;
  assign n48967 = pi10 ? n48878 : n48966;
  assign n48968 = pi09 ? n48827 : n48967;
  assign n48969 = pi15 ? n23730 : n23574;
  assign n48970 = pi14 ? n48969 : n32;
  assign n48971 = pi15 ? n32 : n37197;
  assign n48972 = pi19 ? n349 : ~n1812;
  assign n48973 = pi18 ? n32 : ~n48972;
  assign n48974 = pi17 ? n2736 : ~n48973;
  assign n48975 = pi16 ? n32 : n48974;
  assign n48976 = pi19 ? n236 : ~n1812;
  assign n48977 = pi18 ? n32 : ~n48976;
  assign n48978 = pi17 ? n48834 : ~n48977;
  assign n48979 = pi16 ? n32 : n48978;
  assign n48980 = pi15 ? n48975 : n48979;
  assign n48981 = pi14 ? n48971 : n48980;
  assign n48982 = pi13 ? n48970 : n48981;
  assign n48983 = pi18 ? n48841 : n48972;
  assign n48984 = pi17 ? n32 : n48983;
  assign n48985 = pi16 ? n32 : n48984;
  assign n48986 = pi19 ? n617 : ~n813;
  assign n48987 = pi18 ? n48845 : ~n48986;
  assign n48988 = pi17 ? n32 : ~n48987;
  assign n48989 = pi16 ? n32 : n48988;
  assign n48990 = pi15 ? n48985 : n48989;
  assign n48991 = pi14 ? n48990 : n48854;
  assign n48992 = pi14 ? n48856 : n35384;
  assign n48993 = pi13 ? n48991 : n48992;
  assign n48994 = pi12 ? n48982 : n48993;
  assign n48995 = pi18 ? n936 : n6132;
  assign n48996 = pi17 ? n32 : n48995;
  assign n48997 = pi16 ? n32 : n48996;
  assign n48998 = pi15 ? n48997 : n48867;
  assign n48999 = pi22 ? n34 : n50;
  assign n49000 = pi21 ? n48999 : ~n32;
  assign n49001 = pi20 ? n49000 : ~n32;
  assign n49002 = pi19 ? n349 : ~n49001;
  assign n49003 = pi18 ? n6145 : n49002;
  assign n49004 = pi17 ? n32 : n49003;
  assign n49005 = pi16 ? n32 : n49004;
  assign n49006 = pi15 ? n49005 : n32;
  assign n49007 = pi14 ? n48998 : n49006;
  assign n49008 = pi14 ? n32 : n23326;
  assign n49009 = pi13 ? n49007 : n49008;
  assign n49010 = pi14 ? n23326 : n22540;
  assign n49011 = pi13 ? n49010 : n32;
  assign n49012 = pi12 ? n49009 : n49011;
  assign n49013 = pi11 ? n48994 : n49012;
  assign n49014 = pi20 ? n8943 : ~n20507;
  assign n49015 = pi19 ? n49014 : ~n32;
  assign n49016 = pi18 ? n32 : n49015;
  assign n49017 = pi17 ? n48885 : ~n49016;
  assign n49018 = pi16 ? n32 : n49017;
  assign n49019 = pi15 ? n49018 : n48895;
  assign n49020 = pi14 ? n49019 : n48901;
  assign n49021 = pi13 ? n49020 : n48917;
  assign n49022 = pi12 ? n48884 : n49021;
  assign n49023 = pi17 ? n23052 : n12287;
  assign n49024 = pi16 ? n32 : n49023;
  assign n49025 = pi18 ? n20164 : n520;
  assign n49026 = pi17 ? n48726 : ~n49025;
  assign n49027 = pi16 ? n32 : n49026;
  assign n49028 = pi15 ? n49024 : n49027;
  assign n49029 = pi14 ? n49028 : n48932;
  assign n49030 = pi19 ? n246 : n1324;
  assign n49031 = pi20 ? n310 : ~n13171;
  assign n49032 = pi19 ? n49031 : ~n32;
  assign n49033 = pi18 ? n49030 : n49032;
  assign n49034 = pi17 ? n49033 : ~n35424;
  assign n49035 = pi16 ? n32 : n49034;
  assign n49036 = pi15 ? n49035 : n48952;
  assign n49037 = pi14 ? n48940 : n49036;
  assign n49038 = pi13 ? n49029 : n49037;
  assign n49039 = pi16 ? n129 : n13951;
  assign n49040 = pi15 ? n48961 : n49039;
  assign n49041 = pi14 ? n48757 : n49040;
  assign n49042 = pi13 ? n924 : n49041;
  assign n49043 = pi12 ? n49038 : n49042;
  assign n49044 = pi11 ? n49022 : n49043;
  assign n49045 = pi10 ? n49013 : n49044;
  assign n49046 = pi09 ? n48827 : n49045;
  assign n49047 = pi08 ? n48968 : n49046;
  assign n49048 = pi07 ? n48822 : n49047;
  assign n49049 = pi13 ? n32 : n36873;
  assign n49050 = pi12 ? n32 : n49049;
  assign n49051 = pi11 ? n32 : n49050;
  assign n49052 = pi10 ? n32 : n49051;
  assign n49053 = pi17 ? n1682 : ~n4245;
  assign n49054 = pi16 ? n32 : n49053;
  assign n49055 = pi15 ? n24742 : n49054;
  assign n49056 = pi19 ? n358 : n1812;
  assign n49057 = pi18 ? n32 : n49056;
  assign n49058 = pi17 ? n2519 : ~n49057;
  assign n49059 = pi16 ? n32 : n49058;
  assign n49060 = pi19 ? n32 : ~n18678;
  assign n49061 = pi18 ? n49060 : ~n32;
  assign n49062 = pi17 ? n49061 : ~n4245;
  assign n49063 = pi16 ? n32 : n49062;
  assign n49064 = pi15 ? n49059 : n49063;
  assign n49065 = pi14 ? n49055 : n49064;
  assign n49066 = pi13 ? n16322 : n49065;
  assign n49067 = pi19 ? n322 : n22525;
  assign n49068 = pi18 ? n32 : n49067;
  assign n49069 = pi17 ? n49068 : ~n48977;
  assign n49070 = pi16 ? n32 : n49069;
  assign n49071 = pi18 ? n32 : n8956;
  assign n49072 = pi17 ? n49071 : ~n48835;
  assign n49073 = pi16 ? n32 : n49072;
  assign n49074 = pi15 ? n49070 : n49073;
  assign n49075 = pi19 ? n813 : n5614;
  assign n49076 = pi18 ? n5657 : n49075;
  assign n49077 = pi17 ? n32 : n49076;
  assign n49078 = pi16 ? n32 : n49077;
  assign n49079 = pi19 ? n531 : n5614;
  assign n49080 = pi18 ? n32 : n49079;
  assign n49081 = pi17 ? n32 : n49080;
  assign n49082 = pi16 ? n32 : n49081;
  assign n49083 = pi15 ? n49078 : n49082;
  assign n49084 = pi14 ? n49074 : n49083;
  assign n49085 = pi15 ? n14138 : n32;
  assign n49086 = pi15 ? n25657 : n14339;
  assign n49087 = pi14 ? n49085 : n49086;
  assign n49088 = pi13 ? n49084 : n49087;
  assign n49089 = pi12 ? n49066 : n49088;
  assign n49090 = pi20 ? n246 : ~n1331;
  assign n49091 = pi20 ? n342 : n518;
  assign n49092 = pi19 ? n49090 : ~n49091;
  assign n49093 = pi18 ? n49092 : ~n962;
  assign n49094 = pi17 ? n35241 : n49093;
  assign n49095 = pi16 ? n32 : n49094;
  assign n49096 = pi17 ? n34522 : ~n2724;
  assign n49097 = pi16 ? n32 : n49096;
  assign n49098 = pi15 ? n49095 : n49097;
  assign n49099 = pi20 ? n3523 : ~n6621;
  assign n49100 = pi19 ? n49099 : n5614;
  assign n49101 = pi18 ? n6118 : n49100;
  assign n49102 = pi17 ? n32 : n49101;
  assign n49103 = pi16 ? n32 : n49102;
  assign n49104 = pi15 ? n49103 : n32;
  assign n49105 = pi14 ? n49098 : n49104;
  assign n49106 = pi13 ? n49105 : n32;
  assign n49107 = pi12 ? n49106 : n47581;
  assign n49108 = pi11 ? n49089 : n49107;
  assign n49109 = pi17 ? n2519 : ~n1682;
  assign n49110 = pi16 ? n32 : n49109;
  assign n49111 = pi15 ? n32 : n49110;
  assign n49112 = pi17 ? n1500 : ~n36008;
  assign n49113 = pi16 ? n32 : n49112;
  assign n49114 = pi17 ? n1028 : ~n48166;
  assign n49115 = pi16 ? n17120 : n49114;
  assign n49116 = pi15 ? n49113 : n49115;
  assign n49117 = pi14 ? n49111 : n49116;
  assign n49118 = pi13 ? n22926 : n49117;
  assign n49119 = pi17 ? n1697 : ~n4099;
  assign n49120 = pi16 ? n32 : n49119;
  assign n49121 = pi17 ? n31444 : ~n4099;
  assign n49122 = pi16 ? n32 : n49121;
  assign n49123 = pi15 ? n49120 : n49122;
  assign n49124 = pi17 ? n1215 : ~n4099;
  assign n49125 = pi16 ? n32 : n49124;
  assign n49126 = pi19 ? n462 : n3775;
  assign n49127 = pi18 ? n49126 : ~n32;
  assign n49128 = pi17 ? n49127 : ~n4099;
  assign n49129 = pi16 ? n32 : n49128;
  assign n49130 = pi15 ? n49125 : n49129;
  assign n49131 = pi14 ? n49123 : n49130;
  assign n49132 = pi17 ? n1580 : ~n2618;
  assign n49133 = pi16 ? n32 : n49132;
  assign n49134 = pi17 ? n2325 : ~n2512;
  assign n49135 = pi16 ? n32 : n49134;
  assign n49136 = pi15 ? n49133 : n49135;
  assign n49137 = pi18 ? n6384 : n508;
  assign n49138 = pi17 ? n2959 : ~n49137;
  assign n49139 = pi16 ? n32 : n49138;
  assign n49140 = pi19 ? n236 : ~n33150;
  assign n49141 = pi18 ? n49140 : n35545;
  assign n49142 = pi17 ? n32 : ~n49141;
  assign n49143 = pi16 ? n32 : n49142;
  assign n49144 = pi15 ? n49139 : n49143;
  assign n49145 = pi14 ? n49136 : n49144;
  assign n49146 = pi13 ? n49131 : n49145;
  assign n49147 = pi12 ? n49118 : n49146;
  assign n49148 = pi18 ? n237 : n323;
  assign n49149 = pi17 ? n32 : ~n49148;
  assign n49150 = pi16 ? n337 : n49149;
  assign n49151 = pi18 ? n6163 : n35545;
  assign n49152 = pi17 ? n3164 : ~n49151;
  assign n49153 = pi16 ? n32 : n49152;
  assign n49154 = pi15 ? n49150 : n49153;
  assign n49155 = pi16 ? n2860 : ~n2518;
  assign n49156 = pi17 ? n32 : n5779;
  assign n49157 = pi16 ? n49156 : ~n2518;
  assign n49158 = pi15 ? n49155 : n49157;
  assign n49159 = pi14 ? n49154 : n49158;
  assign n49160 = pi19 ? n22525 : ~n32;
  assign n49161 = pi18 ? n32 : n49160;
  assign n49162 = pi17 ? n32 : n49161;
  assign n49163 = pi16 ? n49162 : ~n2518;
  assign n49164 = pi18 ? n276 : n5372;
  assign n49165 = pi17 ? n32 : n49164;
  assign n49166 = pi16 ? n49165 : ~n2518;
  assign n49167 = pi15 ? n49163 : n49166;
  assign n49168 = pi19 ? n9037 : ~n236;
  assign n49169 = pi18 ? n49168 : n350;
  assign n49170 = pi17 ? n7039 : ~n49169;
  assign n49171 = pi16 ? n32 : n49170;
  assign n49172 = pi20 ? n32 : n309;
  assign n49173 = pi19 ? n32 : n49172;
  assign n49174 = pi18 ? n49173 : n32;
  assign n49175 = pi17 ? n32 : n49174;
  assign n49176 = pi16 ? n49175 : n32;
  assign n49177 = pi15 ? n49171 : n49176;
  assign n49178 = pi14 ? n49167 : n49177;
  assign n49179 = pi13 ? n49159 : n49178;
  assign n49180 = pi18 ? n23194 : n32;
  assign n49181 = pi17 ? n32 : n49180;
  assign n49182 = pi16 ? n49181 : n32;
  assign n49183 = pi15 ? n49182 : n32;
  assign n49184 = pi14 ? n49183 : n32;
  assign n49185 = pi18 ? n37093 : ~n32;
  assign n49186 = pi17 ? n49185 : ~n32;
  assign n49187 = pi16 ? n1233 : ~n49186;
  assign n49188 = pi16 ? n17884 : n32;
  assign n49189 = pi15 ? n49187 : n49188;
  assign n49190 = pi18 ? n41994 : ~n237;
  assign n49191 = pi17 ? n32 : n49190;
  assign n49192 = pi16 ? n49191 : n32;
  assign n49193 = pi18 ? n936 : ~n605;
  assign n49194 = pi17 ? n32 : n49193;
  assign n49195 = pi16 ? n49194 : n32;
  assign n49196 = pi15 ? n49192 : n49195;
  assign n49197 = pi14 ? n49189 : n49196;
  assign n49198 = pi13 ? n49184 : n49197;
  assign n49199 = pi12 ? n49179 : n49198;
  assign n49200 = pi11 ? n49147 : n49199;
  assign n49201 = pi10 ? n49108 : n49200;
  assign n49202 = pi09 ? n49052 : n49201;
  assign n49203 = pi15 ? n24742 : n6985;
  assign n49204 = pi17 ? n2519 : ~n6587;
  assign n49205 = pi16 ? n32 : n49204;
  assign n49206 = pi17 ? n49061 : ~n3067;
  assign n49207 = pi16 ? n32 : n49206;
  assign n49208 = pi15 ? n49205 : n49207;
  assign n49209 = pi14 ? n49203 : n49208;
  assign n49210 = pi13 ? n16322 : n49209;
  assign n49211 = pi19 ? n236 : ~n349;
  assign n49212 = pi18 ? n32 : ~n49211;
  assign n49213 = pi17 ? n49068 : ~n49212;
  assign n49214 = pi16 ? n32 : n49213;
  assign n49215 = pi15 ? n49214 : n49073;
  assign n49216 = pi14 ? n49215 : n49083;
  assign n49217 = pi15 ? n15248 : n14339;
  assign n49218 = pi14 ? n49085 : n49217;
  assign n49219 = pi13 ? n49216 : n49218;
  assign n49220 = pi12 ? n49210 : n49219;
  assign n49221 = pi20 ? n3523 : n309;
  assign n49222 = pi19 ? n49221 : n5614;
  assign n49223 = pi18 ? n6118 : n49222;
  assign n49224 = pi17 ? n32 : n49223;
  assign n49225 = pi16 ? n32 : n49224;
  assign n49226 = pi15 ? n49225 : n32;
  assign n49227 = pi14 ? n49098 : n49226;
  assign n49228 = pi13 ? n49227 : n32;
  assign n49229 = pi12 ? n49228 : n47581;
  assign n49230 = pi11 ? n49220 : n49229;
  assign n49231 = pi17 ? n1697 : ~n2618;
  assign n49232 = pi16 ? n32 : n49231;
  assign n49233 = pi17 ? n31444 : ~n2618;
  assign n49234 = pi16 ? n32 : n49233;
  assign n49235 = pi15 ? n49232 : n49234;
  assign n49236 = pi17 ? n1215 : ~n2618;
  assign n49237 = pi16 ? n32 : n49236;
  assign n49238 = pi17 ? n49127 : ~n2618;
  assign n49239 = pi16 ? n32 : n49238;
  assign n49240 = pi15 ? n49237 : n49239;
  assign n49241 = pi14 ? n49235 : n49240;
  assign n49242 = pi13 ? n49241 : n49145;
  assign n49243 = pi12 ? n49118 : n49242;
  assign n49244 = pi16 ? n17850 : n49149;
  assign n49245 = pi15 ? n49244 : n49153;
  assign n49246 = pi14 ? n49245 : n49158;
  assign n49247 = pi13 ? n49246 : n49178;
  assign n49248 = pi15 ? n49187 : n130;
  assign n49249 = pi18 ? n48958 : ~n237;
  assign n49250 = pi17 ? n32 : n49249;
  assign n49251 = pi16 ? n49250 : n32;
  assign n49252 = pi21 ? n124 : n405;
  assign n49253 = pi20 ? n32 : n49252;
  assign n49254 = pi19 ? n32 : n49253;
  assign n49255 = pi18 ? n49254 : ~n605;
  assign n49256 = pi17 ? n32 : n49255;
  assign n49257 = pi16 ? n49256 : n32;
  assign n49258 = pi15 ? n49251 : n49257;
  assign n49259 = pi14 ? n49248 : n49258;
  assign n49260 = pi13 ? n49184 : n49259;
  assign n49261 = pi12 ? n49247 : n49260;
  assign n49262 = pi11 ? n49243 : n49261;
  assign n49263 = pi10 ? n49230 : n49262;
  assign n49264 = pi09 ? n49052 : n49263;
  assign n49265 = pi08 ? n49202 : n49264;
  assign n49266 = pi15 ? n16377 : n16314;
  assign n49267 = pi14 ? n32 : n49266;
  assign n49268 = pi13 ? n32 : n49267;
  assign n49269 = pi12 ? n32 : n49268;
  assign n49270 = pi11 ? n32 : n49269;
  assign n49271 = pi10 ? n32 : n49270;
  assign n49272 = pi14 ? n27740 : n32;
  assign n49273 = pi18 ? n29418 : ~n32;
  assign n49274 = pi17 ? n49273 : ~n3067;
  assign n49275 = pi16 ? n32 : n49274;
  assign n49276 = pi15 ? n37197 : n49275;
  assign n49277 = pi17 ? n2868 : ~n3067;
  assign n49278 = pi16 ? n32 : n49277;
  assign n49279 = pi17 ? n34251 : ~n3067;
  assign n49280 = pi16 ? n32 : n49279;
  assign n49281 = pi15 ? n49278 : n49280;
  assign n49282 = pi14 ? n49276 : n49281;
  assign n49283 = pi13 ? n49272 : n49282;
  assign n49284 = pi17 ? n48834 : ~n49212;
  assign n49285 = pi16 ? n32 : n49284;
  assign n49286 = pi17 ? n8193 : ~n48977;
  assign n49287 = pi16 ? n32 : n49286;
  assign n49288 = pi15 ? n49285 : n49287;
  assign n49289 = pi19 ? n4391 : n5614;
  assign n49290 = pi18 ? n5657 : n49289;
  assign n49291 = pi17 ? n32 : n49290;
  assign n49292 = pi16 ? n32 : n49291;
  assign n49293 = pi15 ? n49292 : n49082;
  assign n49294 = pi14 ? n49288 : n49293;
  assign n49295 = pi19 ? n32 : n23180;
  assign n49296 = pi18 ? n49295 : n49079;
  assign n49297 = pi17 ? n32 : n49296;
  assign n49298 = pi16 ? n32 : n49297;
  assign n49299 = pi15 ? n49298 : n14917;
  assign n49300 = pi18 ? n32 : n6669;
  assign n49301 = pi17 ? n32 : n49300;
  assign n49302 = pi16 ? n32 : n49301;
  assign n49303 = pi15 ? n14917 : n49302;
  assign n49304 = pi14 ? n49299 : n49303;
  assign n49305 = pi13 ? n49294 : n49304;
  assign n49306 = pi12 ? n49283 : n49305;
  assign n49307 = pi19 ? n4126 : n321;
  assign n49308 = pi18 ? n32 : n49307;
  assign n49309 = pi18 ? n12890 : ~n697;
  assign n49310 = pi17 ? n49308 : n49309;
  assign n49311 = pi16 ? n32 : n49310;
  assign n49312 = pi17 ? n48166 : ~n2736;
  assign n49313 = pi16 ? n32 : n49312;
  assign n49314 = pi15 ? n49311 : n49313;
  assign n49315 = pi14 ? n49314 : n23794;
  assign n49316 = pi13 ? n49315 : n23624;
  assign n49317 = pi12 ? n49316 : n32;
  assign n49318 = pi11 ? n49306 : n49317;
  assign n49319 = pi17 ? n46746 : ~n36008;
  assign n49320 = pi16 ? n32 : n49319;
  assign n49321 = pi15 ? n32 : n49320;
  assign n49322 = pi16 ? n3068 : ~n2860;
  assign n49323 = pi15 ? n49113 : n49322;
  assign n49324 = pi14 ? n49321 : n49323;
  assign n49325 = pi13 ? n22926 : n49324;
  assign n49326 = pi17 ? n1697 : ~n2750;
  assign n49327 = pi16 ? n32 : n49326;
  assign n49328 = pi17 ? n1215 : ~n2750;
  assign n49329 = pi16 ? n32 : n49328;
  assign n49330 = pi15 ? n49329 : n49327;
  assign n49331 = pi14 ? n49327 : n49330;
  assign n49332 = pi19 ? n6398 : n342;
  assign n49333 = pi18 ? n49332 : ~n32;
  assign n49334 = pi17 ? n49333 : ~n2512;
  assign n49335 = pi16 ? n32 : n49334;
  assign n49336 = pi15 ? n49335 : n49135;
  assign n49337 = pi19 ? n349 : ~n9037;
  assign n49338 = pi18 ? n49337 : n25110;
  assign n49339 = pi17 ? n32 : ~n49338;
  assign n49340 = pi16 ? n32 : n49339;
  assign n49341 = pi15 ? n35544 : n49340;
  assign n49342 = pi14 ? n49336 : n49341;
  assign n49343 = pi13 ? n49331 : n49342;
  assign n49344 = pi12 ? n49325 : n49343;
  assign n49345 = pi18 ? n6163 : n28193;
  assign n49346 = pi17 ? n3164 : ~n49345;
  assign n49347 = pi16 ? n32 : n49346;
  assign n49348 = pi15 ? n23892 : n49347;
  assign n49349 = pi16 ? n2860 : ~n2749;
  assign n49350 = pi14 ? n49348 : n49349;
  assign n49351 = pi16 ? n3946 : ~n2749;
  assign n49352 = pi18 ? n32 : n1333;
  assign n49353 = pi17 ? n32 : n49352;
  assign n49354 = pi16 ? n49353 : ~n2749;
  assign n49355 = pi15 ? n49351 : n49354;
  assign n49356 = pi19 ? n267 : n38221;
  assign n49357 = pi18 ? n49356 : n9578;
  assign n49358 = pi17 ? n32 : n49357;
  assign n49359 = pi16 ? n32 : n49358;
  assign n49360 = pi16 ? n17850 : n32;
  assign n49361 = pi15 ? n49359 : n49360;
  assign n49362 = pi14 ? n49355 : n49361;
  assign n49363 = pi13 ? n49350 : n49362;
  assign n49364 = pi15 ? n49360 : n32;
  assign n49365 = pi14 ? n49364 : n32;
  assign n49366 = pi18 ? n12172 : n23302;
  assign n49367 = pi17 ? n32 : n49366;
  assign n49368 = pi16 ? n49367 : n32;
  assign n49369 = pi15 ? n1716 : n49368;
  assign n49370 = pi18 ? n29316 : ~n35818;
  assign n49371 = pi17 ? n32 : n49370;
  assign n49372 = pi16 ? n49371 : n32;
  assign n49373 = pi18 ? n12172 : ~n605;
  assign n49374 = pi17 ? n32 : n49373;
  assign n49375 = pi16 ? n49374 : n32;
  assign n49376 = pi15 ? n49372 : n49375;
  assign n49377 = pi14 ? n49369 : n49376;
  assign n49378 = pi13 ? n49365 : n49377;
  assign n49379 = pi12 ? n49363 : n49378;
  assign n49380 = pi11 ? n49344 : n49379;
  assign n49381 = pi10 ? n49318 : n49380;
  assign n49382 = pi09 ? n49271 : n49381;
  assign n49383 = pi15 ? n16377 : n25070;
  assign n49384 = pi14 ? n32 : n49383;
  assign n49385 = pi13 ? n32 : n49384;
  assign n49386 = pi12 ? n32 : n49385;
  assign n49387 = pi11 ? n32 : n49386;
  assign n49388 = pi10 ? n32 : n49387;
  assign n49389 = pi15 ? n25070 : n32;
  assign n49390 = pi14 ? n49389 : n32;
  assign n49391 = pi17 ? n49273 : ~n2850;
  assign n49392 = pi16 ? n32 : n49391;
  assign n49393 = pi15 ? n14917 : n49392;
  assign n49394 = pi17 ? n2868 : ~n2850;
  assign n49395 = pi16 ? n32 : n49394;
  assign n49396 = pi17 ? n34251 : ~n2850;
  assign n49397 = pi16 ? n32 : n49396;
  assign n49398 = pi15 ? n49395 : n49397;
  assign n49399 = pi14 ? n49393 : n49398;
  assign n49400 = pi13 ? n49390 : n49399;
  assign n49401 = pi19 ? n236 : ~n2848;
  assign n49402 = pi18 ? n32 : ~n49401;
  assign n49403 = pi17 ? n48834 : ~n49402;
  assign n49404 = pi16 ? n32 : n49403;
  assign n49405 = pi17 ? n8193 : ~n49402;
  assign n49406 = pi16 ? n32 : n49405;
  assign n49407 = pi15 ? n49404 : n49406;
  assign n49408 = pi14 ? n49407 : n49293;
  assign n49409 = pi13 ? n49408 : n49304;
  assign n49410 = pi12 ? n49400 : n49409;
  assign n49411 = pi11 ? n49410 : n49317;
  assign n49412 = pi16 ? n3068 : ~n2624;
  assign n49413 = pi15 ? n49113 : n49412;
  assign n49414 = pi14 ? n49321 : n49413;
  assign n49415 = pi13 ? n22926 : n49414;
  assign n49416 = pi18 ? n19232 : n702;
  assign n49417 = pi17 ? n1697 : ~n49416;
  assign n49418 = pi16 ? n32 : n49417;
  assign n49419 = pi15 ? n49418 : n49327;
  assign n49420 = pi14 ? n49419 : n49330;
  assign n49421 = pi13 ? n49420 : n49342;
  assign n49422 = pi12 ? n49415 : n49421;
  assign n49423 = pi14 ? n49348 : n49155;
  assign n49424 = pi20 ? n1817 : ~n266;
  assign n49425 = pi19 ? n49424 : ~n32;
  assign n49426 = pi18 ? n32 : n49425;
  assign n49427 = pi17 ? n32 : n49426;
  assign n49428 = pi16 ? n49427 : ~n2749;
  assign n49429 = pi15 ? n49155 : n49428;
  assign n49430 = pi16 ? n20835 : n49358;
  assign n49431 = pi18 ? n17848 : n5158;
  assign n49432 = pi17 ? n32 : n49431;
  assign n49433 = pi16 ? n49432 : n32;
  assign n49434 = pi15 ? n49430 : n49433;
  assign n49435 = pi14 ? n49429 : n49434;
  assign n49436 = pi13 ? n49423 : n49435;
  assign n49437 = pi15 ? n49433 : n32;
  assign n49438 = pi14 ? n49437 : n32;
  assign n49439 = pi18 ? n29316 : ~n289;
  assign n49440 = pi17 ? n32 : n49439;
  assign n49441 = pi16 ? n49440 : n20830;
  assign n49442 = pi16 ? n49374 : n20830;
  assign n49443 = pi15 ? n49441 : n49442;
  assign n49444 = pi14 ? n49369 : n49443;
  assign n49445 = pi13 ? n49438 : n49444;
  assign n49446 = pi12 ? n49436 : n49445;
  assign n49447 = pi11 ? n49422 : n49446;
  assign n49448 = pi10 ? n49411 : n49447;
  assign n49449 = pi09 ? n49388 : n49448;
  assign n49450 = pi08 ? n49382 : n49449;
  assign n49451 = pi07 ? n49265 : n49450;
  assign n49452 = pi06 ? n49048 : n49451;
  assign n49453 = pi05 ? n48617 : n49452;
  assign n49454 = pi04 ? n47580 : n49453;
  assign n49455 = pi14 ? n32 : n26994;
  assign n49456 = pi13 ? n32 : n49455;
  assign n49457 = pi12 ? n32 : n49456;
  assign n49458 = pi11 ? n32 : n49457;
  assign n49459 = pi10 ? n32 : n49458;
  assign n49460 = pi15 ? n24237 : n33242;
  assign n49461 = pi14 ? n49460 : n32;
  assign n49462 = pi20 ? n1368 : n18261;
  assign n49463 = pi19 ? n49462 : ~n33796;
  assign n49464 = pi18 ? n49463 : n14329;
  assign n49465 = pi17 ? n32 : n49464;
  assign n49466 = pi16 ? n32 : n49465;
  assign n49467 = pi19 ? n18782 : n41496;
  assign n49468 = pi18 ? n32 : n49467;
  assign n49469 = pi20 ? n1324 : n18073;
  assign n49470 = pi19 ? n49469 : n29682;
  assign n49471 = pi19 ? n422 : ~n2848;
  assign n49472 = pi18 ? n49470 : ~n49471;
  assign n49473 = pi17 ? n49468 : ~n49472;
  assign n49474 = pi16 ? n32 : n49473;
  assign n49475 = pi15 ? n49466 : n49474;
  assign n49476 = pi18 ? n32 : n36415;
  assign n49477 = pi20 ? n1611 : n32;
  assign n49478 = pi19 ? n49477 : n41320;
  assign n49479 = pi18 ? n49478 : ~n49471;
  assign n49480 = pi17 ? n49476 : ~n49479;
  assign n49481 = pi16 ? n32 : n49480;
  assign n49482 = pi18 ? n16449 : n39517;
  assign n49483 = pi17 ? n32 : n49482;
  assign n49484 = pi16 ? n32 : n49483;
  assign n49485 = pi15 ? n49481 : n49484;
  assign n49486 = pi14 ? n49475 : n49485;
  assign n49487 = pi13 ? n49461 : n49486;
  assign n49488 = pi19 ? n24055 : n11879;
  assign n49489 = pi19 ? n3524 : ~n2848;
  assign n49490 = pi18 ? n49488 : n49489;
  assign n49491 = pi17 ? n17346 : n49490;
  assign n49492 = pi16 ? n32 : n49491;
  assign n49493 = pi19 ? n507 : ~n2848;
  assign n49494 = pi18 ? n32 : n49493;
  assign n49495 = pi17 ? n32 : n49494;
  assign n49496 = pi16 ? n32 : n49495;
  assign n49497 = pi15 ? n49492 : n49496;
  assign n49498 = pi19 ? n267 : ~n349;
  assign n49499 = pi18 ? n32 : n49498;
  assign n49500 = pi17 ? n32 : n49499;
  assign n49501 = pi16 ? n32 : n49500;
  assign n49502 = pi15 ? n49501 : n24247;
  assign n49503 = pi14 ? n49497 : n49502;
  assign n49504 = pi15 ? n32 : n35889;
  assign n49505 = pi15 ? n35889 : n39520;
  assign n49506 = pi14 ? n49504 : n49505;
  assign n49507 = pi13 ? n49503 : n49506;
  assign n49508 = pi12 ? n49487 : n49507;
  assign n49509 = pi18 ? n32 : n33422;
  assign n49510 = pi18 ? n36866 : n24731;
  assign n49511 = pi17 ? n49509 : n49510;
  assign n49512 = pi16 ? n32 : n49511;
  assign n49513 = pi18 ? n23571 : n38665;
  assign n49514 = pi17 ? n32 : n49513;
  assign n49515 = pi16 ? n32 : n49514;
  assign n49516 = pi15 ? n49512 : n49515;
  assign n49517 = pi14 ? n49516 : n32;
  assign n49518 = pi14 ? n32 : n23726;
  assign n49519 = pi13 ? n49517 : n49518;
  assign n49520 = pi14 ? n32 : n48385;
  assign n49521 = pi13 ? n32 : n49520;
  assign n49522 = pi12 ? n49519 : n49521;
  assign n49523 = pi11 ? n49508 : n49522;
  assign n49524 = pi14 ? n32 : n30209;
  assign n49525 = pi17 ? n1978 : ~n1933;
  assign n49526 = pi16 ? n32 : n49525;
  assign n49527 = pi15 ? n32 : n49526;
  assign n49528 = pi16 ? n2958 : ~n49156;
  assign n49529 = pi17 ? n32 : n4302;
  assign n49530 = pi19 ? n18489 : n32;
  assign n49531 = pi18 ? n20166 : n49530;
  assign n49532 = pi17 ? n49531 : n2623;
  assign n49533 = pi16 ? n49529 : ~n49532;
  assign n49534 = pi15 ? n49528 : n49533;
  assign n49535 = pi14 ? n49527 : n49534;
  assign n49536 = pi13 ? n49524 : n49535;
  assign n49537 = pi17 ? n2750 : ~n2623;
  assign n49538 = pi16 ? n32 : n49537;
  assign n49539 = pi18 ? n880 : n237;
  assign n49540 = pi17 ? n49539 : ~n2623;
  assign n49541 = pi16 ? n32 : n49540;
  assign n49542 = pi15 ? n49538 : n49541;
  assign n49543 = pi18 ? n32 : n1249;
  assign n49544 = pi17 ? n32 : n49543;
  assign n49545 = pi18 ? n36943 : n32;
  assign n49546 = pi17 ? n49545 : n2623;
  assign n49547 = pi16 ? n49544 : ~n49546;
  assign n49548 = pi19 ? n32 : n24055;
  assign n49549 = pi18 ? n49548 : ~n20605;
  assign n49550 = pi17 ? n49549 : ~n2623;
  assign n49551 = pi16 ? n32 : n49550;
  assign n49552 = pi15 ? n49547 : n49551;
  assign n49553 = pi14 ? n49542 : n49552;
  assign n49554 = pi19 ? n37542 : ~n4406;
  assign n49555 = pi18 ? n16389 : ~n49554;
  assign n49556 = pi18 ? n13945 : n702;
  assign n49557 = pi17 ? n49555 : ~n49556;
  assign n49558 = pi16 ? n32 : n49557;
  assign n49559 = pi20 ? n287 : ~n175;
  assign n49560 = pi19 ? n35959 : ~n49559;
  assign n49561 = pi18 ? n49560 : n508;
  assign n49562 = pi17 ? n35958 : ~n49561;
  assign n49563 = pi16 ? n32 : n49562;
  assign n49564 = pi15 ? n49558 : n49563;
  assign n49565 = pi14 ? n49564 : n35974;
  assign n49566 = pi13 ? n49553 : n49565;
  assign n49567 = pi12 ? n49536 : n49566;
  assign n49568 = pi17 ? n32 : n9311;
  assign n49569 = pi19 ? n23644 : n28623;
  assign n49570 = pi18 ? n49569 : n16389;
  assign n49571 = pi17 ? n49570 : n2512;
  assign n49572 = pi16 ? n49568 : ~n49571;
  assign n49573 = pi15 ? n13040 : n49572;
  assign n49574 = pi19 ? n23644 : n1464;
  assign n49575 = pi18 ? n49574 : n32;
  assign n49576 = pi17 ? n49575 : n2512;
  assign n49577 = pi16 ? n49568 : ~n49576;
  assign n49578 = pi16 ? n35982 : ~n2513;
  assign n49579 = pi15 ? n49577 : n49578;
  assign n49580 = pi14 ? n49573 : n49579;
  assign n49581 = pi17 ? n32 : n7039;
  assign n49582 = pi16 ? n49581 : ~n2513;
  assign n49583 = pi15 ? n49582 : n34480;
  assign n49584 = pi14 ? n49583 : n32;
  assign n49585 = pi13 ? n49580 : n49584;
  assign n49586 = pi14 ? n32 : n20969;
  assign n49587 = pi18 ? n366 : ~n36005;
  assign n49588 = pi17 ? n32 : n49587;
  assign n49589 = pi16 ? n49588 : n32;
  assign n49590 = pi15 ? n3254 : n49589;
  assign n49591 = pi18 ? n1012 : n36012;
  assign n49592 = pi17 ? n32 : n49591;
  assign n49593 = pi16 ? n49592 : n32;
  assign n49594 = pi18 ? n1012 : n36018;
  assign n49595 = pi17 ? n32 : n49594;
  assign n49596 = pi16 ? n49595 : n32;
  assign n49597 = pi15 ? n49593 : n49596;
  assign n49598 = pi14 ? n49590 : n49597;
  assign n49599 = pi13 ? n49586 : n49598;
  assign n49600 = pi12 ? n49585 : n49599;
  assign n49601 = pi11 ? n49567 : n49600;
  assign n49602 = pi10 ? n49523 : n49601;
  assign n49603 = pi09 ? n49459 : n49602;
  assign n49604 = pi18 ? n49463 : n24981;
  assign n49605 = pi17 ? n32 : n49604;
  assign n49606 = pi16 ? n32 : n49605;
  assign n49607 = pi19 ? n422 : ~n589;
  assign n49608 = pi18 ? n49470 : ~n49607;
  assign n49609 = pi17 ? n49468 : ~n49608;
  assign n49610 = pi16 ? n32 : n49609;
  assign n49611 = pi15 ? n49606 : n49610;
  assign n49612 = pi18 ? n49478 : ~n49607;
  assign n49613 = pi17 ? n49476 : ~n49612;
  assign n49614 = pi16 ? n32 : n49613;
  assign n49615 = pi18 ? n16449 : n37498;
  assign n49616 = pi17 ? n32 : n49615;
  assign n49617 = pi16 ? n32 : n49616;
  assign n49618 = pi15 ? n49614 : n49617;
  assign n49619 = pi14 ? n49611 : n49618;
  assign n49620 = pi13 ? n49461 : n49619;
  assign n49621 = pi19 ? n3524 : ~n589;
  assign n49622 = pi18 ? n49488 : n49621;
  assign n49623 = pi17 ? n17346 : n49622;
  assign n49624 = pi16 ? n32 : n49623;
  assign n49625 = pi15 ? n49624 : n36100;
  assign n49626 = pi14 ? n49625 : n49502;
  assign n49627 = pi13 ? n49626 : n49506;
  assign n49628 = pi12 ? n49620 : n49627;
  assign n49629 = pi18 ? n32 : n28164;
  assign n49630 = pi17 ? n32 : n49629;
  assign n49631 = pi16 ? n32 : n49630;
  assign n49632 = pi15 ? n49512 : n49631;
  assign n49633 = pi14 ? n49632 : n32;
  assign n49634 = pi13 ? n49633 : n32;
  assign n49635 = pi12 ? n49634 : n49521;
  assign n49636 = pi11 ? n49628 : n49635;
  assign n49637 = pi14 ? n23421 : n30209;
  assign n49638 = pi18 ? n32 : n34621;
  assign n49639 = pi17 ? n32 : n49638;
  assign n49640 = pi16 ? n2958 : ~n49639;
  assign n49641 = pi17 ? n49531 : n2855;
  assign n49642 = pi16 ? n4578 : ~n49641;
  assign n49643 = pi15 ? n49640 : n49642;
  assign n49644 = pi14 ? n49527 : n49643;
  assign n49645 = pi13 ? n49637 : n49644;
  assign n49646 = pi17 ? n2750 : ~n2750;
  assign n49647 = pi16 ? n32 : n49646;
  assign n49648 = pi15 ? n49647 : n49541;
  assign n49649 = pi17 ? n49545 : n2750;
  assign n49650 = pi16 ? n49544 : ~n49649;
  assign n49651 = pi15 ? n49650 : n49551;
  assign n49652 = pi14 ? n49648 : n49651;
  assign n49653 = pi19 ? n2358 : n49559;
  assign n49654 = pi18 ? n49653 : ~n508;
  assign n49655 = pi17 ? n36054 : n49654;
  assign n49656 = pi16 ? n32 : n49655;
  assign n49657 = pi15 ? n49558 : n49656;
  assign n49658 = pi14 ? n49657 : n35974;
  assign n49659 = pi13 ? n49652 : n49658;
  assign n49660 = pi12 ? n49645 : n49659;
  assign n49661 = pi16 ? n2958 : ~n2513;
  assign n49662 = pi15 ? n49577 : n49661;
  assign n49663 = pi14 ? n49573 : n49662;
  assign n49664 = pi16 ? n20835 : n32;
  assign n49665 = pi14 ? n49583 : n49664;
  assign n49666 = pi13 ? n49663 : n49665;
  assign n49667 = pi15 ? n49664 : n32;
  assign n49668 = pi14 ? n49667 : n20969;
  assign n49669 = pi18 ? n366 : ~n36068;
  assign n49670 = pi17 ? n32 : n49669;
  assign n49671 = pi16 ? n49670 : n32;
  assign n49672 = pi15 ? n3254 : n49671;
  assign n49673 = pi18 ? n1012 : n36074;
  assign n49674 = pi17 ? n32 : n49673;
  assign n49675 = pi16 ? n49674 : n32;
  assign n49676 = pi18 ? n1012 : n36078;
  assign n49677 = pi17 ? n32 : n49676;
  assign n49678 = pi16 ? n49677 : n32;
  assign n49679 = pi15 ? n49675 : n49678;
  assign n49680 = pi14 ? n49672 : n49679;
  assign n49681 = pi13 ? n49668 : n49680;
  assign n49682 = pi12 ? n49666 : n49681;
  assign n49683 = pi11 ? n49660 : n49682;
  assign n49684 = pi10 ? n49636 : n49683;
  assign n49685 = pi09 ? n49459 : n49684;
  assign n49686 = pi08 ? n49603 : n49685;
  assign n49687 = pi14 ? n32 : n36807;
  assign n49688 = pi13 ? n32 : n49687;
  assign n49689 = pi12 ? n32 : n49688;
  assign n49690 = pi11 ? n32 : n49689;
  assign n49691 = pi10 ? n32 : n49690;
  assign n49692 = pi14 ? n24573 : n32;
  assign n49693 = pi19 ? n507 : ~n34313;
  assign n49694 = pi18 ? n49693 : n24981;
  assign n49695 = pi17 ? n32 : n49694;
  assign n49696 = pi16 ? n32 : n49695;
  assign n49697 = pi19 ? n22864 : ~n589;
  assign n49698 = pi18 ? n32 : n49697;
  assign n49699 = pi17 ? n32 : n49698;
  assign n49700 = pi16 ? n32 : n49699;
  assign n49701 = pi15 ? n49696 : n49700;
  assign n49702 = pi19 ? n1248 : ~n589;
  assign n49703 = pi18 ? n32 : n49702;
  assign n49704 = pi17 ? n32 : n49703;
  assign n49705 = pi16 ? n32 : n49704;
  assign n49706 = pi19 ? n1490 : ~n589;
  assign n49707 = pi18 ? n32 : n49706;
  assign n49708 = pi17 ? n32 : n49707;
  assign n49709 = pi16 ? n32 : n49708;
  assign n49710 = pi15 ? n49705 : n49709;
  assign n49711 = pi14 ? n49701 : n49710;
  assign n49712 = pi13 ? n49692 : n49711;
  assign n49713 = pi15 ? n37487 : n36100;
  assign n49714 = pi14 ? n49713 : n24247;
  assign n49715 = pi15 ? n32 : n36095;
  assign n49716 = pi15 ? n36100 : n37501;
  assign n49717 = pi14 ? n49715 : n49716;
  assign n49718 = pi13 ? n49714 : n49717;
  assign n49719 = pi12 ? n49712 : n49718;
  assign n49720 = pi18 ? n21287 : n6581;
  assign n49721 = pi17 ? n32 : n49720;
  assign n49722 = pi16 ? n32 : n49721;
  assign n49723 = pi15 ? n49722 : n32;
  assign n49724 = pi14 ? n49723 : n32;
  assign n49725 = pi14 ? n23981 : n35691;
  assign n49726 = pi13 ? n49724 : n49725;
  assign n49727 = pi12 ? n49726 : n49521;
  assign n49728 = pi11 ? n49719 : n49727;
  assign n49729 = pi14 ? n38992 : n36135;
  assign n49730 = pi17 ? n4344 : ~n3509;
  assign n49731 = pi16 ? n32 : n49730;
  assign n49732 = pi15 ? n36139 : n49731;
  assign n49733 = pi18 ? n28164 : ~n4343;
  assign n49734 = pi17 ? n49733 : ~n2855;
  assign n49735 = pi16 ? n32 : n49734;
  assign n49736 = pi19 ? n18390 : ~n32;
  assign n49737 = pi18 ? n32 : n49736;
  assign n49738 = pi17 ? n49737 : ~n2855;
  assign n49739 = pi16 ? n32 : n49738;
  assign n49740 = pi15 ? n49735 : n49739;
  assign n49741 = pi14 ? n49732 : n49740;
  assign n49742 = pi13 ? n49729 : n49741;
  assign n49743 = pi17 ? n6020 : ~n2855;
  assign n49744 = pi16 ? n32 : n49743;
  assign n49745 = pi15 ? n8690 : n49744;
  assign n49746 = pi19 ? n23644 : n18396;
  assign n49747 = pi18 ? n49746 : n6019;
  assign n49748 = pi17 ? n49747 : ~n2855;
  assign n49749 = pi16 ? n32 : n49748;
  assign n49750 = pi19 ? n16002 : ~n30681;
  assign n49751 = pi18 ? n32 : ~n49750;
  assign n49752 = pi19 ? n23895 : ~n4670;
  assign n49753 = pi18 ? n49752 : ~n702;
  assign n49754 = pi17 ? n49751 : n49753;
  assign n49755 = pi16 ? n32 : n49754;
  assign n49756 = pi15 ? n49749 : n49755;
  assign n49757 = pi14 ? n49745 : n49756;
  assign n49758 = pi18 ? n32 : n29140;
  assign n49759 = pi19 ? n1757 : ~n4342;
  assign n49760 = pi18 ? n49759 : ~n702;
  assign n49761 = pi17 ? n49758 : n49760;
  assign n49762 = pi16 ? n32 : n49761;
  assign n49763 = pi18 ? n222 : ~n508;
  assign n49764 = pi17 ? n32 : n49763;
  assign n49765 = pi16 ? n32 : n49764;
  assign n49766 = pi15 ? n49762 : n49765;
  assign n49767 = pi14 ? n49766 : n36173;
  assign n49768 = pi13 ? n49757 : n49767;
  assign n49769 = pi12 ? n49742 : n49768;
  assign n49770 = pi19 ? n9007 : n37324;
  assign n49771 = pi18 ? n49770 : ~n16834;
  assign n49772 = pi17 ? n49771 : ~n2512;
  assign n49773 = pi16 ? n32 : n49772;
  assign n49774 = pi15 ? n13040 : n49773;
  assign n49775 = pi18 ? n28164 : ~n16389;
  assign n49776 = pi17 ? n49775 : ~n2628;
  assign n49777 = pi16 ? n3438 : n49776;
  assign n49778 = pi16 ? n44945 : ~n2629;
  assign n49779 = pi15 ? n49777 : n49778;
  assign n49780 = pi14 ? n49774 : n49779;
  assign n49781 = pi17 ? n32 : n31472;
  assign n49782 = pi16 ? n49781 : ~n2629;
  assign n49783 = pi15 ? n49782 : n32;
  assign n49784 = pi14 ? n49783 : n32;
  assign n49785 = pi13 ? n49780 : n49784;
  assign n49786 = pi18 ? n366 : ~n36209;
  assign n49787 = pi17 ? n32 : n49786;
  assign n49788 = pi16 ? n49787 : n32;
  assign n49789 = pi15 ? n3254 : n49788;
  assign n49790 = pi18 ? n127 : n36216;
  assign n49791 = pi17 ? n32 : n49790;
  assign n49792 = pi16 ? n49791 : n32;
  assign n49793 = pi18 ? n127 : n23571;
  assign n49794 = pi17 ? n32 : n49793;
  assign n49795 = pi16 ? n49794 : n32;
  assign n49796 = pi15 ? n49792 : n49795;
  assign n49797 = pi14 ? n49789 : n49796;
  assign n49798 = pi13 ? n32 : n49797;
  assign n49799 = pi12 ? n49785 : n49798;
  assign n49800 = pi11 ? n49769 : n49799;
  assign n49801 = pi10 ? n49728 : n49800;
  assign n49802 = pi09 ? n49691 : n49801;
  assign n49803 = pi18 ? n49693 : n7216;
  assign n49804 = pi17 ? n32 : n49803;
  assign n49805 = pi16 ? n32 : n49804;
  assign n49806 = pi19 ? n22864 : ~n2317;
  assign n49807 = pi18 ? n32 : n49806;
  assign n49808 = pi17 ? n32 : n49807;
  assign n49809 = pi16 ? n32 : n49808;
  assign n49810 = pi15 ? n49805 : n49809;
  assign n49811 = pi19 ? n1248 : ~n2317;
  assign n49812 = pi18 ? n32 : n49811;
  assign n49813 = pi17 ? n32 : n49812;
  assign n49814 = pi16 ? n32 : n49813;
  assign n49815 = pi19 ? n1490 : ~n2317;
  assign n49816 = pi18 ? n32 : n49815;
  assign n49817 = pi17 ? n32 : n49816;
  assign n49818 = pi16 ? n32 : n49817;
  assign n49819 = pi15 ? n49814 : n49818;
  assign n49820 = pi14 ? n49810 : n49819;
  assign n49821 = pi13 ? n49692 : n49820;
  assign n49822 = pi19 ? n343 : ~n2317;
  assign n49823 = pi18 ? n32 : n49822;
  assign n49824 = pi17 ? n32 : n49823;
  assign n49825 = pi16 ? n32 : n49824;
  assign n49826 = pi15 ? n49825 : n36100;
  assign n49827 = pi14 ? n49826 : n24511;
  assign n49828 = pi13 ? n49827 : n49717;
  assign n49829 = pi12 ? n49821 : n49828;
  assign n49830 = pi15 ? n49722 : n16377;
  assign n49831 = pi14 ? n49830 : n16378;
  assign n49832 = pi14 ? n16319 : n16321;
  assign n49833 = pi13 ? n49831 : n49832;
  assign n49834 = pi15 ? n32 : n23933;
  assign n49835 = pi14 ? n32 : n49834;
  assign n49836 = pi13 ? n32 : n49835;
  assign n49837 = pi12 ? n49833 : n49836;
  assign n49838 = pi11 ? n49829 : n49837;
  assign n49839 = pi15 ? n36257 : n49731;
  assign n49840 = pi14 ? n49839 : n49740;
  assign n49841 = pi13 ? n49729 : n49840;
  assign n49842 = pi12 ? n49841 : n49768;
  assign n49843 = pi17 ? n49771 : ~n2628;
  assign n49844 = pi16 ? n32 : n49843;
  assign n49845 = pi15 ? n13040 : n49844;
  assign n49846 = pi16 ? n3438 : ~n2629;
  assign n49847 = pi15 ? n49777 : n49846;
  assign n49848 = pi14 ? n49845 : n49847;
  assign n49849 = pi13 ? n49848 : n49784;
  assign n49850 = pi18 ? n127 : n36270;
  assign n49851 = pi17 ? n32 : n49850;
  assign n49852 = pi16 ? n49851 : n32;
  assign n49853 = pi15 ? n49852 : n32;
  assign n49854 = pi14 ? n49590 : n49853;
  assign n49855 = pi13 ? n32 : n49854;
  assign n49856 = pi12 ? n49849 : n49855;
  assign n49857 = pi11 ? n49842 : n49856;
  assign n49858 = pi10 ? n49838 : n49857;
  assign n49859 = pi09 ? n49691 : n49858;
  assign n49860 = pi08 ? n49802 : n49859;
  assign n49861 = pi07 ? n49686 : n49860;
  assign n49862 = pi15 ? n24495 : n16452;
  assign n49863 = pi14 ? n32 : n49862;
  assign n49864 = pi13 ? n32 : n49863;
  assign n49865 = pi12 ? n32 : n49864;
  assign n49866 = pi11 ? n32 : n49865;
  assign n49867 = pi10 ? n32 : n49866;
  assign n49868 = pi14 ? n24633 : n22818;
  assign n49869 = pi19 ? n33823 : ~n2317;
  assign n49870 = pi18 ? n20007 : n49869;
  assign n49871 = pi17 ? n32 : n49870;
  assign n49872 = pi16 ? n32 : n49871;
  assign n49873 = pi20 ? n220 : n7939;
  assign n49874 = pi19 ? n32 : ~n49873;
  assign n49875 = pi18 ? n49874 : n37498;
  assign n49876 = pi17 ? n32 : n49875;
  assign n49877 = pi16 ? n32 : n49876;
  assign n49878 = pi15 ? n49872 : n49877;
  assign n49879 = pi19 ? n519 : ~n2317;
  assign n49880 = pi18 ? n16981 : n49879;
  assign n49881 = pi17 ? n32 : n49880;
  assign n49882 = pi16 ? n32 : n49881;
  assign n49883 = pi14 ? n49878 : n49882;
  assign n49884 = pi13 ? n49868 : n49883;
  assign n49885 = pi15 ? n24705 : n24511;
  assign n49886 = pi14 ? n49885 : n24505;
  assign n49887 = pi15 ? n16105 : n24640;
  assign n49888 = pi14 ? n49887 : n24640;
  assign n49889 = pi13 ? n49886 : n49888;
  assign n49890 = pi12 ? n49884 : n49889;
  assign n49891 = pi19 ? n6057 : ~n10890;
  assign n49892 = pi18 ? n32 : n49891;
  assign n49893 = pi17 ? n32 : n49892;
  assign n49894 = pi16 ? n32 : n49893;
  assign n49895 = pi15 ? n49894 : n32;
  assign n49896 = pi14 ? n49895 : n32;
  assign n49897 = pi13 ? n49896 : n32;
  assign n49898 = pi14 ? n23794 : n23574;
  assign n49899 = pi13 ? n32 : n49898;
  assign n49900 = pi12 ? n49897 : n49899;
  assign n49901 = pi11 ? n49890 : n49900;
  assign n49902 = pi18 ? n16449 : n4343;
  assign n49903 = pi17 ? n32 : n49902;
  assign n49904 = pi16 ? n32 : n49903;
  assign n49905 = pi15 ? n23574 : n49904;
  assign n49906 = pi14 ? n49905 : n36333;
  assign n49907 = pi19 ? n6398 : n11879;
  assign n49908 = pi18 ? n49907 : n5005;
  assign n49909 = pi17 ? n32 : n49908;
  assign n49910 = pi16 ? n32 : n49909;
  assign n49911 = pi17 ? n3067 : ~n2855;
  assign n49912 = pi16 ? n32 : n49911;
  assign n49913 = pi15 ? n49910 : n49912;
  assign n49914 = pi17 ? n2959 : ~n2855;
  assign n49915 = pi16 ? n32 : n49914;
  assign n49916 = pi19 ? n3495 : n531;
  assign n49917 = pi18 ? n32 : n49916;
  assign n49918 = pi17 ? n49917 : ~n2616;
  assign n49919 = pi16 ? n32 : n49918;
  assign n49920 = pi15 ? n49915 : n49919;
  assign n49921 = pi14 ? n49913 : n49920;
  assign n49922 = pi13 ? n49906 : n49921;
  assign n49923 = pi19 ? n3495 : ~n32;
  assign n49924 = pi18 ? n32 : n49923;
  assign n49925 = pi17 ? n49924 : ~n2616;
  assign n49926 = pi16 ? n32 : n49925;
  assign n49927 = pi19 ? n32 : ~n4670;
  assign n49928 = pi18 ? n32 : n49927;
  assign n49929 = pi17 ? n49928 : ~n2616;
  assign n49930 = pi16 ? n32 : n49929;
  assign n49931 = pi15 ? n49926 : n49930;
  assign n49932 = pi19 ? n32 : ~n266;
  assign n49933 = pi18 ? n32 : n49932;
  assign n49934 = pi18 ? n268 : n1750;
  assign n49935 = pi17 ? n49933 : ~n49934;
  assign n49936 = pi16 ? n32 : n49935;
  assign n49937 = pi20 ? n260 : n206;
  assign n49938 = pi19 ? n9169 : ~n49937;
  assign n49939 = pi18 ? n32 : n49938;
  assign n49940 = pi19 ? n18728 : ~n38795;
  assign n49941 = pi18 ? n49940 : n702;
  assign n49942 = pi17 ? n49939 : ~n49941;
  assign n49943 = pi16 ? n32 : n49942;
  assign n49944 = pi15 ? n49936 : n49943;
  assign n49945 = pi14 ? n49931 : n49944;
  assign n49946 = pi19 ? n32 : ~n28451;
  assign n49947 = pi18 ? n32 : n49946;
  assign n49948 = pi19 ? n266 : n20923;
  assign n49949 = pi18 ? n49948 : n702;
  assign n49950 = pi17 ? n49947 : ~n49949;
  assign n49951 = pi16 ? n32 : n49950;
  assign n49952 = pi15 ? n49951 : n13040;
  assign n49953 = pi14 ? n49952 : n36368;
  assign n49954 = pi13 ? n49945 : n49953;
  assign n49955 = pi12 ? n49922 : n49954;
  assign n49956 = pi19 ? n246 : n322;
  assign n49957 = pi18 ? n49956 : ~n508;
  assign n49958 = pi17 ? n32 : n49957;
  assign n49959 = pi16 ? n32 : n49958;
  assign n49960 = pi19 ? n176 : ~n5707;
  assign n49961 = pi18 ? n32 : n49960;
  assign n49962 = pi20 ? n357 : ~n342;
  assign n49963 = pi19 ? n49962 : ~n6350;
  assign n49964 = pi18 ? n49963 : ~n508;
  assign n49965 = pi17 ? n49961 : n49964;
  assign n49966 = pi16 ? n32 : n49965;
  assign n49967 = pi15 ? n49959 : n49966;
  assign n49968 = pi20 ? n12882 : n342;
  assign n49969 = pi19 ? n49968 : ~n5614;
  assign n49970 = pi18 ? n209 : ~n49969;
  assign n49971 = pi17 ? n32 : n49970;
  assign n49972 = pi19 ? n6042 : n1757;
  assign n49973 = pi18 ? n702 : ~n49972;
  assign n49974 = pi20 ? n2358 : ~n342;
  assign n49975 = pi19 ? n49974 : ~n6350;
  assign n49976 = pi18 ? n49975 : ~n2627;
  assign n49977 = pi17 ? n49973 : n49976;
  assign n49978 = pi16 ? n49971 : n49977;
  assign n49979 = pi20 ? n1076 : ~n246;
  assign n49980 = pi19 ? n49979 : ~n32;
  assign n49981 = pi18 ? n49980 : ~n32;
  assign n49982 = pi17 ? n49981 : ~n2628;
  assign n49983 = pi16 ? n32 : n49982;
  assign n49984 = pi15 ? n49978 : n49983;
  assign n49985 = pi14 ? n49967 : n49984;
  assign n49986 = pi20 ? n342 : ~n16008;
  assign n49987 = pi19 ? n49986 : n32;
  assign n49988 = pi18 ? n32 : n49987;
  assign n49989 = pi17 ? n32 : n49988;
  assign n49990 = pi16 ? n17347 : n49989;
  assign n49991 = pi15 ? n49990 : n32;
  assign n49992 = pi14 ? n49991 : n32;
  assign n49993 = pi13 ? n49985 : n49992;
  assign n49994 = pi17 ? n33099 : n29699;
  assign n49995 = pi16 ? n32 : n49994;
  assign n49996 = pi15 ? n32 : n49995;
  assign n49997 = pi14 ? n32 : n49996;
  assign n49998 = pi18 ? n1012 : ~n32;
  assign n49999 = pi17 ? n32 : n49998;
  assign n50000 = pi16 ? n49999 : ~n1679;
  assign n50001 = pi18 ? n1012 : ~n940;
  assign n50002 = pi17 ? n32 : n50001;
  assign n50003 = pi18 ? n12135 : n32;
  assign n50004 = pi17 ? n50003 : n14611;
  assign n50005 = pi16 ? n50002 : n50004;
  assign n50006 = pi15 ? n50000 : n50005;
  assign n50007 = pi18 ? n127 : n36415;
  assign n50008 = pi17 ? n32 : n50007;
  assign n50009 = pi16 ? n50008 : n29937;
  assign n50010 = pi16 ? n32 : n29937;
  assign n50011 = pi15 ? n50009 : n50010;
  assign n50012 = pi14 ? n50006 : n50011;
  assign n50013 = pi13 ? n49997 : n50012;
  assign n50014 = pi12 ? n49993 : n50013;
  assign n50015 = pi11 ? n49955 : n50014;
  assign n50016 = pi10 ? n49901 : n50015;
  assign n50017 = pi09 ? n49867 : n50016;
  assign n50018 = pi14 ? n32 : n39563;
  assign n50019 = pi13 ? n32 : n50018;
  assign n50020 = pi12 ? n32 : n50019;
  assign n50021 = pi11 ? n32 : n50020;
  assign n50022 = pi10 ? n32 : n50021;
  assign n50023 = pi19 ? n33823 : ~n343;
  assign n50024 = pi18 ? n20007 : n50023;
  assign n50025 = pi17 ? n32 : n50024;
  assign n50026 = pi16 ? n32 : n50025;
  assign n50027 = pi18 ? n49874 : n14648;
  assign n50028 = pi17 ? n32 : n50027;
  assign n50029 = pi16 ? n32 : n50028;
  assign n50030 = pi15 ? n50026 : n50029;
  assign n50031 = pi18 ? n16981 : n15072;
  assign n50032 = pi17 ? n32 : n50031;
  assign n50033 = pi16 ? n32 : n50032;
  assign n50034 = pi14 ? n50030 : n50033;
  assign n50035 = pi13 ? n49868 : n50034;
  assign n50036 = pi15 ? n15230 : n24640;
  assign n50037 = pi14 ? n50036 : n24505;
  assign n50038 = pi15 ? n16105 : n24511;
  assign n50039 = pi14 ? n50038 : n24640;
  assign n50040 = pi13 ? n50037 : n50039;
  assign n50041 = pi12 ? n50035 : n50040;
  assign n50042 = pi15 ? n24813 : n32;
  assign n50043 = pi14 ? n50042 : n32;
  assign n50044 = pi13 ? n50043 : n32;
  assign n50045 = pi14 ? n32 : n23623;
  assign n50046 = pi13 ? n32 : n50045;
  assign n50047 = pi12 ? n50044 : n50046;
  assign n50048 = pi11 ? n50041 : n50047;
  assign n50049 = pi15 ? n24905 : n49904;
  assign n50050 = pi14 ? n50049 : n36333;
  assign n50051 = pi17 ? n2959 : ~n2616;
  assign n50052 = pi16 ? n32 : n50051;
  assign n50053 = pi15 ? n50052 : n49919;
  assign n50054 = pi14 ? n49913 : n50053;
  assign n50055 = pi13 ? n50050 : n50054;
  assign n50056 = pi18 ? n49940 : n1750;
  assign n50057 = pi17 ? n49939 : ~n50056;
  assign n50058 = pi16 ? n32 : n50057;
  assign n50059 = pi15 ? n49936 : n50058;
  assign n50060 = pi14 ? n49931 : n50059;
  assign n50061 = pi14 ? n49952 : n36453;
  assign n50062 = pi13 ? n50060 : n50061;
  assign n50063 = pi12 ? n50055 : n50062;
  assign n50064 = pi18 ? n49956 : ~n595;
  assign n50065 = pi17 ? n32 : n50064;
  assign n50066 = pi16 ? n32 : n50065;
  assign n50067 = pi18 ? n49963 : ~n595;
  assign n50068 = pi17 ? n49961 : n50067;
  assign n50069 = pi16 ? n32 : n50068;
  assign n50070 = pi15 ? n50066 : n50069;
  assign n50071 = pi20 ? n11107 : n428;
  assign n50072 = pi19 ? n50071 : ~n43838;
  assign n50073 = pi18 ? n1395 : ~n50072;
  assign n50074 = pi17 ? n32 : n50073;
  assign n50075 = pi18 ? n49975 : ~n595;
  assign n50076 = pi17 ? n49973 : n50075;
  assign n50077 = pi16 ? n50074 : n50076;
  assign n50078 = pi18 ? n49160 : ~n32;
  assign n50079 = pi17 ? n50078 : ~n2618;
  assign n50080 = pi16 ? n32 : n50079;
  assign n50081 = pi15 ? n50077 : n50080;
  assign n50082 = pi14 ? n50070 : n50081;
  assign n50083 = pi16 ? n17347 : n21345;
  assign n50084 = pi15 ? n50083 : n32;
  assign n50085 = pi14 ? n50084 : n32;
  assign n50086 = pi13 ? n50082 : n50085;
  assign n50087 = pi19 ? n502 : ~n322;
  assign n50088 = pi18 ? n50087 : n32;
  assign n50089 = pi17 ? n50088 : n32;
  assign n50090 = pi16 ? n50002 : n50089;
  assign n50091 = pi15 ? n50000 : n50090;
  assign n50092 = pi17 ? n32 : n49476;
  assign n50093 = pi17 ? n19432 : n20658;
  assign n50094 = pi16 ? n50092 : n50093;
  assign n50095 = pi15 ? n50094 : n50010;
  assign n50096 = pi14 ? n50091 : n50095;
  assign n50097 = pi13 ? n49997 : n50096;
  assign n50098 = pi12 ? n50086 : n50097;
  assign n50099 = pi11 ? n50063 : n50098;
  assign n50100 = pi10 ? n50048 : n50099;
  assign n50101 = pi09 ? n50022 : n50100;
  assign n50102 = pi08 ? n50017 : n50101;
  assign n50103 = pi14 ? n32 : n24880;
  assign n50104 = pi13 ? n32 : n50103;
  assign n50105 = pi12 ? n32 : n50104;
  assign n50106 = pi11 ? n32 : n50105;
  assign n50107 = pi10 ? n32 : n50106;
  assign n50108 = pi14 ? n25965 : n22818;
  assign n50109 = pi19 ? n9037 : ~n589;
  assign n50110 = pi18 ? n1249 : n50109;
  assign n50111 = pi17 ? n32 : n50110;
  assign n50112 = pi16 ? n32 : n50111;
  assign n50113 = pi19 ? n32 : ~n18728;
  assign n50114 = pi19 ? n2359 : ~n589;
  assign n50115 = pi18 ? n50113 : n50114;
  assign n50116 = pi17 ? n32 : n50115;
  assign n50117 = pi16 ? n32 : n50116;
  assign n50118 = pi15 ? n50112 : n50117;
  assign n50119 = pi14 ? n50118 : n14651;
  assign n50120 = pi13 ? n50108 : n50119;
  assign n50121 = pi15 ? n15230 : n24511;
  assign n50122 = pi14 ? n50121 : n24505;
  assign n50123 = pi15 ? n24511 : n24700;
  assign n50124 = pi14 ? n50123 : n24700;
  assign n50125 = pi13 ? n50122 : n50124;
  assign n50126 = pi12 ? n50120 : n50125;
  assign n50127 = pi13 ? n32 : n36030;
  assign n50128 = pi14 ? n32 : n23924;
  assign n50129 = pi13 ? n50128 : n32;
  assign n50130 = pi12 ? n50127 : n50129;
  assign n50131 = pi11 ? n50126 : n50130;
  assign n50132 = pi19 ? n594 : n18728;
  assign n50133 = pi18 ? n50132 : n36511;
  assign n50134 = pi17 ? n32 : n50133;
  assign n50135 = pi16 ? n32 : n50134;
  assign n50136 = pi15 ? n32 : n50135;
  assign n50137 = pi14 ? n50136 : n36520;
  assign n50138 = pi20 ? n14286 : ~n206;
  assign n50139 = pi19 ? n50138 : ~n236;
  assign n50140 = pi18 ? n36522 : n50139;
  assign n50141 = pi17 ? n32 : n50140;
  assign n50142 = pi16 ? n32 : n50141;
  assign n50143 = pi15 ? n50142 : n7124;
  assign n50144 = pi15 ? n49915 : n9408;
  assign n50145 = pi14 ? n50143 : n50144;
  assign n50146 = pi13 ? n50137 : n50145;
  assign n50147 = pi19 ? n32 : ~n4491;
  assign n50148 = pi18 ? n32 : n50147;
  assign n50149 = pi17 ? n50148 : ~n2616;
  assign n50150 = pi16 ? n32 : n50149;
  assign n50151 = pi15 ? n8688 : n50150;
  assign n50152 = pi19 ? n32 : n2358;
  assign n50153 = pi18 ? n32 : n50152;
  assign n50154 = pi19 ? n1844 : n9591;
  assign n50155 = pi18 ? n50154 : n2615;
  assign n50156 = pi17 ? n50153 : ~n50155;
  assign n50157 = pi16 ? n32 : n50156;
  assign n50158 = pi19 ? n10485 : n507;
  assign n50159 = pi18 ? n50158 : ~n1750;
  assign n50160 = pi17 ? n32 : n50159;
  assign n50161 = pi16 ? n32 : n50160;
  assign n50162 = pi15 ? n50157 : n50161;
  assign n50163 = pi14 ? n50151 : n50162;
  assign n50164 = pi19 ? n32331 : ~n18678;
  assign n50165 = pi18 ? n50164 : n702;
  assign n50166 = pi17 ? n15845 : ~n50165;
  assign n50167 = pi16 ? n32 : n50166;
  assign n50168 = pi15 ? n50167 : n23892;
  assign n50169 = pi14 ? n50168 : n36543;
  assign n50170 = pi13 ? n50163 : n50169;
  assign n50171 = pi12 ? n50146 : n50170;
  assign n50172 = pi18 ? n21274 : ~n595;
  assign n50173 = pi17 ? n8617 : n50172;
  assign n50174 = pi16 ? n32 : n50173;
  assign n50175 = pi15 ? n36542 : n50174;
  assign n50176 = pi19 ? n5356 : n1757;
  assign n50177 = pi18 ? n702 : ~n50176;
  assign n50178 = pi19 ? n18489 : n4342;
  assign n50179 = pi18 ? n50178 : n595;
  assign n50180 = pi17 ? n50177 : ~n50179;
  assign n50181 = pi16 ? n32 : n50180;
  assign n50182 = pi17 ? n1994 : ~n2618;
  assign n50183 = pi16 ? n32 : n50182;
  assign n50184 = pi15 ? n50181 : n50183;
  assign n50185 = pi14 ? n50175 : n50184;
  assign n50186 = pi17 ? n29220 : n32;
  assign n50187 = pi16 ? n32 : n50186;
  assign n50188 = pi15 ? n50187 : n32;
  assign n50189 = pi14 ? n50188 : n32;
  assign n50190 = pi13 ? n50185 : n50189;
  assign n50191 = pi20 ? n1331 : ~n173;
  assign n50192 = pi19 ? n175 : n50191;
  assign n50193 = pi18 ? n32 : n50192;
  assign n50194 = pi17 ? n32 : n50193;
  assign n50195 = pi18 ? n359 : n36578;
  assign n50196 = pi18 ? n36580 : n32;
  assign n50197 = pi17 ? n50195 : ~n50196;
  assign n50198 = pi16 ? n50194 : ~n50197;
  assign n50199 = pi15 ? n32 : n50198;
  assign n50200 = pi14 ? n32 : n50199;
  assign n50201 = pi16 ? n45307 : ~n1679;
  assign n50202 = pi18 ? n127 : ~n940;
  assign n50203 = pi17 ? n32 : n50202;
  assign n50204 = pi19 ? n36588 : ~n322;
  assign n50205 = pi18 ? n50204 : n32;
  assign n50206 = pi17 ? n50205 : n32;
  assign n50207 = pi16 ? n50203 : n50206;
  assign n50208 = pi15 ? n50201 : n50207;
  assign n50209 = pi18 ? n1012 : n16847;
  assign n50210 = pi17 ? n32 : n50209;
  assign n50211 = pi17 ? n36598 : n32;
  assign n50212 = pi16 ? n50210 : n50211;
  assign n50213 = pi18 ? n21316 : n32;
  assign n50214 = pi17 ? n50213 : n664;
  assign n50215 = pi16 ? n32 : n50214;
  assign n50216 = pi15 ? n50212 : n50215;
  assign n50217 = pi14 ? n50208 : n50216;
  assign n50218 = pi13 ? n50200 : n50217;
  assign n50219 = pi12 ? n50190 : n50218;
  assign n50220 = pi11 ? n50171 : n50219;
  assign n50221 = pi10 ? n50131 : n50220;
  assign n50222 = pi09 ? n50107 : n50221;
  assign n50223 = pi14 ? n16607 : n22818;
  assign n50224 = pi19 ? n9037 : ~n2303;
  assign n50225 = pi18 ? n1249 : n50224;
  assign n50226 = pi17 ? n32 : n50225;
  assign n50227 = pi16 ? n32 : n50226;
  assign n50228 = pi19 ? n2359 : ~n2303;
  assign n50229 = pi18 ? n50113 : n50228;
  assign n50230 = pi17 ? n32 : n50229;
  assign n50231 = pi16 ? n32 : n50230;
  assign n50232 = pi15 ? n50227 : n50231;
  assign n50233 = pi19 ? n322 : ~n2303;
  assign n50234 = pi18 ? n32 : n50233;
  assign n50235 = pi17 ? n32 : n50234;
  assign n50236 = pi16 ? n32 : n50235;
  assign n50237 = pi14 ? n50232 : n50236;
  assign n50238 = pi13 ? n50223 : n50237;
  assign n50239 = pi15 ? n37923 : n24700;
  assign n50240 = pi14 ? n50239 : n24505;
  assign n50241 = pi13 ? n50240 : n50124;
  assign n50242 = pi12 ? n50238 : n50241;
  assign n50243 = pi14 ? n24368 : n24370;
  assign n50244 = pi13 ? n50243 : n36030;
  assign n50245 = pi12 ? n50244 : n32;
  assign n50246 = pi11 ? n50242 : n50245;
  assign n50247 = pi19 ? n50138 : ~n1941;
  assign n50248 = pi18 ? n36522 : n50247;
  assign n50249 = pi17 ? n32 : n50248;
  assign n50250 = pi16 ? n32 : n50249;
  assign n50251 = pi17 ? n3067 : ~n3070;
  assign n50252 = pi16 ? n32 : n50251;
  assign n50253 = pi15 ? n50250 : n50252;
  assign n50254 = pi15 ? n9681 : n9403;
  assign n50255 = pi14 ? n50253 : n50254;
  assign n50256 = pi13 ? n50137 : n50255;
  assign n50257 = pi17 ? n2750 : ~n2736;
  assign n50258 = pi16 ? n32 : n50257;
  assign n50259 = pi17 ? n50148 : ~n2736;
  assign n50260 = pi16 ? n32 : n50259;
  assign n50261 = pi15 ? n50258 : n50260;
  assign n50262 = pi18 ? n50154 : n1750;
  assign n50263 = pi17 ? n50153 : ~n50262;
  assign n50264 = pi16 ? n32 : n50263;
  assign n50265 = pi18 ? n42558 : ~n1750;
  assign n50266 = pi17 ? n32 : n50265;
  assign n50267 = pi16 ? n32 : n50266;
  assign n50268 = pi15 ? n50264 : n50267;
  assign n50269 = pi14 ? n50261 : n50268;
  assign n50270 = pi13 ? n50269 : n50169;
  assign n50271 = pi12 ? n50256 : n50270;
  assign n50272 = pi18 ? n50178 : n4098;
  assign n50273 = pi17 ? n50177 : ~n50272;
  assign n50274 = pi16 ? n32 : n50273;
  assign n50275 = pi17 ? n1718 : ~n2618;
  assign n50276 = pi16 ? n32 : n50275;
  assign n50277 = pi15 ? n50274 : n50276;
  assign n50278 = pi14 ? n50175 : n50277;
  assign n50279 = pi18 ? n9578 : n32;
  assign n50280 = pi17 ? n50279 : n32;
  assign n50281 = pi16 ? n32 : n50280;
  assign n50282 = pi14 ? n50188 : n50281;
  assign n50283 = pi13 ? n50278 : n50282;
  assign n50284 = pi15 ? n50281 : n32;
  assign n50285 = pi21 ? n140 : n405;
  assign n50286 = pi20 ? n32 : n50285;
  assign n50287 = pi19 ? n32 : n50286;
  assign n50288 = pi18 ? n50287 : ~n32;
  assign n50289 = pi17 ? n32 : n50288;
  assign n50290 = pi17 ? n36579 : ~n50196;
  assign n50291 = pi16 ? n50289 : ~n50290;
  assign n50292 = pi15 ? n32 : n50291;
  assign n50293 = pi14 ? n50284 : n50292;
  assign n50294 = pi19 ? n5688 : ~n322;
  assign n50295 = pi18 ? n50294 : n32;
  assign n50296 = pi17 ? n50295 : n32;
  assign n50297 = pi16 ? n50203 : n50296;
  assign n50298 = pi15 ? n50201 : n50297;
  assign n50299 = pi17 ? n36651 : n32;
  assign n50300 = pi16 ? n50210 : n50299;
  assign n50301 = pi17 ? n50213 : n20658;
  assign n50302 = pi16 ? n32 : n50301;
  assign n50303 = pi15 ? n50300 : n50302;
  assign n50304 = pi14 ? n50298 : n50303;
  assign n50305 = pi13 ? n50293 : n50304;
  assign n50306 = pi12 ? n50283 : n50305;
  assign n50307 = pi11 ? n50271 : n50306;
  assign n50308 = pi10 ? n50246 : n50307;
  assign n50309 = pi09 ? n50107 : n50308;
  assign n50310 = pi08 ? n50222 : n50309;
  assign n50311 = pi07 ? n50102 : n50310;
  assign n50312 = pi06 ? n49861 : n50311;
  assign n50313 = pi14 ? n32 : n16837;
  assign n50314 = pi13 ? n32 : n50313;
  assign n50315 = pi12 ? n32 : n50314;
  assign n50316 = pi11 ? n32 : n50315;
  assign n50317 = pi10 ? n32 : n50316;
  assign n50318 = pi19 ? n342 : ~n343;
  assign n50319 = pi18 ? n4380 : n50318;
  assign n50320 = pi17 ? n32 : n50319;
  assign n50321 = pi16 ? n32 : n50320;
  assign n50322 = pi15 ? n16452 : n50321;
  assign n50323 = pi14 ? n37470 : n50322;
  assign n50324 = pi18 ? n209 : ~n684;
  assign n50325 = pi17 ? n32 : n50324;
  assign n50326 = pi16 ? n32 : n50325;
  assign n50327 = pi19 ? n4391 : ~n2303;
  assign n50328 = pi18 ? n32 : n50327;
  assign n50329 = pi17 ? n32 : n50328;
  assign n50330 = pi16 ? n32 : n50329;
  assign n50331 = pi15 ? n50326 : n50330;
  assign n50332 = pi19 ? n321 : ~n2303;
  assign n50333 = pi18 ? n32 : n50332;
  assign n50334 = pi17 ? n32 : n50333;
  assign n50335 = pi16 ? n32 : n50334;
  assign n50336 = pi14 ? n50331 : n50335;
  assign n50337 = pi13 ? n50323 : n50336;
  assign n50338 = pi19 ? n32 : ~n2303;
  assign n50339 = pi18 ? n32 : n50338;
  assign n50340 = pi17 ? n32 : n50339;
  assign n50341 = pi16 ? n32 : n50340;
  assign n50342 = pi15 ? n50341 : n16452;
  assign n50343 = pi18 ? n49295 : n24697;
  assign n50344 = pi17 ? n32 : n50343;
  assign n50345 = pi16 ? n32 : n50344;
  assign n50346 = pi18 ? n49295 : n14648;
  assign n50347 = pi17 ? n32 : n50346;
  assign n50348 = pi16 ? n32 : n50347;
  assign n50349 = pi15 ? n50345 : n50348;
  assign n50350 = pi14 ? n50342 : n50349;
  assign n50351 = pi15 ? n24700 : n25044;
  assign n50352 = pi19 ? n32 : ~n16431;
  assign n50353 = pi19 ? n462 : ~n2303;
  assign n50354 = pi18 ? n50352 : n50353;
  assign n50355 = pi17 ? n32 : n50354;
  assign n50356 = pi16 ? n32 : n50355;
  assign n50357 = pi15 ? n50356 : n16786;
  assign n50358 = pi14 ? n50351 : n50357;
  assign n50359 = pi13 ? n50350 : n50358;
  assign n50360 = pi12 ? n50337 : n50359;
  assign n50361 = pi14 ? n23924 : n32;
  assign n50362 = pi13 ? n32 : n50361;
  assign n50363 = pi12 ? n32 : n50362;
  assign n50364 = pi11 ? n50360 : n50363;
  assign n50365 = pi18 ? n29140 : n24015;
  assign n50366 = pi17 ? n32 : n50365;
  assign n50367 = pi16 ? n32 : n50366;
  assign n50368 = pi15 ? n50367 : n9141;
  assign n50369 = pi15 ? n9403 : n8476;
  assign n50370 = pi14 ? n50368 : n50369;
  assign n50371 = pi13 ? n36705 : n50370;
  assign n50372 = pi20 ? n342 : n915;
  assign n50373 = pi19 ? n32 : n50372;
  assign n50374 = pi18 ? n32 : ~n50373;
  assign n50375 = pi18 ? n359 : n697;
  assign n50376 = pi17 ? n50374 : ~n50375;
  assign n50377 = pi16 ? n32 : n50376;
  assign n50378 = pi15 ? n9403 : n50377;
  assign n50379 = pi18 ? n24306 : n6163;
  assign n50380 = pi17 ? n32 : n50379;
  assign n50381 = pi16 ? n32 : n50380;
  assign n50382 = pi19 ? n322 : n37542;
  assign n50383 = pi18 ? n50382 : n6163;
  assign n50384 = pi17 ? n32 : n50383;
  assign n50385 = pi16 ? n32 : n50384;
  assign n50386 = pi15 ? n50381 : n50385;
  assign n50387 = pi14 ? n50378 : n50386;
  assign n50388 = pi18 ? n36720 : n13335;
  assign n50389 = pi17 ? n32 : n50388;
  assign n50390 = pi16 ? n32 : n50389;
  assign n50391 = pi15 ? n50390 : n36729;
  assign n50392 = pi18 ? n16041 : n36732;
  assign n50393 = pi17 ? n32 : n50392;
  assign n50394 = pi16 ? n32 : n50393;
  assign n50395 = pi15 ? n36735 : n50394;
  assign n50396 = pi14 ? n50391 : n50395;
  assign n50397 = pi13 ? n50387 : n50396;
  assign n50398 = pi12 ? n50371 : n50397;
  assign n50399 = pi18 ? n15844 : n5742;
  assign n50400 = pi17 ? n32 : n50399;
  assign n50401 = pi16 ? n32 : n50400;
  assign n50402 = pi17 ? n1807 : ~n2512;
  assign n50403 = pi16 ? n32 : n50402;
  assign n50404 = pi15 ? n50401 : n50403;
  assign n50405 = pi17 ? n1682 : ~n4099;
  assign n50406 = pi16 ? n32 : n50405;
  assign n50407 = pi15 ? n50406 : n32;
  assign n50408 = pi14 ? n50404 : n50407;
  assign n50409 = pi13 ? n50408 : n32;
  assign n50410 = pi18 ? n127 : n532;
  assign n50411 = pi17 ? n32 : n50410;
  assign n50412 = pi16 ? n50411 : ~n2727;
  assign n50413 = pi15 ? n32 : n50412;
  assign n50414 = pi14 ? n32 : n50413;
  assign n50415 = pi18 ? n1012 : n532;
  assign n50416 = pi17 ? n32 : n50415;
  assign n50417 = pi19 ? n18497 : n32;
  assign n50418 = pi18 ? n50417 : n32;
  assign n50419 = pi17 ? n24781 : ~n50418;
  assign n50420 = pi16 ? n50416 : ~n50419;
  assign n50421 = pi18 ? n6645 : n23073;
  assign n50422 = pi17 ? n50421 : ~n32;
  assign n50423 = pi16 ? n50411 : ~n50422;
  assign n50424 = pi15 ? n50420 : n50423;
  assign n50425 = pi17 ? n36794 : n32;
  assign n50426 = pi16 ? n129 : n50425;
  assign n50427 = pi17 ? n50213 : n32;
  assign n50428 = pi16 ? n32 : n50427;
  assign n50429 = pi15 ? n50426 : n50428;
  assign n50430 = pi14 ? n50424 : n50429;
  assign n50431 = pi13 ? n50414 : n50430;
  assign n50432 = pi12 ? n50409 : n50431;
  assign n50433 = pi11 ? n50398 : n50432;
  assign n50434 = pi10 ? n50364 : n50433;
  assign n50435 = pi09 ? n50317 : n50434;
  assign n50436 = pi18 ? n209 : ~n1965;
  assign n50437 = pi17 ? n32 : n50436;
  assign n50438 = pi16 ? n32 : n50437;
  assign n50439 = pi19 ? n4391 : ~n429;
  assign n50440 = pi18 ? n32 : n50439;
  assign n50441 = pi17 ? n32 : n50440;
  assign n50442 = pi16 ? n32 : n50441;
  assign n50443 = pi15 ? n50438 : n50442;
  assign n50444 = pi19 ? n321 : ~n429;
  assign n50445 = pi18 ? n32 : n50444;
  assign n50446 = pi17 ? n32 : n50445;
  assign n50447 = pi16 ? n32 : n50446;
  assign n50448 = pi14 ? n50443 : n50447;
  assign n50449 = pi13 ? n50323 : n50448;
  assign n50450 = pi14 ? n27529 : n50349;
  assign n50451 = pi13 ? n50450 : n50358;
  assign n50452 = pi12 ? n50449 : n50451;
  assign n50453 = pi14 ? n32 : n24368;
  assign n50454 = pi13 ? n50453 : n32;
  assign n50455 = pi12 ? n50454 : n50362;
  assign n50456 = pi11 ? n50452 : n50455;
  assign n50457 = pi17 ? n2519 : ~n2731;
  assign n50458 = pi16 ? n32 : n50457;
  assign n50459 = pi15 ? n9403 : n50458;
  assign n50460 = pi14 ? n50368 : n50459;
  assign n50461 = pi13 ? n36705 : n50460;
  assign n50462 = pi17 ? n2726 : ~n2731;
  assign n50463 = pi16 ? n32 : n50462;
  assign n50464 = pi15 ? n50463 : n50377;
  assign n50465 = pi14 ? n50464 : n50386;
  assign n50466 = pi13 ? n50465 : n50396;
  assign n50467 = pi12 ? n50461 : n50466;
  assign n50468 = pi17 ? n1682 : ~n2618;
  assign n50469 = pi16 ? n32 : n50468;
  assign n50470 = pi15 ? n50469 : n32;
  assign n50471 = pi14 ? n50404 : n50470;
  assign n50472 = pi14 ? n32 : n50281;
  assign n50473 = pi13 ? n50471 : n50472;
  assign n50474 = pi14 ? n50284 : n50413;
  assign n50475 = pi18 ? n25595 : n23073;
  assign n50476 = pi17 ? n50475 : ~n32;
  assign n50477 = pi16 ? n50411 : ~n50476;
  assign n50478 = pi15 ? n50420 : n50477;
  assign n50479 = pi17 ? n36837 : n32;
  assign n50480 = pi16 ? n129 : n50479;
  assign n50481 = pi15 ? n50480 : n50302;
  assign n50482 = pi14 ? n50478 : n50481;
  assign n50483 = pi13 ? n50474 : n50482;
  assign n50484 = pi12 ? n50473 : n50483;
  assign n50485 = pi11 ? n50467 : n50484;
  assign n50486 = pi10 ? n50456 : n50485;
  assign n50487 = pi09 ? n50317 : n50486;
  assign n50488 = pi08 ? n50435 : n50487;
  assign n50489 = pi14 ? n32 : n25823;
  assign n50490 = pi13 ? n32 : n50489;
  assign n50491 = pi12 ? n32 : n50490;
  assign n50492 = pi11 ? n32 : n50491;
  assign n50493 = pi10 ? n32 : n50492;
  assign n50494 = pi19 ? n6057 : n2303;
  assign n50495 = pi18 ? n222 : ~n50494;
  assign n50496 = pi17 ? n32 : n50495;
  assign n50497 = pi16 ? n32 : n50496;
  assign n50498 = pi15 ? n16101 : n50497;
  assign n50499 = pi14 ? n26770 : n50498;
  assign n50500 = pi18 ? n684 : ~n2830;
  assign n50501 = pi17 ? n32 : n50500;
  assign n50502 = pi16 ? n32 : n50501;
  assign n50503 = pi18 ? n936 : n50444;
  assign n50504 = pi17 ? n32 : n50503;
  assign n50505 = pi16 ? n32 : n50504;
  assign n50506 = pi15 ? n50502 : n50505;
  assign n50507 = pi14 ? n50506 : n50505;
  assign n50508 = pi13 ? n50499 : n50507;
  assign n50509 = pi15 ? n27528 : n24874;
  assign n50510 = pi19 ? n1464 : ~n429;
  assign n50511 = pi18 ? n32 : n50510;
  assign n50512 = pi17 ? n32 : n50511;
  assign n50513 = pi16 ? n32 : n50512;
  assign n50514 = pi15 ? n50513 : n14895;
  assign n50515 = pi14 ? n50509 : n50514;
  assign n50516 = pi15 ? n27528 : n25211;
  assign n50517 = pi18 ? n32 : n35966;
  assign n50518 = pi17 ? n32 : n50517;
  assign n50519 = pi16 ? n32 : n50518;
  assign n50520 = pi15 ? n50519 : n32;
  assign n50521 = pi14 ? n50516 : n50520;
  assign n50522 = pi13 ? n50515 : n50521;
  assign n50523 = pi12 ? n50508 : n50522;
  assign n50524 = pi14 ? n32 : n24498;
  assign n50525 = pi13 ? n50524 : n32;
  assign n50526 = pi14 ? n32 : n35688;
  assign n50527 = pi13 ? n32 : n50526;
  assign n50528 = pi12 ? n50525 : n50527;
  assign n50529 = pi11 ? n50523 : n50528;
  assign n50530 = pi19 ? n32 : ~n23895;
  assign n50531 = pi19 ? n8611 : ~n236;
  assign n50532 = pi18 ? n50530 : n50531;
  assign n50533 = pi17 ? n32 : n50532;
  assign n50534 = pi16 ? n32 : n50533;
  assign n50535 = pi15 ? n32 : n50534;
  assign n50536 = pi14 ? n36893 : n50535;
  assign n50537 = pi19 ? n15527 : n236;
  assign n50538 = pi18 ? n605 : ~n50537;
  assign n50539 = pi17 ? n32 : n50538;
  assign n50540 = pi16 ? n32 : n50539;
  assign n50541 = pi15 ? n50540 : n9141;
  assign n50542 = pi17 ? n2531 : ~n2731;
  assign n50543 = pi16 ? n32 : n50542;
  assign n50544 = pi15 ? n50463 : n50543;
  assign n50545 = pi14 ? n50541 : n50544;
  assign n50546 = pi13 ? n50536 : n50545;
  assign n50547 = pi19 ? n247 : n531;
  assign n50548 = pi18 ? n32 : n50547;
  assign n50549 = pi17 ? n50548 : ~n2731;
  assign n50550 = pi16 ? n32 : n50549;
  assign n50551 = pi18 ? n32 : ~n16847;
  assign n50552 = pi18 ? n24647 : ~n48314;
  assign n50553 = pi17 ? n50551 : ~n50552;
  assign n50554 = pi16 ? n32 : n50553;
  assign n50555 = pi15 ? n50550 : n50554;
  assign n50556 = pi18 ? n20020 : n6163;
  assign n50557 = pi17 ? n32 : n50556;
  assign n50558 = pi16 ? n32 : n50557;
  assign n50559 = pi19 ? n322 : n36903;
  assign n50560 = pi18 ? n50559 : ~n35719;
  assign n50561 = pi17 ? n32 : n50560;
  assign n50562 = pi16 ? n32 : n50561;
  assign n50563 = pi15 ? n50558 : n50562;
  assign n50564 = pi14 ? n50555 : n50563;
  assign n50565 = pi18 ? n36911 : ~n47647;
  assign n50566 = pi17 ? n32 : n50565;
  assign n50567 = pi16 ? n32 : n50566;
  assign n50568 = pi18 ? n36917 : ~n32928;
  assign n50569 = pi17 ? n32 : n50568;
  assign n50570 = pi16 ? n32 : n50569;
  assign n50571 = pi15 ? n50567 : n50570;
  assign n50572 = pi18 ? n15844 : n34401;
  assign n50573 = pi17 ? n32 : n50572;
  assign n50574 = pi16 ? n32 : n50573;
  assign n50575 = pi14 ? n50571 : n50574;
  assign n50576 = pi13 ? n50564 : n50575;
  assign n50577 = pi12 ? n50546 : n50576;
  assign n50578 = pi18 ? n15844 : n13901;
  assign n50579 = pi17 ? n32 : n50578;
  assign n50580 = pi16 ? n32 : n50579;
  assign n50581 = pi15 ? n50580 : n7355;
  assign n50582 = pi17 ? n1682 : ~n2512;
  assign n50583 = pi16 ? n32 : n50582;
  assign n50584 = pi17 ? n36981 : n32;
  assign n50585 = pi16 ? n32 : n50584;
  assign n50586 = pi15 ? n50583 : n50585;
  assign n50587 = pi14 ? n50581 : n50586;
  assign n50588 = pi17 ? n28638 : n32;
  assign n50589 = pi16 ? n32 : n50588;
  assign n50590 = pi14 ? n32 : n50589;
  assign n50591 = pi13 ? n50587 : n50590;
  assign n50592 = pi18 ? n24942 : n32;
  assign n50593 = pi17 ? n2726 : ~n50592;
  assign n50594 = pi16 ? n3625 : ~n50593;
  assign n50595 = pi15 ? n32 : n50594;
  assign n50596 = pi14 ? n50589 : n50595;
  assign n50597 = pi19 ? n28854 : n23644;
  assign n50598 = pi18 ? n50597 : n248;
  assign n50599 = pi17 ? n24948 : ~n50598;
  assign n50600 = pi16 ? n3625 : ~n50599;
  assign n50601 = pi18 ? n36959 : n605;
  assign n50602 = pi17 ? n50601 : ~n32;
  assign n50603 = pi16 ? n3625 : ~n50602;
  assign n50604 = pi15 ? n50600 : n50603;
  assign n50605 = pi17 ? n36965 : n32;
  assign n50606 = pi16 ? n129 : n50605;
  assign n50607 = pi15 ? n50606 : n20660;
  assign n50608 = pi14 ? n50604 : n50607;
  assign n50609 = pi13 ? n50596 : n50608;
  assign n50610 = pi12 ? n50591 : n50609;
  assign n50611 = pi11 ? n50577 : n50610;
  assign n50612 = pi10 ? n50529 : n50611;
  assign n50613 = pi09 ? n50493 : n50612;
  assign n50614 = pi14 ? n32 : n26063;
  assign n50615 = pi13 ? n32 : n50614;
  assign n50616 = pi12 ? n32 : n50615;
  assign n50617 = pi11 ? n32 : n50616;
  assign n50618 = pi10 ? n32 : n50617;
  assign n50619 = pi19 ? n6057 : n429;
  assign n50620 = pi18 ? n222 : ~n50619;
  assign n50621 = pi17 ? n32 : n50620;
  assign n50622 = pi16 ? n32 : n50621;
  assign n50623 = pi15 ? n25211 : n50622;
  assign n50624 = pi14 ? n26770 : n50623;
  assign n50625 = pi18 ? n684 : ~n2962;
  assign n50626 = pi17 ? n32 : n50625;
  assign n50627 = pi16 ? n32 : n50626;
  assign n50628 = pi19 ? n321 : ~n2297;
  assign n50629 = pi18 ? n936 : n50628;
  assign n50630 = pi17 ? n32 : n50629;
  assign n50631 = pi16 ? n32 : n50630;
  assign n50632 = pi15 ? n50627 : n50631;
  assign n50633 = pi14 ? n50632 : n50631;
  assign n50634 = pi13 ? n50624 : n50633;
  assign n50635 = pi19 ? n32 : ~n2297;
  assign n50636 = pi18 ? n32 : n50635;
  assign n50637 = pi17 ? n32 : n50636;
  assign n50638 = pi16 ? n32 : n50637;
  assign n50639 = pi15 ? n50638 : n24874;
  assign n50640 = pi14 ? n50639 : n50514;
  assign n50641 = pi13 ? n50640 : n50521;
  assign n50642 = pi12 ? n50634 : n50641;
  assign n50643 = pi11 ? n50642 : n32;
  assign n50644 = pi17 ? n2726 : ~n2724;
  assign n50645 = pi16 ? n32 : n50644;
  assign n50646 = pi17 ? n2531 : ~n2724;
  assign n50647 = pi16 ? n32 : n50646;
  assign n50648 = pi15 ? n50645 : n50647;
  assign n50649 = pi14 ? n50541 : n50648;
  assign n50650 = pi13 ? n50536 : n50649;
  assign n50651 = pi17 ? n50548 : ~n2736;
  assign n50652 = pi16 ? n32 : n50651;
  assign n50653 = pi19 ? n32 : n30461;
  assign n50654 = pi18 ? n50653 : ~n48314;
  assign n50655 = pi17 ? n50551 : ~n50654;
  assign n50656 = pi16 ? n32 : n50655;
  assign n50657 = pi15 ? n50652 : n50656;
  assign n50658 = pi14 ? n50657 : n50563;
  assign n50659 = pi18 ? n15844 : n34613;
  assign n50660 = pi17 ? n32 : n50659;
  assign n50661 = pi16 ? n32 : n50660;
  assign n50662 = pi14 ? n50571 : n50661;
  assign n50663 = pi13 ? n50658 : n50662;
  assign n50664 = pi12 ? n50650 : n50663;
  assign n50665 = pi15 ? n50589 : n32;
  assign n50666 = pi16 ? n50411 : ~n50593;
  assign n50667 = pi15 ? n32 : n50666;
  assign n50668 = pi14 ? n50665 : n50667;
  assign n50669 = pi19 ? n28854 : n39054;
  assign n50670 = pi18 ? n50669 : n248;
  assign n50671 = pi17 ? n32 : ~n50670;
  assign n50672 = pi16 ? n50411 : ~n50671;
  assign n50673 = pi18 ? n37013 : n605;
  assign n50674 = pi17 ? n50673 : ~n32;
  assign n50675 = pi16 ? n50411 : ~n50674;
  assign n50676 = pi15 ? n50672 : n50675;
  assign n50677 = pi17 ? n37019 : n32;
  assign n50678 = pi16 ? n32 : n50677;
  assign n50679 = pi15 ? n50678 : n20660;
  assign n50680 = pi14 ? n50676 : n50679;
  assign n50681 = pi13 ? n50668 : n50680;
  assign n50682 = pi12 ? n50591 : n50681;
  assign n50683 = pi11 ? n50664 : n50682;
  assign n50684 = pi10 ? n50643 : n50683;
  assign n50685 = pi09 ? n50618 : n50684;
  assign n50686 = pi08 ? n50613 : n50685;
  assign n50687 = pi07 ? n50488 : n50686;
  assign n50688 = pi15 ? n17039 : n15847;
  assign n50689 = pi14 ? n32 : n50688;
  assign n50690 = pi13 ? n32 : n50689;
  assign n50691 = pi12 ? n32 : n50690;
  assign n50692 = pi11 ? n32 : n50691;
  assign n50693 = pi10 ? n32 : n50692;
  assign n50694 = pi19 ? n267 : ~n343;
  assign n50695 = pi18 ? n32 : n50694;
  assign n50696 = pi17 ? n32 : n50695;
  assign n50697 = pi16 ? n32 : n50696;
  assign n50698 = pi15 ? n17039 : n50697;
  assign n50699 = pi19 ? n18390 : n429;
  assign n50700 = pi18 ? n858 : ~n50699;
  assign n50701 = pi17 ? n32 : n50700;
  assign n50702 = pi16 ? n32 : n50701;
  assign n50703 = pi15 ? n27528 : n50702;
  assign n50704 = pi14 ? n50698 : n50703;
  assign n50705 = pi18 ? n702 : ~n2962;
  assign n50706 = pi17 ? n32 : n50705;
  assign n50707 = pi16 ? n32 : n50706;
  assign n50708 = pi18 ? n1741 : ~n2962;
  assign n50709 = pi17 ? n32 : n50708;
  assign n50710 = pi16 ? n32 : n50709;
  assign n50711 = pi15 ? n50707 : n50710;
  assign n50712 = pi20 ? n428 : n6822;
  assign n50713 = pi19 ? n32 : n50712;
  assign n50714 = pi20 ? n18408 : ~n32;
  assign n50715 = pi19 ? n50714 : ~n13085;
  assign n50716 = pi18 ? n50713 : ~n50715;
  assign n50717 = pi17 ? n32 : n50716;
  assign n50718 = pi16 ? n32 : n50717;
  assign n50719 = pi15 ? n50718 : n25384;
  assign n50720 = pi14 ? n50711 : n50719;
  assign n50721 = pi13 ? n50704 : n50720;
  assign n50722 = pi20 ? n428 : n1324;
  assign n50723 = pi19 ? n32 : n50722;
  assign n50724 = pi19 ? n5694 : n429;
  assign n50725 = pi18 ? n50723 : ~n50724;
  assign n50726 = pi17 ? n32 : n50725;
  assign n50727 = pi16 ? n32 : n50726;
  assign n50728 = pi15 ? n25211 : n50727;
  assign n50729 = pi14 ? n25385 : n50728;
  assign n50730 = pi15 ? n27528 : n27304;
  assign n50731 = pi21 ? n405 : n2076;
  assign n50732 = pi20 ? n50731 : n32;
  assign n50733 = pi19 ? n1818 : n50732;
  assign n50734 = pi18 ? n32 : n50733;
  assign n50735 = pi17 ? n32 : n50734;
  assign n50736 = pi16 ? n32 : n50735;
  assign n50737 = pi15 ? n50736 : n32;
  assign n50738 = pi14 ? n50730 : n50737;
  assign n50739 = pi13 ? n50729 : n50738;
  assign n50740 = pi12 ? n50721 : n50739;
  assign n50741 = pi19 ? n4126 : n3495;
  assign n50742 = pi18 ? n32 : n50741;
  assign n50743 = pi17 ? n32 : n50742;
  assign n50744 = pi16 ? n32 : n50743;
  assign n50745 = pi15 ? n32 : n50744;
  assign n50746 = pi14 ? n32 : n50745;
  assign n50747 = pi13 ? n32 : n50746;
  assign n50748 = pi12 ? n32 : n50747;
  assign n50749 = pi11 ? n50740 : n50748;
  assign n50750 = pi19 ? n2386 : n236;
  assign n50751 = pi18 ? n16847 : ~n50750;
  assign n50752 = pi17 ? n32 : n50751;
  assign n50753 = pi16 ? n32 : n50752;
  assign n50754 = pi19 ? n32 : n34092;
  assign n50755 = pi19 ? n4670 : n1812;
  assign n50756 = pi18 ? n50754 : ~n50755;
  assign n50757 = pi17 ? n32 : n50756;
  assign n50758 = pi16 ? n32 : n50757;
  assign n50759 = pi15 ? n50753 : n50758;
  assign n50760 = pi14 ? n37072 : n50759;
  assign n50761 = pi18 ? n350 : ~n4244;
  assign n50762 = pi17 ? n32 : n50761;
  assign n50763 = pi16 ? n32 : n50762;
  assign n50764 = pi17 ? n3164 : ~n2724;
  assign n50765 = pi16 ? n32 : n50764;
  assign n50766 = pi15 ? n50763 : n50765;
  assign n50767 = pi17 ? n7396 : ~n2724;
  assign n50768 = pi16 ? n32 : n50767;
  assign n50769 = pi15 ? n9663 : n50768;
  assign n50770 = pi14 ? n50766 : n50769;
  assign n50771 = pi13 ? n50760 : n50770;
  assign n50772 = pi19 ? n208 : n18502;
  assign n50773 = pi18 ? n32 : n50772;
  assign n50774 = pi17 ? n50773 : ~n2724;
  assign n50775 = pi16 ? n32 : n50774;
  assign n50776 = pi20 ? n3523 : ~n266;
  assign n50777 = pi19 ? n50776 : ~n32;
  assign n50778 = pi18 ? n32 : n50777;
  assign n50779 = pi17 ? n50778 : ~n2736;
  assign n50780 = pi16 ? n32 : n50779;
  assign n50781 = pi15 ? n50775 : n50780;
  assign n50782 = pi18 ? n34208 : ~n702;
  assign n50783 = pi17 ? n32 : n50782;
  assign n50784 = pi16 ? n32 : n50783;
  assign n50785 = pi15 ? n12056 : n50784;
  assign n50786 = pi14 ? n50781 : n50785;
  assign n50787 = pi18 ? n7647 : ~n702;
  assign n50788 = pi17 ? n32 : n50787;
  assign n50789 = pi16 ? n32 : n50788;
  assign n50790 = pi15 ? n50789 : n37099;
  assign n50791 = pi18 ? n9346 : ~n702;
  assign n50792 = pi17 ? n32 : n50791;
  assign n50793 = pi16 ? n32 : n50792;
  assign n50794 = pi18 ? n7038 : n25787;
  assign n50795 = pi17 ? n32 : n50794;
  assign n50796 = pi16 ? n32 : n50795;
  assign n50797 = pi15 ? n50793 : n50796;
  assign n50798 = pi14 ? n50790 : n50797;
  assign n50799 = pi13 ? n50786 : n50798;
  assign n50800 = pi12 ? n50771 : n50799;
  assign n50801 = pi20 ? n3523 : n1331;
  assign n50802 = pi19 ? n32 : n50801;
  assign n50803 = pi18 ? n209 : ~n50802;
  assign n50804 = pi17 ? n32 : n50803;
  assign n50805 = pi20 ? n6050 : n220;
  assign n50806 = pi19 ? n50805 : n3524;
  assign n50807 = pi18 ? n50806 : ~n32;
  assign n50808 = pi18 ? n17118 : ~n32928;
  assign n50809 = pi17 ? n50807 : ~n50808;
  assign n50810 = pi16 ? n50804 : ~n50809;
  assign n50811 = pi17 ? n35572 : ~n2750;
  assign n50812 = pi16 ? n32 : n50811;
  assign n50813 = pi15 ? n50810 : n50812;
  assign n50814 = pi14 ? n50813 : n32;
  assign n50815 = pi18 ? n16981 : n359;
  assign n50816 = pi17 ? n50815 : n32;
  assign n50817 = pi16 ? n32 : n50816;
  assign n50818 = pi14 ? n32 : n50817;
  assign n50819 = pi13 ? n50814 : n50818;
  assign n50820 = pi18 ? n25109 : ~n32;
  assign n50821 = pi17 ? n32 : n50820;
  assign n50822 = pi16 ? n3061 : ~n50821;
  assign n50823 = pi15 ? n32 : n50822;
  assign n50824 = pi14 ? n50817 : n50823;
  assign n50825 = pi19 ? n32 : ~n19749;
  assign n50826 = pi18 ? n50825 : ~n32;
  assign n50827 = pi17 ? n32 : n50826;
  assign n50828 = pi16 ? n3061 : ~n50827;
  assign n50829 = pi18 ? n31959 : ~n32;
  assign n50830 = pi17 ? n19071 : n50829;
  assign n50831 = pi16 ? n2958 : ~n50830;
  assign n50832 = pi15 ? n50828 : n50831;
  assign n50833 = pi17 ? n20065 : n22085;
  assign n50834 = pi16 ? n32 : n50833;
  assign n50835 = pi15 ? n50834 : n32;
  assign n50836 = pi14 ? n50832 : n50835;
  assign n50837 = pi13 ? n50824 : n50836;
  assign n50838 = pi12 ? n50819 : n50837;
  assign n50839 = pi11 ? n50800 : n50838;
  assign n50840 = pi10 ? n50749 : n50839;
  assign n50841 = pi09 ? n50693 : n50840;
  assign n50842 = pi19 ? n18390 : n531;
  assign n50843 = pi18 ? n858 : ~n50842;
  assign n50844 = pi17 ? n32 : n50843;
  assign n50845 = pi16 ? n32 : n50844;
  assign n50846 = pi15 ? n27528 : n50845;
  assign n50847 = pi14 ? n50698 : n50846;
  assign n50848 = pi18 ? n1741 : ~n880;
  assign n50849 = pi17 ? n32 : n50848;
  assign n50850 = pi16 ? n32 : n50849;
  assign n50851 = pi15 ? n10291 : n50850;
  assign n50852 = pi20 ? n18173 : ~n32;
  assign n50853 = pi19 ? n50852 : ~n5707;
  assign n50854 = pi18 ? n17848 : ~n50853;
  assign n50855 = pi17 ? n32 : n50854;
  assign n50856 = pi16 ? n32 : n50855;
  assign n50857 = pi15 ? n50856 : n15847;
  assign n50858 = pi14 ? n50851 : n50857;
  assign n50859 = pi13 ? n50847 : n50858;
  assign n50860 = pi14 ? n25640 : n50728;
  assign n50861 = pi14 ? n50730 : n16974;
  assign n50862 = pi13 ? n50860 : n50861;
  assign n50863 = pi12 ? n50859 : n50862;
  assign n50864 = pi14 ? n16786 : n16840;
  assign n50865 = pi13 ? n32 : n50864;
  assign n50866 = pi12 ? n50865 : n50747;
  assign n50867 = pi11 ? n50863 : n50866;
  assign n50868 = pi18 ? n50754 : ~n38127;
  assign n50869 = pi17 ? n32 : n50868;
  assign n50870 = pi16 ? n32 : n50869;
  assign n50871 = pi15 ? n50753 : n50870;
  assign n50872 = pi14 ? n37072 : n50871;
  assign n50873 = pi18 ? n350 : ~n496;
  assign n50874 = pi17 ? n32 : n50873;
  assign n50875 = pi16 ? n32 : n50874;
  assign n50876 = pi15 ? n50875 : n50765;
  assign n50877 = pi17 ? n7396 : ~n4245;
  assign n50878 = pi16 ? n32 : n50877;
  assign n50879 = pi15 ? n9663 : n50878;
  assign n50880 = pi14 ? n50876 : n50879;
  assign n50881 = pi13 ? n50872 : n50880;
  assign n50882 = pi17 ? n36742 : ~n2736;
  assign n50883 = pi16 ? n32 : n50882;
  assign n50884 = pi15 ? n50775 : n50883;
  assign n50885 = pi14 ? n50884 : n50785;
  assign n50886 = pi13 ? n50885 : n50798;
  assign n50887 = pi12 ? n50881 : n50886;
  assign n50888 = pi18 ? n245 : ~n19082;
  assign n50889 = pi17 ? n32 : n50888;
  assign n50890 = pi20 ? n8943 : n5854;
  assign n50891 = pi19 ? n50890 : n804;
  assign n50892 = pi18 ? n50891 : ~n32;
  assign n50893 = pi17 ? n50892 : ~n50808;
  assign n50894 = pi16 ? n50889 : ~n50893;
  assign n50895 = pi15 ? n50894 : n50812;
  assign n50896 = pi14 ? n50895 : n32;
  assign n50897 = pi13 ? n50896 : n50590;
  assign n50898 = pi14 ? n50589 : n50823;
  assign n50899 = pi17 ? n37213 : n21317;
  assign n50900 = pi16 ? n32 : n50899;
  assign n50901 = pi15 ? n50900 : n32;
  assign n50902 = pi14 ? n50832 : n50901;
  assign n50903 = pi13 ? n50898 : n50902;
  assign n50904 = pi12 ? n50897 : n50903;
  assign n50905 = pi11 ? n50887 : n50904;
  assign n50906 = pi10 ? n50867 : n50905;
  assign n50907 = pi09 ? n50693 : n50906;
  assign n50908 = pi08 ? n50841 : n50907;
  assign n50909 = pi20 ? n18834 : ~n207;
  assign n50910 = pi19 ? n50909 : n365;
  assign n50911 = pi18 ? n32 : ~n50910;
  assign n50912 = pi17 ? n32 : n50911;
  assign n50913 = pi16 ? n32 : n50912;
  assign n50914 = pi15 ? n50913 : n16485;
  assign n50915 = pi14 ? n17273 : n50914;
  assign n50916 = pi13 ? n32 : n50915;
  assign n50917 = pi12 ? n32 : n50916;
  assign n50918 = pi11 ? n32 : n50917;
  assign n50919 = pi10 ? n32 : n50918;
  assign n50920 = pi19 ? n275 : ~n429;
  assign n50921 = pi18 ? n32 : n50920;
  assign n50922 = pi17 ? n32 : n50921;
  assign n50923 = pi16 ? n32 : n50922;
  assign n50924 = pi18 ? n863 : ~n50842;
  assign n50925 = pi17 ? n32 : n50924;
  assign n50926 = pi16 ? n32 : n50925;
  assign n50927 = pi15 ? n50923 : n50926;
  assign n50928 = pi14 ? n50698 : n50927;
  assign n50929 = pi20 ? n5854 : n1817;
  assign n50930 = pi19 ? n50929 : n531;
  assign n50931 = pi18 ? n42108 : ~n50930;
  assign n50932 = pi17 ? n32 : n50931;
  assign n50933 = pi16 ? n32 : n50932;
  assign n50934 = pi20 ? n3523 : ~n831;
  assign n50935 = pi19 ? n50934 : n5707;
  assign n50936 = pi18 ? n32 : n50935;
  assign n50937 = pi17 ? n32 : n50936;
  assign n50938 = pi16 ? n32 : n50937;
  assign n50939 = pi15 ? n50933 : n50938;
  assign n50940 = pi19 ? n32 : n6171;
  assign n50941 = pi18 ? n32 : n50940;
  assign n50942 = pi17 ? n32 : n50941;
  assign n50943 = pi16 ? n32 : n50942;
  assign n50944 = pi15 ? n15847 : n50943;
  assign n50945 = pi14 ? n50939 : n50944;
  assign n50946 = pi13 ? n50928 : n50945;
  assign n50947 = pi18 ? n32 : n22889;
  assign n50948 = pi17 ? n32 : n50947;
  assign n50949 = pi16 ? n32 : n50948;
  assign n50950 = pi15 ? n22817 : n50949;
  assign n50951 = pi20 ? n9194 : n6026;
  assign n50952 = pi19 ? n50951 : ~n11108;
  assign n50953 = pi18 ? n1819 : n50952;
  assign n50954 = pi17 ? n32 : n50953;
  assign n50955 = pi16 ? n32 : n50954;
  assign n50956 = pi20 ? n9194 : n3897;
  assign n50957 = pi19 ? n50956 : ~n11108;
  assign n50958 = pi18 ? n32 : n50957;
  assign n50959 = pi17 ? n32 : n50958;
  assign n50960 = pi16 ? n32 : n50959;
  assign n50961 = pi15 ? n50955 : n50960;
  assign n50962 = pi14 ? n50950 : n50961;
  assign n50963 = pi19 ? n6398 : ~n11108;
  assign n50964 = pi18 ? n32 : n50963;
  assign n50965 = pi17 ? n32 : n50964;
  assign n50966 = pi16 ? n32 : n50965;
  assign n50967 = pi15 ? n50966 : n15403;
  assign n50968 = pi15 ? n16973 : n16606;
  assign n50969 = pi14 ? n50967 : n50968;
  assign n50970 = pi13 ? n50962 : n50969;
  assign n50971 = pi12 ? n50946 : n50970;
  assign n50972 = pi15 ? n24572 : n37258;
  assign n50973 = pi14 ? n24368 : n50972;
  assign n50974 = pi13 ? n32 : n50973;
  assign n50975 = pi12 ? n32 : n50974;
  assign n50976 = pi11 ? n50971 : n50975;
  assign n50977 = pi18 ? n16847 : ~n496;
  assign n50978 = pi17 ? n32 : n50977;
  assign n50979 = pi16 ? n32 : n50978;
  assign n50980 = pi18 ? n222 : ~n496;
  assign n50981 = pi17 ? n32 : n50980;
  assign n50982 = pi16 ? n32 : n50981;
  assign n50983 = pi15 ? n50979 : n50982;
  assign n50984 = pi14 ? n30921 : n50983;
  assign n50985 = pi17 ? n3067 : ~n4245;
  assign n50986 = pi16 ? n32 : n50985;
  assign n50987 = pi15 ? n50765 : n50986;
  assign n50988 = pi14 ? n50876 : n50987;
  assign n50989 = pi13 ? n50984 : n50988;
  assign n50990 = pi20 ? n3843 : ~n9863;
  assign n50991 = pi19 ? n32 : n50990;
  assign n50992 = pi18 ? n32 : n50991;
  assign n50993 = pi17 ? n50992 : ~n4245;
  assign n50994 = pi16 ? n32 : n50993;
  assign n50995 = pi17 ? n6236 : ~n2724;
  assign n50996 = pi16 ? n32 : n50995;
  assign n50997 = pi15 ? n50994 : n50996;
  assign n50998 = pi18 ? n496 : ~n962;
  assign n50999 = pi17 ? n32 : n50998;
  assign n51000 = pi16 ? n32 : n50999;
  assign n51001 = pi18 ? n34208 : ~n697;
  assign n51002 = pi17 ? n32 : n51001;
  assign n51003 = pi16 ? n32 : n51002;
  assign n51004 = pi15 ? n51000 : n51003;
  assign n51005 = pi14 ? n50997 : n51004;
  assign n51006 = pi15 ? n12261 : n37296;
  assign n51007 = pi18 ? n880 : ~n1750;
  assign n51008 = pi17 ? n32 : n51007;
  assign n51009 = pi16 ? n32 : n51008;
  assign n51010 = pi15 ? n51009 : n50796;
  assign n51011 = pi14 ? n51006 : n51010;
  assign n51012 = pi13 ? n51005 : n51011;
  assign n51013 = pi12 ? n50989 : n51012;
  assign n51014 = pi18 ? n1464 : ~n32;
  assign n51015 = pi18 ? n22885 : ~n37298;
  assign n51016 = pi17 ? n51014 : ~n51015;
  assign n51017 = pi16 ? n1323 : ~n51016;
  assign n51018 = pi17 ? n2750 : ~n7922;
  assign n51019 = pi16 ? n32 : n51018;
  assign n51020 = pi15 ? n51017 : n51019;
  assign n51021 = pi14 ? n51020 : n32;
  assign n51022 = pi17 ? n28818 : n32;
  assign n51023 = pi16 ? n32 : n51022;
  assign n51024 = pi14 ? n32 : n51023;
  assign n51025 = pi13 ? n51021 : n51024;
  assign n51026 = pi17 ? n18292 : n32;
  assign n51027 = pi16 ? n32 : n51026;
  assign n51028 = pi15 ? n51023 : n51027;
  assign n51029 = pi18 ? n25266 : n46870;
  assign n51030 = pi17 ? n32 : n51029;
  assign n51031 = pi16 ? n2958 : ~n51030;
  assign n51032 = pi15 ? n32 : n51031;
  assign n51033 = pi14 ? n51028 : n51032;
  assign n51034 = pi18 ? n20193 : n237;
  assign n51035 = pi17 ? n32 : n51034;
  assign n51036 = pi16 ? n2958 : ~n51035;
  assign n51037 = pi18 ? n20788 : ~n32;
  assign n51038 = pi17 ? n19071 : n51037;
  assign n51039 = pi16 ? n2958 : ~n51038;
  assign n51040 = pi15 ? n51036 : n51039;
  assign n51041 = pi17 ? n37353 : n21317;
  assign n51042 = pi16 ? n32 : n51041;
  assign n51043 = pi19 ? n507 : ~n5707;
  assign n51044 = pi18 ? n1575 : ~n51043;
  assign n51045 = pi17 ? n32 : n51044;
  assign n51046 = pi16 ? n51045 : n32;
  assign n51047 = pi15 ? n51042 : n51046;
  assign n51048 = pi14 ? n51040 : n51047;
  assign n51049 = pi13 ? n51033 : n51048;
  assign n51050 = pi12 ? n51025 : n51049;
  assign n51051 = pi11 ? n51013 : n51050;
  assign n51052 = pi10 ? n50976 : n51051;
  assign n51053 = pi09 ? n50919 : n51052;
  assign n51054 = pi20 ? n7839 : n207;
  assign n51055 = pi19 ? n51054 : ~n365;
  assign n51056 = pi18 ? n32 : n51055;
  assign n51057 = pi17 ? n32 : n51056;
  assign n51058 = pi16 ? n32 : n51057;
  assign n51059 = pi15 ? n51058 : n16485;
  assign n51060 = pi14 ? n17273 : n51059;
  assign n51061 = pi13 ? n32 : n51060;
  assign n51062 = pi12 ? n32 : n51061;
  assign n51063 = pi11 ? n32 : n51062;
  assign n51064 = pi10 ? n32 : n51063;
  assign n51065 = pi19 ? n18390 : n365;
  assign n51066 = pi18 ? n863 : ~n51065;
  assign n51067 = pi17 ? n32 : n51066;
  assign n51068 = pi16 ? n32 : n51067;
  assign n51069 = pi15 ? n50923 : n51068;
  assign n51070 = pi14 ? n50698 : n51069;
  assign n51071 = pi19 ? n50934 : n13074;
  assign n51072 = pi18 ? n32 : n51071;
  assign n51073 = pi17 ? n32 : n51072;
  assign n51074 = pi16 ? n32 : n51073;
  assign n51075 = pi15 ? n50933 : n51074;
  assign n51076 = pi15 ? n16485 : n50943;
  assign n51077 = pi14 ? n51075 : n51076;
  assign n51078 = pi13 ? n51070 : n51077;
  assign n51079 = pi19 ? n507 : n4491;
  assign n51080 = pi18 ? n32 : n51079;
  assign n51081 = pi17 ? n32 : n51080;
  assign n51082 = pi16 ? n32 : n51081;
  assign n51083 = pi19 ? n507 : n6171;
  assign n51084 = pi18 ? n32 : n51083;
  assign n51085 = pi17 ? n32 : n51084;
  assign n51086 = pi16 ? n32 : n51085;
  assign n51087 = pi15 ? n51082 : n51086;
  assign n51088 = pi19 ? n50951 : ~n8818;
  assign n51089 = pi18 ? n1819 : n51088;
  assign n51090 = pi17 ? n32 : n51089;
  assign n51091 = pi16 ? n32 : n51090;
  assign n51092 = pi19 ? n50956 : ~n8818;
  assign n51093 = pi18 ? n32 : n51092;
  assign n51094 = pi17 ? n32 : n51093;
  assign n51095 = pi16 ? n32 : n51094;
  assign n51096 = pi15 ? n51091 : n51095;
  assign n51097 = pi14 ? n51087 : n51096;
  assign n51098 = pi19 ? n6398 : ~n8818;
  assign n51099 = pi18 ? n32 : n51098;
  assign n51100 = pi17 ? n32 : n51099;
  assign n51101 = pi16 ? n32 : n51100;
  assign n51102 = pi15 ? n51101 : n15403;
  assign n51103 = pi14 ? n51102 : n32;
  assign n51104 = pi13 ? n51097 : n51103;
  assign n51105 = pi12 ? n51078 : n51104;
  assign n51106 = pi15 ? n24237 : n37383;
  assign n51107 = pi14 ? n32 : n51106;
  assign n51108 = pi13 ? n32 : n51107;
  assign n51109 = pi12 ? n32 : n51108;
  assign n51110 = pi11 ? n51105 : n51109;
  assign n51111 = pi18 ? n16847 : ~n590;
  assign n51112 = pi17 ? n32 : n51111;
  assign n51113 = pi16 ? n32 : n51112;
  assign n51114 = pi18 ? n222 : ~n2849;
  assign n51115 = pi17 ? n32 : n51114;
  assign n51116 = pi16 ? n32 : n51115;
  assign n51117 = pi15 ? n51113 : n51116;
  assign n51118 = pi14 ? n30921 : n51117;
  assign n51119 = pi18 ? n350 : ~n2849;
  assign n51120 = pi17 ? n32 : n51119;
  assign n51121 = pi16 ? n32 : n51120;
  assign n51122 = pi15 ? n51121 : n7743;
  assign n51123 = pi15 ? n7743 : n50986;
  assign n51124 = pi14 ? n51122 : n51123;
  assign n51125 = pi13 ? n51118 : n51124;
  assign n51126 = pi20 ? n1331 : ~n1685;
  assign n51127 = pi19 ? n32 : n51126;
  assign n51128 = pi18 ? n32 : n51127;
  assign n51129 = pi17 ? n51128 : ~n4245;
  assign n51130 = pi16 ? n32 : n51129;
  assign n51131 = pi17 ? n6236 : ~n4245;
  assign n51132 = pi16 ? n32 : n51131;
  assign n51133 = pi15 ? n51130 : n51132;
  assign n51134 = pi18 ? n496 : ~n4244;
  assign n51135 = pi17 ? n32 : n51134;
  assign n51136 = pi16 ? n32 : n51135;
  assign n51137 = pi18 ? n34208 : ~n2730;
  assign n51138 = pi17 ? n32 : n51137;
  assign n51139 = pi16 ? n32 : n51138;
  assign n51140 = pi15 ? n51136 : n51139;
  assign n51141 = pi14 ? n51133 : n51140;
  assign n51142 = pi18 ? n684 : ~n2730;
  assign n51143 = pi17 ? n32 : n51142;
  assign n51144 = pi16 ? n32 : n51143;
  assign n51145 = pi15 ? n51144 : n37296;
  assign n51146 = pi18 ? n880 : ~n697;
  assign n51147 = pi17 ? n32 : n51146;
  assign n51148 = pi16 ? n32 : n51147;
  assign n51149 = pi18 ? n32 : n19065;
  assign n51150 = pi17 ? n32 : n51149;
  assign n51151 = pi16 ? n51150 : n50795;
  assign n51152 = pi15 ? n51148 : n51151;
  assign n51153 = pi14 ? n51145 : n51152;
  assign n51154 = pi13 ? n51141 : n51153;
  assign n51155 = pi12 ? n51125 : n51154;
  assign n51156 = pi18 ? n1464 : ~n359;
  assign n51157 = pi17 ? n51156 : ~n51015;
  assign n51158 = pi16 ? n1683 : ~n51157;
  assign n51159 = pi19 ? n2141 : n617;
  assign n51160 = pi18 ? n32 : n51159;
  assign n51161 = pi17 ? n2750 : ~n51160;
  assign n51162 = pi16 ? n32 : n51161;
  assign n51163 = pi15 ? n51158 : n51162;
  assign n51164 = pi14 ? n51163 : n32;
  assign n51165 = pi17 ? n20658 : n32;
  assign n51166 = pi16 ? n32 : n51165;
  assign n51167 = pi14 ? n32 : n51166;
  assign n51168 = pi13 ? n51164 : n51167;
  assign n51169 = pi15 ? n51166 : n32;
  assign n51170 = pi18 ? n25357 : n532;
  assign n51171 = pi17 ? n32 : n51170;
  assign n51172 = pi16 ? n2958 : ~n51171;
  assign n51173 = pi15 ? n32 : n51172;
  assign n51174 = pi14 ? n51169 : n51173;
  assign n51175 = pi19 ? n5446 : n531;
  assign n51176 = pi18 ? n32 : n51175;
  assign n51177 = pi17 ? n32 : n51176;
  assign n51178 = pi16 ? n51177 : ~n51038;
  assign n51179 = pi15 ? n51036 : n51178;
  assign n51180 = pi17 ? n37443 : n21317;
  assign n51181 = pi16 ? n32 : n51180;
  assign n51182 = pi20 ? n749 : ~n342;
  assign n51183 = pi19 ? n51182 : n5707;
  assign n51184 = pi18 ? n32 : n51183;
  assign n51185 = pi17 ? n32 : n51184;
  assign n51186 = pi16 ? n51185 : n32;
  assign n51187 = pi15 ? n51181 : n51186;
  assign n51188 = pi14 ? n51179 : n51187;
  assign n51189 = pi13 ? n51174 : n51188;
  assign n51190 = pi12 ? n51168 : n51189;
  assign n51191 = pi11 ? n51155 : n51190;
  assign n51192 = pi10 ? n51110 : n51191;
  assign n51193 = pi09 ? n51064 : n51192;
  assign n51194 = pi08 ? n51053 : n51193;
  assign n51195 = pi07 ? n50908 : n51194;
  assign n51196 = pi06 ? n50687 : n51195;
  assign n51197 = pi05 ? n50312 : n51196;
  assign n51198 = pi14 ? n17112 : n37719;
  assign n51199 = pi13 ? n32 : n51198;
  assign n51200 = pi12 ? n32 : n51199;
  assign n51201 = pi11 ? n32 : n51200;
  assign n51202 = pi10 ? n32 : n51201;
  assign n51203 = pi19 ? n1464 : n5707;
  assign n51204 = pi18 ? n32 : n51203;
  assign n51205 = pi17 ? n32 : n51204;
  assign n51206 = pi16 ? n32 : n51205;
  assign n51207 = pi15 ? n16832 : n51206;
  assign n51208 = pi19 ? n32 : ~n9345;
  assign n51209 = pi18 ? n32 : n51208;
  assign n51210 = pi17 ? n32 : n51209;
  assign n51211 = pi16 ? n32 : n51210;
  assign n51212 = pi15 ? n14985 : n51211;
  assign n51213 = pi14 ? n51207 : n51212;
  assign n51214 = pi19 ? n507 : n13074;
  assign n51215 = pi18 ? n32 : n51214;
  assign n51216 = pi17 ? n32 : n51215;
  assign n51217 = pi16 ? n32 : n51216;
  assign n51218 = pi15 ? n51217 : n16485;
  assign n51219 = pi15 ? n16485 : n16392;
  assign n51220 = pi14 ? n51218 : n51219;
  assign n51221 = pi13 ? n51213 : n51220;
  assign n51222 = pi15 ? n16392 : n24874;
  assign n51223 = pi19 ? n594 : n10645;
  assign n51224 = pi18 ? n32 : n51223;
  assign n51225 = pi17 ? n32 : n51224;
  assign n51226 = pi16 ? n32 : n51225;
  assign n51227 = pi19 ? n594 : n5707;
  assign n51228 = pi18 ? n32 : n51227;
  assign n51229 = pi17 ? n32 : n51228;
  assign n51230 = pi16 ? n32 : n51229;
  assign n51231 = pi15 ? n51226 : n51230;
  assign n51232 = pi14 ? n51222 : n51231;
  assign n51233 = pi15 ? n16392 : n17036;
  assign n51234 = pi14 ? n51233 : n32;
  assign n51235 = pi13 ? n51232 : n51234;
  assign n51236 = pi12 ? n51221 : n51235;
  assign n51237 = pi15 ? n37644 : n36296;
  assign n51238 = pi14 ? n32 : n51237;
  assign n51239 = pi13 ? n32 : n51238;
  assign n51240 = pi12 ? n32 : n51239;
  assign n51241 = pi11 ? n51236 : n51240;
  assign n51242 = pi15 ? n23933 : n14696;
  assign n51243 = pi19 ? n1757 : n4342;
  assign n51244 = pi18 ? n51243 : ~n496;
  assign n51245 = pi17 ? n3282 : n51244;
  assign n51246 = pi16 ? n32 : n51245;
  assign n51247 = pi18 ? n32 : n5747;
  assign n51248 = pi17 ? n32 : n51247;
  assign n51249 = pi16 ? n32 : n51248;
  assign n51250 = pi15 ? n51246 : n51249;
  assign n51251 = pi14 ? n51242 : n51250;
  assign n51252 = pi18 ? n863 : ~n496;
  assign n51253 = pi17 ? n26267 : n51252;
  assign n51254 = pi16 ? n32 : n51253;
  assign n51255 = pi21 ? n174 : ~n173;
  assign n51256 = pi20 ? n32 : n51255;
  assign n51257 = pi19 ? n32 : n51256;
  assign n51258 = pi18 ? n32 : n51257;
  assign n51259 = pi18 ? n32255 : ~n496;
  assign n51260 = pi17 ? n51258 : n51259;
  assign n51261 = pi16 ? n32 : n51260;
  assign n51262 = pi15 ? n51254 : n51261;
  assign n51263 = pi19 ? n6298 : n236;
  assign n51264 = pi18 ? n51263 : ~n496;
  assign n51265 = pi17 ? n32 : n51264;
  assign n51266 = pi16 ? n32 : n51265;
  assign n51267 = pi18 ? n359 : n496;
  assign n51268 = pi17 ? n32 : ~n51267;
  assign n51269 = pi16 ? n32 : n51268;
  assign n51270 = pi15 ? n51266 : n51269;
  assign n51271 = pi14 ? n51262 : n51270;
  assign n51272 = pi13 ? n51251 : n51271;
  assign n51273 = pi17 ? n3292 : ~n2736;
  assign n51274 = pi16 ? n32 : n51273;
  assign n51275 = pi20 ? n18253 : n18261;
  assign n51276 = pi19 ? n51275 : ~n501;
  assign n51277 = pi18 ? n51276 : n37418;
  assign n51278 = pi17 ? n19886 : ~n51277;
  assign n51279 = pi16 ? n32 : n51278;
  assign n51280 = pi15 ? n51274 : n51279;
  assign n51281 = pi19 ? n32 : n31941;
  assign n51282 = pi19 ? n24218 : ~n236;
  assign n51283 = pi18 ? n51281 : n51282;
  assign n51284 = pi17 ? n32 : n51283;
  assign n51285 = pi16 ? n32 : n51284;
  assign n51286 = pi18 ? n4380 : n5725;
  assign n51287 = pi17 ? n32 : n51286;
  assign n51288 = pi16 ? n32 : n51287;
  assign n51289 = pi15 ? n51285 : n51288;
  assign n51290 = pi14 ? n51280 : n51289;
  assign n51291 = pi18 ? n1819 : n6132;
  assign n51292 = pi17 ? n32 : n51291;
  assign n51293 = pi16 ? n32 : n51292;
  assign n51294 = pi18 ? n12368 : ~n37510;
  assign n51295 = pi17 ? n32 : n51294;
  assign n51296 = pi16 ? n32 : n51295;
  assign n51297 = pi15 ? n51293 : n51296;
  assign n51298 = pi19 ? n28926 : ~n4721;
  assign n51299 = pi18 ? n32 : n51298;
  assign n51300 = pi17 ? n32 : n51299;
  assign n51301 = pi18 ? n4127 : n6405;
  assign n51302 = pi17 ? n32 : n51301;
  assign n51303 = pi16 ? n51300 : n51302;
  assign n51304 = pi15 ? n24018 : n51303;
  assign n51305 = pi14 ? n51297 : n51304;
  assign n51306 = pi13 ? n51290 : n51305;
  assign n51307 = pi12 ? n51272 : n51306;
  assign n51308 = pi18 ? n863 : n9012;
  assign n51309 = pi17 ? n32 : n51308;
  assign n51310 = pi16 ? n32 : n51309;
  assign n51311 = pi15 ? n51310 : n32;
  assign n51312 = pi14 ? n51311 : n22543;
  assign n51313 = pi13 ? n51312 : n51167;
  assign n51314 = pi18 ? n12368 : n237;
  assign n51315 = pi17 ? n32 : n51314;
  assign n51316 = pi16 ? n32 : ~n51315;
  assign n51317 = pi15 ? n32 : n51316;
  assign n51318 = pi14 ? n51166 : n51317;
  assign n51319 = pi16 ? n32 : ~n4394;
  assign n51320 = pi16 ? n2530 : ~n4060;
  assign n51321 = pi15 ? n51319 : n51320;
  assign n51322 = pi17 ? n32 : n45911;
  assign n51323 = pi16 ? n51322 : n21318;
  assign n51324 = pi16 ? n2320 : n21318;
  assign n51325 = pi15 ? n51323 : n51324;
  assign n51326 = pi14 ? n51321 : n51325;
  assign n51327 = pi13 ? n51318 : n51326;
  assign n51328 = pi12 ? n51313 : n51327;
  assign n51329 = pi11 ? n51307 : n51328;
  assign n51330 = pi10 ? n51241 : n51329;
  assign n51331 = pi09 ? n51202 : n51330;
  assign n51332 = pi14 ? n16985 : n37719;
  assign n51333 = pi13 ? n32 : n51332;
  assign n51334 = pi12 ? n32 : n51333;
  assign n51335 = pi11 ? n32 : n51334;
  assign n51336 = pi10 ? n32 : n51335;
  assign n51337 = pi15 ? n16392 : n51206;
  assign n51338 = pi19 ? n32 : ~n33215;
  assign n51339 = pi18 ? n32 : n51338;
  assign n51340 = pi17 ? n32 : n51339;
  assign n51341 = pi16 ? n32 : n51340;
  assign n51342 = pi15 ? n14985 : n51341;
  assign n51343 = pi14 ? n51337 : n51342;
  assign n51344 = pi15 ? n51217 : n25708;
  assign n51345 = pi15 ? n25708 : n16832;
  assign n51346 = pi14 ? n51344 : n51345;
  assign n51347 = pi13 ? n51343 : n51346;
  assign n51348 = pi15 ? n16832 : n24874;
  assign n51349 = pi14 ? n51348 : n51231;
  assign n51350 = pi14 ? n51233 : n17189;
  assign n51351 = pi13 ? n51349 : n51350;
  assign n51352 = pi12 ? n51347 : n51351;
  assign n51353 = pi11 ? n51352 : n51240;
  assign n51354 = pi18 ? n51243 : ~n590;
  assign n51355 = pi17 ? n32 : n51354;
  assign n51356 = pi16 ? n32 : n51355;
  assign n51357 = pi18 ? n32 : n37376;
  assign n51358 = pi17 ? n32 : n51357;
  assign n51359 = pi16 ? n32 : n51358;
  assign n51360 = pi15 ? n51356 : n51359;
  assign n51361 = pi14 ? n51242 : n51360;
  assign n51362 = pi18 ? n863 : ~n590;
  assign n51363 = pi17 ? n32 : n51362;
  assign n51364 = pi16 ? n32 : n51363;
  assign n51365 = pi18 ? n32 : n44259;
  assign n51366 = pi17 ? n51365 : n51259;
  assign n51367 = pi16 ? n32 : n51366;
  assign n51368 = pi15 ? n51364 : n51367;
  assign n51369 = pi15 ? n51266 : n10424;
  assign n51370 = pi14 ? n51368 : n51369;
  assign n51371 = pi13 ? n51361 : n51370;
  assign n51372 = pi20 ? n3843 : ~n18261;
  assign n51373 = pi19 ? n51372 : n501;
  assign n51374 = pi18 ? n51373 : ~n37418;
  assign n51375 = pi17 ? n19886 : n51374;
  assign n51376 = pi16 ? n32 : n51375;
  assign n51377 = pi15 ? n9952 : n51376;
  assign n51378 = pi19 ? n24218 : ~n813;
  assign n51379 = pi18 ? n51281 : n51378;
  assign n51380 = pi17 ? n32 : n51379;
  assign n51381 = pi16 ? n32 : n51380;
  assign n51382 = pi15 ? n51381 : n51288;
  assign n51383 = pi14 ? n51377 : n51382;
  assign n51384 = pi18 ? n1819 : n37589;
  assign n51385 = pi17 ? n32 : n51384;
  assign n51386 = pi16 ? n32 : n51385;
  assign n51387 = pi18 ? n12368 : ~n37593;
  assign n51388 = pi17 ? n32 : n51387;
  assign n51389 = pi16 ? n32 : n51388;
  assign n51390 = pi15 ? n51386 : n51389;
  assign n51391 = pi20 ? n2140 : n342;
  assign n51392 = pi19 ? n51391 : ~n4721;
  assign n51393 = pi18 ? n32 : n51392;
  assign n51394 = pi17 ? n32 : n51393;
  assign n51395 = pi16 ? n51394 : n51302;
  assign n51396 = pi15 ? n24018 : n51395;
  assign n51397 = pi14 ? n51390 : n51396;
  assign n51398 = pi13 ? n51383 : n51397;
  assign n51399 = pi12 ? n51371 : n51398;
  assign n51400 = pi16 ? n2426 : ~n4060;
  assign n51401 = pi15 ? n51319 : n51400;
  assign n51402 = pi16 ? n2654 : n21318;
  assign n51403 = pi15 ? n51323 : n51402;
  assign n51404 = pi14 ? n51401 : n51403;
  assign n51405 = pi13 ? n51318 : n51404;
  assign n51406 = pi12 ? n51313 : n51405;
  assign n51407 = pi11 ? n51399 : n51406;
  assign n51408 = pi10 ? n51353 : n51407;
  assign n51409 = pi09 ? n51336 : n51408;
  assign n51410 = pi08 ? n51331 : n51409;
  assign n51411 = pi14 ? n25557 : n26684;
  assign n51412 = pi13 ? n32 : n51411;
  assign n51413 = pi12 ? n32 : n51412;
  assign n51414 = pi11 ? n32 : n51413;
  assign n51415 = pi10 ? n32 : n51414;
  assign n51416 = pi15 ? n16984 : n15139;
  assign n51417 = pi14 ? n51416 : n25291;
  assign n51418 = pi20 ? n518 : n125;
  assign n51419 = pi19 ? n32 : n51418;
  assign n51420 = pi18 ? n32 : n51419;
  assign n51421 = pi17 ? n32 : n51420;
  assign n51422 = pi16 ? n32 : n51421;
  assign n51423 = pi15 ? n51422 : n25704;
  assign n51424 = pi14 ? n51423 : n26330;
  assign n51425 = pi13 ? n51417 : n51424;
  assign n51426 = pi15 ? n15847 : n16485;
  assign n51427 = pi14 ? n32 : n51426;
  assign n51428 = pi15 ? n16832 : n32;
  assign n51429 = pi15 ? n32 : n36851;
  assign n51430 = pi14 ? n51428 : n51429;
  assign n51431 = pi13 ? n51427 : n51430;
  assign n51432 = pi12 ? n51425 : n51431;
  assign n51433 = pi14 ? n24627 : n37644;
  assign n51434 = pi13 ? n32 : n51433;
  assign n51435 = pi12 ? n32 : n51434;
  assign n51436 = pi11 ? n51432 : n51435;
  assign n51437 = pi18 ? n15844 : ~n590;
  assign n51438 = pi17 ? n32 : n51437;
  assign n51439 = pi16 ? n32 : n51438;
  assign n51440 = pi15 ? n51439 : n51359;
  assign n51441 = pi14 ? n37649 : n51440;
  assign n51442 = pi18 ? n32 : ~n496;
  assign n51443 = pi17 ? n32 : n51442;
  assign n51444 = pi16 ? n32 : n51443;
  assign n51445 = pi18 ? n7889 : ~n496;
  assign n51446 = pi17 ? n32 : n51445;
  assign n51447 = pi16 ? n32 : n51446;
  assign n51448 = pi15 ? n51444 : n51447;
  assign n51449 = pi19 ? n1464 : n343;
  assign n51450 = pi18 ? n51449 : ~n496;
  assign n51451 = pi17 ? n32 : n51450;
  assign n51452 = pi16 ? n32 : n51451;
  assign n51453 = pi18 ? n323 : ~n2849;
  assign n51454 = pi17 ? n32 : n51453;
  assign n51455 = pi16 ? n32 : n51454;
  assign n51456 = pi15 ? n51452 : n51455;
  assign n51457 = pi14 ? n51448 : n51456;
  assign n51458 = pi13 ? n51441 : n51457;
  assign n51459 = pi17 ? n23052 : n36495;
  assign n51460 = pi16 ? n32 : n51459;
  assign n51461 = pi19 ? n8818 : ~n236;
  assign n51462 = pi18 ? n32 : n51461;
  assign n51463 = pi17 ? n32 : n51462;
  assign n51464 = pi16 ? n32 : n51463;
  assign n51465 = pi15 ? n51460 : n51464;
  assign n51466 = pi19 ? n5688 : ~n813;
  assign n51467 = pi18 ? n940 : n51466;
  assign n51468 = pi17 ? n32 : n51467;
  assign n51469 = pi16 ? n32 : n51468;
  assign n51470 = pi15 ? n51469 : n35701;
  assign n51471 = pi14 ? n51465 : n51470;
  assign n51472 = pi18 ? n4380 : n6132;
  assign n51473 = pi17 ? n32 : n51472;
  assign n51474 = pi16 ? n32 : n51473;
  assign n51475 = pi15 ? n35393 : n51474;
  assign n51476 = pi19 ? n519 : ~n5694;
  assign n51477 = pi18 ? n32 : n51476;
  assign n51478 = pi17 ? n32 : n51477;
  assign n51479 = pi18 ? n863 : n6405;
  assign n51480 = pi17 ? n32 : n51479;
  assign n51481 = pi16 ? n51478 : n51480;
  assign n51482 = pi15 ? n35452 : n51481;
  assign n51483 = pi14 ? n51475 : n51482;
  assign n51484 = pi13 ? n51471 : n51483;
  assign n51485 = pi12 ? n51458 : n51484;
  assign n51486 = pi13 ? n36305 : n32;
  assign n51487 = pi17 ? n1028 : ~n31073;
  assign n51488 = pi16 ? n32 : n51487;
  assign n51489 = pi15 ? n32 : n51488;
  assign n51490 = pi14 ? n32 : n51489;
  assign n51491 = pi17 ? n1028 : ~n4393;
  assign n51492 = pi16 ? n32 : n51491;
  assign n51493 = pi16 ? n2518 : ~n4060;
  assign n51494 = pi15 ? n51492 : n51493;
  assign n51495 = pi16 ? n2513 : ~n1029;
  assign n51496 = pi16 ? n2293 : n14396;
  assign n51497 = pi15 ? n51495 : n51496;
  assign n51498 = pi14 ? n51494 : n51497;
  assign n51499 = pi13 ? n51490 : n51498;
  assign n51500 = pi12 ? n51486 : n51499;
  assign n51501 = pi11 ? n51485 : n51500;
  assign n51502 = pi10 ? n51436 : n51501;
  assign n51503 = pi09 ? n51415 : n51502;
  assign n51504 = pi15 ? n16485 : n16832;
  assign n51505 = pi14 ? n51416 : n51504;
  assign n51506 = pi20 ? n518 : ~n243;
  assign n51507 = pi19 ? n32 : n51506;
  assign n51508 = pi18 ? n32 : n51507;
  assign n51509 = pi17 ? n32 : n51508;
  assign n51510 = pi16 ? n32 : n51509;
  assign n51511 = pi15 ? n25704 : n51510;
  assign n51512 = pi14 ? n51511 : n25815;
  assign n51513 = pi13 ? n51505 : n51512;
  assign n51514 = pi14 ? n32 : n15847;
  assign n51515 = pi15 ? n25763 : n16984;
  assign n51516 = pi14 ? n51515 : n17412;
  assign n51517 = pi13 ? n51514 : n51516;
  assign n51518 = pi12 ? n51513 : n51517;
  assign n51519 = pi14 ? n32 : n37644;
  assign n51520 = pi13 ? n32 : n51519;
  assign n51521 = pi12 ? n32 : n51520;
  assign n51522 = pi11 ? n51518 : n51521;
  assign n51523 = pi14 ? n37735 : n51440;
  assign n51524 = pi18 ? n323 : ~n496;
  assign n51525 = pi17 ? n32 : n51524;
  assign n51526 = pi16 ? n32 : n51525;
  assign n51527 = pi15 ? n51452 : n51526;
  assign n51528 = pi14 ? n51448 : n51527;
  assign n51529 = pi13 ? n51523 : n51528;
  assign n51530 = pi19 ? n1840 : ~n5694;
  assign n51531 = pi18 ? n32 : n51530;
  assign n51532 = pi17 ? n32 : n51531;
  assign n51533 = pi16 ? n51532 : n51480;
  assign n51534 = pi15 ? n35452 : n51533;
  assign n51535 = pi14 ? n51475 : n51534;
  assign n51536 = pi13 ? n51471 : n51535;
  assign n51537 = pi12 ? n51529 : n51536;
  assign n51538 = pi16 ? n4100 : ~n4060;
  assign n51539 = pi15 ? n51492 : n51538;
  assign n51540 = pi16 ? n2860 : n14396;
  assign n51541 = pi15 ? n51495 : n51540;
  assign n51542 = pi14 ? n51539 : n51541;
  assign n51543 = pi13 ? n51490 : n51542;
  assign n51544 = pi12 ? n51486 : n51543;
  assign n51545 = pi11 ? n51537 : n51544;
  assign n51546 = pi10 ? n51522 : n51545;
  assign n51547 = pi09 ? n51415 : n51546;
  assign n51548 = pi08 ? n51503 : n51547;
  assign n51549 = pi07 ? n51410 : n51548;
  assign n51550 = pi13 ? n32 : n25755;
  assign n51551 = pi12 ? n32 : n51550;
  assign n51552 = pi11 ? n32 : n51551;
  assign n51553 = pi10 ? n32 : n51552;
  assign n51554 = pi14 ? n15848 : n25291;
  assign n51555 = pi19 ? n32 : n23406;
  assign n51556 = pi18 ? n32 : n51555;
  assign n51557 = pi17 ? n32 : n51556;
  assign n51558 = pi16 ? n32 : n51557;
  assign n51559 = pi15 ? n51558 : n25563;
  assign n51560 = pi15 ? n25563 : n25763;
  assign n51561 = pi14 ? n51559 : n51560;
  assign n51562 = pi13 ? n51554 : n51561;
  assign n51563 = pi18 ? n32 : n28987;
  assign n51564 = pi17 ? n32 : n51563;
  assign n51565 = pi16 ? n32 : n51564;
  assign n51566 = pi15 ? n16546 : n51565;
  assign n51567 = pi14 ? n16392 : n51566;
  assign n51568 = pi14 ? n16984 : n32;
  assign n51569 = pi13 ? n51567 : n51568;
  assign n51570 = pi12 ? n51562 : n51569;
  assign n51571 = pi13 ? n32 : n17375;
  assign n51572 = pi14 ? n32 : n37781;
  assign n51573 = pi13 ? n32 : n51572;
  assign n51574 = pi12 ? n51571 : n51573;
  assign n51575 = pi11 ? n51570 : n51574;
  assign n51576 = pi19 ? n18478 : ~n349;
  assign n51577 = pi18 ? n32 : n51576;
  assign n51578 = pi17 ? n32 : n51577;
  assign n51579 = pi16 ? n32 : n51578;
  assign n51580 = pi15 ? n15244 : n51579;
  assign n51581 = pi14 ? n37786 : n51580;
  assign n51582 = pi19 ? n1757 : n589;
  assign n51583 = pi18 ? n32 : ~n51582;
  assign n51584 = pi17 ? n32 : n51583;
  assign n51585 = pi16 ? n32 : n51584;
  assign n51586 = pi15 ? n12556 : n51585;
  assign n51587 = pi15 ? n51359 : n51249;
  assign n51588 = pi14 ? n51586 : n51587;
  assign n51589 = pi13 ? n51581 : n51588;
  assign n51590 = pi18 ? n13945 : n28433;
  assign n51591 = pi17 ? n32 : n51590;
  assign n51592 = pi16 ? n32 : n51591;
  assign n51593 = pi15 ? n51592 : n14917;
  assign n51594 = pi15 ? n14570 : n24659;
  assign n51595 = pi14 ? n51593 : n51594;
  assign n51596 = pi15 ? n24659 : n35030;
  assign n51597 = pi19 ? n32 : n51182;
  assign n51598 = pi18 ? n32 : n51597;
  assign n51599 = pi17 ? n32 : n51598;
  assign n51600 = pi17 ? n1227 : ~n25596;
  assign n51601 = pi16 ? n51599 : ~n51600;
  assign n51602 = pi15 ? n51601 : n24742;
  assign n51603 = pi14 ? n51596 : n51602;
  assign n51604 = pi13 ? n51595 : n51603;
  assign n51605 = pi12 ? n51589 : n51604;
  assign n51606 = pi19 ? n4126 : n1757;
  assign n51607 = pi18 ? n51606 : n32;
  assign n51608 = pi17 ? n32 : n51607;
  assign n51609 = pi16 ? n32 : n51608;
  assign n51610 = pi15 ? n32 : n51609;
  assign n51611 = pi14 ? n51610 : n32;
  assign n51612 = pi13 ? n32 : n51611;
  assign n51613 = pi20 ? n17652 : n17665;
  assign n51614 = pi19 ? n975 : n51613;
  assign n51615 = pi18 ? n51614 : n21194;
  assign n51616 = pi17 ? n32 : n51615;
  assign n51617 = pi16 ? n32 : n51616;
  assign n51618 = pi18 ? n32 : n21350;
  assign n51619 = pi17 ? n2355 : ~n51618;
  assign n51620 = pi16 ? n32 : n51619;
  assign n51621 = pi15 ? n51617 : n51620;
  assign n51622 = pi14 ? n32 : n51621;
  assign n51623 = pi17 ? n37834 : n34522;
  assign n51624 = pi16 ? n3165 : ~n51623;
  assign n51625 = pi18 ? n32 : n31959;
  assign n51626 = pi17 ? n32 : n51625;
  assign n51627 = pi16 ? n2745 : ~n51626;
  assign n51628 = pi15 ? n51624 : n51627;
  assign n51629 = pi17 ? n37834 : n32;
  assign n51630 = pi16 ? n15408 : n51629;
  assign n51631 = pi17 ? n1215 : ~n21317;
  assign n51632 = pi16 ? n2745 : ~n51631;
  assign n51633 = pi15 ? n51630 : n51632;
  assign n51634 = pi14 ? n51628 : n51633;
  assign n51635 = pi13 ? n51622 : n51634;
  assign n51636 = pi12 ? n51612 : n51635;
  assign n51637 = pi11 ? n51605 : n51636;
  assign n51638 = pi10 ? n51575 : n51637;
  assign n51639 = pi09 ? n51553 : n51638;
  assign n51640 = pi15 ? n25556 : n15847;
  assign n51641 = pi19 ? n32 : n21723;
  assign n51642 = pi18 ? n32 : n51641;
  assign n51643 = pi17 ? n32 : n51642;
  assign n51644 = pi16 ? n32 : n51643;
  assign n51645 = pi15 ? n15847 : n51644;
  assign n51646 = pi14 ? n51640 : n51645;
  assign n51647 = pi15 ? n51558 : n17121;
  assign n51648 = pi15 ? n17121 : n25763;
  assign n51649 = pi14 ? n51647 : n51648;
  assign n51650 = pi13 ? n51646 : n51649;
  assign n51651 = pi14 ? n25630 : n32;
  assign n51652 = pi13 ? n51567 : n51651;
  assign n51653 = pi12 ? n51650 : n51652;
  assign n51654 = pi12 ? n32 : n51573;
  assign n51655 = pi11 ? n51653 : n51654;
  assign n51656 = pi15 ? n51601 : n25657;
  assign n51657 = pi14 ? n51596 : n51656;
  assign n51658 = pi13 ? n51595 : n51657;
  assign n51659 = pi12 ? n51589 : n51658;
  assign n51660 = pi20 ? n339 : ~n4279;
  assign n51661 = pi19 ? n975 : n51660;
  assign n51662 = pi18 ? n51661 : ~n18891;
  assign n51663 = pi17 ? n32 : n51662;
  assign n51664 = pi16 ? n32 : n51663;
  assign n51665 = pi15 ? n51664 : n51620;
  assign n51666 = pi14 ? n32 : n51665;
  assign n51667 = pi17 ? n37886 : n34522;
  assign n51668 = pi16 ? n3165 : ~n51667;
  assign n51669 = pi16 ? n2851 : ~n51626;
  assign n51670 = pi15 ? n51668 : n51669;
  assign n51671 = pi17 ? n37886 : n32;
  assign n51672 = pi16 ? n16396 : n51671;
  assign n51673 = pi16 ? n2837 : ~n51631;
  assign n51674 = pi15 ? n51672 : n51673;
  assign n51675 = pi14 ? n51670 : n51674;
  assign n51676 = pi13 ? n51666 : n51675;
  assign n51677 = pi12 ? n51612 : n51676;
  assign n51678 = pi11 ? n51659 : n51677;
  assign n51679 = pi10 ? n51655 : n51678;
  assign n51680 = pi09 ? n51553 : n51679;
  assign n51681 = pi08 ? n51639 : n51680;
  assign n51682 = pi13 ? n32 : n26048;
  assign n51683 = pi12 ? n32 : n51682;
  assign n51684 = pi11 ? n32 : n51683;
  assign n51685 = pi10 ? n32 : n51684;
  assign n51686 = pi15 ? n16392 : n17435;
  assign n51687 = pi14 ? n38060 : n51686;
  assign n51688 = pi15 ? n17435 : n17121;
  assign n51689 = pi15 ? n17121 : n25814;
  assign n51690 = pi14 ? n51688 : n51689;
  assign n51691 = pi13 ? n51687 : n51690;
  assign n51692 = pi15 ? n25708 : n25763;
  assign n51693 = pi14 ? n51692 : n25763;
  assign n51694 = pi14 ? n25625 : n32;
  assign n51695 = pi13 ? n51693 : n51694;
  assign n51696 = pi12 ? n51691 : n51695;
  assign n51697 = pi13 ? n38696 : n32;
  assign n51698 = pi14 ? n24498 : n37915;
  assign n51699 = pi13 ? n24564 : n51698;
  assign n51700 = pi12 ? n51697 : n51699;
  assign n51701 = pi11 ? n51696 : n51700;
  assign n51702 = pi19 ? n321 : ~n343;
  assign n51703 = pi18 ? n32 : n51702;
  assign n51704 = pi17 ? n32 : n51703;
  assign n51705 = pi16 ? n32 : n51704;
  assign n51706 = pi15 ? n15230 : n51705;
  assign n51707 = pi14 ? n37924 : n51706;
  assign n51708 = pi15 ? n14016 : n51359;
  assign n51709 = pi19 ? n4391 : ~n589;
  assign n51710 = pi18 ? n32 : n51709;
  assign n51711 = pi17 ? n32 : n51710;
  assign n51712 = pi16 ? n32 : n51711;
  assign n51713 = pi15 ? n51359 : n51712;
  assign n51714 = pi14 ? n51708 : n51713;
  assign n51715 = pi13 ? n51707 : n51714;
  assign n51716 = pi15 ? n37190 : n14917;
  assign n51717 = pi15 ? n37190 : n24659;
  assign n51718 = pi14 ? n51716 : n51717;
  assign n51719 = pi15 ? n23443 : n24659;
  assign n51720 = pi15 ? n24659 : n22817;
  assign n51721 = pi14 ? n51719 : n51720;
  assign n51722 = pi13 ? n51718 : n51721;
  assign n51723 = pi12 ? n51715 : n51722;
  assign n51724 = pi18 ? n37954 : ~n6059;
  assign n51725 = pi17 ? n37953 : ~n51724;
  assign n51726 = pi16 ? n32 : n51725;
  assign n51727 = pi17 ? n1718 : ~n2119;
  assign n51728 = pi16 ? n32 : n51727;
  assign n51729 = pi15 ? n51726 : n51728;
  assign n51730 = pi14 ? n32 : n51729;
  assign n51731 = pi16 ? n4578 : ~n1934;
  assign n51732 = pi16 ? n2958 : ~n3625;
  assign n51733 = pi15 ? n51731 : n51732;
  assign n51734 = pi15 ? n32 : n37959;
  assign n51735 = pi14 ? n51733 : n51734;
  assign n51736 = pi13 ? n51730 : n51735;
  assign n51737 = pi12 ? n51612 : n51736;
  assign n51738 = pi11 ? n51723 : n51737;
  assign n51739 = pi10 ? n51701 : n51738;
  assign n51740 = pi09 ? n51685 : n51739;
  assign n51741 = pi15 ? n17298 : n17261;
  assign n51742 = pi15 ? n17261 : n25997;
  assign n51743 = pi14 ? n51741 : n51742;
  assign n51744 = pi13 ? n51687 : n51743;
  assign n51745 = pi15 ? n16237 : n25763;
  assign n51746 = pi14 ? n51745 : n25763;
  assign n51747 = pi14 ? n25693 : n32;
  assign n51748 = pi13 ? n51746 : n51747;
  assign n51749 = pi12 ? n51744 : n51748;
  assign n51750 = pi14 ? n32 : n24563;
  assign n51751 = pi14 ? n24498 : n37990;
  assign n51752 = pi13 ? n51750 : n51751;
  assign n51753 = pi12 ? n32 : n51752;
  assign n51754 = pi11 ? n51749 : n51753;
  assign n51755 = pi14 ? n37999 : n51706;
  assign n51756 = pi19 ? n4391 : ~n2317;
  assign n51757 = pi18 ? n32 : n51756;
  assign n51758 = pi17 ? n32 : n51757;
  assign n51759 = pi16 ? n32 : n51758;
  assign n51760 = pi15 ? n51359 : n51759;
  assign n51761 = pi14 ? n51708 : n51760;
  assign n51762 = pi13 ? n51755 : n51761;
  assign n51763 = pi18 ? n16603 : n14553;
  assign n51764 = pi17 ? n32 : n51763;
  assign n51765 = pi16 ? n32 : n51764;
  assign n51766 = pi15 ? n51765 : n14917;
  assign n51767 = pi14 ? n51766 : n51717;
  assign n51768 = pi13 ? n51767 : n51721;
  assign n51769 = pi12 ? n51762 : n51768;
  assign n51770 = pi19 ? n4126 : n39001;
  assign n51771 = pi18 ? n51770 : n32;
  assign n51772 = pi17 ? n32 : n51771;
  assign n51773 = pi16 ? n32 : n51772;
  assign n51774 = pi15 ? n32 : n51773;
  assign n51775 = pi14 ? n51774 : n32;
  assign n51776 = pi13 ? n32 : n51775;
  assign n51777 = pi18 ? n4127 : ~n6059;
  assign n51778 = pi17 ? n37953 : ~n51777;
  assign n51779 = pi16 ? n32 : n51778;
  assign n51780 = pi15 ? n51779 : n51728;
  assign n51781 = pi14 ? n32 : n51780;
  assign n51782 = pi16 ? n3588 : ~n1934;
  assign n51783 = pi16 ? n3165 : ~n3625;
  assign n51784 = pi15 ? n51782 : n51783;
  assign n51785 = pi16 ? n3047 : ~n37958;
  assign n51786 = pi15 ? n32 : n51785;
  assign n51787 = pi14 ? n51784 : n51786;
  assign n51788 = pi13 ? n51781 : n51787;
  assign n51789 = pi12 ? n51776 : n51788;
  assign n51790 = pi11 ? n51769 : n51789;
  assign n51791 = pi10 ? n51754 : n51790;
  assign n51792 = pi09 ? n51685 : n51791;
  assign n51793 = pi08 ? n51740 : n51792;
  assign n51794 = pi07 ? n51681 : n51793;
  assign n51795 = pi06 ? n51549 : n51794;
  assign n51796 = pi15 ? n26479 : n25948;
  assign n51797 = pi14 ? n26147 : n51796;
  assign n51798 = pi13 ? n32 : n51797;
  assign n51799 = pi12 ? n32 : n51798;
  assign n51800 = pi11 ? n32 : n51799;
  assign n51801 = pi10 ? n32 : n51800;
  assign n51802 = pi19 ? n32 : n22019;
  assign n51803 = pi18 ? n32 : n51802;
  assign n51804 = pi17 ? n32 : n51803;
  assign n51805 = pi16 ? n32 : n51804;
  assign n51806 = pi20 ? n1076 : ~n207;
  assign n51807 = pi19 ? n32 : n51806;
  assign n51808 = pi18 ? n32 : n51807;
  assign n51809 = pi17 ? n32 : n51808;
  assign n51810 = pi16 ? n32 : n51809;
  assign n51811 = pi15 ? n51805 : n51810;
  assign n51812 = pi14 ? n51811 : n25133;
  assign n51813 = pi15 ? n17336 : n17261;
  assign n51814 = pi14 ? n51813 : n51742;
  assign n51815 = pi13 ? n51812 : n51814;
  assign n51816 = pi14 ? n27734 : n27678;
  assign n51817 = pi14 ? n38620 : n32;
  assign n51818 = pi13 ? n51816 : n51817;
  assign n51819 = pi12 ? n51815 : n51818;
  assign n51820 = pi15 ? n25563 : n26115;
  assign n51821 = pi14 ? n51820 : n37565;
  assign n51822 = pi13 ? n25558 : n51821;
  assign n51823 = pi15 ? n24874 : n27528;
  assign n51824 = pi14 ? n32 : n51823;
  assign n51825 = pi13 ? n32 : n51824;
  assign n51826 = pi12 ? n51822 : n51825;
  assign n51827 = pi11 ? n51819 : n51826;
  assign n51828 = pi15 ? n27528 : n14651;
  assign n51829 = pi15 ? n14651 : n15230;
  assign n51830 = pi14 ? n51828 : n51829;
  assign n51831 = pi15 ? n50236 : n14207;
  assign n51832 = pi15 ? n14488 : n14917;
  assign n51833 = pi14 ? n51831 : n51832;
  assign n51834 = pi13 ? n51830 : n51833;
  assign n51835 = pi18 ? n268 : n24637;
  assign n51836 = pi17 ? n32 : n51835;
  assign n51837 = pi16 ? n32 : n51836;
  assign n51838 = pi15 ? n51837 : n24511;
  assign n51839 = pi15 ? n15244 : n49496;
  assign n51840 = pi14 ? n51838 : n51839;
  assign n51841 = pi20 ? n3523 : ~n354;
  assign n51842 = pi19 ? n51841 : n6085;
  assign n51843 = pi19 ? n28483 : n38539;
  assign n51844 = pi18 ? n51842 : n51843;
  assign n51845 = pi17 ? n51844 : n25655;
  assign n51846 = pi16 ? n32 : n51845;
  assign n51847 = pi15 ? n14917 : n51846;
  assign n51848 = pi14 ? n51847 : n48187;
  assign n51849 = pi13 ? n51840 : n51848;
  assign n51850 = pi12 ? n51834 : n51849;
  assign n51851 = pi19 ? n32 : ~n5356;
  assign n51852 = pi18 ? n51851 : n32;
  assign n51853 = pi17 ? n32 : n51852;
  assign n51854 = pi16 ? n32 : n51853;
  assign n51855 = pi15 ? n32 : n51854;
  assign n51856 = pi14 ? n51855 : n32;
  assign n51857 = pi13 ? n32 : n51856;
  assign n51858 = pi18 ? n36119 : ~n605;
  assign n51859 = pi17 ? n32 : n51858;
  assign n51860 = pi16 ? n32 : n51859;
  assign n51861 = pi17 ? n38122 : ~n2119;
  assign n51862 = pi16 ? n32 : n51861;
  assign n51863 = pi15 ? n51860 : n51862;
  assign n51864 = pi14 ? n47688 : n51863;
  assign n51865 = pi16 ? n3438 : ~n49156;
  assign n51866 = pi16 ? n32 : ~n49156;
  assign n51867 = pi15 ? n51865 : n51866;
  assign n51868 = pi17 ? n38128 : ~n14154;
  assign n51869 = pi16 ? n3438 : ~n51868;
  assign n51870 = pi15 ? n32 : n51869;
  assign n51871 = pi14 ? n51867 : n51870;
  assign n51872 = pi13 ? n51864 : n51871;
  assign n51873 = pi12 ? n51857 : n51872;
  assign n51874 = pi11 ? n51850 : n51873;
  assign n51875 = pi10 ? n51827 : n51874;
  assign n51876 = pi09 ? n51801 : n51875;
  assign n51877 = pi20 ? n428 : n52;
  assign n51878 = pi19 ? n32 : n51877;
  assign n51879 = pi18 ? n32 : n51878;
  assign n51880 = pi17 ? n32 : n51879;
  assign n51881 = pi16 ? n32 : n51880;
  assign n51882 = pi15 ? n51881 : n17298;
  assign n51883 = pi14 ? n16893 : n51882;
  assign n51884 = pi15 ? n25948 : n26479;
  assign n51885 = pi14 ? n26318 : n51884;
  assign n51886 = pi13 ? n51883 : n51885;
  assign n51887 = pi15 ? n26201 : n16392;
  assign n51888 = pi14 ? n51887 : n27678;
  assign n51889 = pi15 ? n17261 : n17454;
  assign n51890 = pi14 ? n51889 : n25805;
  assign n51891 = pi13 ? n51888 : n51890;
  assign n51892 = pi12 ? n51886 : n51891;
  assign n51893 = pi14 ? n25563 : n17412;
  assign n51894 = pi13 ? n25558 : n51893;
  assign n51895 = pi15 ? n15847 : n14985;
  assign n51896 = pi14 ? n32 : n51895;
  assign n51897 = pi13 ? n32 : n51896;
  assign n51898 = pi12 ? n51894 : n51897;
  assign n51899 = pi11 ? n51892 : n51898;
  assign n51900 = pi15 ? n14985 : n14651;
  assign n51901 = pi14 ? n51900 : n51829;
  assign n51902 = pi15 ? n14651 : n14207;
  assign n51903 = pi15 ? n14207 : n14917;
  assign n51904 = pi14 ? n51902 : n51903;
  assign n51905 = pi13 ? n51901 : n51904;
  assign n51906 = pi18 ? n268 : n24508;
  assign n51907 = pi17 ? n32 : n51906;
  assign n51908 = pi16 ? n32 : n51907;
  assign n51909 = pi15 ? n51908 : n24511;
  assign n51910 = pi15 ? n15244 : n36100;
  assign n51911 = pi14 ? n51909 : n51910;
  assign n51912 = pi20 ? n7839 : ~n9491;
  assign n51913 = pi19 ? n275 : n51912;
  assign n51914 = pi20 ? n1331 : ~n260;
  assign n51915 = pi20 ? n18840 : n309;
  assign n51916 = pi19 ? n51914 : n51915;
  assign n51917 = pi18 ? n51913 : ~n51916;
  assign n51918 = pi17 ? n51917 : ~n25655;
  assign n51919 = pi16 ? n3283 : ~n51918;
  assign n51920 = pi15 ? n14917 : n51919;
  assign n51921 = pi20 ? n974 : ~n518;
  assign n51922 = pi19 ? n51921 : ~n32;
  assign n51923 = pi18 ? n51922 : ~n32;
  assign n51924 = pi17 ? n51923 : ~n19886;
  assign n51925 = pi16 ? n3283 : ~n51924;
  assign n51926 = pi15 ? n51925 : n32;
  assign n51927 = pi14 ? n51920 : n51926;
  assign n51928 = pi13 ? n51911 : n51927;
  assign n51929 = pi12 ? n51905 : n51928;
  assign n51930 = pi20 ? n321 : ~n4279;
  assign n51931 = pi19 ? n32 : ~n51930;
  assign n51932 = pi18 ? n51931 : n32;
  assign n51933 = pi17 ? n32 : n51932;
  assign n51934 = pi16 ? n32 : n51933;
  assign n51935 = pi15 ? n32 : n51934;
  assign n51936 = pi14 ? n51935 : n32;
  assign n51937 = pi13 ? n32 : n51936;
  assign n51938 = pi17 ? n3557 : ~n5779;
  assign n51939 = pi16 ? n32 : n51938;
  assign n51940 = pi17 ? n3719 : ~n5779;
  assign n51941 = pi16 ? n32 : n51940;
  assign n51942 = pi15 ? n51939 : n51941;
  assign n51943 = pi18 ? n41071 : n32;
  assign n51944 = pi17 ? n51943 : n14154;
  assign n51945 = pi16 ? n32 : n51944;
  assign n51946 = pi15 ? n32 : n51945;
  assign n51947 = pi14 ? n51942 : n51946;
  assign n51948 = pi13 ? n51864 : n51947;
  assign n51949 = pi12 ? n51937 : n51948;
  assign n51950 = pi11 ? n51929 : n51949;
  assign n51951 = pi10 ? n51899 : n51950;
  assign n51952 = pi09 ? n51801 : n51951;
  assign n51953 = pi08 ? n51876 : n51952;
  assign n51954 = pi15 ? n32 : n17216;
  assign n51955 = pi15 ? n17056 : n17216;
  assign n51956 = pi14 ? n51954 : n51955;
  assign n51957 = pi13 ? n32 : n51956;
  assign n51958 = pi12 ? n32 : n51957;
  assign n51959 = pi11 ? n32 : n51958;
  assign n51960 = pi10 ? n32 : n51959;
  assign n51961 = pi15 ? n38750 : n16804;
  assign n51962 = pi14 ? n51961 : n26034;
  assign n51963 = pi13 ? n51962 : n51885;
  assign n51964 = pi15 ? n17121 : n16392;
  assign n51965 = pi15 ? n16804 : n32;
  assign n51966 = pi14 ? n51964 : n51965;
  assign n51967 = pi15 ? n17336 : n16984;
  assign n51968 = pi14 ? n51967 : n32;
  assign n51969 = pi13 ? n51966 : n51968;
  assign n51970 = pi12 ? n51963 : n51969;
  assign n51971 = pi14 ? n32 : n38620;
  assign n51972 = pi14 ? n17178 : n32;
  assign n51973 = pi13 ? n51971 : n51972;
  assign n51974 = pi14 ? n17188 : n51895;
  assign n51975 = pi13 ? n32 : n51974;
  assign n51976 = pi12 ? n51973 : n51975;
  assign n51977 = pi11 ? n51970 : n51976;
  assign n51978 = pi15 ? n15403 : n14895;
  assign n51979 = pi15 ? n14895 : n37998;
  assign n51980 = pi14 ? n51978 : n51979;
  assign n51981 = pi15 ? n37998 : n14651;
  assign n51982 = pi15 ? n14651 : n37501;
  assign n51983 = pi14 ? n51981 : n51982;
  assign n51984 = pi13 ? n51980 : n51983;
  assign n51985 = pi15 ? n24640 : n24504;
  assign n51986 = pi14 ? n51985 : n36100;
  assign n51987 = pi19 ? n275 : n1844;
  assign n51988 = pi18 ? n51987 : n32;
  assign n51989 = pi17 ? n51988 : n15242;
  assign n51990 = pi16 ? n32 : n51989;
  assign n51991 = pi18 ? n237 : ~n34006;
  assign n51992 = pi18 ? n20605 : n15359;
  assign n51993 = pi17 ? n51991 : n51992;
  assign n51994 = pi16 ? n32 : n51993;
  assign n51995 = pi15 ? n51990 : n51994;
  assign n51996 = pi14 ? n51995 : n22543;
  assign n51997 = pi13 ? n51986 : n51996;
  assign n51998 = pi12 ? n51984 : n51997;
  assign n51999 = pi19 ? n1785 : n358;
  assign n52000 = pi18 ? n32 : n51999;
  assign n52001 = pi17 ? n32 : n52000;
  assign n52002 = pi16 ? n32 : n52001;
  assign n52003 = pi15 ? n32 : n52002;
  assign n52004 = pi14 ? n22541 : n52003;
  assign n52005 = pi18 ? n51851 : n1541;
  assign n52006 = pi17 ? n32 : n52005;
  assign n52007 = pi16 ? n32 : n52006;
  assign n52008 = pi15 ? n15123 : n52007;
  assign n52009 = pi15 ? n22817 : n38257;
  assign n52010 = pi14 ? n52008 : n52009;
  assign n52011 = pi13 ? n52004 : n52010;
  assign n52012 = pi19 ? n4867 : n32;
  assign n52013 = pi18 ? n32 : n52012;
  assign n52014 = pi17 ? n32 : n52013;
  assign n52015 = pi16 ? n32 : n52014;
  assign n52016 = pi19 ? n28926 : n32;
  assign n52017 = pi18 ? n32 : n52016;
  assign n52018 = pi17 ? n32 : n52017;
  assign n52019 = pi16 ? n32 : n52018;
  assign n52020 = pi15 ? n52015 : n52019;
  assign n52021 = pi19 ? n589 : ~n1844;
  assign n52022 = pi18 ? n52021 : ~n32;
  assign n52023 = pi17 ? n52022 : ~n2119;
  assign n52024 = pi16 ? n32 : n52023;
  assign n52025 = pi15 ? n51860 : n52024;
  assign n52026 = pi14 ? n52020 : n52025;
  assign n52027 = pi17 ? n3704 : ~n2512;
  assign n52028 = pi16 ? n32 : n52027;
  assign n52029 = pi20 ? n1368 : n206;
  assign n52030 = pi19 ? n52029 : ~n32;
  assign n52031 = pi18 ? n32 : n52030;
  assign n52032 = pi17 ? n52022 : ~n52031;
  assign n52033 = pi16 ? n32 : n52032;
  assign n52034 = pi15 ? n52028 : n52033;
  assign n52035 = pi17 ? n38265 : n32;
  assign n52036 = pi16 ? n32 : n52035;
  assign n52037 = pi19 ? n349 : ~n6298;
  assign n52038 = pi18 ? n52037 : n32;
  assign n52039 = pi17 ? n52038 : n14154;
  assign n52040 = pi16 ? n32 : n52039;
  assign n52041 = pi15 ? n52036 : n52040;
  assign n52042 = pi14 ? n52034 : n52041;
  assign n52043 = pi13 ? n52026 : n52042;
  assign n52044 = pi12 ? n52011 : n52043;
  assign n52045 = pi11 ? n51998 : n52044;
  assign n52046 = pi10 ? n51977 : n52045;
  assign n52047 = pi09 ? n51960 : n52046;
  assign n52048 = pi14 ? n51954 : n17216;
  assign n52049 = pi13 ? n32 : n52048;
  assign n52050 = pi12 ? n32 : n52049;
  assign n52051 = pi11 ? n32 : n52050;
  assign n52052 = pi10 ? n32 : n52051;
  assign n52053 = pi15 ? n17039 : n16804;
  assign n52054 = pi14 ? n52053 : n25990;
  assign n52055 = pi15 ? n17216 : n16824;
  assign n52056 = pi14 ? n26761 : n52055;
  assign n52057 = pi13 ? n52054 : n52056;
  assign n52058 = pi14 ? n25905 : n32;
  assign n52059 = pi13 ? n51966 : n52058;
  assign n52060 = pi12 ? n52057 : n52059;
  assign n52061 = pi15 ? n16485 : n14985;
  assign n52062 = pi14 ? n32 : n52061;
  assign n52063 = pi13 ? n32 : n52062;
  assign n52064 = pi12 ? n51973 : n52063;
  assign n52065 = pi11 ? n52060 : n52064;
  assign n52066 = pi15 ? n15403 : n14909;
  assign n52067 = pi19 ? n507 : ~n30701;
  assign n52068 = pi18 ? n32 : n52067;
  assign n52069 = pi17 ? n32 : n52068;
  assign n52070 = pi16 ? n32 : n52069;
  assign n52071 = pi15 ? n14895 : n52070;
  assign n52072 = pi14 ? n52066 : n52071;
  assign n52073 = pi13 ? n52072 : n51983;
  assign n52074 = pi15 ? n24700 : n24504;
  assign n52075 = pi14 ? n52074 : n36100;
  assign n52076 = pi20 ? n518 : ~n820;
  assign n52077 = pi19 ? n52076 : n16304;
  assign n52078 = pi18 ? n52077 : n32;
  assign n52079 = pi17 ? n52078 : n15242;
  assign n52080 = pi16 ? n32 : n52079;
  assign n52081 = pi18 ? n1548 : ~n34006;
  assign n52082 = pi19 ? n7642 : n594;
  assign n52083 = pi18 ? n52082 : n15359;
  assign n52084 = pi17 ? n52081 : n52083;
  assign n52085 = pi16 ? n32 : n52084;
  assign n52086 = pi15 ? n52080 : n52085;
  assign n52087 = pi14 ? n52086 : n22543;
  assign n52088 = pi13 ? n52075 : n52087;
  assign n52089 = pi12 ? n52073 : n52088;
  assign n52090 = pi18 ? n32 : n28317;
  assign n52091 = pi17 ? n32 : n52090;
  assign n52092 = pi16 ? n32 : n52091;
  assign n52093 = pi15 ? n32 : n52092;
  assign n52094 = pi14 ? n22541 : n52093;
  assign n52095 = pi13 ? n52094 : n52010;
  assign n52096 = pi15 ? n52015 : n22817;
  assign n52097 = pi17 ? n3855 : ~n2119;
  assign n52098 = pi16 ? n32 : n52097;
  assign n52099 = pi15 ? n51860 : n52098;
  assign n52100 = pi14 ? n52096 : n52099;
  assign n52101 = pi20 ? n175 : n206;
  assign n52102 = pi19 ? n52101 : ~n32;
  assign n52103 = pi18 ? n32 : n52102;
  assign n52104 = pi17 ? n1219 : ~n52103;
  assign n52105 = pi16 ? n32 : n52104;
  assign n52106 = pi15 ? n5814 : n52105;
  assign n52107 = pi17 ? n38322 : n32;
  assign n52108 = pi16 ? n32 : n52107;
  assign n52109 = pi19 ? n429 : ~n6298;
  assign n52110 = pi18 ? n52109 : n32;
  assign n52111 = pi17 ? n52110 : n14154;
  assign n52112 = pi16 ? n32 : n52111;
  assign n52113 = pi15 ? n52108 : n52112;
  assign n52114 = pi14 ? n52106 : n52113;
  assign n52115 = pi13 ? n52100 : n52114;
  assign n52116 = pi12 ? n52095 : n52115;
  assign n52117 = pi11 ? n52089 : n52116;
  assign n52118 = pi10 ? n52065 : n52117;
  assign n52119 = pi09 ? n52052 : n52118;
  assign n52120 = pi08 ? n52047 : n52119;
  assign n52121 = pi07 ? n51953 : n52120;
  assign n52122 = pi14 ? n26133 : n16850;
  assign n52123 = pi13 ? n32 : n52122;
  assign n52124 = pi12 ? n32 : n52123;
  assign n52125 = pi11 ? n32 : n52124;
  assign n52126 = pi10 ? n32 : n52125;
  assign n52127 = pi14 ? n16804 : n38491;
  assign n52128 = pi15 ? n17056 : n25948;
  assign n52129 = pi14 ? n26824 : n52128;
  assign n52130 = pi13 ? n52127 : n52129;
  assign n52131 = pi13 ? n51971 : n52058;
  assign n52132 = pi12 ? n52130 : n52131;
  assign n52133 = pi14 ? n32 : n25861;
  assign n52134 = pi14 ? n25805 : n32;
  assign n52135 = pi13 ? n52133 : n52134;
  assign n52136 = pi15 ? n16984 : n36851;
  assign n52137 = pi14 ? n32 : n52136;
  assign n52138 = pi15 ? n32 : n16965;
  assign n52139 = pi15 ? n15847 : n15403;
  assign n52140 = pi14 ? n52138 : n52139;
  assign n52141 = pi13 ? n52137 : n52140;
  assign n52142 = pi12 ? n52135 : n52141;
  assign n52143 = pi11 ? n52132 : n52142;
  assign n52144 = pi15 ? n15531 : n27528;
  assign n52145 = pi14 ? n52144 : n50516;
  assign n52146 = pi15 ? n27304 : n15637;
  assign n52147 = pi14 ? n52146 : n15637;
  assign n52148 = pi13 ? n52145 : n52147;
  assign n52149 = pi19 ? n267 : ~n589;
  assign n52150 = pi18 ? n32 : n52149;
  assign n52151 = pi17 ? n32 : n52150;
  assign n52152 = pi16 ? n32 : n52151;
  assign n52153 = pi15 ? n52152 : n24572;
  assign n52154 = pi15 ? n26074 : n24237;
  assign n52155 = pi14 ? n52153 : n52154;
  assign n52156 = pi19 ? n531 : ~n24218;
  assign n52157 = pi18 ? n52156 : n32;
  assign n52158 = pi19 ? n32 : ~n766;
  assign n52159 = pi18 ? n32 : n52158;
  assign n52160 = pi17 ? n52157 : n52159;
  assign n52161 = pi16 ? n32 : n52160;
  assign n52162 = pi18 ? n532 : ~n5657;
  assign n52163 = pi19 ? n4342 : ~n589;
  assign n52164 = pi18 ? n34905 : ~n52163;
  assign n52165 = pi17 ? n52162 : ~n52164;
  assign n52166 = pi16 ? n32 : n52165;
  assign n52167 = pi15 ? n52161 : n52166;
  assign n52168 = pi21 ? n10182 : n32;
  assign n52169 = pi20 ? n52168 : n32;
  assign n52170 = pi19 ? n32 : n52169;
  assign n52171 = pi18 ? n32 : n52170;
  assign n52172 = pi17 ? n32 : n52171;
  assign n52173 = pi16 ? n32 : n52172;
  assign n52174 = pi15 ? n16319 : n52173;
  assign n52175 = pi14 ? n52167 : n52174;
  assign n52176 = pi13 ? n52155 : n52175;
  assign n52177 = pi12 ? n52148 : n52176;
  assign n52178 = pi16 ? n32 : n34080;
  assign n52179 = pi15 ? n52178 : n23250;
  assign n52180 = pi14 ? n24329 : n52179;
  assign n52181 = pi15 ? n21853 : n23443;
  assign n52182 = pi14 ? n23485 : n52181;
  assign n52183 = pi13 ? n52180 : n52182;
  assign n52184 = pi19 ? n46184 : n32;
  assign n52185 = pi18 ? n32 : n52184;
  assign n52186 = pi17 ? n32 : n52185;
  assign n52187 = pi16 ? n32 : n52186;
  assign n52188 = pi15 ? n32 : n52187;
  assign n52189 = pi18 ? n32 : n21888;
  assign n52190 = pi18 ? n23073 : ~n323;
  assign n52191 = pi17 ? n52189 : n52190;
  assign n52192 = pi16 ? n32 : n52191;
  assign n52193 = pi15 ? n52192 : n5803;
  assign n52194 = pi14 ? n52188 : n52193;
  assign n52195 = pi19 ? n750 : ~n28976;
  assign n52196 = pi18 ? n52195 : n38402;
  assign n52197 = pi20 ? n11107 : ~n207;
  assign n52198 = pi19 ? n52197 : n32;
  assign n52199 = pi18 ? n38406 : n52198;
  assign n52200 = pi17 ? n52196 : n52199;
  assign n52201 = pi16 ? n32 : n52200;
  assign n52202 = pi15 ? n5803 : n52201;
  assign n52203 = pi17 ? n464 : n32;
  assign n52204 = pi16 ? n32 : n52203;
  assign n52205 = pi20 ? n749 : ~n206;
  assign n52206 = pi19 ? n208 : n52205;
  assign n52207 = pi18 ? n52206 : n6059;
  assign n52208 = pi17 ? n52207 : n14154;
  assign n52209 = pi16 ? n32 : n52208;
  assign n52210 = pi15 ? n52204 : n52209;
  assign n52211 = pi14 ? n52202 : n52210;
  assign n52212 = pi13 ? n52194 : n52211;
  assign n52213 = pi12 ? n52183 : n52212;
  assign n52214 = pi11 ? n52177 : n52213;
  assign n52215 = pi10 ? n52143 : n52214;
  assign n52216 = pi09 ? n52126 : n52215;
  assign n52217 = pi15 ? n17428 : n32;
  assign n52218 = pi14 ? n16804 : n52217;
  assign n52219 = pi15 ? n17428 : n16736;
  assign n52220 = pi20 ? n175 : ~n749;
  assign n52221 = pi19 ? n32 : n52220;
  assign n52222 = pi18 ? n32 : n52221;
  assign n52223 = pi17 ? n32 : n52222;
  assign n52224 = pi16 ? n32 : n52223;
  assign n52225 = pi15 ? n16736 : n52224;
  assign n52226 = pi14 ? n52219 : n52225;
  assign n52227 = pi13 ? n52218 : n52226;
  assign n52228 = pi14 ? n25989 : n26034;
  assign n52229 = pi13 ? n51971 : n52228;
  assign n52230 = pi12 ? n52227 : n52229;
  assign n52231 = pi15 ? n17111 : n16837;
  assign n52232 = pi14 ? n32 : n52231;
  assign n52233 = pi15 ? n16837 : n16832;
  assign n52234 = pi15 ? n16485 : n25713;
  assign n52235 = pi14 ? n52233 : n52234;
  assign n52236 = pi13 ? n52232 : n52235;
  assign n52237 = pi12 ? n52135 : n52236;
  assign n52238 = pi11 ? n52230 : n52237;
  assign n52239 = pi15 ? n25384 : n50638;
  assign n52240 = pi15 ? n50638 : n27304;
  assign n52241 = pi14 ? n52239 : n52240;
  assign n52242 = pi15 ? n27304 : n27528;
  assign n52243 = pi15 ? n27528 : n15633;
  assign n52244 = pi14 ? n52242 : n52243;
  assign n52245 = pi13 ? n52241 : n52244;
  assign n52246 = pi19 ? n267 : ~n2848;
  assign n52247 = pi18 ? n32 : n52246;
  assign n52248 = pi17 ? n32 : n52247;
  assign n52249 = pi16 ? n32 : n52248;
  assign n52250 = pi15 ? n52249 : n32;
  assign n52251 = pi15 ? n24504 : n24237;
  assign n52252 = pi14 ? n52250 : n52251;
  assign n52253 = pi19 ? n750 : ~n24218;
  assign n52254 = pi18 ? n52253 : n32;
  assign n52255 = pi17 ? n52254 : n52159;
  assign n52256 = pi16 ? n32 : n52255;
  assign n52257 = pi18 ? n797 : ~n5657;
  assign n52258 = pi19 ? n4342 : ~n349;
  assign n52259 = pi18 ? n34905 : ~n52258;
  assign n52260 = pi17 ? n52257 : ~n52259;
  assign n52261 = pi16 ? n32 : n52260;
  assign n52262 = pi15 ? n52256 : n52261;
  assign n52263 = pi15 ? n32 : n52173;
  assign n52264 = pi14 ? n52262 : n52263;
  assign n52265 = pi13 ? n52252 : n52264;
  assign n52266 = pi12 ? n52245 : n52265;
  assign n52267 = pi14 ? n15119 : n52179;
  assign n52268 = pi13 ? n52267 : n52182;
  assign n52269 = pi15 ? n52192 : n5961;
  assign n52270 = pi14 ? n33991 : n52269;
  assign n52271 = pi19 ? n519 : ~n28686;
  assign n52272 = pi18 ? n52271 : n38402;
  assign n52273 = pi17 ? n52272 : n52199;
  assign n52274 = pi16 ? n32 : n52273;
  assign n52275 = pi15 ? n5961 : n52274;
  assign n52276 = pi18 ? n473 : n32;
  assign n52277 = pi17 ? n52276 : n32;
  assign n52278 = pi16 ? n32 : n52277;
  assign n52279 = pi19 ? n519 : n30681;
  assign n52280 = pi18 ? n52279 : n6059;
  assign n52281 = pi17 ? n52280 : n14154;
  assign n52282 = pi16 ? n32 : n52281;
  assign n52283 = pi15 ? n52278 : n52282;
  assign n52284 = pi14 ? n52275 : n52283;
  assign n52285 = pi13 ? n52270 : n52284;
  assign n52286 = pi12 ? n52268 : n52285;
  assign n52287 = pi11 ? n52266 : n52286;
  assign n52288 = pi10 ? n52238 : n52287;
  assign n52289 = pi09 ? n52126 : n52288;
  assign n52290 = pi08 ? n52216 : n52289;
  assign n52291 = pi14 ? n26184 : n26183;
  assign n52292 = pi13 ? n32 : n52291;
  assign n52293 = pi12 ? n32 : n52292;
  assign n52294 = pi11 ? n32 : n52293;
  assign n52295 = pi10 ? n32 : n52294;
  assign n52296 = pi15 ? n16804 : n25948;
  assign n52297 = pi15 ? n26225 : n25904;
  assign n52298 = pi14 ? n52296 : n52297;
  assign n52299 = pi15 ? n16850 : n17428;
  assign n52300 = pi15 ? n17428 : n17121;
  assign n52301 = pi14 ? n52299 : n52300;
  assign n52302 = pi13 ? n52298 : n52301;
  assign n52303 = pi14 ? n26034 : n32;
  assign n52304 = pi13 ? n52058 : n52303;
  assign n52305 = pi12 ? n52302 : n52304;
  assign n52306 = pi14 ? n32 : n25905;
  assign n52307 = pi13 ? n52306 : n52058;
  assign n52308 = pi14 ? n32 : n17412;
  assign n52309 = pi13 ? n52308 : n38506;
  assign n52310 = pi12 ? n52307 : n52309;
  assign n52311 = pi11 ? n52305 : n52310;
  assign n52312 = pi19 ? n32 : ~n6042;
  assign n52313 = pi18 ? n32 : n52312;
  assign n52314 = pi17 ? n32 : n52313;
  assign n52315 = pi16 ? n32 : n52314;
  assign n52316 = pi15 ? n52315 : n16515;
  assign n52317 = pi14 ? n24882 : n52316;
  assign n52318 = pi20 ? n8630 : n32;
  assign n52319 = pi19 ? n32 : n52318;
  assign n52320 = pi18 ? n32 : n52319;
  assign n52321 = pi17 ? n32 : n52320;
  assign n52322 = pi16 ? n32 : n52321;
  assign n52323 = pi21 ? n32 : ~n631;
  assign n52324 = pi20 ? n52323 : ~n32;
  assign n52325 = pi19 ? n32 : ~n52324;
  assign n52326 = pi18 ? n32 : n52325;
  assign n52327 = pi17 ? n32 : n52326;
  assign n52328 = pi16 ? n32 : n52327;
  assign n52329 = pi15 ? n52322 : n52328;
  assign n52330 = pi21 ? n206 : n10182;
  assign n52331 = pi20 ? n52330 : ~n32;
  assign n52332 = pi19 ? n32 : ~n52331;
  assign n52333 = pi18 ? n32 : n52332;
  assign n52334 = pi17 ? n32 : n52333;
  assign n52335 = pi16 ? n32 : n52334;
  assign n52336 = pi15 ? n52335 : n15633;
  assign n52337 = pi14 ? n52329 : n52336;
  assign n52338 = pi13 ? n52317 : n52337;
  assign n52339 = pi19 ? n267 : ~n1077;
  assign n52340 = pi18 ? n32 : n52339;
  assign n52341 = pi17 ? n32 : n52340;
  assign n52342 = pi16 ? n32 : n52341;
  assign n52343 = pi15 ? n52342 : n16606;
  assign n52344 = pi15 ? n16101 : n52278;
  assign n52345 = pi14 ? n52343 : n52344;
  assign n52346 = pi20 ? n260 : ~n11107;
  assign n52347 = pi19 ? n507 : n52346;
  assign n52348 = pi18 ? n52347 : ~n618;
  assign n52349 = pi17 ? n52348 : n20173;
  assign n52350 = pi16 ? n32 : n52349;
  assign n52351 = pi20 ? n28761 : ~n13171;
  assign n52352 = pi19 ? n507 : ~n52351;
  assign n52353 = pi20 ? n18255 : n29452;
  assign n52354 = pi20 ? n246 : ~n1368;
  assign n52355 = pi19 ? n52353 : ~n52354;
  assign n52356 = pi18 ? n52352 : ~n52355;
  assign n52357 = pi20 ? n18832 : ~n2358;
  assign n52358 = pi19 ? n52357 : ~n32;
  assign n52359 = pi19 ? n4342 : ~n236;
  assign n52360 = pi18 ? n52358 : ~n52359;
  assign n52361 = pi17 ? n52356 : ~n52360;
  assign n52362 = pi16 ? n32 : n52361;
  assign n52363 = pi15 ? n52350 : n52362;
  assign n52364 = pi20 ? n30456 : n32;
  assign n52365 = pi19 ? n32 : n52364;
  assign n52366 = pi18 ? n32 : n52365;
  assign n52367 = pi17 ? n32 : n52366;
  assign n52368 = pi16 ? n32 : n52367;
  assign n52369 = pi15 ? n32 : n52368;
  assign n52370 = pi14 ? n52363 : n52369;
  assign n52371 = pi13 ? n52345 : n52370;
  assign n52372 = pi12 ? n52338 : n52371;
  assign n52373 = pi18 ? n6118 : n38521;
  assign n52374 = pi18 ? n22159 : ~n323;
  assign n52375 = pi17 ? n52373 : n52374;
  assign n52376 = pi16 ? n32 : n52375;
  assign n52377 = pi15 ? n52376 : n5377;
  assign n52378 = pi14 ? n21320 : n52377;
  assign n52379 = pi19 ? n32 : n34093;
  assign n52380 = pi18 ? n52379 : n38541;
  assign n52381 = pi19 ? n6504 : n32;
  assign n52382 = pi18 ? n38544 : n52381;
  assign n52383 = pi17 ? n52380 : n52382;
  assign n52384 = pi16 ? n32 : n52383;
  assign n52385 = pi15 ? n5377 : n52384;
  assign n52386 = pi17 ? n17883 : n32;
  assign n52387 = pi16 ? n32 : n52386;
  assign n52388 = pi18 ? n24932 : ~n350;
  assign n52389 = pi18 ? n4671 : n5731;
  assign n52390 = pi17 ? n52388 : n52389;
  assign n52391 = pi16 ? n32 : n52390;
  assign n52392 = pi15 ? n52387 : n52391;
  assign n52393 = pi14 ? n52385 : n52392;
  assign n52394 = pi13 ? n52378 : n52393;
  assign n52395 = pi12 ? n52183 : n52394;
  assign n52396 = pi11 ? n52372 : n52395;
  assign n52397 = pi10 ? n52311 : n52396;
  assign n52398 = pi09 ? n52295 : n52397;
  assign n52399 = pi20 ? n32 : n29949;
  assign n52400 = pi19 ? n32 : n52399;
  assign n52401 = pi18 ? n32 : n52400;
  assign n52402 = pi17 ? n32 : n52401;
  assign n52403 = pi16 ? n32 : n52402;
  assign n52404 = pi15 ? n26400 : n52403;
  assign n52405 = pi15 ? n52403 : n17121;
  assign n52406 = pi14 ? n52404 : n52405;
  assign n52407 = pi13 ? n52298 : n52406;
  assign n52408 = pi13 ? n52058 : n32;
  assign n52409 = pi12 ? n52407 : n52408;
  assign n52410 = pi13 ? n32 : n38567;
  assign n52411 = pi12 ? n52307 : n52410;
  assign n52412 = pi11 ? n52409 : n52411;
  assign n52413 = pi15 ? n52335 : n52315;
  assign n52414 = pi14 ? n52329 : n52413;
  assign n52415 = pi13 ? n52317 : n52414;
  assign n52416 = pi19 ? n267 : ~n7206;
  assign n52417 = pi18 ? n32 : n52416;
  assign n52418 = pi17 ? n32 : n52417;
  assign n52419 = pi16 ? n32 : n52418;
  assign n52420 = pi15 ? n52419 : n16606;
  assign n52421 = pi15 ? n16101 : n32;
  assign n52422 = pi14 ? n52420 : n52421;
  assign n52423 = pi20 ? n831 : ~n266;
  assign n52424 = pi19 ? n32 : n52423;
  assign n52425 = pi18 ? n52424 : ~n618;
  assign n52426 = pi18 ? n19232 : n20172;
  assign n52427 = pi17 ? n52425 : n52426;
  assign n52428 = pi16 ? n32 : n52427;
  assign n52429 = pi20 ? n785 : n7939;
  assign n52430 = pi19 ? n52429 : ~n36199;
  assign n52431 = pi18 ? n38747 : ~n52430;
  assign n52432 = pi20 ? n18173 : ~n321;
  assign n52433 = pi19 ? n52432 : ~n32;
  assign n52434 = pi18 ? n52433 : ~n52359;
  assign n52435 = pi17 ? n52431 : ~n52434;
  assign n52436 = pi16 ? n32 : n52435;
  assign n52437 = pi15 ? n52428 : n52436;
  assign n52438 = pi14 ? n52437 : n52369;
  assign n52439 = pi13 ? n52422 : n52438;
  assign n52440 = pi12 ? n52415 : n52439;
  assign n52441 = pi18 ? n32 : n38572;
  assign n52442 = pi18 ? n38575 : ~n323;
  assign n52443 = pi17 ? n52441 : n52442;
  assign n52444 = pi16 ? n32 : n52443;
  assign n52445 = pi15 ? n52444 : n5522;
  assign n52446 = pi14 ? n21320 : n52445;
  assign n52447 = pi17 ? n4497 : ~n2408;
  assign n52448 = pi16 ? n32 : n52447;
  assign n52449 = pi18 ? n16316 : n32;
  assign n52450 = pi17 ? n52449 : n32;
  assign n52451 = pi16 ? n32 : n52450;
  assign n52452 = pi15 ? n52448 : n52451;
  assign n52453 = pi20 ? n653 : n428;
  assign n52454 = pi19 ? n32 : n52453;
  assign n52455 = pi18 ? n52454 : n32;
  assign n52456 = pi17 ? n52455 : n32;
  assign n52457 = pi16 ? n32 : n52456;
  assign n52458 = pi20 ? n749 : ~n266;
  assign n52459 = pi19 ? n32 : n52458;
  assign n52460 = pi18 ? n52459 : ~n350;
  assign n52461 = pi17 ? n52460 : n52389;
  assign n52462 = pi16 ? n32 : n52461;
  assign n52463 = pi15 ? n52457 : n52462;
  assign n52464 = pi14 ? n52452 : n52463;
  assign n52465 = pi13 ? n52446 : n52464;
  assign n52466 = pi12 ? n52183 : n52465;
  assign n52467 = pi11 ? n52440 : n52466;
  assign n52468 = pi10 ? n52412 : n52467;
  assign n52469 = pi09 ? n52295 : n52468;
  assign n52470 = pi08 ? n52398 : n52469;
  assign n52471 = pi07 ? n52290 : n52470;
  assign n52472 = pi06 ? n52121 : n52471;
  assign n52473 = pi05 ? n51795 : n52472;
  assign n52474 = pi04 ? n51197 : n52473;
  assign n52475 = pi03 ? n49454 : n52474;
  assign n52476 = pi02 ? n45884 : n52475;
  assign n52477 = pi01 ? n32 : n52476;
  assign n52478 = pi15 ? n32 : n26272;
  assign n52479 = pi14 ? n52478 : n26269;
  assign n52480 = pi13 ? n32 : n52479;
  assign n52481 = pi12 ? n32 : n52480;
  assign n52482 = pi11 ? n32 : n52481;
  assign n52483 = pi10 ? n32 : n52482;
  assign n52484 = pi14 ? n17348 : n26303;
  assign n52485 = pi14 ? n26400 : n26235;
  assign n52486 = pi13 ? n52484 : n52485;
  assign n52487 = pi14 ? n38491 : n32;
  assign n52488 = pi13 ? n52487 : n32;
  assign n52489 = pi12 ? n52486 : n52488;
  assign n52490 = pi14 ? n32 : n25984;
  assign n52491 = pi13 ? n52490 : n52058;
  assign n52492 = pi14 ? n25861 : n24797;
  assign n52493 = pi14 ? n27557 : n16392;
  assign n52494 = pi13 ? n52492 : n52493;
  assign n52495 = pi12 ? n52491 : n52494;
  assign n52496 = pi11 ? n52489 : n52495;
  assign n52497 = pi15 ? n15847 : n25704;
  assign n52498 = pi15 ? n16546 : n16333;
  assign n52499 = pi14 ? n52497 : n52498;
  assign n52500 = pi15 ? n52322 : n26885;
  assign n52501 = pi15 ? n16377 : n22817;
  assign n52502 = pi14 ? n52500 : n52501;
  assign n52503 = pi13 ? n52499 : n52502;
  assign n52504 = pi19 ? n507 : ~n7206;
  assign n52505 = pi18 ? n32 : n52504;
  assign n52506 = pi17 ? n32 : n52505;
  assign n52507 = pi16 ? n32 : n52506;
  assign n52508 = pi18 ? n23978 : n32;
  assign n52509 = pi17 ? n52508 : n32;
  assign n52510 = pi16 ? n32 : n52509;
  assign n52511 = pi15 ? n16452 : n52510;
  assign n52512 = pi14 ? n52507 : n52511;
  assign n52513 = pi20 ? n9641 : ~n1076;
  assign n52514 = pi19 ? n32 : n52513;
  assign n52515 = pi21 ? n14158 : ~n173;
  assign n52516 = pi20 ? n52515 : n1331;
  assign n52517 = pi19 ? n52516 : ~n617;
  assign n52518 = pi18 ? n52514 : n52517;
  assign n52519 = pi18 ? n17650 : n32;
  assign n52520 = pi17 ? n52518 : n52519;
  assign n52521 = pi16 ? n32 : n52520;
  assign n52522 = pi15 ? n52521 : n32;
  assign n52523 = pi15 ? n24247 : n52368;
  assign n52524 = pi14 ? n52522 : n52523;
  assign n52525 = pi13 ? n52512 : n52524;
  assign n52526 = pi12 ? n52503 : n52525;
  assign n52527 = pi19 ? n507 : ~n6683;
  assign n52528 = pi18 ? n32 : n52527;
  assign n52529 = pi17 ? n32 : n52528;
  assign n52530 = pi16 ? n32 : n52529;
  assign n52531 = pi15 ? n52530 : n23011;
  assign n52532 = pi15 ? n52178 : n39812;
  assign n52533 = pi14 ? n52531 : n52532;
  assign n52534 = pi14 ? n23485 : n32;
  assign n52535 = pi13 ? n52533 : n52534;
  assign n52536 = pi15 ? n22817 : n33901;
  assign n52537 = pi19 ? n4964 : ~n16431;
  assign n52538 = pi18 ? n16603 : ~n52537;
  assign n52539 = pi19 ? n4964 : n5688;
  assign n52540 = pi18 ? n52539 : n4428;
  assign n52541 = pi17 ? n52538 : ~n52540;
  assign n52542 = pi16 ? n32 : n52541;
  assign n52543 = pi19 ? n9536 : ~n32;
  assign n52544 = pi18 ? n2835 : n52543;
  assign n52545 = pi17 ? n52544 : ~n49638;
  assign n52546 = pi16 ? n32 : n52545;
  assign n52547 = pi15 ? n52542 : n52546;
  assign n52548 = pi14 ? n52536 : n52547;
  assign n52549 = pi19 ? n2386 : ~n32;
  assign n52550 = pi18 ? n32 : n52549;
  assign n52551 = pi17 ? n4656 : ~n52550;
  assign n52552 = pi16 ? n32 : n52551;
  assign n52553 = pi17 ? n464 : n20021;
  assign n52554 = pi16 ? n32 : n52553;
  assign n52555 = pi15 ? n52552 : n52554;
  assign n52556 = pi18 ? n19082 : n9170;
  assign n52557 = pi17 ? n52556 : n385;
  assign n52558 = pi16 ? n32 : n52557;
  assign n52559 = pi20 ? n342 : n260;
  assign n52560 = pi19 ? n32 : n52559;
  assign n52561 = pi19 ? n1248 : n349;
  assign n52562 = pi18 ? n52560 : ~n52561;
  assign n52563 = pi17 ? n52562 : n5731;
  assign n52564 = pi16 ? n32 : n52563;
  assign n52565 = pi15 ? n52558 : n52564;
  assign n52566 = pi14 ? n52555 : n52565;
  assign n52567 = pi13 ? n52548 : n52566;
  assign n52568 = pi12 ? n52535 : n52567;
  assign n52569 = pi11 ? n52526 : n52568;
  assign n52570 = pi10 ? n52496 : n52569;
  assign n52571 = pi09 ? n52483 : n52570;
  assign n52572 = pi14 ? n17286 : n26272;
  assign n52573 = pi13 ? n52484 : n52572;
  assign n52574 = pi14 ? n26225 : n32;
  assign n52575 = pi13 ? n52487 : n52574;
  assign n52576 = pi12 ? n52573 : n52575;
  assign n52577 = pi14 ? n32 : n24797;
  assign n52578 = pi13 ? n52577 : n52493;
  assign n52579 = pi12 ? n52491 : n52578;
  assign n52580 = pi11 ? n52576 : n52579;
  assign n52581 = pi19 ? n6398 : n161;
  assign n52582 = pi18 ? n32 : n52581;
  assign n52583 = pi17 ? n32 : n52582;
  assign n52584 = pi16 ? n32 : n52583;
  assign n52585 = pi15 ? n52584 : n22817;
  assign n52586 = pi14 ? n52500 : n52585;
  assign n52587 = pi13 ? n52499 : n52586;
  assign n52588 = pi19 ? n507 : ~n1077;
  assign n52589 = pi18 ? n32 : n52588;
  assign n52590 = pi17 ? n32 : n52589;
  assign n52591 = pi16 ? n32 : n52590;
  assign n52592 = pi15 ? n52507 : n52591;
  assign n52593 = pi14 ? n52592 : n24633;
  assign n52594 = pi20 ? n428 : ~n342;
  assign n52595 = pi19 ? n32 : n52594;
  assign n52596 = pi20 ? n20396 : n1331;
  assign n52597 = pi19 ? n52596 : ~n617;
  assign n52598 = pi18 ? n52595 : n52597;
  assign n52599 = pi17 ? n52598 : n52519;
  assign n52600 = pi16 ? n32 : n52599;
  assign n52601 = pi15 ? n52600 : n32;
  assign n52602 = pi14 ? n52601 : n52523;
  assign n52603 = pi13 ? n52593 : n52602;
  assign n52604 = pi12 ? n52587 : n52603;
  assign n52605 = pi15 ? n23250 : n22923;
  assign n52606 = pi14 ? n52605 : n32;
  assign n52607 = pi13 ? n52533 : n52606;
  assign n52608 = pi18 ? n32 : ~n52537;
  assign n52609 = pi17 ? n52608 : ~n52540;
  assign n52610 = pi16 ? n32 : n52609;
  assign n52611 = pi18 ? n366 : n52543;
  assign n52612 = pi17 ? n52611 : ~n49638;
  assign n52613 = pi16 ? n32 : n52612;
  assign n52614 = pi15 ? n52610 : n52613;
  assign n52615 = pi14 ? n52536 : n52614;
  assign n52616 = pi17 ? n1232 : ~n52550;
  assign n52617 = pi16 ? n32 : n52616;
  assign n52618 = pi15 ? n52617 : n52554;
  assign n52619 = pi18 ? n25746 : n32;
  assign n52620 = pi17 ? n52619 : n21541;
  assign n52621 = pi16 ? n32 : n52620;
  assign n52622 = pi19 ? n32847 : n349;
  assign n52623 = pi18 ? n356 : ~n52622;
  assign n52624 = pi17 ? n52623 : n5731;
  assign n52625 = pi16 ? n32 : n52624;
  assign n52626 = pi15 ? n52621 : n52625;
  assign n52627 = pi14 ? n52618 : n52626;
  assign n52628 = pi13 ? n52615 : n52627;
  assign n52629 = pi12 ? n52607 : n52628;
  assign n52630 = pi11 ? n52604 : n52629;
  assign n52631 = pi10 ? n52580 : n52630;
  assign n52632 = pi09 ? n52483 : n52631;
  assign n52633 = pi08 ? n52571 : n52632;
  assign n52634 = pi15 ? n32 : n38847;
  assign n52635 = pi14 ? n52634 : n26354;
  assign n52636 = pi13 ? n32 : n52635;
  assign n52637 = pi12 ? n32 : n52636;
  assign n52638 = pi11 ? n32 : n52637;
  assign n52639 = pi10 ? n32 : n52638;
  assign n52640 = pi14 ? n26303 : n17515;
  assign n52641 = pi15 ? n17286 : n17152;
  assign n52642 = pi14 ? n52641 : n26272;
  assign n52643 = pi13 ? n52640 : n52642;
  assign n52644 = pi12 ? n52643 : n52488;
  assign n52645 = pi18 ? n32 : n46185;
  assign n52646 = pi17 ? n32 : n52645;
  assign n52647 = pi16 ? n32 : n52646;
  assign n52648 = pi15 ? n17348 : n52647;
  assign n52649 = pi14 ? n32 : n52648;
  assign n52650 = pi15 ? n52647 : n17039;
  assign n52651 = pi14 ? n52650 : n25133;
  assign n52652 = pi13 ? n52649 : n52651;
  assign n52653 = pi15 ? n40426 : n16804;
  assign n52654 = pi14 ? n38431 : n52653;
  assign n52655 = pi14 ? n27557 : n32;
  assign n52656 = pi13 ? n52654 : n52655;
  assign n52657 = pi12 ? n52652 : n52656;
  assign n52658 = pi11 ? n52644 : n52657;
  assign n52659 = pi15 ? n25704 : n16333;
  assign n52660 = pi14 ? n25387 : n52659;
  assign n52661 = pi13 ? n52660 : n52502;
  assign n52662 = pi19 ? n32 : n21412;
  assign n52663 = pi21 ? n85 : ~n259;
  assign n52664 = pi20 ? n428 : n52663;
  assign n52665 = pi19 ? n52664 : n32;
  assign n52666 = pi18 ? n52662 : n52665;
  assign n52667 = pi17 ? n52666 : n32;
  assign n52668 = pi16 ? n32 : n52667;
  assign n52669 = pi15 ? n52668 : n32;
  assign n52670 = pi14 ? n52669 : n24719;
  assign n52671 = pi13 ? n52593 : n52670;
  assign n52672 = pi12 ? n52661 : n52671;
  assign n52673 = pi20 ? n14318 : ~n32;
  assign n52674 = pi19 ? n594 : ~n52673;
  assign n52675 = pi18 ? n32 : n52674;
  assign n52676 = pi17 ? n32 : n52675;
  assign n52677 = pi16 ? n32 : n52676;
  assign n52678 = pi15 ? n16105 : n52677;
  assign n52679 = pi19 ? n507 : n440;
  assign n52680 = pi18 ? n32 : n52679;
  assign n52681 = pi17 ? n32 : n52680;
  assign n52682 = pi16 ? n32 : n52681;
  assign n52683 = pi19 ? n322 : n358;
  assign n52684 = pi18 ? n32 : n52683;
  assign n52685 = pi17 ? n32 : n52684;
  assign n52686 = pi16 ? n32 : n52685;
  assign n52687 = pi15 ? n52682 : n52686;
  assign n52688 = pi14 ? n52678 : n52687;
  assign n52689 = pi19 ? n857 : n5635;
  assign n52690 = pi18 ? n32 : n52689;
  assign n52691 = pi17 ? n32 : n52690;
  assign n52692 = pi16 ? n32 : n52691;
  assign n52693 = pi15 ? n52692 : n24274;
  assign n52694 = pi14 ? n52693 : n22925;
  assign n52695 = pi13 ? n52688 : n52694;
  assign n52696 = pi15 ? n22540 : n33970;
  assign n52697 = pi19 ? n6988 : ~n22501;
  assign n52698 = pi18 ? n2387 : ~n52697;
  assign n52699 = pi18 ? n4965 : n4428;
  assign n52700 = pi17 ? n52698 : ~n52699;
  assign n52701 = pi16 ? n32 : n52700;
  assign n52702 = pi21 ? n100 : ~n309;
  assign n52703 = pi20 ? n32 : n52702;
  assign n52704 = pi19 ? n32 : n52703;
  assign n52705 = pi18 ? n52704 : ~n32;
  assign n52706 = pi17 ? n52705 : ~n5779;
  assign n52707 = pi16 ? n32 : n52706;
  assign n52708 = pi15 ? n52701 : n52707;
  assign n52709 = pi14 ? n52696 : n52708;
  assign n52710 = pi18 ? n52704 : ~n863;
  assign n52711 = pi18 ? n16389 : n5778;
  assign n52712 = pi17 ? n52710 : ~n52711;
  assign n52713 = pi16 ? n32 : n52712;
  assign n52714 = pi20 ? n32 : n10183;
  assign n52715 = pi19 ? n32 : n52714;
  assign n52716 = pi18 ? n52715 : n9012;
  assign n52717 = pi17 ? n52716 : n20021;
  assign n52718 = pi16 ? n32 : n52717;
  assign n52719 = pi15 ? n52713 : n52718;
  assign n52720 = pi20 ? n357 : n266;
  assign n52721 = pi19 ? n52720 : n32;
  assign n52722 = pi18 ? n32 : n52721;
  assign n52723 = pi17 ? n52722 : n32;
  assign n52724 = pi16 ? n32 : n52723;
  assign n52725 = pi18 ? n52715 : ~n52561;
  assign n52726 = pi18 ? n14153 : n5731;
  assign n52727 = pi17 ? n52725 : n52726;
  assign n52728 = pi16 ? n32 : n52727;
  assign n52729 = pi15 ? n52724 : n52728;
  assign n52730 = pi14 ? n52719 : n52729;
  assign n52731 = pi13 ? n52709 : n52730;
  assign n52732 = pi12 ? n52695 : n52731;
  assign n52733 = pi11 ? n52672 : n52732;
  assign n52734 = pi10 ? n52658 : n52733;
  assign n52735 = pi09 ? n52639 : n52734;
  assign n52736 = pi15 ? n38847 : n17152;
  assign n52737 = pi14 ? n26303 : n52736;
  assign n52738 = pi15 ? n38847 : n26272;
  assign n52739 = pi14 ? n26390 : n52738;
  assign n52740 = pi13 ? n52737 : n52739;
  assign n52741 = pi12 ? n52740 : n52488;
  assign n52742 = pi11 ? n52741 : n52657;
  assign n52743 = pi17 ? n17849 : n32;
  assign n52744 = pi16 ? n32 : n52743;
  assign n52745 = pi15 ? n16452 : n52744;
  assign n52746 = pi14 ? n52507 : n52745;
  assign n52747 = pi20 ? n17671 : n9863;
  assign n52748 = pi19 ? n52747 : n32;
  assign n52749 = pi18 ? n17819 : n52748;
  assign n52750 = pi17 ? n52749 : n32;
  assign n52751 = pi16 ? n32 : n52750;
  assign n52752 = pi15 ? n52751 : n32;
  assign n52753 = pi14 ? n52752 : n24719;
  assign n52754 = pi13 ? n52746 : n52753;
  assign n52755 = pi12 ? n52661 : n52754;
  assign n52756 = pi19 ? n594 : n5614;
  assign n52757 = pi18 ? n32 : n52756;
  assign n52758 = pi17 ? n32 : n52757;
  assign n52759 = pi16 ? n32 : n52758;
  assign n52760 = pi15 ? n16105 : n52759;
  assign n52761 = pi14 ? n52760 : n52687;
  assign n52762 = pi15 ? n37312 : n22923;
  assign n52763 = pi14 ? n52762 : n22925;
  assign n52764 = pi13 ? n52761 : n52763;
  assign n52765 = pi18 ? n2142 : ~n52697;
  assign n52766 = pi17 ? n52765 : ~n52699;
  assign n52767 = pi16 ? n32 : n52766;
  assign n52768 = pi17 ? n2143 : ~n5779;
  assign n52769 = pi16 ? n32 : n52768;
  assign n52770 = pi15 ? n52767 : n52769;
  assign n52771 = pi14 ? n52696 : n52770;
  assign n52772 = pi18 ? n936 : ~n863;
  assign n52773 = pi17 ? n52772 : ~n52711;
  assign n52774 = pi16 ? n32 : n52773;
  assign n52775 = pi18 ? n936 : n9012;
  assign n52776 = pi17 ? n52775 : n20021;
  assign n52777 = pi16 ? n32 : n52776;
  assign n52778 = pi15 ? n52774 : n52777;
  assign n52779 = pi17 ? n20834 : n32;
  assign n52780 = pi16 ? n32 : n52779;
  assign n52781 = pi18 ? n936 : ~n52561;
  assign n52782 = pi17 ? n52781 : n52726;
  assign n52783 = pi16 ? n32 : n52782;
  assign n52784 = pi15 ? n52780 : n52783;
  assign n52785 = pi14 ? n52778 : n52784;
  assign n52786 = pi13 ? n52771 : n52785;
  assign n52787 = pi12 ? n52764 : n52786;
  assign n52788 = pi11 ? n52755 : n52787;
  assign n52789 = pi10 ? n52742 : n52788;
  assign n52790 = pi09 ? n52639 : n52789;
  assign n52791 = pi08 ? n52735 : n52790;
  assign n52792 = pi07 ? n52633 : n52791;
  assign n52793 = pi14 ? n17466 : n26462;
  assign n52794 = pi13 ? n32 : n52793;
  assign n52795 = pi12 ? n32 : n52794;
  assign n52796 = pi11 ? n32 : n52795;
  assign n52797 = pi10 ? n32 : n52796;
  assign n52798 = pi15 ? n26462 : n17316;
  assign n52799 = pi14 ? n32 : n52798;
  assign n52800 = pi20 ? n32 : n38008;
  assign n52801 = pi19 ? n32 : n52800;
  assign n52802 = pi18 ? n32 : n52801;
  assign n52803 = pi17 ? n32 : n52802;
  assign n52804 = pi16 ? n32 : n52803;
  assign n52805 = pi15 ? n52804 : n17435;
  assign n52806 = pi14 ? n26390 : n52805;
  assign n52807 = pi13 ? n52799 : n52806;
  assign n52808 = pi15 ? n17435 : n26269;
  assign n52809 = pi14 ? n52808 : n26269;
  assign n52810 = pi13 ? n52809 : n32;
  assign n52811 = pi12 ? n52807 : n52810;
  assign n52812 = pi14 ? n17043 : n25133;
  assign n52813 = pi13 ? n40816 : n52812;
  assign n52814 = pi20 ? n175 : n274;
  assign n52815 = pi19 ? n32 : n52814;
  assign n52816 = pi18 ? n32 : n52815;
  assign n52817 = pi17 ? n32 : n52816;
  assign n52818 = pi16 ? n32 : n52817;
  assign n52819 = pi15 ? n52818 : n26479;
  assign n52820 = pi14 ? n32 : n52819;
  assign n52821 = pi14 ? n16804 : n24799;
  assign n52822 = pi13 ? n52820 : n52821;
  assign n52823 = pi12 ? n52813 : n52822;
  assign n52824 = pi11 ? n52811 : n52823;
  assign n52825 = pi20 ? n1839 : ~n339;
  assign n52826 = pi19 ? n32 : n52825;
  assign n52827 = pi18 ? n32 : n52826;
  assign n52828 = pi17 ? n32 : n52827;
  assign n52829 = pi16 ? n32 : n52828;
  assign n52830 = pi15 ? n52829 : n16333;
  assign n52831 = pi14 ? n25387 : n52830;
  assign n52832 = pi15 ? n15847 : n24237;
  assign n52833 = pi15 ? n16314 : n16105;
  assign n52834 = pi14 ? n52832 : n52833;
  assign n52835 = pi13 ? n52831 : n52834;
  assign n52836 = pi21 ? n206 : n35;
  assign n52837 = pi20 ? n52836 : n32;
  assign n52838 = pi19 ? n32 : n52837;
  assign n52839 = pi18 ? n32 : n52838;
  assign n52840 = pi17 ? n32 : n52839;
  assign n52841 = pi16 ? n32 : n52840;
  assign n52842 = pi20 ? n1817 : n18158;
  assign n52843 = pi19 ? n52842 : n32;
  assign n52844 = pi18 ? n32 : n52843;
  assign n52845 = pi17 ? n52844 : n16450;
  assign n52846 = pi16 ? n32 : n52845;
  assign n52847 = pi21 ? n32 : n30090;
  assign n52848 = pi20 ? n1817 : n52847;
  assign n52849 = pi19 ? n52848 : n32;
  assign n52850 = pi18 ? n32 : n52849;
  assign n52851 = pi17 ? n52850 : n20173;
  assign n52852 = pi16 ? n32 : n52851;
  assign n52853 = pi15 ? n52846 : n52852;
  assign n52854 = pi14 ? n52841 : n52853;
  assign n52855 = pi15 ? n24582 : n24247;
  assign n52856 = pi14 ? n38992 : n52855;
  assign n52857 = pi13 ? n52854 : n52856;
  assign n52858 = pi12 ? n52835 : n52857;
  assign n52859 = pi15 ? n15244 : n23443;
  assign n52860 = pi14 ? n52859 : n34408;
  assign n52861 = pi15 ? n21853 : n25247;
  assign n52862 = pi14 ? n52861 : n38175;
  assign n52863 = pi13 ? n52860 : n52862;
  assign n52864 = pi19 ? n9037 : ~n322;
  assign n52865 = pi18 ? n32 : n52864;
  assign n52866 = pi18 ? n16847 : n28602;
  assign n52867 = pi17 ? n52865 : n52866;
  assign n52868 = pi16 ? n32 : n52867;
  assign n52869 = pi15 ? n32 : n52868;
  assign n52870 = pi19 ? n6683 : ~n18678;
  assign n52871 = pi18 ? n32 : n52870;
  assign n52872 = pi18 ? n4380 : ~n5357;
  assign n52873 = pi17 ? n52871 : ~n52872;
  assign n52874 = pi16 ? n32 : n52873;
  assign n52875 = pi18 ? n20164 : ~n5357;
  assign n52876 = pi17 ? n5437 : ~n52875;
  assign n52877 = pi16 ? n32 : n52876;
  assign n52878 = pi15 ? n52874 : n52877;
  assign n52879 = pi14 ? n52869 : n52878;
  assign n52880 = pi21 ? n7659 : ~n32;
  assign n52881 = pi20 ? n52880 : ~n32;
  assign n52882 = pi19 ? n52881 : ~n32;
  assign n52883 = pi18 ? n32 : n52882;
  assign n52884 = pi17 ? n52883 : ~n2519;
  assign n52885 = pi16 ? n32 : n52884;
  assign n52886 = pi17 ? n18533 : n14395;
  assign n52887 = pi16 ? n32 : n52886;
  assign n52888 = pi15 ? n52885 : n52887;
  assign n52889 = pi17 ? n16317 : n21317;
  assign n52890 = pi16 ? n32 : n52889;
  assign n52891 = pi17 ? n46740 : n14395;
  assign n52892 = pi16 ? n32 : n52891;
  assign n52893 = pi15 ? n52890 : n52892;
  assign n52894 = pi14 ? n52888 : n52893;
  assign n52895 = pi13 ? n52879 : n52894;
  assign n52896 = pi12 ? n52863 : n52895;
  assign n52897 = pi11 ? n52858 : n52896;
  assign n52898 = pi10 ? n52824 : n52897;
  assign n52899 = pi09 ? n52797 : n52898;
  assign n52900 = pi15 ? n17428 : n17435;
  assign n52901 = pi14 ? n17316 : n52900;
  assign n52902 = pi13 ? n26507 : n52901;
  assign n52903 = pi15 ? n17367 : n26269;
  assign n52904 = pi14 ? n52903 : n26269;
  assign n52905 = pi14 ? n26349 : n38814;
  assign n52906 = pi13 ? n52904 : n52905;
  assign n52907 = pi12 ? n52902 : n52906;
  assign n52908 = pi15 ? n32 : n17066;
  assign n52909 = pi14 ? n32 : n52908;
  assign n52910 = pi14 ? n38505 : n25133;
  assign n52911 = pi13 ? n52909 : n52910;
  assign n52912 = pi12 ? n52911 : n52822;
  assign n52913 = pi11 ? n52907 : n52912;
  assign n52914 = pi20 ? n1324 : ~n339;
  assign n52915 = pi19 ? n32 : n52914;
  assign n52916 = pi18 ? n32 : n52915;
  assign n52917 = pi17 ? n32 : n52916;
  assign n52918 = pi16 ? n32 : n52917;
  assign n52919 = pi15 ? n52918 : n15847;
  assign n52920 = pi14 ? n25387 : n52919;
  assign n52921 = pi13 ? n52920 : n52834;
  assign n52922 = pi20 ? n1817 : n3523;
  assign n52923 = pi19 ? n52922 : n32;
  assign n52924 = pi18 ? n32 : n52923;
  assign n52925 = pi17 ? n52924 : n16450;
  assign n52926 = pi16 ? n32 : n52925;
  assign n52927 = pi20 ? n26832 : n3523;
  assign n52928 = pi19 ? n52927 : n32;
  assign n52929 = pi18 ? n32 : n52928;
  assign n52930 = pi17 ? n52929 : n20173;
  assign n52931 = pi16 ? n32 : n52930;
  assign n52932 = pi15 ? n52926 : n52931;
  assign n52933 = pi14 ? n52841 : n52932;
  assign n52934 = pi14 ? n38992 : n39249;
  assign n52935 = pi13 ? n52933 : n52934;
  assign n52936 = pi12 ? n52921 : n52935;
  assign n52937 = pi15 ? n21853 : n22923;
  assign n52938 = pi14 ? n52859 : n52937;
  assign n52939 = pi13 ? n52938 : n52862;
  assign n52940 = pi19 ? n1812 : ~n18678;
  assign n52941 = pi18 ? n32 : n52940;
  assign n52942 = pi17 ? n52941 : ~n52872;
  assign n52943 = pi16 ? n32 : n52942;
  assign n52944 = pi15 ? n52943 : n52877;
  assign n52945 = pi14 ? n52869 : n52944;
  assign n52946 = pi15 ? n38958 : n14397;
  assign n52947 = pi19 ? n462 : n7693;
  assign n52948 = pi18 ? n32 : n52947;
  assign n52949 = pi17 ? n52948 : n21317;
  assign n52950 = pi16 ? n32 : n52949;
  assign n52951 = pi15 ? n52950 : n52892;
  assign n52952 = pi14 ? n52946 : n52951;
  assign n52953 = pi13 ? n52945 : n52952;
  assign n52954 = pi12 ? n52939 : n52953;
  assign n52955 = pi11 ? n52936 : n52954;
  assign n52956 = pi10 ? n52913 : n52955;
  assign n52957 = pi09 ? n52797 : n52956;
  assign n52958 = pi08 ? n52899 : n52957;
  assign n52959 = pi19 ? n32 : n14382;
  assign n52960 = pi18 ? n32 : n52959;
  assign n52961 = pi17 ? n32 : n52960;
  assign n52962 = pi16 ? n32 : n52961;
  assign n52963 = pi15 ? n32 : n52962;
  assign n52964 = pi14 ? n52963 : n38973;
  assign n52965 = pi13 ? n32 : n52964;
  assign n52966 = pi12 ? n32 : n52965;
  assign n52967 = pi11 ? n32 : n52966;
  assign n52968 = pi10 ? n32 : n52967;
  assign n52969 = pi15 ? n38913 : n17465;
  assign n52970 = pi14 ? n32 : n52969;
  assign n52971 = pi13 ? n52970 : n38975;
  assign n52972 = pi15 ? n17111 : n38937;
  assign n52973 = pi15 ? n38937 : n16984;
  assign n52974 = pi14 ? n52972 : n52973;
  assign n52975 = pi13 ? n52905 : n52974;
  assign n52976 = pi12 ? n52971 : n52975;
  assign n52977 = pi20 ? n428 : ~n287;
  assign n52978 = pi19 ? n32 : n52977;
  assign n52979 = pi18 ? n32 : n52978;
  assign n52980 = pi17 ? n32 : n52979;
  assign n52981 = pi16 ? n32 : n52980;
  assign n52982 = pi15 ? n32 : n52981;
  assign n52983 = pi14 ? n32 : n52982;
  assign n52984 = pi14 ? n38628 : n25133;
  assign n52985 = pi13 ? n52983 : n52984;
  assign n52986 = pi14 ? n32 : n16893;
  assign n52987 = pi14 ? n16804 : n32;
  assign n52988 = pi13 ? n52986 : n52987;
  assign n52989 = pi12 ? n52985 : n52988;
  assign n52990 = pi11 ? n52976 : n52989;
  assign n52991 = pi14 ? n16452 : n15847;
  assign n52992 = pi15 ? n24289 : n52841;
  assign n52993 = pi14 ? n52832 : n52992;
  assign n52994 = pi13 ? n52991 : n52993;
  assign n52995 = pi20 ? n39817 : n32;
  assign n52996 = pi19 ? n32 : n52995;
  assign n52997 = pi18 ? n32 : n52996;
  assign n52998 = pi17 ? n32 : n52997;
  assign n52999 = pi16 ? n32 : n52998;
  assign n53000 = pi15 ? n52999 : n16101;
  assign n53001 = pi20 ? n151 : n1817;
  assign n53002 = pi19 ? n53001 : n32;
  assign n53003 = pi18 ? n32 : n53002;
  assign n53004 = pi18 ? n17118 : n16449;
  assign n53005 = pi17 ? n53003 : n53004;
  assign n53006 = pi16 ? n32 : n53005;
  assign n53007 = pi19 ? n29363 : n7853;
  assign n53008 = pi18 ? n32 : n53007;
  assign n53009 = pi17 ? n53008 : n20173;
  assign n53010 = pi16 ? n32 : n53009;
  assign n53011 = pi15 ? n53006 : n53010;
  assign n53012 = pi14 ? n53000 : n53011;
  assign n53013 = pi14 ? n24719 : n39249;
  assign n53014 = pi13 ? n53012 : n53013;
  assign n53015 = pi12 ? n52994 : n53014;
  assign n53016 = pi15 ? n24742 : n23443;
  assign n53017 = pi14 ? n53016 : n34408;
  assign n53018 = pi13 ? n53017 : n52862;
  assign n53019 = pi19 ? n2033 : ~n322;
  assign n53020 = pi18 ? n32 : n53019;
  assign n53021 = pi17 ? n53020 : n52866;
  assign n53022 = pi16 ? n32 : n53021;
  assign n53023 = pi15 ? n32 : n53022;
  assign n53024 = pi20 ? n428 : ~n17665;
  assign n53025 = pi19 ? n53024 : ~n4342;
  assign n53026 = pi18 ? n32 : n53025;
  assign n53027 = pi18 ? n6057 : ~n5357;
  assign n53028 = pi17 ? n53026 : ~n53027;
  assign n53029 = pi16 ? n32 : n53028;
  assign n53030 = pi17 ? n2644 : ~n52875;
  assign n53031 = pi16 ? n32 : n53030;
  assign n53032 = pi15 ? n53029 : n53031;
  assign n53033 = pi14 ? n53023 : n53032;
  assign n53034 = pi19 ? n28036 : ~n322;
  assign n53035 = pi18 ? n53034 : ~n14153;
  assign n53036 = pi17 ? n14395 : ~n53035;
  assign n53037 = pi16 ? n32 : n53036;
  assign n53038 = pi15 ? n39066 : n53037;
  assign n53039 = pi18 ? n858 : n21316;
  assign n53040 = pi17 ? n20834 : n53039;
  assign n53041 = pi16 ? n32 : n53040;
  assign n53042 = pi17 ? n46740 : n20834;
  assign n53043 = pi16 ? n32 : n53042;
  assign n53044 = pi15 ? n53041 : n53043;
  assign n53045 = pi14 ? n53038 : n53044;
  assign n53046 = pi13 ? n53033 : n53045;
  assign n53047 = pi12 ? n53018 : n53046;
  assign n53048 = pi11 ? n53015 : n53047;
  assign n53049 = pi10 ? n52990 : n53048;
  assign n53050 = pi09 ? n52968 : n53049;
  assign n53051 = pi14 ? n26591 : n38973;
  assign n53052 = pi13 ? n32 : n53051;
  assign n53053 = pi12 ? n32 : n53052;
  assign n53054 = pi11 ? n32 : n53053;
  assign n53055 = pi10 ? n32 : n53054;
  assign n53056 = pi13 ? n52970 : n39034;
  assign n53057 = pi12 ? n53056 : n32;
  assign n53058 = pi11 ? n53057 : n52989;
  assign n53059 = pi15 ? n15847 : n16319;
  assign n53060 = pi15 ? n24289 : n25301;
  assign n53061 = pi14 ? n53059 : n53060;
  assign n53062 = pi13 ? n52991 : n53061;
  assign n53063 = pi15 ? n52999 : n27686;
  assign n53064 = pi20 ? n974 : n32;
  assign n53065 = pi19 ? n1818 : n53064;
  assign n53066 = pi18 ? n32 : n53065;
  assign n53067 = pi17 ? n53066 : n53004;
  assign n53068 = pi16 ? n32 : n53067;
  assign n53069 = pi21 ? n174 : ~n13784;
  assign n53070 = pi20 ? n32 : n53069;
  assign n53071 = pi19 ? n53070 : n6136;
  assign n53072 = pi18 ? n32 : n53071;
  assign n53073 = pi17 ? n53072 : n20173;
  assign n53074 = pi16 ? n32 : n53073;
  assign n53075 = pi15 ? n53068 : n53074;
  assign n53076 = pi14 ? n53063 : n53075;
  assign n53077 = pi13 ? n53076 : n53013;
  assign n53078 = pi12 ? n53062 : n53077;
  assign n53079 = pi17 ? n14430 : n52866;
  assign n53080 = pi16 ? n32 : n53079;
  assign n53081 = pi15 ? n32 : n53080;
  assign n53082 = pi19 ? n35361 : ~n3495;
  assign n53083 = pi18 ? n32 : n53082;
  assign n53084 = pi17 ? n53083 : ~n5358;
  assign n53085 = pi16 ? n32 : n53084;
  assign n53086 = pi17 ? n2425 : ~n52875;
  assign n53087 = pi16 ? n32 : n53086;
  assign n53088 = pi15 ? n53085 : n53087;
  assign n53089 = pi14 ? n53081 : n53088;
  assign n53090 = pi17 ? n2425 : ~n2519;
  assign n53091 = pi16 ? n32 : n53090;
  assign n53092 = pi15 ? n53091 : n53037;
  assign n53093 = pi18 ? n858 : n9012;
  assign n53094 = pi17 ? n20834 : n53093;
  assign n53095 = pi16 ? n32 : n53094;
  assign n53096 = pi15 ? n53095 : n53043;
  assign n53097 = pi14 ? n53092 : n53096;
  assign n53098 = pi13 ? n53089 : n53097;
  assign n53099 = pi12 ? n53018 : n53098;
  assign n53100 = pi11 ? n53078 : n53099;
  assign n53101 = pi10 ? n53058 : n53100;
  assign n53102 = pi09 ? n53055 : n53101;
  assign n53103 = pi08 ? n53050 : n53102;
  assign n53104 = pi07 ? n52958 : n53103;
  assign n53105 = pi06 ? n52792 : n53104;
  assign n53106 = pi14 ? n17608 : n17607;
  assign n53107 = pi13 ? n32 : n53106;
  assign n53108 = pi12 ? n32 : n53107;
  assign n53109 = pi11 ? n32 : n53108;
  assign n53110 = pi10 ? n32 : n53109;
  assign n53111 = pi15 ? n17607 : n17618;
  assign n53112 = pi14 ? n17316 : n53111;
  assign n53113 = pi13 ? n53112 : n17278;
  assign n53114 = pi12 ? n53113 : n39227;
  assign n53115 = pi20 ? n428 : ~n518;
  assign n53116 = pi19 ? n32 : n53115;
  assign n53117 = pi18 ? n32 : n53116;
  assign n53118 = pi17 ? n32 : n53117;
  assign n53119 = pi16 ? n32 : n53118;
  assign n53120 = pi15 ? n32 : n53119;
  assign n53121 = pi14 ? n32 : n53120;
  assign n53122 = pi14 ? n16736 : n25133;
  assign n53123 = pi13 ? n53121 : n53122;
  assign n53124 = pi15 ? n26479 : n16804;
  assign n53125 = pi14 ? n32 : n53124;
  assign n53126 = pi13 ? n53125 : n52987;
  assign n53127 = pi12 ? n53123 : n53126;
  assign n53128 = pi11 ? n53114 : n53127;
  assign n53129 = pi15 ? n16452 : n25708;
  assign n53130 = pi18 ? n32 : n48472;
  assign n53131 = pi17 ? n32 : n53130;
  assign n53132 = pi16 ? n32 : n53131;
  assign n53133 = pi15 ? n53132 : n15847;
  assign n53134 = pi14 ? n53129 : n53133;
  assign n53135 = pi15 ? n16319 : n15244;
  assign n53136 = pi21 ? n32 : ~n1009;
  assign n53137 = pi20 ? n53136 : ~n32;
  assign n53138 = pi19 ? n507 : ~n53137;
  assign n53139 = pi18 ? n32 : n53138;
  assign n53140 = pi17 ? n32 : n53139;
  assign n53141 = pi16 ? n32 : n53140;
  assign n53142 = pi15 ? n39520 : n53141;
  assign n53143 = pi14 ? n53135 : n53142;
  assign n53144 = pi13 ? n53134 : n53143;
  assign n53145 = pi19 ? n6398 : n18390;
  assign n53146 = pi18 ? n32 : n53145;
  assign n53147 = pi19 ? n531 : ~n16511;
  assign n53148 = pi18 ? n32 : ~n53147;
  assign n53149 = pi17 ? n53146 : n53148;
  assign n53150 = pi16 ? n32 : n53149;
  assign n53151 = pi19 ? n358 : n16511;
  assign n53152 = pi18 ? n32 : n53151;
  assign n53153 = pi17 ? n21926 : n53152;
  assign n53154 = pi16 ? n32 : n53153;
  assign n53155 = pi15 ? n53150 : n53154;
  assign n53156 = pi19 ? n358 : n247;
  assign n53157 = pi18 ? n32 : n53156;
  assign n53158 = pi17 ? n21926 : n53157;
  assign n53159 = pi16 ? n32 : n53158;
  assign n53160 = pi15 ? n53159 : n24247;
  assign n53161 = pi14 ? n53155 : n53160;
  assign n53162 = pi15 ? n24247 : n15244;
  assign n53163 = pi15 ? n15244 : n22817;
  assign n53164 = pi14 ? n53162 : n53163;
  assign n53165 = pi13 ? n53161 : n53164;
  assign n53166 = pi12 ? n53144 : n53165;
  assign n53167 = pi15 ? n24742 : n21853;
  assign n53168 = pi14 ? n53167 : n21853;
  assign n53169 = pi15 ? n23443 : n15119;
  assign n53170 = pi15 ? n38175 : n14156;
  assign n53171 = pi14 ? n53169 : n53170;
  assign n53172 = pi13 ? n53168 : n53171;
  assign n53173 = pi21 ? n100 : n259;
  assign n53174 = pi20 ? n32 : n53173;
  assign n53175 = pi19 ? n53174 : ~n4342;
  assign n53176 = pi18 ? n32 : n53175;
  assign n53177 = pi19 ? n266 : n1757;
  assign n53178 = pi18 ? n53177 : n508;
  assign n53179 = pi17 ? n53176 : ~n53178;
  assign n53180 = pi16 ? n32 : n53179;
  assign n53181 = pi15 ? n14147 : n53180;
  assign n53182 = pi17 ? n2292 : ~n2512;
  assign n53183 = pi16 ? n32 : n53182;
  assign n53184 = pi18 ? n32 : n1712;
  assign n53185 = pi18 ? n16847 : n508;
  assign n53186 = pi17 ? n53184 : ~n53185;
  assign n53187 = pi16 ? n32 : n53186;
  assign n53188 = pi15 ? n53183 : n53187;
  assign n53189 = pi14 ? n53181 : n53188;
  assign n53190 = pi17 ? n53184 : ~n2868;
  assign n53191 = pi16 ? n32 : n53190;
  assign n53192 = pi17 ? n2750 : ~n2119;
  assign n53193 = pi16 ? n32 : n53192;
  assign n53194 = pi15 ? n53191 : n53193;
  assign n53195 = pi20 ? n357 : n7388;
  assign n53196 = pi19 ? n32 : n53195;
  assign n53197 = pi18 ? n32 : n53196;
  assign n53198 = pi17 ? n53197 : n32;
  assign n53199 = pi16 ? n32 : n53198;
  assign n53200 = pi19 ? n32 : ~n25120;
  assign n53201 = pi18 ? n32 : n53200;
  assign n53202 = pi18 ? n350 : ~n5005;
  assign n53203 = pi17 ? n53201 : ~n53202;
  assign n53204 = pi16 ? n32 : n53203;
  assign n53205 = pi15 ? n53199 : n53204;
  assign n53206 = pi14 ? n53194 : n53205;
  assign n53207 = pi13 ? n53189 : n53206;
  assign n53208 = pi12 ? n53172 : n53207;
  assign n53209 = pi11 ? n53166 : n53208;
  assign n53210 = pi10 ? n53128 : n53209;
  assign n53211 = pi09 ? n53110 : n53210;
  assign n53212 = pi15 ? n17316 : n17278;
  assign n53213 = pi14 ? n53212 : n17278;
  assign n53214 = pi13 ? n17316 : n53213;
  assign n53215 = pi12 ? n53214 : n39287;
  assign n53216 = pi11 ? n53215 : n53127;
  assign n53217 = pi19 ? n507 : ~n4342;
  assign n53218 = pi18 ? n32 : n53217;
  assign n53219 = pi17 ? n53218 : ~n53178;
  assign n53220 = pi16 ? n32 : n53219;
  assign n53221 = pi15 ? n14147 : n53220;
  assign n53222 = pi17 ? n2736 : ~n53185;
  assign n53223 = pi16 ? n32 : n53222;
  assign n53224 = pi15 ? n8331 : n53223;
  assign n53225 = pi14 ? n53221 : n53224;
  assign n53226 = pi15 ? n39192 : n39146;
  assign n53227 = pi20 ? n357 : n274;
  assign n53228 = pi19 ? n32 : n53227;
  assign n53229 = pi18 ? n32 : n53228;
  assign n53230 = pi17 ? n53229 : n32;
  assign n53231 = pi16 ? n32 : n53230;
  assign n53232 = pi19 ? n1574 : ~n25120;
  assign n53233 = pi18 ? n32 : n53232;
  assign n53234 = pi17 ? n53233 : ~n53202;
  assign n53235 = pi16 ? n32 : n53234;
  assign n53236 = pi15 ? n53231 : n53235;
  assign n53237 = pi14 ? n53226 : n53236;
  assign n53238 = pi13 ? n53225 : n53237;
  assign n53239 = pi12 ? n53172 : n53238;
  assign n53240 = pi11 ? n53166 : n53239;
  assign n53241 = pi10 ? n53216 : n53240;
  assign n53242 = pi09 ? n53110 : n53241;
  assign n53243 = pi08 ? n53211 : n53242;
  assign n53244 = pi14 ? n17466 : n17465;
  assign n53245 = pi13 ? n32 : n53244;
  assign n53246 = pi12 ? n32 : n53245;
  assign n53247 = pi11 ? n32 : n53246;
  assign n53248 = pi10 ? n32 : n53247;
  assign n53249 = pi13 ? n32 : n39156;
  assign n53250 = pi12 ? n17465 : n53249;
  assign n53251 = pi14 ? n16736 : n32;
  assign n53252 = pi13 ? n53121 : n53251;
  assign n53253 = pi13 ? n53125 : n38864;
  assign n53254 = pi12 ? n53252 : n53253;
  assign n53255 = pi11 ? n53250 : n53254;
  assign n53256 = pi19 ? n4721 : ~n16511;
  assign n53257 = pi18 ? n32 : ~n53256;
  assign n53258 = pi17 ? n8193 : n53257;
  assign n53259 = pi16 ? n32 : n53258;
  assign n53260 = pi19 ? n32 : n52842;
  assign n53261 = pi18 ? n32 : n53260;
  assign n53262 = pi21 ? n174 : n1009;
  assign n53263 = pi20 ? n53262 : n32;
  assign n53264 = pi19 ? n1464 : n53263;
  assign n53265 = pi18 ? n32 : n53264;
  assign n53266 = pi17 ? n53261 : n53265;
  assign n53267 = pi16 ? n32 : n53266;
  assign n53268 = pi15 ? n53259 : n53267;
  assign n53269 = pi19 ? n1757 : n247;
  assign n53270 = pi18 ? n32 : n53269;
  assign n53271 = pi17 ? n53261 : n53270;
  assign n53272 = pi16 ? n32 : n53271;
  assign n53273 = pi15 ? n53272 : n24247;
  assign n53274 = pi14 ? n53268 : n53273;
  assign n53275 = pi14 ? n15362 : n53163;
  assign n53276 = pi13 ? n53274 : n53275;
  assign n53277 = pi12 ? n53144 : n53276;
  assign n53278 = pi15 ? n27355 : n22437;
  assign n53279 = pi14 ? n53278 : n21853;
  assign n53280 = pi15 ? n23443 : n22817;
  assign n53281 = pi14 ? n53280 : n53170;
  assign n53282 = pi13 ? n53279 : n53281;
  assign n53283 = pi19 ? n52720 : n6314;
  assign n53284 = pi18 ? n53283 : n33476;
  assign n53285 = pi17 ? n2852 : ~n53284;
  assign n53286 = pi16 ? n32 : n53285;
  assign n53287 = pi15 ? n14147 : n53286;
  assign n53288 = pi19 ? n32 : n52881;
  assign n53289 = pi18 ? n32 : n53288;
  assign n53290 = pi17 ? n53289 : ~n53185;
  assign n53291 = pi16 ? n32 : n53290;
  assign n53292 = pi15 ? n8701 : n53291;
  assign n53293 = pi14 ? n53287 : n53292;
  assign n53294 = pi17 ? n53289 : ~n2517;
  assign n53295 = pi16 ? n32 : n53294;
  assign n53296 = pi17 ? n8653 : ~n2119;
  assign n53297 = pi16 ? n32 : n53296;
  assign n53298 = pi15 ? n53295 : n53297;
  assign n53299 = pi20 ? n17671 : n6303;
  assign n53300 = pi19 ? n32 : n53299;
  assign n53301 = pi18 ? n32 : n53300;
  assign n53302 = pi20 ? n3843 : n17671;
  assign n53303 = pi19 ? n53302 : n462;
  assign n53304 = pi19 ? n29270 : n32;
  assign n53305 = pi18 ? n53303 : n53304;
  assign n53306 = pi17 ? n53301 : n53305;
  assign n53307 = pi16 ? n32 : n53306;
  assign n53308 = pi17 ? n16395 : ~n53202;
  assign n53309 = pi16 ? n32 : n53308;
  assign n53310 = pi15 ? n53307 : n53309;
  assign n53311 = pi14 ? n53298 : n53310;
  assign n53312 = pi13 ? n53293 : n53311;
  assign n53313 = pi12 ? n53282 : n53312;
  assign n53314 = pi11 ? n53277 : n53313;
  assign n53315 = pi10 ? n53255 : n53314;
  assign n53316 = pi09 ? n53248 : n53315;
  assign n53317 = pi17 ? n26423 : n53265;
  assign n53318 = pi16 ? n32 : n53317;
  assign n53319 = pi15 ? n53259 : n53318;
  assign n53320 = pi17 ? n26423 : n53270;
  assign n53321 = pi16 ? n32 : n53320;
  assign n53322 = pi15 ? n53321 : n24247;
  assign n53323 = pi14 ? n53319 : n53322;
  assign n53324 = pi15 ? n40538 : n22817;
  assign n53325 = pi14 ? n15362 : n53324;
  assign n53326 = pi13 ? n53323 : n53325;
  assign n53327 = pi12 ? n53144 : n53326;
  assign n53328 = pi19 ? n1785 : ~n813;
  assign n53329 = pi18 ? n32 : n53328;
  assign n53330 = pi17 ? n32 : n53329;
  assign n53331 = pi16 ? n32 : n53330;
  assign n53332 = pi15 ? n53331 : n22437;
  assign n53333 = pi14 ? n53332 : n21853;
  assign n53334 = pi13 ? n53333 : n53281;
  assign n53335 = pi19 ? n267 : n6314;
  assign n53336 = pi18 ? n53335 : n33476;
  assign n53337 = pi17 ? n4245 : ~n53336;
  assign n53338 = pi16 ? n32 : n53337;
  assign n53339 = pi15 ? n14147 : n53338;
  assign n53340 = pi17 ? n3067 : ~n24861;
  assign n53341 = pi16 ? n32 : n53340;
  assign n53342 = pi15 ? n8899 : n53341;
  assign n53343 = pi14 ? n53339 : n53342;
  assign n53344 = pi20 ? n13792 : n1091;
  assign n53345 = pi19 ? n32 : n53344;
  assign n53346 = pi18 ? n32 : n53345;
  assign n53347 = pi20 ? n220 : n17671;
  assign n53348 = pi20 ? n174 : n357;
  assign n53349 = pi19 ? n53347 : n53348;
  assign n53350 = pi18 ? n53349 : n53304;
  assign n53351 = pi17 ? n53346 : n53350;
  assign n53352 = pi16 ? n32 : n53351;
  assign n53353 = pi15 ? n53352 : n53309;
  assign n53354 = pi14 ? n39218 : n53353;
  assign n53355 = pi13 ? n53343 : n53354;
  assign n53356 = pi12 ? n53334 : n53355;
  assign n53357 = pi11 ? n53327 : n53356;
  assign n53358 = pi10 ? n53255 : n53357;
  assign n53359 = pi09 ? n53248 : n53358;
  assign n53360 = pi08 ? n53316 : n53359;
  assign n53361 = pi07 ? n53243 : n53360;
  assign n53362 = pi15 ? n16392 : n16397;
  assign n53363 = pi14 ? n32 : n53362;
  assign n53364 = pi13 ? n53363 : n53251;
  assign n53365 = pi14 ? n32 : n16804;
  assign n53366 = pi14 ? n25133 : n24691;
  assign n53367 = pi13 ? n53365 : n53366;
  assign n53368 = pi12 ? n53364 : n53367;
  assign n53369 = pi11 ? n39228 : n53368;
  assign n53370 = pi15 ? n16452 : n15847;
  assign n53371 = pi18 ? n19232 : n32;
  assign n53372 = pi17 ? n32 : n53371;
  assign n53373 = pi16 ? n32 : n53372;
  assign n53374 = pi15 ? n32 : n53373;
  assign n53375 = pi14 ? n53370 : n53374;
  assign n53376 = pi18 ? n19232 : n16316;
  assign n53377 = pi17 ? n32 : n53376;
  assign n53378 = pi16 ? n32 : n53377;
  assign n53379 = pi15 ? n53378 : n39243;
  assign n53380 = pi20 ? n428 : ~n266;
  assign n53381 = pi20 ? n5854 : ~n266;
  assign n53382 = pi19 ? n53380 : n53381;
  assign n53383 = pi19 ? n5688 : n53263;
  assign n53384 = pi18 ? n53382 : n53383;
  assign n53385 = pi17 ? n4319 : n53384;
  assign n53386 = pi16 ? n32 : n53385;
  assign n53387 = pi15 ? n39243 : n53386;
  assign n53388 = pi14 ? n53379 : n53387;
  assign n53389 = pi13 ? n53375 : n53388;
  assign n53390 = pi20 ? n14286 : n207;
  assign n53391 = pi19 ? n32 : n53390;
  assign n53392 = pi18 ? n32 : n53391;
  assign n53393 = pi19 ? n5356 : n28685;
  assign n53394 = pi20 ? n7861 : ~n32;
  assign n53395 = pi19 ? n267 : ~n53394;
  assign n53396 = pi18 ? n53393 : n53395;
  assign n53397 = pi17 ? n53392 : n53396;
  assign n53398 = pi16 ? n32 : n53397;
  assign n53399 = pi19 ? n6057 : ~n6652;
  assign n53400 = pi18 ? n32 : n53399;
  assign n53401 = pi17 ? n32 : n53400;
  assign n53402 = pi16 ? n32 : n53401;
  assign n53403 = pi15 ? n53398 : n53402;
  assign n53404 = pi19 ? n449 : ~n502;
  assign n53405 = pi18 ? n32 : n53404;
  assign n53406 = pi17 ? n32 : n53405;
  assign n53407 = pi16 ? n32 : n53406;
  assign n53408 = pi15 ? n53407 : n16105;
  assign n53409 = pi14 ? n53403 : n53408;
  assign n53410 = pi15 ? n16105 : n23574;
  assign n53411 = pi19 ? n2141 : n5614;
  assign n53412 = pi18 ? n32 : n53411;
  assign n53413 = pi17 ? n32 : n53412;
  assign n53414 = pi16 ? n32 : n53413;
  assign n53415 = pi15 ? n53414 : n23933;
  assign n53416 = pi14 ? n53410 : n53415;
  assign n53417 = pi13 ? n53409 : n53416;
  assign n53418 = pi12 ? n53389 : n53417;
  assign n53419 = pi18 ? n32 : n29556;
  assign n53420 = pi17 ? n32 : n53419;
  assign n53421 = pi16 ? n32 : n53420;
  assign n53422 = pi15 ? n53421 : n14790;
  assign n53423 = pi15 ? n21853 : n22540;
  assign n53424 = pi14 ? n53422 : n53423;
  assign n53425 = pi14 ? n23264 : n22856;
  assign n53426 = pi13 ? n53424 : n53425;
  assign n53427 = pi17 ? n2733 : ~n2517;
  assign n53428 = pi16 ? n32 : n53427;
  assign n53429 = pi15 ? n14147 : n53428;
  assign n53430 = pi19 ? n49091 : ~n32;
  assign n53431 = pi18 ? n9012 : n53430;
  assign n53432 = pi17 ? n2733 : ~n53431;
  assign n53433 = pi16 ? n32 : n53432;
  assign n53434 = pi19 ? n32 : n39006;
  assign n53435 = pi18 ? n32 : n53434;
  assign n53436 = pi19 ? n14688 : ~n32;
  assign n53437 = pi18 ? n32 : n53436;
  assign n53438 = pi17 ? n53435 : ~n53437;
  assign n53439 = pi16 ? n32 : n53438;
  assign n53440 = pi15 ? n53433 : n53439;
  assign n53441 = pi14 ? n53429 : n53440;
  assign n53442 = pi17 ? n53435 : ~n34900;
  assign n53443 = pi16 ? n32 : n53442;
  assign n53444 = pi17 ? n4128 : ~n2292;
  assign n53445 = pi16 ? n32 : n53444;
  assign n53446 = pi15 ? n53443 : n53445;
  assign n53447 = pi18 ? n4343 : ~n4343;
  assign n53448 = pi17 ? n49543 : ~n53447;
  assign n53449 = pi16 ? n32 : n53448;
  assign n53450 = pi20 ? n101 : ~n18762;
  assign n53451 = pi19 ? n32 : n53450;
  assign n53452 = pi18 ? n32 : n53451;
  assign n53453 = pi18 ? n20729 : ~n5005;
  assign n53454 = pi17 ? n53452 : ~n53453;
  assign n53455 = pi16 ? n32 : n53454;
  assign n53456 = pi15 ? n53449 : n53455;
  assign n53457 = pi14 ? n53446 : n53456;
  assign n53458 = pi13 ? n53441 : n53457;
  assign n53459 = pi12 ? n53426 : n53458;
  assign n53460 = pi11 ? n53418 : n53459;
  assign n53461 = pi10 ? n53369 : n53460;
  assign n53462 = pi09 ? n32 : n53461;
  assign n53463 = pi11 ? n39288 : n53368;
  assign n53464 = pi18 ? n19232 : n23978;
  assign n53465 = pi17 ? n32 : n53464;
  assign n53466 = pi16 ? n32 : n53465;
  assign n53467 = pi15 ? n32 : n53466;
  assign n53468 = pi14 ? n53370 : n53467;
  assign n53469 = pi21 ? n7107 : ~n206;
  assign n53470 = pi20 ? n53469 : n32;
  assign n53471 = pi19 ? n322 : n53470;
  assign n53472 = pi18 ? n32 : n53471;
  assign n53473 = pi17 ? n32 : n53472;
  assign n53474 = pi16 ? n32 : n53473;
  assign n53475 = pi21 ? n454 : ~n32;
  assign n53476 = pi20 ? n32 : n53475;
  assign n53477 = pi19 ? n32 : n53476;
  assign n53478 = pi18 ? n32 : n53477;
  assign n53479 = pi20 ? n518 : ~n266;
  assign n53480 = pi19 ? n53479 : n53381;
  assign n53481 = pi18 ? n53480 : n53383;
  assign n53482 = pi17 ? n53478 : n53481;
  assign n53483 = pi16 ? n32 : n53482;
  assign n53484 = pi15 ? n53474 : n53483;
  assign n53485 = pi14 ? n53379 : n53484;
  assign n53486 = pi13 ? n53468 : n53485;
  assign n53487 = pi18 ? n32 : n1395;
  assign n53488 = pi17 ? n53487 : n53396;
  assign n53489 = pi16 ? n32 : n53488;
  assign n53490 = pi18 ? n19774 : n53399;
  assign n53491 = pi17 ? n32 : n53490;
  assign n53492 = pi16 ? n32 : n53491;
  assign n53493 = pi15 ? n53489 : n53492;
  assign n53494 = pi14 ? n53493 : n53408;
  assign n53495 = pi19 ? n507 : n5614;
  assign n53496 = pi18 ? n32 : n53495;
  assign n53497 = pi17 ? n32 : n53496;
  assign n53498 = pi16 ? n32 : n53497;
  assign n53499 = pi15 ? n53498 : n23933;
  assign n53500 = pi14 ? n53410 : n53499;
  assign n53501 = pi13 ? n53494 : n53500;
  assign n53502 = pi12 ? n53486 : n53501;
  assign n53503 = pi17 ? n3050 : ~n2517;
  assign n53504 = pi16 ? n32 : n53503;
  assign n53505 = pi15 ? n14147 : n53504;
  assign n53506 = pi17 ? n3050 : ~n53431;
  assign n53507 = pi16 ? n32 : n53506;
  assign n53508 = pi17 ? n2959 : ~n53437;
  assign n53509 = pi16 ? n32 : n53508;
  assign n53510 = pi15 ? n53507 : n53509;
  assign n53511 = pi14 ? n53505 : n53510;
  assign n53512 = pi17 ? n2959 : ~n2868;
  assign n53513 = pi16 ? n32 : n53512;
  assign n53514 = pi17 ? n4128 : ~n2408;
  assign n53515 = pi16 ? n32 : n53514;
  assign n53516 = pi15 ? n53513 : n53515;
  assign n53517 = pi17 ? n3046 : ~n53447;
  assign n53518 = pi16 ? n32 : n53517;
  assign n53519 = pi18 ? n21316 : ~n5005;
  assign n53520 = pi17 ? n2959 : ~n53519;
  assign n53521 = pi16 ? n32 : n53520;
  assign n53522 = pi15 ? n53518 : n53521;
  assign n53523 = pi14 ? n53516 : n53522;
  assign n53524 = pi13 ? n53511 : n53523;
  assign n53525 = pi12 ? n53426 : n53524;
  assign n53526 = pi11 ? n53502 : n53525;
  assign n53527 = pi10 ? n53463 : n53526;
  assign n53528 = pi09 ? n32 : n53527;
  assign n53529 = pi08 ? n53462 : n53528;
  assign n53530 = pi15 ? n16397 : n16850;
  assign n53531 = pi14 ? n53530 : n32;
  assign n53532 = pi13 ? n53363 : n53531;
  assign n53533 = pi15 ? n17061 : n16804;
  assign n53534 = pi14 ? n26163 : n53533;
  assign n53535 = pi13 ? n53534 : n24876;
  assign n53536 = pi12 ? n53532 : n53535;
  assign n53537 = pi11 ? n39288 : n53536;
  assign n53538 = pi14 ? n53370 : n23982;
  assign n53539 = pi15 ? n16319 : n39243;
  assign n53540 = pi19 ? n1248 : n5371;
  assign n53541 = pi18 ? n53540 : n53383;
  assign n53542 = pi17 ? n32 : n53541;
  assign n53543 = pi16 ? n32 : n53542;
  assign n53544 = pi15 ? n53474 : n53543;
  assign n53545 = pi14 ? n53539 : n53544;
  assign n53546 = pi13 ? n53538 : n53545;
  assign n53547 = pi19 ? n267 : ~n6652;
  assign n53548 = pi18 ? n45386 : n53547;
  assign n53549 = pi17 ? n32 : n53548;
  assign n53550 = pi16 ? n32 : n53549;
  assign n53551 = pi21 ? n174 : ~n124;
  assign n53552 = pi20 ? n53551 : ~n32;
  assign n53553 = pi19 ? n267 : ~n53552;
  assign n53554 = pi18 ? n9578 : n53553;
  assign n53555 = pi17 ? n32 : n53554;
  assign n53556 = pi16 ? n32 : n53555;
  assign n53557 = pi15 ? n53550 : n53556;
  assign n53558 = pi15 ? n38371 : n16319;
  assign n53559 = pi14 ? n53557 : n53558;
  assign n53560 = pi19 ? n472 : ~n236;
  assign n53561 = pi18 ? n32 : n53560;
  assign n53562 = pi17 ? n32 : n53561;
  assign n53563 = pi16 ? n32 : n53562;
  assign n53564 = pi15 ? n23574 : n53563;
  assign n53565 = pi14 ? n23574 : n53564;
  assign n53566 = pi13 ? n53559 : n53565;
  assign n53567 = pi12 ? n53546 : n53566;
  assign n53568 = pi21 ? n32 : ~n42173;
  assign n53569 = pi20 ? n32 : n53568;
  assign n53570 = pi19 ? n53569 : n32;
  assign n53571 = pi18 ? n32 : n53570;
  assign n53572 = pi17 ? n32 : n53571;
  assign n53573 = pi16 ? n32 : n53572;
  assign n53574 = pi15 ? n53421 : n53573;
  assign n53575 = pi15 ? n21543 : n14397;
  assign n53576 = pi14 ? n53574 : n53575;
  assign n53577 = pi14 ? n21217 : n23679;
  assign n53578 = pi13 ? n53576 : n53577;
  assign n53579 = pi17 ? n3164 : ~n2517;
  assign n53580 = pi16 ? n32 : n53579;
  assign n53581 = pi15 ? n14147 : n53580;
  assign n53582 = pi20 ? n175 : n266;
  assign n53583 = pi19 ? n267 : n53582;
  assign n53584 = pi18 ? n53583 : n1491;
  assign n53585 = pi17 ? n3164 : ~n53584;
  assign n53586 = pi16 ? n32 : n53585;
  assign n53587 = pi17 ? n46383 : ~n38897;
  assign n53588 = pi16 ? n32 : n53587;
  assign n53589 = pi15 ? n53586 : n53588;
  assign n53590 = pi14 ? n53581 : n53589;
  assign n53591 = pi20 ? n32 : n13792;
  assign n53592 = pi19 ? n32 : n53591;
  assign n53593 = pi18 ? n32 : n53592;
  assign n53594 = pi17 ? n53593 : ~n2119;
  assign n53595 = pi16 ? n32 : n53594;
  assign n53596 = pi18 ? n4343 : ~n13080;
  assign n53597 = pi17 ? n32 : ~n53596;
  assign n53598 = pi16 ? n32 : n53597;
  assign n53599 = pi20 ? n357 : ~n321;
  assign n53600 = pi19 ? n53599 : n32;
  assign n53601 = pi18 ? n53600 : ~n13372;
  assign n53602 = pi17 ? n32 : ~n53601;
  assign n53603 = pi16 ? n32 : n53602;
  assign n53604 = pi15 ? n53598 : n53603;
  assign n53605 = pi14 ? n53595 : n53604;
  assign n53606 = pi13 ? n53590 : n53605;
  assign n53607 = pi12 ? n53578 : n53606;
  assign n53608 = pi11 ? n53567 : n53607;
  assign n53609 = pi10 ? n53537 : n53608;
  assign n53610 = pi09 ? n32 : n53609;
  assign n53611 = pi15 ? n23981 : n39243;
  assign n53612 = pi14 ? n53611 : n53544;
  assign n53613 = pi13 ? n53538 : n53612;
  assign n53614 = pi18 ? n248 : n53547;
  assign n53615 = pi17 ? n32 : n53614;
  assign n53616 = pi16 ? n32 : n53615;
  assign n53617 = pi20 ? n274 : n17712;
  assign n53618 = pi19 ? n53617 : n32;
  assign n53619 = pi19 ? n267 : ~n10890;
  assign n53620 = pi18 ? n53618 : n53619;
  assign n53621 = pi17 ? n32 : n53620;
  assign n53622 = pi16 ? n32 : n53621;
  assign n53623 = pi15 ? n53616 : n53622;
  assign n53624 = pi15 ? n38371 : n16105;
  assign n53625 = pi14 ? n53623 : n53624;
  assign n53626 = pi15 ? n32 : n53421;
  assign n53627 = pi14 ? n23574 : n53626;
  assign n53628 = pi13 ? n53625 : n53627;
  assign n53629 = pi12 ? n53613 : n53628;
  assign n53630 = pi15 ? n37644 : n14790;
  assign n53631 = pi14 ? n53630 : n53575;
  assign n53632 = pi15 ? n14397 : n15263;
  assign n53633 = pi14 ? n53632 : n22437;
  assign n53634 = pi13 ? n53631 : n53633;
  assign n53635 = pi17 ? n2954 : ~n2517;
  assign n53636 = pi16 ? n32 : n53635;
  assign n53637 = pi15 ? n14147 : n53636;
  assign n53638 = pi17 ? n3569 : ~n53584;
  assign n53639 = pi16 ? n32 : n53638;
  assign n53640 = pi17 ? n3569 : ~n38897;
  assign n53641 = pi16 ? n32 : n53640;
  assign n53642 = pi15 ? n53639 : n53641;
  assign n53643 = pi14 ? n53637 : n53642;
  assign n53644 = pi14 ? n39370 : n53604;
  assign n53645 = pi13 ? n53643 : n53644;
  assign n53646 = pi12 ? n53634 : n53645;
  assign n53647 = pi11 ? n53629 : n53646;
  assign n53648 = pi10 ? n53537 : n53647;
  assign n53649 = pi09 ? n32 : n53648;
  assign n53650 = pi08 ? n53610 : n53649;
  assign n53651 = pi07 ? n53529 : n53650;
  assign n53652 = pi06 ? n53361 : n53651;
  assign n53653 = pi05 ? n53105 : n53652;
  assign n53654 = pi14 ? n16392 : n53362;
  assign n53655 = pi13 ? n53654 : n32;
  assign n53656 = pi15 ? n32 : n26322;
  assign n53657 = pi19 ? n32 : n52197;
  assign n53658 = pi18 ? n32 : n53657;
  assign n53659 = pi17 ? n32 : n53658;
  assign n53660 = pi16 ? n32 : n53659;
  assign n53661 = pi15 ? n53660 : n17039;
  assign n53662 = pi14 ? n53656 : n53661;
  assign n53663 = pi15 ? n16101 : n16452;
  assign n53664 = pi15 ? n16101 : n24874;
  assign n53665 = pi14 ? n53663 : n53664;
  assign n53666 = pi13 ? n53662 : n53665;
  assign n53667 = pi12 ? n53655 : n53666;
  assign n53668 = pi11 ? n39288 : n53667;
  assign n53669 = pi19 ? n322 : n4670;
  assign n53670 = pi18 ? n32 : n53669;
  assign n53671 = pi17 ? n32 : n53670;
  assign n53672 = pi16 ? n32 : n53671;
  assign n53673 = pi15 ? n53672 : n24659;
  assign n53674 = pi15 ? n38371 : n16293;
  assign n53675 = pi14 ? n53673 : n53674;
  assign n53676 = pi15 ? n16101 : n27686;
  assign n53677 = pi18 ? n268 : n53471;
  assign n53678 = pi17 ? n32 : n53677;
  assign n53679 = pi16 ? n32 : n53678;
  assign n53680 = pi18 ? n16847 : n6645;
  assign n53681 = pi17 ? n32 : n53680;
  assign n53682 = pi16 ? n32 : n53681;
  assign n53683 = pi15 ? n53679 : n53682;
  assign n53684 = pi14 ? n53676 : n53683;
  assign n53685 = pi13 ? n53675 : n53684;
  assign n53686 = pi19 ? n322 : ~n6652;
  assign n53687 = pi18 ? n32 : n53686;
  assign n53688 = pi17 ? n32 : n53687;
  assign n53689 = pi16 ? n32 : n53688;
  assign n53690 = pi15 ? n53689 : n37501;
  assign n53691 = pi14 ? n53690 : n16105;
  assign n53692 = pi19 ? n8662 : n358;
  assign n53693 = pi18 ? n32 : n53692;
  assign n53694 = pi17 ? n32 : n53693;
  assign n53695 = pi16 ? n32 : n53694;
  assign n53696 = pi15 ? n21543 : n53695;
  assign n53697 = pi14 ? n32 : n53696;
  assign n53698 = pi13 ? n53691 : n53697;
  assign n53699 = pi12 ? n53685 : n53698;
  assign n53700 = pi19 ? n6398 : ~n2614;
  assign n53701 = pi18 ? n32 : n53700;
  assign n53702 = pi17 ? n32 : n53701;
  assign n53703 = pi16 ? n32 : n53702;
  assign n53704 = pi15 ? n24659 : n53703;
  assign n53705 = pi18 ? n32 : n29718;
  assign n53706 = pi17 ? n32 : n53705;
  assign n53707 = pi16 ? n32 : n53706;
  assign n53708 = pi15 ? n53707 : n13948;
  assign n53709 = pi14 ? n53704 : n53708;
  assign n53710 = pi15 ? n40063 : n14967;
  assign n53711 = pi15 ? n14967 : n21853;
  assign n53712 = pi14 ? n53710 : n53711;
  assign n53713 = pi13 ? n53709 : n53712;
  assign n53714 = pi19 ? n28177 : ~n32;
  assign n53715 = pi18 ? n350 : ~n53714;
  assign n53716 = pi17 ? n32 : n53715;
  assign n53717 = pi16 ? n32 : n53716;
  assign n53718 = pi18 ? n3350 : ~n532;
  assign n53719 = pi17 ? n32 : n53718;
  assign n53720 = pi16 ? n32 : n53719;
  assign n53721 = pi15 ? n53717 : n53720;
  assign n53722 = pi18 ? n5436 : ~n28193;
  assign n53723 = pi17 ? n32 : n53722;
  assign n53724 = pi16 ? n32 : n53723;
  assign n53725 = pi19 ? n1686 : ~n32;
  assign n53726 = pi18 ? n53725 : ~n323;
  assign n53727 = pi17 ? n32 : n53726;
  assign n53728 = pi16 ? n32 : n53727;
  assign n53729 = pi15 ? n53724 : n53728;
  assign n53730 = pi14 ? n53721 : n53729;
  assign n53731 = pi18 ? n31385 : ~n532;
  assign n53732 = pi17 ? n32 : n53731;
  assign n53733 = pi16 ? n32 : n53732;
  assign n53734 = pi20 ? n53173 : ~n32;
  assign n53735 = pi19 ? n53734 : ~n32;
  assign n53736 = pi18 ? n53735 : ~n20788;
  assign n53737 = pi17 ? n32 : n53736;
  assign n53738 = pi16 ? n32 : n53737;
  assign n53739 = pi15 ? n53733 : n53738;
  assign n53740 = pi18 ? n53735 : ~n532;
  assign n53741 = pi17 ? n32 : n53740;
  assign n53742 = pi16 ? n32 : n53741;
  assign n53743 = pi15 ? n53742 : n29701;
  assign n53744 = pi14 ? n53739 : n53743;
  assign n53745 = pi13 ? n53730 : n53744;
  assign n53746 = pi12 ? n53713 : n53745;
  assign n53747 = pi11 ? n53699 : n53746;
  assign n53748 = pi10 ? n53668 : n53747;
  assign n53749 = pi09 ? n32 : n53748;
  assign n53750 = pi15 ? n16832 : n16397;
  assign n53751 = pi14 ? n16392 : n53750;
  assign n53752 = pi13 ? n53751 : n32;
  assign n53753 = pi12 ? n53752 : n53666;
  assign n53754 = pi11 ? n39288 : n53753;
  assign n53755 = pi15 ? n38371 : n16298;
  assign n53756 = pi14 ? n53673 : n53755;
  assign n53757 = pi15 ? n16101 : n40632;
  assign n53758 = pi14 ? n53757 : n53683;
  assign n53759 = pi13 ? n53756 : n53758;
  assign n53760 = pi19 ? n1464 : n15651;
  assign n53761 = pi18 ? n32 : n53760;
  assign n53762 = pi17 ? n32 : n53761;
  assign n53763 = pi16 ? n32 : n53762;
  assign n53764 = pi15 ? n21853 : n53763;
  assign n53765 = pi14 ? n32 : n53764;
  assign n53766 = pi13 ? n53691 : n53765;
  assign n53767 = pi12 ? n53759 : n53766;
  assign n53768 = pi15 ? n24659 : n22923;
  assign n53769 = pi15 ? n22540 : n13948;
  assign n53770 = pi14 ? n53768 : n53769;
  assign n53771 = pi15 ? n40063 : n22437;
  assign n53772 = pi14 ? n53771 : n26788;
  assign n53773 = pi13 ? n53770 : n53772;
  assign n53774 = pi17 ? n32 : n45327;
  assign n53775 = pi16 ? n32 : n53774;
  assign n53776 = pi15 ? n53775 : n46562;
  assign n53777 = pi20 ? n151 : ~n32;
  assign n53778 = pi19 ? n53777 : ~n32;
  assign n53779 = pi18 ? n53778 : ~n323;
  assign n53780 = pi17 ? n32 : n53779;
  assign n53781 = pi16 ? n32 : n53780;
  assign n53782 = pi15 ? n53724 : n53781;
  assign n53783 = pi14 ? n53776 : n53782;
  assign n53784 = pi18 ? n344 : ~n20788;
  assign n53785 = pi17 ? n32 : n53784;
  assign n53786 = pi16 ? n32 : n53785;
  assign n53787 = pi15 ? n39449 : n53786;
  assign n53788 = pi18 ? n1541 : n4492;
  assign n53789 = pi17 ? n32 : n53788;
  assign n53790 = pi16 ? n32 : n53789;
  assign n53791 = pi15 ? n39449 : n53790;
  assign n53792 = pi14 ? n53787 : n53791;
  assign n53793 = pi13 ? n53783 : n53792;
  assign n53794 = pi12 ? n53773 : n53793;
  assign n53795 = pi11 ? n53767 : n53794;
  assign n53796 = pi10 ? n53754 : n53795;
  assign n53797 = pi09 ? n32 : n53796;
  assign n53798 = pi08 ? n53749 : n53797;
  assign n53799 = pi13 ? n53751 : n38860;
  assign n53800 = pi19 ? n32 : n28179;
  assign n53801 = pi18 ? n32 : n53800;
  assign n53802 = pi17 ? n32 : n53801;
  assign n53803 = pi16 ? n32 : n53802;
  assign n53804 = pi15 ? n53803 : n16837;
  assign n53805 = pi14 ? n39388 : n53804;
  assign n53806 = pi15 ? n25211 : n15403;
  assign n53807 = pi14 ? n53664 : n53806;
  assign n53808 = pi13 ? n53805 : n53807;
  assign n53809 = pi12 ? n53799 : n53808;
  assign n53810 = pi11 ? n39288 : n53809;
  assign n53811 = pi19 ? n322 : n7642;
  assign n53812 = pi18 ? n32 : n53811;
  assign n53813 = pi17 ? n32 : n53812;
  assign n53814 = pi16 ? n32 : n53813;
  assign n53815 = pi15 ? n53814 : n14917;
  assign n53816 = pi15 ? n39474 : n16204;
  assign n53817 = pi14 ? n53815 : n53816;
  assign n53818 = pi19 ? n19773 : n267;
  assign n53819 = pi19 ? n2359 : ~n11117;
  assign n53820 = pi18 ? n53818 : n53819;
  assign n53821 = pi17 ? n32 : n53820;
  assign n53822 = pi16 ? n32 : n53821;
  assign n53823 = pi19 ? n19773 : n5694;
  assign n53824 = pi18 ? n53823 : n6645;
  assign n53825 = pi17 ? n32 : n53824;
  assign n53826 = pi16 ? n32 : n53825;
  assign n53827 = pi15 ? n53822 : n53826;
  assign n53828 = pi14 ? n40632 : n53827;
  assign n53829 = pi13 ? n53817 : n53828;
  assign n53830 = pi21 ? n14399 : ~n32;
  assign n53831 = pi20 ? n53830 : ~n32;
  assign n53832 = pi19 ? n322 : ~n53831;
  assign n53833 = pi18 ? n9170 : n53832;
  assign n53834 = pi17 ? n32 : n53833;
  assign n53835 = pi16 ? n32 : n53834;
  assign n53836 = pi19 ? n16597 : n6057;
  assign n53837 = pi18 ? n53836 : n6600;
  assign n53838 = pi17 ? n32 : n53837;
  assign n53839 = pi16 ? n32 : n53838;
  assign n53840 = pi15 ? n53835 : n53839;
  assign n53841 = pi14 ? n53840 : n16218;
  assign n53842 = pi15 ? n21853 : n23169;
  assign n53843 = pi15 ? n23169 : n24659;
  assign n53844 = pi14 ? n53842 : n53843;
  assign n53845 = pi13 ? n53841 : n53844;
  assign n53846 = pi12 ? n53829 : n53845;
  assign n53847 = pi14 ? n48187 : n24555;
  assign n53848 = pi15 ? n14397 : n22437;
  assign n53849 = pi14 ? n53848 : n32;
  assign n53850 = pi13 ? n53847 : n53849;
  assign n53851 = pi17 ? n32 : n21894;
  assign n53852 = pi16 ? n32 : n53851;
  assign n53853 = pi19 ? n14022 : ~n32;
  assign n53854 = pi18 ? n344 : ~n53853;
  assign n53855 = pi17 ? n32 : n53854;
  assign n53856 = pi16 ? n32 : n53855;
  assign n53857 = pi15 ? n53852 : n53856;
  assign n53858 = pi20 ? n101 : ~n357;
  assign n53859 = pi19 ? n53858 : ~n32;
  assign n53860 = pi18 ? n53859 : ~n323;
  assign n53861 = pi17 ? n32 : n53860;
  assign n53862 = pi16 ? n32 : n53861;
  assign n53863 = pi18 ? n418 : ~n22159;
  assign n53864 = pi17 ? n32 : n53863;
  assign n53865 = pi16 ? n32 : n53864;
  assign n53866 = pi15 ? n53862 : n53865;
  assign n53867 = pi14 ? n53857 : n53866;
  assign n53868 = pi18 ? n1405 : ~n20788;
  assign n53869 = pi17 ? n32 : n53868;
  assign n53870 = pi16 ? n32 : n53869;
  assign n53871 = pi15 ? n39540 : n53870;
  assign n53872 = pi19 ? n8622 : n462;
  assign n53873 = pi18 ? n53872 : n20298;
  assign n53874 = pi17 ? n32 : n53873;
  assign n53875 = pi16 ? n32 : n53874;
  assign n53876 = pi15 ? n39540 : n53875;
  assign n53877 = pi14 ? n53871 : n53876;
  assign n53878 = pi13 ? n53867 : n53877;
  assign n53879 = pi12 ? n53850 : n53878;
  assign n53880 = pi11 ? n53846 : n53879;
  assign n53881 = pi10 ? n53810 : n53880;
  assign n53882 = pi09 ? n32 : n53881;
  assign n53883 = pi15 ? n25763 : n16397;
  assign n53884 = pi14 ? n16832 : n53883;
  assign n53885 = pi13 ? n53884 : n38860;
  assign n53886 = pi12 ? n53885 : n53808;
  assign n53887 = pi11 ? n39288 : n53886;
  assign n53888 = pi15 ? n24247 : n16204;
  assign n53889 = pi14 ? n53815 : n53888;
  assign n53890 = pi21 ? n7500 : ~n206;
  assign n53891 = pi20 ? n53890 : n32;
  assign n53892 = pi19 ? n32 : n53891;
  assign n53893 = pi18 ? n32 : n53892;
  assign n53894 = pi17 ? n32 : n53893;
  assign n53895 = pi16 ? n32 : n53894;
  assign n53896 = pi15 ? n40632 : n53895;
  assign n53897 = pi18 ? n268 : n53819;
  assign n53898 = pi17 ? n32 : n53897;
  assign n53899 = pi16 ? n32 : n53898;
  assign n53900 = pi19 ? n1138 : ~n12245;
  assign n53901 = pi18 ? n16847 : n53900;
  assign n53902 = pi17 ? n32 : n53901;
  assign n53903 = pi16 ? n32 : n53902;
  assign n53904 = pi15 ? n53899 : n53903;
  assign n53905 = pi14 ? n53896 : n53904;
  assign n53906 = pi13 ? n53889 : n53905;
  assign n53907 = pi19 ? n1138 : ~n813;
  assign n53908 = pi18 ? n32 : n53907;
  assign n53909 = pi17 ? n32 : n53908;
  assign n53910 = pi16 ? n32 : n53909;
  assign n53911 = pi19 ? n322 : n7488;
  assign n53912 = pi18 ? n32 : n53911;
  assign n53913 = pi17 ? n32 : n53912;
  assign n53914 = pi16 ? n32 : n53913;
  assign n53915 = pi15 ? n53910 : n53914;
  assign n53916 = pi15 ? n24289 : n23574;
  assign n53917 = pi14 ? n53915 : n53916;
  assign n53918 = pi15 ? n39812 : n37644;
  assign n53919 = pi15 ? n37644 : n24659;
  assign n53920 = pi14 ? n53918 : n53919;
  assign n53921 = pi13 ? n53917 : n53920;
  assign n53922 = pi12 ? n53906 : n53921;
  assign n53923 = pi15 ? n22817 : n658;
  assign n53924 = pi19 ? n21065 : n32;
  assign n53925 = pi18 ? n32 : n53924;
  assign n53926 = pi17 ? n32 : n53925;
  assign n53927 = pi16 ? n32 : n53926;
  assign n53928 = pi15 ? n21954 : n53927;
  assign n53929 = pi14 ? n53923 : n53928;
  assign n53930 = pi19 ? n334 : n32;
  assign n53931 = pi18 ? n32 : n53930;
  assign n53932 = pi17 ? n32 : n53931;
  assign n53933 = pi16 ? n32 : n53932;
  assign n53934 = pi15 ? n53933 : n21853;
  assign n53935 = pi14 ? n53934 : n32;
  assign n53936 = pi13 ? n53929 : n53935;
  assign n53937 = pi18 ? n2424 : ~n323;
  assign n53938 = pi17 ? n32 : n53937;
  assign n53939 = pi16 ? n32 : n53938;
  assign n53940 = pi15 ? n10721 : n53939;
  assign n53941 = pi14 ? n53940 : n39536;
  assign n53942 = pi18 ? n605 : ~n20788;
  assign n53943 = pi17 ? n32 : n53942;
  assign n53944 = pi16 ? n32 : n53943;
  assign n53945 = pi15 ? n39540 : n53944;
  assign n53946 = pi20 ? n141 : ~n439;
  assign n53947 = pi19 ? n594 : ~n53946;
  assign n53948 = pi18 ? n53947 : n20298;
  assign n53949 = pi17 ? n32 : n53948;
  assign n53950 = pi16 ? n32 : n53949;
  assign n53951 = pi15 ? n39540 : n53950;
  assign n53952 = pi14 ? n53945 : n53951;
  assign n53953 = pi13 ? n53941 : n53952;
  assign n53954 = pi12 ? n53936 : n53953;
  assign n53955 = pi11 ? n53922 : n53954;
  assign n53956 = pi10 ? n53887 : n53955;
  assign n53957 = pi09 ? n32 : n53956;
  assign n53958 = pi08 ? n53882 : n53957;
  assign n53959 = pi07 ? n53798 : n53958;
  assign n53960 = pi19 ? n32 : n13916;
  assign n53961 = pi18 ? n32 : n53960;
  assign n53962 = pi17 ? n32 : n53961;
  assign n53963 = pi16 ? n32 : n53962;
  assign n53964 = pi15 ? n53963 : n16397;
  assign n53965 = pi14 ? n16832 : n53964;
  assign n53966 = pi19 ? n32 : n6342;
  assign n53967 = pi18 ? n32 : n53966;
  assign n53968 = pi17 ? n32 : n53967;
  assign n53969 = pi16 ? n32 : n53968;
  assign n53970 = pi15 ? n16452 : n53969;
  assign n53971 = pi14 ? n32 : n53970;
  assign n53972 = pi13 ? n53965 : n53971;
  assign n53973 = pi15 ? n16804 : n24874;
  assign n53974 = pi14 ? n39556 : n53973;
  assign n53975 = pi15 ? n38065 : n16193;
  assign n53976 = pi14 ? n40109 : n53975;
  assign n53977 = pi13 ? n53974 : n53976;
  assign n53978 = pi12 ? n53972 : n53977;
  assign n53979 = pi11 ? n39288 : n53978;
  assign n53980 = pi15 ? n16193 : n24504;
  assign n53981 = pi21 ? n1939 : n309;
  assign n53982 = pi20 ? n53981 : n32;
  assign n53983 = pi19 ? n32 : n53982;
  assign n53984 = pi18 ? n32 : n53983;
  assign n53985 = pi17 ? n32 : n53984;
  assign n53986 = pi16 ? n32 : n53985;
  assign n53987 = pi15 ? n39243 : n53986;
  assign n53988 = pi14 ? n53980 : n53987;
  assign n53989 = pi21 ? n66 : n14158;
  assign n53990 = pi20 ? n53989 : n32;
  assign n53991 = pi19 ? n32 : n53990;
  assign n53992 = pi18 ? n32 : n53991;
  assign n53993 = pi17 ? n32 : n53992;
  assign n53994 = pi16 ? n32 : n53993;
  assign n53995 = pi19 ? n267 : ~n1941;
  assign n53996 = pi18 ? n32 : n53995;
  assign n53997 = pi17 ? n32 : n53996;
  assign n53998 = pi16 ? n32 : n53997;
  assign n53999 = pi15 ? n53994 : n53998;
  assign n54000 = pi19 ? n4391 : ~n1941;
  assign n54001 = pi18 ? n16847 : n54000;
  assign n54002 = pi17 ? n32 : n54001;
  assign n54003 = pi16 ? n32 : n54002;
  assign n54004 = pi18 ? n15849 : ~n496;
  assign n54005 = pi17 ? n32 : n54004;
  assign n54006 = pi16 ? n32 : n54005;
  assign n54007 = pi15 ? n54003 : n54006;
  assign n54008 = pi14 ? n53999 : n54007;
  assign n54009 = pi13 ? n53988 : n54008;
  assign n54010 = pi18 ? n17063 : n24981;
  assign n54011 = pi17 ? n32 : n54010;
  assign n54012 = pi16 ? n32 : n54011;
  assign n54013 = pi19 ? n322 : n26833;
  assign n54014 = pi18 ? n32 : n54013;
  assign n54015 = pi17 ? n32 : n54014;
  assign n54016 = pi16 ? n32 : n54015;
  assign n54017 = pi15 ? n54012 : n54016;
  assign n54018 = pi14 ? n54017 : n32;
  assign n54019 = pi14 ? n23484 : n23749;
  assign n54020 = pi13 ? n54018 : n54019;
  assign n54021 = pi12 ? n54009 : n54020;
  assign n54022 = pi20 ? n32 : n9628;
  assign n54023 = pi19 ? n54022 : n32;
  assign n54024 = pi18 ? n32 : n54023;
  assign n54025 = pi17 ? n32 : n54024;
  assign n54026 = pi16 ? n32 : n54025;
  assign n54027 = pi15 ? n54026 : n21801;
  assign n54028 = pi20 ? n32 : ~n8630;
  assign n54029 = pi19 ? n54028 : n32;
  assign n54030 = pi18 ? n32 : n54029;
  assign n54031 = pi17 ? n32 : n54030;
  assign n54032 = pi16 ? n32 : n54031;
  assign n54033 = pi15 ? n54032 : n39887;
  assign n54034 = pi14 ? n54027 : n54033;
  assign n54035 = pi22 ? n65 : n84;
  assign n54036 = pi21 ? n174 : n54035;
  assign n54037 = pi20 ? n32 : n54036;
  assign n54038 = pi19 ? n54037 : n32;
  assign n54039 = pi18 ? n32 : n54038;
  assign n54040 = pi17 ? n32 : n54039;
  assign n54041 = pi16 ? n32 : n54040;
  assign n54042 = pi15 ? n54041 : n39582;
  assign n54043 = pi20 ? n32 : n9367;
  assign n54044 = pi19 ? n54043 : ~n32;
  assign n54045 = pi18 ? n508 : ~n54044;
  assign n54046 = pi17 ? n32 : n54045;
  assign n54047 = pi16 ? n32 : n54046;
  assign n54048 = pi15 ? n13369 : n54047;
  assign n54049 = pi14 ? n54042 : n54048;
  assign n54050 = pi13 ? n54034 : n54049;
  assign n54051 = pi18 ? n1712 : ~n39598;
  assign n54052 = pi17 ? n32 : n54051;
  assign n54053 = pi16 ? n32 : n54052;
  assign n54054 = pi19 ? n4518 : ~n32;
  assign n54055 = pi18 ? n54054 : ~n22159;
  assign n54056 = pi17 ? n32 : n54055;
  assign n54057 = pi16 ? n32 : n54056;
  assign n54058 = pi15 ? n54053 : n54057;
  assign n54059 = pi14 ? n11194 : n54058;
  assign n54060 = pi19 ? n32 : ~n17766;
  assign n54061 = pi18 ? n54060 : n13080;
  assign n54062 = pi17 ? n32 : n54061;
  assign n54063 = pi16 ? n32 : n54062;
  assign n54064 = pi15 ? n54063 : n44497;
  assign n54065 = pi18 ? n595 : ~n532;
  assign n54066 = pi17 ? n32 : n54065;
  assign n54067 = pi16 ? n32 : n54066;
  assign n54068 = pi15 ? n54067 : n39613;
  assign n54069 = pi14 ? n54064 : n54068;
  assign n54070 = pi13 ? n54059 : n54069;
  assign n54071 = pi12 ? n54050 : n54070;
  assign n54072 = pi11 ? n54021 : n54071;
  assign n54073 = pi10 ? n53979 : n54072;
  assign n54074 = pi09 ? n32 : n54073;
  assign n54075 = pi11 ? n39623 : n53978;
  assign n54076 = pi15 ? n39243 : n25301;
  assign n54077 = pi14 ? n53980 : n54076;
  assign n54078 = pi15 ? n26990 : n53998;
  assign n54079 = pi14 ? n54078 : n54007;
  assign n54080 = pi13 ? n54077 : n54079;
  assign n54081 = pi18 ? n6071 : n24981;
  assign n54082 = pi17 ? n32 : n54081;
  assign n54083 = pi16 ? n32 : n54082;
  assign n54084 = pi15 ? n54083 : n54016;
  assign n54085 = pi14 ? n54084 : n32;
  assign n54086 = pi14 ? n23484 : n24909;
  assign n54087 = pi13 ? n54085 : n54086;
  assign n54088 = pi12 ? n54080 : n54087;
  assign n54089 = pi15 ? n54026 : n14156;
  assign n54090 = pi15 ? n14147 : n34846;
  assign n54091 = pi14 ? n54089 : n54090;
  assign n54092 = pi21 ? n174 : ~n6898;
  assign n54093 = pi20 ? n32 : n54092;
  assign n54094 = pi19 ? n54093 : n32;
  assign n54095 = pi18 ? n32 : n54094;
  assign n54096 = pi17 ? n32 : n54095;
  assign n54097 = pi16 ? n32 : n54096;
  assign n54098 = pi15 ? n54097 : n14798;
  assign n54099 = pi18 ? n508 : ~n1405;
  assign n54100 = pi17 ? n32 : n54099;
  assign n54101 = pi16 ? n32 : n54100;
  assign n54102 = pi15 ? n13369 : n54101;
  assign n54103 = pi14 ? n54098 : n54102;
  assign n54104 = pi13 ? n54091 : n54103;
  assign n54105 = pi15 ? n11202 : n11198;
  assign n54106 = pi18 ? n6235 : ~n532;
  assign n54107 = pi17 ? n32 : n54106;
  assign n54108 = pi16 ? n32 : n54107;
  assign n54109 = pi15 ? n54108 : n33135;
  assign n54110 = pi14 ? n54105 : n54109;
  assign n54111 = pi15 ? n54063 : n33135;
  assign n54112 = pi14 ? n54111 : n39653;
  assign n54113 = pi13 ? n54110 : n54112;
  assign n54114 = pi12 ? n54104 : n54113;
  assign n54115 = pi11 ? n54088 : n54114;
  assign n54116 = pi10 ? n54075 : n54115;
  assign n54117 = pi09 ? n32 : n54116;
  assign n54118 = pi08 ? n54074 : n54117;
  assign n54119 = pi15 ? n53119 : n16736;
  assign n54120 = pi14 ? n17036 : n54119;
  assign n54121 = pi13 ? n54120 : n53971;
  assign n54122 = pi19 ? n32 : n7427;
  assign n54123 = pi18 ? n32 : n54122;
  assign n54124 = pi17 ? n32 : n54123;
  assign n54125 = pi16 ? n32 : n54124;
  assign n54126 = pi15 ? n38065 : n54125;
  assign n54127 = pi14 ? n40109 : n54126;
  assign n54128 = pi13 ? n53974 : n54127;
  assign n54129 = pi12 ? n54121 : n54128;
  assign n54130 = pi11 ? n39623 : n54129;
  assign n54131 = pi19 ? n32 : n7661;
  assign n54132 = pi18 ? n32 : n54131;
  assign n54133 = pi17 ? n32 : n54132;
  assign n54134 = pi16 ? n32 : n54133;
  assign n54135 = pi15 ? n54134 : n24712;
  assign n54136 = pi19 ? n322 : n7412;
  assign n54137 = pi18 ? n32 : n54136;
  assign n54138 = pi17 ? n32 : n54137;
  assign n54139 = pi16 ? n32 : n54138;
  assign n54140 = pi15 ? n54139 : n27304;
  assign n54141 = pi14 ? n54135 : n54140;
  assign n54142 = pi19 ? n358 : n19847;
  assign n54143 = pi18 ? n32 : n54142;
  assign n54144 = pi17 ? n32 : n54143;
  assign n54145 = pi16 ? n32 : n54144;
  assign n54146 = pi19 ? n36073 : ~n1941;
  assign n54147 = pi18 ? n16834 : n54146;
  assign n54148 = pi17 ? n32 : n54147;
  assign n54149 = pi16 ? n32 : n54148;
  assign n54150 = pi15 ? n54145 : n54149;
  assign n54151 = pi20 ? n175 : ~n321;
  assign n54152 = pi19 ? n32 : n54151;
  assign n54153 = pi21 ? n66 : n259;
  assign n54154 = pi20 ? n54153 : ~n32;
  assign n54155 = pi19 ? n47028 : ~n54154;
  assign n54156 = pi18 ? n54152 : n54155;
  assign n54157 = pi17 ? n32 : n54156;
  assign n54158 = pi16 ? n32 : n54157;
  assign n54159 = pi20 ? n915 : n321;
  assign n54160 = pi19 ? n594 : ~n54159;
  assign n54161 = pi18 ? n54160 : ~n590;
  assign n54162 = pi17 ? n32 : n54161;
  assign n54163 = pi16 ? n32 : n54162;
  assign n54164 = pi15 ? n54158 : n54163;
  assign n54165 = pi14 ? n54150 : n54164;
  assign n54166 = pi13 ? n54141 : n54165;
  assign n54167 = pi19 ? n531 : ~n39789;
  assign n54168 = pi18 ? n32 : n54167;
  assign n54169 = pi17 ? n32 : n54168;
  assign n54170 = pi16 ? n32 : n54169;
  assign n54171 = pi19 ? n322 : n15696;
  assign n54172 = pi18 ? n32 : n54171;
  assign n54173 = pi17 ? n32 : n54172;
  assign n54174 = pi16 ? n32 : n54173;
  assign n54175 = pi15 ? n54170 : n54174;
  assign n54176 = pi14 ? n54175 : n32;
  assign n54177 = pi19 ? n275 : ~n236;
  assign n54178 = pi18 ? n32 : n54177;
  assign n54179 = pi17 ? n32 : n54178;
  assign n54180 = pi16 ? n32 : n54179;
  assign n54181 = pi15 ? n23749 : n54180;
  assign n54182 = pi14 ? n23484 : n54181;
  assign n54183 = pi13 ? n54176 : n54182;
  assign n54184 = pi12 ? n54166 : n54183;
  assign n54185 = pi20 ? n32 : n100;
  assign n54186 = pi19 ? n54185 : n32;
  assign n54187 = pi18 ? n32 : n54186;
  assign n54188 = pi17 ? n32 : n54187;
  assign n54189 = pi16 ? n32 : n54188;
  assign n54190 = pi15 ? n54189 : n14156;
  assign n54191 = pi21 ? n174 : ~n100;
  assign n54192 = pi20 ? n32 : n54191;
  assign n54193 = pi19 ? n54192 : n32;
  assign n54194 = pi18 ? n32 : n54193;
  assign n54195 = pi17 ? n32 : n54194;
  assign n54196 = pi16 ? n32 : n54195;
  assign n54197 = pi15 ? n13948 : n54196;
  assign n54198 = pi14 ? n54190 : n54197;
  assign n54199 = pi21 ? n405 : ~n10445;
  assign n54200 = pi20 ? n32 : n54199;
  assign n54201 = pi19 ? n54200 : n32;
  assign n54202 = pi18 ? n32 : n54201;
  assign n54203 = pi17 ? n32 : n54202;
  assign n54204 = pi16 ? n32 : n54203;
  assign n54205 = pi15 ? n22347 : n54204;
  assign n54206 = pi15 ? n33939 : n11650;
  assign n54207 = pi14 ? n54205 : n54206;
  assign n54208 = pi13 ? n54198 : n54207;
  assign n54209 = pi20 ? n32 : n7013;
  assign n54210 = pi19 ? n54209 : ~n32;
  assign n54211 = pi18 ? n702 : ~n54210;
  assign n54212 = pi17 ? n32 : n54211;
  assign n54213 = pi16 ? n32 : n54212;
  assign n54214 = pi15 ? n11423 : n54213;
  assign n54215 = pi18 ? n962 : ~n532;
  assign n54216 = pi17 ? n32 : n54215;
  assign n54217 = pi16 ? n32 : n54216;
  assign n54218 = pi14 ? n54214 : n54217;
  assign n54219 = pi20 ? n915 : ~n32;
  assign n54220 = pi19 ? n54219 : ~n32;
  assign n54221 = pi18 ? n9038 : ~n54220;
  assign n54222 = pi17 ? n32 : n54221;
  assign n54223 = pi16 ? n32 : n54222;
  assign n54224 = pi15 ? n54223 : n33618;
  assign n54225 = pi18 ? n4407 : ~n418;
  assign n54226 = pi17 ? n32 : n54225;
  assign n54227 = pi16 ? n32 : n54226;
  assign n54228 = pi15 ? n54227 : n39713;
  assign n54229 = pi14 ? n54224 : n54228;
  assign n54230 = pi13 ? n54218 : n54229;
  assign n54231 = pi12 ? n54208 : n54230;
  assign n54232 = pi11 ? n54184 : n54231;
  assign n54233 = pi10 ? n54130 : n54232;
  assign n54234 = pi09 ? n32 : n54233;
  assign n54235 = pi12 ? n54121 : n53977;
  assign n54236 = pi11 ? n39623 : n54235;
  assign n54237 = pi15 ? n24504 : n25044;
  assign n54238 = pi19 ? n322 : n7443;
  assign n54239 = pi18 ? n32 : n54238;
  assign n54240 = pi17 ? n32 : n54239;
  assign n54241 = pi16 ? n32 : n54240;
  assign n54242 = pi15 ? n54241 : n27304;
  assign n54243 = pi14 ? n54237 : n54242;
  assign n54244 = pi19 ? n358 : n19749;
  assign n54245 = pi18 ? n16962 : n54244;
  assign n54246 = pi17 ? n32 : n54245;
  assign n54247 = pi16 ? n32 : n54246;
  assign n54248 = pi19 ? n5371 : n1941;
  assign n54249 = pi18 ? n16389 : ~n54248;
  assign n54250 = pi17 ? n32 : n54249;
  assign n54251 = pi16 ? n32 : n54250;
  assign n54252 = pi15 ? n54247 : n54251;
  assign n54253 = pi19 ? n9007 : n589;
  assign n54254 = pi18 ? n16394 : ~n54253;
  assign n54255 = pi17 ? n32 : n54254;
  assign n54256 = pi16 ? n32 : n54255;
  assign n54257 = pi18 ? n15849 : ~n590;
  assign n54258 = pi17 ? n32 : n54257;
  assign n54259 = pi16 ? n32 : n54258;
  assign n54260 = pi15 ? n54256 : n54259;
  assign n54261 = pi14 ? n54252 : n54260;
  assign n54262 = pi13 ? n54243 : n54261;
  assign n54263 = pi14 ? n35176 : n54181;
  assign n54264 = pi13 ? n54176 : n54263;
  assign n54265 = pi12 ? n54262 : n54264;
  assign n54266 = pi21 ? n1939 : n405;
  assign n54267 = pi20 ? n32 : n54266;
  assign n54268 = pi19 ? n54267 : n32;
  assign n54269 = pi18 ? n32 : n54268;
  assign n54270 = pi17 ? n32 : n54269;
  assign n54271 = pi16 ? n32 : n54270;
  assign n54272 = pi15 ? n54271 : n14156;
  assign n54273 = pi14 ? n54272 : n54197;
  assign n54274 = pi15 ? n15123 : n22381;
  assign n54275 = pi14 ? n54274 : n54206;
  assign n54276 = pi13 ? n54273 : n54275;
  assign n54277 = pi18 ? n496 : ~n54210;
  assign n54278 = pi17 ? n32 : n54277;
  assign n54279 = pi16 ? n32 : n54278;
  assign n54280 = pi15 ? n45941 : n54279;
  assign n54281 = pi14 ? n54280 : n33448;
  assign n54282 = pi20 ? n1324 : n501;
  assign n54283 = pi19 ? n32 : n54282;
  assign n54284 = pi18 ? n54283 : ~n44347;
  assign n54285 = pi17 ? n32 : n54284;
  assign n54286 = pi16 ? n32 : n54285;
  assign n54287 = pi15 ? n54286 : n33448;
  assign n54288 = pi14 ? n54287 : n39747;
  assign n54289 = pi13 ? n54281 : n54288;
  assign n54290 = pi12 ? n54276 : n54289;
  assign n54291 = pi11 ? n54265 : n54290;
  assign n54292 = pi10 ? n54236 : n54291;
  assign n54293 = pi09 ? n32 : n54292;
  assign n54294 = pi08 ? n54234 : n54293;
  assign n54295 = pi07 ? n54118 : n54294;
  assign n54296 = pi06 ? n53959 : n54295;
  assign n54297 = pi15 ? n16736 : n16850;
  assign n54298 = pi14 ? n26161 : n54297;
  assign n54299 = pi14 ? n24247 : n26163;
  assign n54300 = pi13 ? n54298 : n54299;
  assign n54301 = pi14 ? n39762 : n24874;
  assign n54302 = pi20 ? n206 : n481;
  assign n54303 = pi19 ? n32 : n54302;
  assign n54304 = pi18 ? n32 : n54303;
  assign n54305 = pi17 ? n32 : n54304;
  assign n54306 = pi16 ? n32 : n54305;
  assign n54307 = pi15 ? n54306 : n51565;
  assign n54308 = pi14 ? n52315 : n54307;
  assign n54309 = pi13 ? n54301 : n54308;
  assign n54310 = pi12 ? n54300 : n54309;
  assign n54311 = pi11 ? n39759 : n54310;
  assign n54312 = pi15 ? n16101 : n14651;
  assign n54313 = pi19 ? n322 : ~n8286;
  assign n54314 = pi18 ? n32 : n54313;
  assign n54315 = pi17 ? n32 : n54314;
  assign n54316 = pi16 ? n32 : n54315;
  assign n54317 = pi19 ? n32 : ~n11783;
  assign n54318 = pi18 ? n32 : n54317;
  assign n54319 = pi17 ? n32 : n54318;
  assign n54320 = pi16 ? n32 : n54319;
  assign n54321 = pi15 ? n54316 : n54320;
  assign n54322 = pi14 ? n54312 : n54321;
  assign n54323 = pi19 ? n5614 : n7435;
  assign n54324 = pi18 ? n32 : n54323;
  assign n54325 = pi17 ? n32 : n54324;
  assign n54326 = pi16 ? n32 : n54325;
  assign n54327 = pi20 ? n321 : n2358;
  assign n54328 = pi19 ? n54327 : ~n1941;
  assign n54329 = pi18 ? n32 : n54328;
  assign n54330 = pi17 ? n32 : n54329;
  assign n54331 = pi16 ? n32 : n54330;
  assign n54332 = pi15 ? n54326 : n54331;
  assign n54333 = pi20 ? n428 : ~n220;
  assign n54334 = pi19 ? n32 : n54333;
  assign n54335 = pi19 ? n8622 : n349;
  assign n54336 = pi18 ? n54334 : ~n54335;
  assign n54337 = pi17 ? n32 : n54336;
  assign n54338 = pi16 ? n32 : n54337;
  assign n54339 = pi20 ? n342 : ~n915;
  assign n54340 = pi19 ? n54339 : ~n9724;
  assign n54341 = pi18 ? n54334 : ~n54340;
  assign n54342 = pi17 ? n32 : n54341;
  assign n54343 = pi16 ? n32 : n54342;
  assign n54344 = pi15 ? n54338 : n54343;
  assign n54345 = pi14 ? n54332 : n54344;
  assign n54346 = pi13 ? n54322 : n54345;
  assign n54347 = pi15 ? n26837 : n15700;
  assign n54348 = pi14 ? n54347 : n38992;
  assign n54349 = pi19 ? n32 : ~n10447;
  assign n54350 = pi18 ? n32 : n54349;
  assign n54351 = pi17 ? n32 : n54350;
  assign n54352 = pi16 ? n32 : n54351;
  assign n54353 = pi15 ? n32 : n54352;
  assign n54354 = pi19 ? n267 : n53;
  assign n54355 = pi18 ? n32 : n54354;
  assign n54356 = pi17 ? n32 : n54355;
  assign n54357 = pi16 ? n32 : n54356;
  assign n54358 = pi19 ? n267 : n358;
  assign n54359 = pi18 ? n32 : n54358;
  assign n54360 = pi17 ? n32 : n54359;
  assign n54361 = pi16 ? n32 : n54360;
  assign n54362 = pi15 ? n54357 : n54361;
  assign n54363 = pi14 ? n54353 : n54362;
  assign n54364 = pi13 ? n54348 : n54363;
  assign n54365 = pi12 ? n54346 : n54364;
  assign n54366 = pi15 ? n22087 : n14156;
  assign n54367 = pi21 ? n206 : ~n27422;
  assign n54368 = pi20 ? n32 : ~n54367;
  assign n54369 = pi19 ? n54368 : n32;
  assign n54370 = pi18 ? n32 : n54369;
  assign n54371 = pi17 ? n32 : n54370;
  assign n54372 = pi16 ? n32 : n54371;
  assign n54373 = pi15 ? n35939 : n54372;
  assign n54374 = pi14 ? n54366 : n54373;
  assign n54375 = pi20 ? n32 : ~n6651;
  assign n54376 = pi19 ? n54375 : n32;
  assign n54377 = pi18 ? n32 : n54376;
  assign n54378 = pi17 ? n32 : n54377;
  assign n54379 = pi16 ? n32 : n54378;
  assign n54380 = pi15 ? n54379 : n39835;
  assign n54381 = pi18 ? n4722 : ~n323;
  assign n54382 = pi17 ? n32 : n54381;
  assign n54383 = pi16 ? n32 : n54382;
  assign n54384 = pi15 ? n39840 : n54383;
  assign n54385 = pi14 ? n54380 : n54384;
  assign n54386 = pi13 ? n54374 : n54385;
  assign n54387 = pi15 ? n32468 : n11860;
  assign n54388 = pi18 ? n42416 : ~n20788;
  assign n54389 = pi17 ? n32 : n54388;
  assign n54390 = pi16 ? n32 : n54389;
  assign n54391 = pi15 ? n11860 : n54390;
  assign n54392 = pi14 ? n54387 : n54391;
  assign n54393 = pi18 ? n1741 : ~n418;
  assign n54394 = pi17 ? n32 : n54393;
  assign n54395 = pi16 ? n32 : n54394;
  assign n54396 = pi18 ? n222 : ~n532;
  assign n54397 = pi17 ? n32 : n54396;
  assign n54398 = pi16 ? n32 : n54397;
  assign n54399 = pi15 ? n54395 : n54398;
  assign n54400 = pi16 ? n32 : n432;
  assign n54401 = pi15 ? n54400 : n20319;
  assign n54402 = pi14 ? n54399 : n54401;
  assign n54403 = pi13 ? n54392 : n54402;
  assign n54404 = pi12 ? n54386 : n54403;
  assign n54405 = pi11 ? n54365 : n54404;
  assign n54406 = pi10 ? n54311 : n54405;
  assign n54407 = pi09 ? n32 : n54406;
  assign n54408 = pi14 ? n32 : n16913;
  assign n54409 = pi13 ? n54408 : n39858;
  assign n54410 = pi12 ? n32 : n54409;
  assign n54411 = pi14 ? n39861 : n24874;
  assign n54412 = pi19 ? n32 : ~n11986;
  assign n54413 = pi18 ? n32 : n54412;
  assign n54414 = pi17 ? n32 : n54413;
  assign n54415 = pi16 ? n32 : n54414;
  assign n54416 = pi15 ? n52315 : n54415;
  assign n54417 = pi14 ? n54416 : n51565;
  assign n54418 = pi13 ? n54411 : n54417;
  assign n54419 = pi12 ? n54300 : n54418;
  assign n54420 = pi11 ? n54410 : n54419;
  assign n54421 = pi19 ? n322 : ~n11561;
  assign n54422 = pi18 ? n32 : n54421;
  assign n54423 = pi17 ? n32 : n54422;
  assign n54424 = pi16 ? n32 : n54423;
  assign n54425 = pi15 ? n54424 : n54320;
  assign n54426 = pi14 ? n54312 : n54425;
  assign n54427 = pi19 ? n54339 : ~n26833;
  assign n54428 = pi18 ? n54334 : ~n54427;
  assign n54429 = pi17 ? n32 : n54428;
  assign n54430 = pi16 ? n32 : n54429;
  assign n54431 = pi15 ? n54338 : n54430;
  assign n54432 = pi14 ? n54332 : n54431;
  assign n54433 = pi13 ? n54426 : n54432;
  assign n54434 = pi15 ? n26837 : n16105;
  assign n54435 = pi14 ? n54434 : n38992;
  assign n54436 = pi14 ? n24327 : n14397;
  assign n54437 = pi13 ? n54435 : n54436;
  assign n54438 = pi12 ? n54433 : n54437;
  assign n54439 = pi15 ? n39487 : n54372;
  assign n54440 = pi14 ? n24555 : n54439;
  assign n54441 = pi15 ? n13948 : n39835;
  assign n54442 = pi15 ? n39594 : n54383;
  assign n54443 = pi14 ? n54441 : n54442;
  assign n54444 = pi13 ? n54440 : n54443;
  assign n54445 = pi18 ? n222 : ~n20628;
  assign n54446 = pi17 ? n32 : n54445;
  assign n54447 = pi16 ? n32 : n54446;
  assign n54448 = pi15 ? n12304 : n54447;
  assign n54449 = pi14 ? n34259 : n54448;
  assign n54450 = pi18 ? n222 : ~n2298;
  assign n54451 = pi17 ? n32 : n54450;
  assign n54452 = pi16 ? n32 : n54451;
  assign n54453 = pi15 ? n39906 : n54452;
  assign n54454 = pi14 ? n54453 : n39909;
  assign n54455 = pi13 ? n54449 : n54454;
  assign n54456 = pi12 ? n54444 : n54455;
  assign n54457 = pi11 ? n54438 : n54456;
  assign n54458 = pi10 ? n54420 : n54457;
  assign n54459 = pi09 ? n32 : n54458;
  assign n54460 = pi08 ? n54407 : n54459;
  assign n54461 = pi14 ? n16393 : n32;
  assign n54462 = pi14 ? n17278 : n16393;
  assign n54463 = pi13 ? n54461 : n54462;
  assign n54464 = pi12 ? n32 : n54463;
  assign n54465 = pi14 ? n16832 : n16850;
  assign n54466 = pi14 ? n24247 : n17039;
  assign n54467 = pi13 ? n54465 : n54466;
  assign n54468 = pi14 ? n39917 : n24874;
  assign n54469 = pi19 ? n32 : ~n21179;
  assign n54470 = pi18 ? n32 : n54469;
  assign n54471 = pi17 ? n32 : n54470;
  assign n54472 = pi16 ? n32 : n54471;
  assign n54473 = pi15 ? n24247 : n54472;
  assign n54474 = pi14 ? n54473 : n16105;
  assign n54475 = pi13 ? n54468 : n54474;
  assign n54476 = pi12 ? n54467 : n54475;
  assign n54477 = pi11 ? n54464 : n54476;
  assign n54478 = pi15 ? n16101 : n39243;
  assign n54479 = pi19 ? n322 : n19749;
  assign n54480 = pi18 ? n32 : n54479;
  assign n54481 = pi17 ? n32 : n54480;
  assign n54482 = pi16 ? n32 : n54481;
  assign n54483 = pi15 ? n54482 : n32;
  assign n54484 = pi14 ? n54478 : n54483;
  assign n54485 = pi19 ? n5371 : ~n349;
  assign n54486 = pi18 ? n32 : n54485;
  assign n54487 = pi17 ? n32 : n54486;
  assign n54488 = pi16 ? n32 : n54487;
  assign n54489 = pi15 ? n15650 : n54488;
  assign n54490 = pi17 ? n32 : n51252;
  assign n54491 = pi16 ? n32 : n54490;
  assign n54492 = pi15 ? n54491 : n12773;
  assign n54493 = pi14 ? n54489 : n54492;
  assign n54494 = pi13 ? n54484 : n54493;
  assign n54495 = pi15 ? n23484 : n22923;
  assign n54496 = pi21 ? n174 : n9326;
  assign n54497 = pi20 ? n32 : n54496;
  assign n54498 = pi19 ? n54497 : n32;
  assign n54499 = pi18 ? n32 : n54498;
  assign n54500 = pi17 ? n32 : n54499;
  assign n54501 = pi16 ? n32 : n54500;
  assign n54502 = pi15 ? n32 : n54501;
  assign n54503 = pi14 ? n54495 : n54502;
  assign n54504 = pi13 ? n49520 : n54503;
  assign n54505 = pi12 ? n54494 : n54504;
  assign n54506 = pi19 ? n1138 : n32;
  assign n54507 = pi18 ? n32 : n54506;
  assign n54508 = pi17 ? n32 : n54507;
  assign n54509 = pi16 ? n32 : n54508;
  assign n54510 = pi15 ? n54509 : n666;
  assign n54511 = pi21 ? n35 : ~n206;
  assign n54512 = pi20 ? n32 : n54511;
  assign n54513 = pi19 ? n54512 : n32;
  assign n54514 = pi18 ? n32 : n54513;
  assign n54515 = pi17 ? n32 : n54514;
  assign n54516 = pi16 ? n32 : n54515;
  assign n54517 = pi15 ? n54516 : n32;
  assign n54518 = pi14 ? n54510 : n54517;
  assign n54519 = pi19 ? n565 : n32;
  assign n54520 = pi18 ? n32 : n54519;
  assign n54521 = pi17 ? n32 : n54520;
  assign n54522 = pi16 ? n32 : n54521;
  assign n54523 = pi15 ? n54522 : n32685;
  assign n54524 = pi18 ? n268 : n13058;
  assign n54525 = pi17 ? n32 : n54524;
  assign n54526 = pi16 ? n32 : n54525;
  assign n54527 = pi18 ? n4127 : ~n605;
  assign n54528 = pi17 ? n32 : n54527;
  assign n54529 = pi16 ? n32 : n54528;
  assign n54530 = pi15 ? n54526 : n54529;
  assign n54531 = pi14 ? n54523 : n54530;
  assign n54532 = pi13 ? n54518 : n54531;
  assign n54533 = pi18 ? n1592 : ~n418;
  assign n54534 = pi17 ? n32 : n54533;
  assign n54535 = pi16 ? n32 : n54534;
  assign n54536 = pi15 ? n54535 : n20997;
  assign n54537 = pi14 ? n12538 : n54536;
  assign n54538 = pi15 ? n20072 : n39952;
  assign n54539 = pi14 ? n20543 : n54538;
  assign n54540 = pi13 ? n54537 : n54539;
  assign n54541 = pi12 ? n54532 : n54540;
  assign n54542 = pi11 ? n54505 : n54541;
  assign n54543 = pi10 ? n54477 : n54542;
  assign n54544 = pi09 ? n32 : n54543;
  assign n54545 = pi15 ? n32 : n16832;
  assign n54546 = pi14 ? n17278 : n54545;
  assign n54547 = pi13 ? n54461 : n54546;
  assign n54548 = pi12 ? n32 : n54547;
  assign n54549 = pi15 ? n26322 : n26009;
  assign n54550 = pi14 ? n54549 : n24874;
  assign n54551 = pi13 ? n54550 : n54474;
  assign n54552 = pi12 ? n54467 : n54551;
  assign n54553 = pi11 ? n54548 : n54552;
  assign n54554 = pi19 ? n15651 : n15646;
  assign n54555 = pi18 ? n32 : n54554;
  assign n54556 = pi17 ? n32 : n54555;
  assign n54557 = pi16 ? n32 : n54556;
  assign n54558 = pi19 ? n36202 : ~n349;
  assign n54559 = pi18 ? n32 : n54558;
  assign n54560 = pi17 ? n32 : n54559;
  assign n54561 = pi16 ? n32 : n54560;
  assign n54562 = pi15 ? n54557 : n54561;
  assign n54563 = pi19 ? n4491 : n349;
  assign n54564 = pi18 ? n863 : ~n54563;
  assign n54565 = pi17 ? n32 : n54564;
  assign n54566 = pi16 ? n32 : n54565;
  assign n54567 = pi18 ? n863 : ~n10486;
  assign n54568 = pi17 ? n32 : n54567;
  assign n54569 = pi16 ? n32 : n54568;
  assign n54570 = pi15 ? n54566 : n54569;
  assign n54571 = pi14 ? n54562 : n54570;
  assign n54572 = pi13 ? n54484 : n54571;
  assign n54573 = pi15 ? n32 : n15655;
  assign n54574 = pi14 ? n32 : n54573;
  assign n54575 = pi20 ? n32 : n11116;
  assign n54576 = pi19 ? n54575 : n32;
  assign n54577 = pi18 ? n32 : n54576;
  assign n54578 = pi17 ? n32 : n54577;
  assign n54579 = pi16 ? n32 : n54578;
  assign n54580 = pi15 ? n32 : n54579;
  assign n54581 = pi14 ? n54495 : n54580;
  assign n54582 = pi13 ? n54574 : n54581;
  assign n54583 = pi12 ? n54572 : n54582;
  assign n54584 = pi20 ? n32 : n12244;
  assign n54585 = pi19 ? n54584 : n32;
  assign n54586 = pi18 ? n32 : n54585;
  assign n54587 = pi17 ? n32 : n54586;
  assign n54588 = pi16 ? n32 : n54587;
  assign n54589 = pi15 ? n54588 : n32;
  assign n54590 = pi19 ? n37233 : n32;
  assign n54591 = pi18 ? n32 : n54590;
  assign n54592 = pi17 ? n32 : n54591;
  assign n54593 = pi16 ? n32 : n54592;
  assign n54594 = pi15 ? n54593 : n21319;
  assign n54595 = pi14 ? n54589 : n54594;
  assign n54596 = pi19 ? n50372 : n32;
  assign n54597 = pi18 ? n32 : n54596;
  assign n54598 = pi17 ? n32 : n54597;
  assign n54599 = pi16 ? n32 : n54598;
  assign n54600 = pi15 ? n21954 : n54599;
  assign n54601 = pi18 ? n863 : ~n605;
  assign n54602 = pi17 ? n32 : n54601;
  assign n54603 = pi16 ? n32 : n54602;
  assign n54604 = pi15 ? n13061 : n54603;
  assign n54605 = pi14 ? n54600 : n54604;
  assign n54606 = pi13 ? n54595 : n54605;
  assign n54607 = pi14 ? n54603 : n12542;
  assign n54608 = pi13 ? n54607 : n39988;
  assign n54609 = pi12 ? n54606 : n54608;
  assign n54610 = pi11 ? n54583 : n54609;
  assign n54611 = pi10 ? n54553 : n54610;
  assign n54612 = pi09 ? n32 : n54611;
  assign n54613 = pi08 ? n54544 : n54612;
  assign n54614 = pi07 ? n54460 : n54613;
  assign n54615 = pi13 ? n32 : n54546;
  assign n54616 = pi12 ? n32 : n54615;
  assign n54617 = pi14 ? n16832 : n17364;
  assign n54618 = pi19 ? n32 : n21588;
  assign n54619 = pi18 ? n32 : n54618;
  assign n54620 = pi17 ? n32 : n54619;
  assign n54621 = pi16 ? n32 : n54620;
  assign n54622 = pi19 ? n1818 : n13926;
  assign n54623 = pi18 ? n32 : n54622;
  assign n54624 = pi17 ? n32 : n54623;
  assign n54625 = pi16 ? n32 : n54624;
  assign n54626 = pi15 ? n54621 : n54625;
  assign n54627 = pi14 ? n53162 : n54626;
  assign n54628 = pi13 ? n54617 : n54627;
  assign n54629 = pi15 ? n17039 : n26009;
  assign n54630 = pi15 ? n16546 : n27528;
  assign n54631 = pi14 ? n54629 : n54630;
  assign n54632 = pi20 ? n1385 : n243;
  assign n54633 = pi19 ? n32 : ~n54632;
  assign n54634 = pi18 ? n32 : n54633;
  assign n54635 = pi17 ? n32 : n54634;
  assign n54636 = pi16 ? n32 : n54635;
  assign n54637 = pi15 ? n54636 : n24247;
  assign n54638 = pi14 ? n54637 : n36481;
  assign n54639 = pi13 ? n54631 : n54638;
  assign n54640 = pi12 ? n54628 : n54639;
  assign n54641 = pi11 ? n54616 : n54640;
  assign n54642 = pi15 ? n16452 : n25384;
  assign n54643 = pi20 ? n20944 : n32;
  assign n54644 = pi19 ? n18396 : n54643;
  assign n54645 = pi18 ? n32 : n54644;
  assign n54646 = pi17 ? n32 : n54645;
  assign n54647 = pi16 ? n32 : n54646;
  assign n54648 = pi15 ? n54647 : n15834;
  assign n54649 = pi14 ? n54642 : n54648;
  assign n54650 = pi19 ? n1757 : ~n6683;
  assign n54651 = pi18 ? n936 : n54650;
  assign n54652 = pi17 ? n32 : n54651;
  assign n54653 = pi16 ? n32 : n54652;
  assign n54654 = pi15 ? n24511 : n54653;
  assign n54655 = pi20 ? n259 : ~n32;
  assign n54656 = pi19 ? n6173 : n54655;
  assign n54657 = pi18 ? n936 : ~n54656;
  assign n54658 = pi17 ? n32 : n54657;
  assign n54659 = pi16 ? n32 : n54658;
  assign n54660 = pi18 ? n936 : n38172;
  assign n54661 = pi17 ? n32 : n54660;
  assign n54662 = pi16 ? n32 : n54661;
  assign n54663 = pi15 ? n54659 : n54662;
  assign n54664 = pi14 ? n54654 : n54663;
  assign n54665 = pi13 ? n54649 : n54664;
  assign n54666 = pi15 ? n23443 : n37801;
  assign n54667 = pi15 ? n39812 : n32;
  assign n54668 = pi14 ? n54666 : n54667;
  assign n54669 = pi15 ? n15123 : n22817;
  assign n54670 = pi14 ? n22252 : n54669;
  assign n54671 = pi13 ? n54668 : n54670;
  assign n54672 = pi12 ? n54665 : n54671;
  assign n54673 = pi15 ? n40196 : n13948;
  assign n54674 = pi14 ? n54673 : n31120;
  assign n54675 = pi15 ? n14397 : n20836;
  assign n54676 = pi20 ? n785 : ~n749;
  assign n54677 = pi19 ? n54676 : n32;
  assign n54678 = pi18 ? n32 : n54677;
  assign n54679 = pi17 ? n32 : n54678;
  assign n54680 = pi16 ? n32 : n54679;
  assign n54681 = pi20 ? n820 : ~n207;
  assign n54682 = pi19 ? n54681 : n32;
  assign n54683 = pi18 ? n32 : n54682;
  assign n54684 = pi17 ? n32 : n54683;
  assign n54685 = pi16 ? n32 : n54684;
  assign n54686 = pi15 ? n54680 : n54685;
  assign n54687 = pi14 ? n54675 : n54686;
  assign n54688 = pi13 ? n54674 : n54687;
  assign n54689 = pi19 ? n9321 : ~n32;
  assign n54690 = pi18 ? n32 : ~n54689;
  assign n54691 = pi17 ? n32 : n54690;
  assign n54692 = pi16 ? n32 : n54691;
  assign n54693 = pi18 ? n32 : ~n20680;
  assign n54694 = pi17 ? n32 : n54693;
  assign n54695 = pi16 ? n32 : n54694;
  assign n54696 = pi15 ? n54692 : n54695;
  assign n54697 = pi14 ? n54696 : n20692;
  assign n54698 = pi19 ? n10879 : n32;
  assign n54699 = pi18 ? n32 : n54698;
  assign n54700 = pi17 ? n32 : n54699;
  assign n54701 = pi16 ? n32 : n54700;
  assign n54702 = pi15 ? n54701 : n20067;
  assign n54703 = pi14 ? n54702 : n19814;
  assign n54704 = pi13 ? n54697 : n54703;
  assign n54705 = pi12 ? n54688 : n54704;
  assign n54706 = pi11 ? n54672 : n54705;
  assign n54707 = pi10 ? n54641 : n54706;
  assign n54708 = pi09 ? n17493 : n54707;
  assign n54709 = pi14 ? n25633 : n17364;
  assign n54710 = pi19 ? n1818 : n21637;
  assign n54711 = pi18 ? n32 : n54710;
  assign n54712 = pi17 ? n32 : n54711;
  assign n54713 = pi16 ? n32 : n54712;
  assign n54714 = pi15 ? n54621 : n54713;
  assign n54715 = pi14 ? n53162 : n54714;
  assign n54716 = pi13 ? n54709 : n54715;
  assign n54717 = pi15 ? n54472 : n24247;
  assign n54718 = pi14 ? n54717 : n36481;
  assign n54719 = pi13 ? n54631 : n54718;
  assign n54720 = pi12 ? n54716 : n54719;
  assign n54721 = pi11 ? n54616 : n54720;
  assign n54722 = pi15 ? n54647 : n24247;
  assign n54723 = pi14 ? n54642 : n54722;
  assign n54724 = pi20 ? n1445 : n32;
  assign n54725 = pi19 ? n37 : n54724;
  assign n54726 = pi18 ? n32 : n54725;
  assign n54727 = pi17 ? n32 : n54726;
  assign n54728 = pi16 ? n32 : n54727;
  assign n54729 = pi21 ? n242 : n309;
  assign n54730 = pi20 ? n54729 : n32;
  assign n54731 = pi19 ? n54730 : ~n6683;
  assign n54732 = pi18 ? n32 : n54731;
  assign n54733 = pi17 ? n32 : n54732;
  assign n54734 = pi16 ? n32 : n54733;
  assign n54735 = pi15 ? n54728 : n54734;
  assign n54736 = pi20 ? n371 : ~n220;
  assign n54737 = pi20 ? n15732 : ~n32;
  assign n54738 = pi19 ? n54736 : ~n54737;
  assign n54739 = pi18 ? n32 : n54738;
  assign n54740 = pi17 ? n32 : n54739;
  assign n54741 = pi16 ? n32 : n54740;
  assign n54742 = pi15 ? n54741 : n38175;
  assign n54743 = pi14 ? n54735 : n54742;
  assign n54744 = pi13 ? n54723 : n54743;
  assign n54745 = pi15 ? n37644 : n32;
  assign n54746 = pi14 ? n54666 : n54745;
  assign n54747 = pi14 ? n22818 : n22931;
  assign n54748 = pi13 ? n54746 : n54747;
  assign n54749 = pi12 ? n54744 : n54748;
  assign n54750 = pi14 ? n54673 : n32;
  assign n54751 = pi19 ? n41923 : n32;
  assign n54752 = pi18 ? n32 : n54751;
  assign n54753 = pi17 ? n32 : n54752;
  assign n54754 = pi16 ? n32 : n54753;
  assign n54755 = pi15 ? n20836 : n54754;
  assign n54756 = pi15 ? n54680 : n40074;
  assign n54757 = pi14 ? n54755 : n54756;
  assign n54758 = pi13 ? n54750 : n54757;
  assign n54759 = pi20 ? n9628 : n32;
  assign n54760 = pi19 ? n54759 : n32;
  assign n54761 = pi18 ? n32 : n54760;
  assign n54762 = pi17 ? n32 : n54761;
  assign n54763 = pi16 ? n32 : n54762;
  assign n54764 = pi15 ? n54763 : n19972;
  assign n54765 = pi14 ? n54764 : n40087;
  assign n54766 = pi13 ? n54765 : n40090;
  assign n54767 = pi12 ? n54758 : n54766;
  assign n54768 = pi11 ? n54749 : n54767;
  assign n54769 = pi10 ? n54721 : n54768;
  assign n54770 = pi09 ? n17493 : n54769;
  assign n54771 = pi08 ? n54708 : n54770;
  assign n54772 = pi15 ? n17188 : n16832;
  assign n54773 = pi14 ? n17278 : n54772;
  assign n54774 = pi13 ? n32 : n54773;
  assign n54775 = pi12 ? n32 : n54774;
  assign n54776 = pi15 ? n17363 : n17039;
  assign n54777 = pi14 ? n25633 : n54776;
  assign n54778 = pi19 ? n507 : ~n1386;
  assign n54779 = pi18 ? n32 : n54778;
  assign n54780 = pi17 ? n32 : n54779;
  assign n54781 = pi16 ? n32 : n54780;
  assign n54782 = pi15 ? n24247 : n54781;
  assign n54783 = pi14 ? n54782 : n38294;
  assign n54784 = pi13 ? n54777 : n54783;
  assign n54785 = pi15 ? n16546 : n25306;
  assign n54786 = pi14 ? n40305 : n54785;
  assign n54787 = pi19 ? n6398 : ~n589;
  assign n54788 = pi18 ? n32 : n54787;
  assign n54789 = pi17 ? n32 : n54788;
  assign n54790 = pi16 ? n32 : n54789;
  assign n54791 = pi15 ? n54472 : n54790;
  assign n54792 = pi15 ? n24247 : n27528;
  assign n54793 = pi14 ? n54791 : n54792;
  assign n54794 = pi13 ? n54786 : n54793;
  assign n54795 = pi12 ? n54784 : n54794;
  assign n54796 = pi11 ? n54775 : n54795;
  assign n54797 = pi20 ? n18256 : ~n32;
  assign n54798 = pi19 ? n32 : ~n54797;
  assign n54799 = pi18 ? n32 : n54798;
  assign n54800 = pi17 ? n32 : n54799;
  assign n54801 = pi16 ? n32 : n54800;
  assign n54802 = pi15 ? n16606 : n54801;
  assign n54803 = pi20 ? n342 : n1385;
  assign n54804 = pi19 ? n54803 : ~n349;
  assign n54805 = pi18 ? n32 : n54804;
  assign n54806 = pi17 ? n32 : n54805;
  assign n54807 = pi16 ? n32 : n54806;
  assign n54808 = pi15 ? n54807 : n32;
  assign n54809 = pi14 ? n54802 : n54808;
  assign n54810 = pi19 ? n52453 : n5635;
  assign n54811 = pi18 ? n32 : n54810;
  assign n54812 = pi17 ? n32 : n54811;
  assign n54813 = pi16 ? n32 : n54812;
  assign n54814 = pi19 ? n52453 : ~n6683;
  assign n54815 = pi18 ? n32 : n54814;
  assign n54816 = pi17 ? n32 : n54815;
  assign n54817 = pi16 ? n32 : n54816;
  assign n54818 = pi15 ? n54813 : n54817;
  assign n54819 = pi19 ? n18113 : ~n1105;
  assign n54820 = pi18 ? n32 : n54819;
  assign n54821 = pi17 ? n32 : n54820;
  assign n54822 = pi16 ? n32 : n54821;
  assign n54823 = pi15 ? n54822 : n54361;
  assign n54824 = pi14 ? n54818 : n54823;
  assign n54825 = pi13 ? n54809 : n54824;
  assign n54826 = pi19 ? n1464 : n440;
  assign n54827 = pi18 ? n32 : n54826;
  assign n54828 = pi17 ? n32 : n54827;
  assign n54829 = pi16 ? n32 : n54828;
  assign n54830 = pi15 ? n54829 : n37801;
  assign n54831 = pi15 ? n23169 : n22540;
  assign n54832 = pi14 ? n54830 : n54831;
  assign n54833 = pi15 ? n22540 : n13952;
  assign n54834 = pi14 ? n54833 : n32;
  assign n54835 = pi13 ? n54832 : n54834;
  assign n54836 = pi12 ? n54825 : n54835;
  assign n54837 = pi15 ? n20048 : n13952;
  assign n54838 = pi14 ? n34020 : n54837;
  assign n54839 = pi19 ? n51806 : n32;
  assign n54840 = pi18 ? n32 : n54839;
  assign n54841 = pi17 ? n32 : n54840;
  assign n54842 = pi16 ? n32 : n54841;
  assign n54843 = pi15 ? n13943 : n54842;
  assign n54844 = pi19 ? n53064 : n32;
  assign n54845 = pi18 ? n32 : n54844;
  assign n54846 = pi17 ? n32 : n54845;
  assign n54847 = pi16 ? n32 : n54846;
  assign n54848 = pi15 ? n13952 : n54847;
  assign n54849 = pi14 ? n54843 : n54848;
  assign n54850 = pi13 ? n54838 : n54849;
  assign n54851 = pi15 ? n156 : n20048;
  assign n54852 = pi14 ? n54851 : n40141;
  assign n54853 = pi13 ? n54852 : n40142;
  assign n54854 = pi12 ? n54850 : n54853;
  assign n54855 = pi11 ? n54836 : n54854;
  assign n54856 = pi10 ? n54796 : n54855;
  assign n54857 = pi09 ? n17493 : n54856;
  assign n54858 = pi20 ? n342 : n125;
  assign n54859 = pi19 ? n32 : n54858;
  assign n54860 = pi18 ? n32 : n54859;
  assign n54861 = pi17 ? n32 : n54860;
  assign n54862 = pi16 ? n32 : n54861;
  assign n54863 = pi15 ? n16832 : n54862;
  assign n54864 = pi14 ? n54863 : n54776;
  assign n54865 = pi19 ? n1785 : n14609;
  assign n54866 = pi18 ? n32 : n54865;
  assign n54867 = pi17 ? n32 : n54866;
  assign n54868 = pi16 ? n32 : n54867;
  assign n54869 = pi19 ? n32 : n32694;
  assign n54870 = pi18 ? n32 : n54869;
  assign n54871 = pi17 ? n32 : n54870;
  assign n54872 = pi16 ? n32 : n54871;
  assign n54873 = pi15 ? n54868 : n54872;
  assign n54874 = pi14 ? n54782 : n54873;
  assign n54875 = pi13 ? n54864 : n54874;
  assign n54876 = pi19 ? n6398 : ~n12680;
  assign n54877 = pi18 ? n32 : n54876;
  assign n54878 = pi17 ? n32 : n54877;
  assign n54879 = pi16 ? n32 : n54878;
  assign n54880 = pi15 ? n16467 : n54879;
  assign n54881 = pi14 ? n39670 : n54880;
  assign n54882 = pi19 ? n32 : ~n14287;
  assign n54883 = pi18 ? n32 : n54882;
  assign n54884 = pi17 ? n32 : n54883;
  assign n54885 = pi16 ? n32 : n54884;
  assign n54886 = pi15 ? n54885 : n24511;
  assign n54887 = pi15 ? n24247 : n15633;
  assign n54888 = pi14 ? n54886 : n54887;
  assign n54889 = pi13 ? n54881 : n54888;
  assign n54890 = pi12 ? n54875 : n54889;
  assign n54891 = pi11 ? n54775 : n54890;
  assign n54892 = pi21 ? n259 : ~n66;
  assign n54893 = pi20 ? n32 : ~n54892;
  assign n54894 = pi19 ? n54893 : n32;
  assign n54895 = pi18 ? n32 : n54894;
  assign n54896 = pi17 ? n32 : n54895;
  assign n54897 = pi16 ? n32 : n54896;
  assign n54898 = pi15 ? n54807 : n54897;
  assign n54899 = pi14 ? n54802 : n54898;
  assign n54900 = pi20 ? n151 : n17134;
  assign n54901 = pi19 ? n54900 : ~n617;
  assign n54902 = pi18 ? n32 : n54901;
  assign n54903 = pi17 ? n32 : n54902;
  assign n54904 = pi16 ? n32 : n54903;
  assign n54905 = pi20 ? n151 : ~n831;
  assign n54906 = pi19 ? n54905 : n1757;
  assign n54907 = pi18 ? n32 : n54906;
  assign n54908 = pi17 ? n32 : n54907;
  assign n54909 = pi16 ? n32 : n54908;
  assign n54910 = pi15 ? n54904 : n54909;
  assign n54911 = pi20 ? n3523 : ~n9000;
  assign n54912 = pi19 ? n54911 : n32;
  assign n54913 = pi18 ? n32 : n54912;
  assign n54914 = pi17 ? n32 : n54913;
  assign n54915 = pi16 ? n32 : n54914;
  assign n54916 = pi15 ? n54915 : n54361;
  assign n54917 = pi14 ? n54910 : n54916;
  assign n54918 = pi13 ? n54899 : n54917;
  assign n54919 = pi15 ? n23169 : n22817;
  assign n54920 = pi14 ? n54830 : n54919;
  assign n54921 = pi14 ? n22543 : n31301;
  assign n54922 = pi13 ? n54920 : n54921;
  assign n54923 = pi12 ? n54918 : n54922;
  assign n54924 = pi15 ? n671 : n14156;
  assign n54925 = pi15 ? n13684 : n21226;
  assign n54926 = pi14 ? n54924 : n54925;
  assign n54927 = pi15 ? n13952 : n20048;
  assign n54928 = pi14 ? n21407 : n54927;
  assign n54929 = pi13 ? n54926 : n54928;
  assign n54930 = pi12 ? n54929 : n32;
  assign n54931 = pi11 ? n54923 : n54930;
  assign n54932 = pi10 ? n54891 : n54931;
  assign n54933 = pi09 ? n17493 : n54932;
  assign n54934 = pi08 ? n54857 : n54933;
  assign n54935 = pi07 ? n54771 : n54934;
  assign n54936 = pi06 ? n54614 : n54935;
  assign n54937 = pi05 ? n54296 : n54936;
  assign n54938 = pi04 ? n53653 : n54937;
  assign n54939 = pi15 ? n16832 : n17188;
  assign n54940 = pi14 ? n17278 : n54939;
  assign n54941 = pi13 ? n32 : n54940;
  assign n54942 = pi12 ? n32 : n54941;
  assign n54943 = pi15 ? n16832 : n17205;
  assign n54944 = pi15 ? n16850 : n16392;
  assign n54945 = pi14 ? n54943 : n54944;
  assign n54946 = pi19 ? n142 : n17212;
  assign n54947 = pi18 ? n32 : n54946;
  assign n54948 = pi17 ? n32 : n54947;
  assign n54949 = pi16 ? n32 : n54948;
  assign n54950 = pi19 ? n142 : n5163;
  assign n54951 = pi18 ? n32 : n54950;
  assign n54952 = pi17 ? n32 : n54951;
  assign n54953 = pi16 ? n32 : n54952;
  assign n54954 = pi15 ? n54949 : n54953;
  assign n54955 = pi14 ? n17039 : n54954;
  assign n54956 = pi13 ? n54945 : n54955;
  assign n54957 = pi20 ? n86 : ~n32;
  assign n54958 = pi19 ? n2386 : ~n54957;
  assign n54959 = pi18 ? n32 : n54958;
  assign n54960 = pi17 ? n32 : n54959;
  assign n54961 = pi16 ? n32 : n54960;
  assign n54962 = pi19 ? n4126 : ~n14275;
  assign n54963 = pi18 ? n32 : n54962;
  assign n54964 = pi17 ? n32 : n54963;
  assign n54965 = pi16 ? n32 : n54964;
  assign n54966 = pi15 ? n54961 : n54965;
  assign n54967 = pi14 ? n39670 : n54966;
  assign n54968 = pi19 ? n2386 : ~n14287;
  assign n54969 = pi18 ? n32 : n54968;
  assign n54970 = pi17 ? n32 : n54969;
  assign n54971 = pi16 ? n32 : n54970;
  assign n54972 = pi15 ? n54971 : n15225;
  assign n54973 = pi14 ? n54972 : n52243;
  assign n54974 = pi13 ? n54967 : n54973;
  assign n54975 = pi12 ? n54956 : n54974;
  assign n54976 = pi11 ? n54942 : n54975;
  assign n54977 = pi15 ? n26990 : n16452;
  assign n54978 = pi19 ? n6622 : n3495;
  assign n54979 = pi18 ? n32 : n54978;
  assign n54980 = pi17 ? n32 : n54979;
  assign n54981 = pi16 ? n32 : n54980;
  assign n54982 = pi19 ? n4126 : ~n349;
  assign n54983 = pi18 ? n32 : n54982;
  assign n54984 = pi17 ? n32 : n54983;
  assign n54985 = pi16 ? n32 : n54984;
  assign n54986 = pi15 ? n54981 : n54985;
  assign n54987 = pi14 ? n54977 : n54986;
  assign n54988 = pi19 ? n4280 : n19317;
  assign n54989 = pi18 ? n32 : n54988;
  assign n54990 = pi17 ? n32 : n54989;
  assign n54991 = pi16 ? n32 : n54990;
  assign n54992 = pi20 ? n428 : n354;
  assign n54993 = pi19 ? n54992 : n32;
  assign n54994 = pi18 ? n32 : n54993;
  assign n54995 = pi17 ? n32 : n54994;
  assign n54996 = pi16 ? n32 : n54995;
  assign n54997 = pi15 ? n54991 : n54996;
  assign n54998 = pi19 ? n1348 : ~n236;
  assign n54999 = pi18 ? n32 : n54998;
  assign n55000 = pi17 ? n32 : n54999;
  assign n55001 = pi16 ? n32 : n55000;
  assign n55002 = pi15 ? n55001 : n23250;
  assign n55003 = pi14 ? n54997 : n55002;
  assign n55004 = pi13 ? n54987 : n55003;
  assign n55005 = pi15 ? n15655 : n22923;
  assign n55006 = pi14 ? n55005 : n24747;
  assign n55007 = pi19 ? n11929 : n32;
  assign n55008 = pi18 ? n32 : n55007;
  assign n55009 = pi17 ? n32 : n55008;
  assign n55010 = pi16 ? n32 : n55009;
  assign n55011 = pi20 ? n32 : ~n12882;
  assign n55012 = pi19 ? n55011 : n32;
  assign n55013 = pi18 ? n32 : n55012;
  assign n55014 = pi17 ? n32 : n55013;
  assign n55015 = pi16 ? n32 : n55014;
  assign n55016 = pi15 ? n55010 : n55015;
  assign n55017 = pi14 ? n55016 : n33991;
  assign n55018 = pi13 ? n55006 : n55017;
  assign n55019 = pi12 ? n55004 : n55018;
  assign n55020 = pi15 ? n14397 : n13948;
  assign n55021 = pi15 ? n13952 : n20660;
  assign n55022 = pi14 ? n55020 : n55021;
  assign n55023 = pi13 ? n55022 : n40247;
  assign n55024 = pi12 ? n55023 : n32;
  assign n55025 = pi11 ? n55019 : n55024;
  assign n55026 = pi10 ? n54976 : n55025;
  assign n55027 = pi09 ? n17493 : n55026;
  assign n55028 = pi15 ? n17363 : n16392;
  assign n55029 = pi14 ? n54943 : n55028;
  assign n55030 = pi20 ? n175 : ~n1475;
  assign n55031 = pi19 ? n32 : n55030;
  assign n55032 = pi18 ? n32 : n55031;
  assign n55033 = pi17 ? n32 : n55032;
  assign n55034 = pi16 ? n32 : n55033;
  assign n55035 = pi15 ? n55034 : n16352;
  assign n55036 = pi14 ? n17039 : n55035;
  assign n55037 = pi13 ? n55029 : n55036;
  assign n55038 = pi19 ? n2386 : ~n422;
  assign n55039 = pi18 ? n32 : n55038;
  assign n55040 = pi17 ? n32 : n55039;
  assign n55041 = pi16 ? n32 : n55040;
  assign n55042 = pi19 ? n18198 : ~n14275;
  assign n55043 = pi18 ? n32 : n55042;
  assign n55044 = pi17 ? n32 : n55043;
  assign n55045 = pi16 ? n32 : n55044;
  assign n55046 = pi15 ? n55041 : n55045;
  assign n55047 = pi14 ? n39670 : n55046;
  assign n55048 = pi21 ? n10182 : n206;
  assign n55049 = pi20 ? n32 : n55048;
  assign n55050 = pi19 ? n55049 : ~n14287;
  assign n55051 = pi18 ? n32 : n55050;
  assign n55052 = pi17 ? n32 : n55051;
  assign n55053 = pi16 ? n32 : n55052;
  assign n55054 = pi21 ? n54035 : n206;
  assign n55055 = pi20 ? n32 : n55054;
  assign n55056 = pi19 ? n55055 : ~n13793;
  assign n55057 = pi18 ? n32 : n55056;
  assign n55058 = pi17 ? n32 : n55057;
  assign n55059 = pi16 ? n32 : n55058;
  assign n55060 = pi15 ? n55053 : n55059;
  assign n55061 = pi21 ? n32 : n14513;
  assign n55062 = pi20 ? n55061 : ~n32;
  assign n55063 = pi19 ? n32 : ~n55062;
  assign n55064 = pi18 ? n32 : n55063;
  assign n55065 = pi17 ? n32 : n55064;
  assign n55066 = pi16 ? n32 : n55065;
  assign n55067 = pi15 ? n55066 : n15633;
  assign n55068 = pi14 ? n55060 : n55067;
  assign n55069 = pi13 ? n55047 : n55068;
  assign n55070 = pi12 ? n55037 : n55069;
  assign n55071 = pi11 ? n54942 : n55070;
  assign n55072 = pi15 ? n27410 : n16452;
  assign n55073 = pi19 ? n267 : n19317;
  assign n55074 = pi18 ? n32 : n55073;
  assign n55075 = pi17 ? n32 : n55074;
  assign n55076 = pi16 ? n32 : n55075;
  assign n55077 = pi19 ? n18198 : ~n349;
  assign n55078 = pi18 ? n32 : n55077;
  assign n55079 = pi17 ? n32 : n55078;
  assign n55080 = pi16 ? n32 : n55079;
  assign n55081 = pi15 ? n55076 : n55080;
  assign n55082 = pi14 ? n55072 : n55081;
  assign n55083 = pi19 ? n507 : n19317;
  assign n55084 = pi18 ? n32 : n55083;
  assign n55085 = pi17 ? n32 : n55084;
  assign n55086 = pi16 ? n32 : n55085;
  assign n55087 = pi15 ? n55086 : n40025;
  assign n55088 = pi19 ? n365 : ~n236;
  assign n55089 = pi18 ? n32 : n55088;
  assign n55090 = pi17 ? n32 : n55089;
  assign n55091 = pi16 ? n32 : n55090;
  assign n55092 = pi15 ? n55091 : n23250;
  assign n55093 = pi14 ? n55087 : n55092;
  assign n55094 = pi13 ? n55082 : n55093;
  assign n55095 = pi14 ? n52605 : n24747;
  assign n55096 = pi14 ? n23025 : n33991;
  assign n55097 = pi13 ? n55095 : n55096;
  assign n55098 = pi12 ? n55094 : n55097;
  assign n55099 = pi15 ? n14397 : n20660;
  assign n55100 = pi14 ? n55099 : n40292;
  assign n55101 = pi13 ? n55100 : n32;
  assign n55102 = pi12 ? n55101 : n32;
  assign n55103 = pi11 ? n55098 : n55102;
  assign n55104 = pi10 ? n55071 : n55103;
  assign n55105 = pi09 ? n17493 : n55104;
  assign n55106 = pi08 ? n55027 : n55105;
  assign n55107 = pi15 ? n17216 : n16352;
  assign n55108 = pi14 ? n16392 : n55107;
  assign n55109 = pi13 ? n55029 : n55108;
  assign n55110 = pi19 ? n507 : ~n14275;
  assign n55111 = pi18 ? n32 : n55110;
  assign n55112 = pi17 ? n32 : n55111;
  assign n55113 = pi16 ? n32 : n55112;
  assign n55114 = pi15 ? n15230 : n55113;
  assign n55115 = pi14 ? n16467 : n55114;
  assign n55116 = pi19 ? n507 : ~n13793;
  assign n55117 = pi18 ? n32 : n55116;
  assign n55118 = pi17 ? n32 : n55117;
  assign n55119 = pi16 ? n32 : n55118;
  assign n55120 = pi15 ? n36100 : n55119;
  assign n55121 = pi21 ? n32 : ~n13784;
  assign n55122 = pi20 ? n55121 : ~n32;
  assign n55123 = pi19 ? n40320 : ~n55122;
  assign n55124 = pi18 ? n32 : n55123;
  assign n55125 = pi17 ? n32 : n55124;
  assign n55126 = pi16 ? n32 : n55125;
  assign n55127 = pi14 ? n55120 : n55126;
  assign n55128 = pi13 ? n55115 : n55127;
  assign n55129 = pi12 ? n55109 : n55128;
  assign n55130 = pi11 ? n54942 : n55129;
  assign n55131 = pi19 ? n40320 : n27066;
  assign n55132 = pi18 ? n32 : n55131;
  assign n55133 = pi17 ? n32 : n55132;
  assign n55134 = pi16 ? n32 : n55133;
  assign n55135 = pi19 ? n662 : n247;
  assign n55136 = pi18 ? n32 : n55135;
  assign n55137 = pi17 ? n32 : n55136;
  assign n55138 = pi16 ? n32 : n55137;
  assign n55139 = pi15 ? n55134 : n55138;
  assign n55140 = pi19 ? n41320 : n19317;
  assign n55141 = pi18 ? n32 : n55140;
  assign n55142 = pi17 ? n32 : n55141;
  assign n55143 = pi16 ? n32 : n55142;
  assign n55144 = pi20 ? n32 : n16008;
  assign n55145 = pi19 ? n55144 : ~n589;
  assign n55146 = pi18 ? n32 : n55145;
  assign n55147 = pi17 ? n32 : n55146;
  assign n55148 = pi16 ? n32 : n55147;
  assign n55149 = pi15 ? n55143 : n55148;
  assign n55150 = pi14 ? n55139 : n55149;
  assign n55151 = pi19 ? n2386 : n32;
  assign n55152 = pi18 ? n32 : n55151;
  assign n55153 = pi17 ? n32 : n55152;
  assign n55154 = pi16 ? n32 : n55153;
  assign n55155 = pi15 ? n22817 : n55154;
  assign n55156 = pi19 ? n4518 : ~n813;
  assign n55157 = pi18 ? n32 : n55156;
  assign n55158 = pi17 ? n32 : n55157;
  assign n55159 = pi16 ? n32 : n55158;
  assign n55160 = pi15 ? n55159 : n23484;
  assign n55161 = pi14 ? n55155 : n55160;
  assign n55162 = pi13 ? n55150 : n55161;
  assign n55163 = pi19 ? n18330 : ~n617;
  assign n55164 = pi18 ? n32 : n55163;
  assign n55165 = pi17 ? n32 : n55164;
  assign n55166 = pi16 ? n32 : n55165;
  assign n55167 = pi15 ? n21928 : n55166;
  assign n55168 = pi19 ? n2201 : ~n617;
  assign n55169 = pi18 ? n32 : n55168;
  assign n55170 = pi17 ? n32 : n55169;
  assign n55171 = pi16 ? n32 : n55170;
  assign n55172 = pi19 ? n786 : ~n617;
  assign n55173 = pi18 ? n32 : n55172;
  assign n55174 = pi17 ? n32 : n55173;
  assign n55175 = pi16 ? n32 : n55174;
  assign n55176 = pi15 ? n55171 : n55175;
  assign n55177 = pi14 ? n55167 : n55176;
  assign n55178 = pi15 ? n55154 : n15123;
  assign n55179 = pi14 ? n55178 : n32;
  assign n55180 = pi13 ? n55177 : n55179;
  assign n55181 = pi12 ? n55162 : n55180;
  assign n55182 = pi11 ? n55181 : n40356;
  assign n55183 = pi10 ? n55130 : n55182;
  assign n55184 = pi09 ? n17493 : n55183;
  assign n55185 = pi19 ? n472 : n5163;
  assign n55186 = pi18 ? n32 : n55185;
  assign n55187 = pi17 ? n32 : n55186;
  assign n55188 = pi16 ? n32 : n55187;
  assign n55189 = pi15 ? n17216 : n55188;
  assign n55190 = pi14 ? n16392 : n55189;
  assign n55191 = pi13 ? n55029 : n55190;
  assign n55192 = pi14 ? n16546 : n55114;
  assign n55193 = pi15 ? n55119 : n15225;
  assign n55194 = pi19 ? n32 : ~n55122;
  assign n55195 = pi18 ? n32 : n55194;
  assign n55196 = pi17 ? n32 : n55195;
  assign n55197 = pi16 ? n32 : n55196;
  assign n55198 = pi15 ? n55197 : n15633;
  assign n55199 = pi14 ? n55193 : n55198;
  assign n55200 = pi13 ? n55192 : n55199;
  assign n55201 = pi12 ? n55191 : n55200;
  assign n55202 = pi11 ? n54942 : n55201;
  assign n55203 = pi21 ? n1939 : n173;
  assign n55204 = pi20 ? n32 : n55203;
  assign n55205 = pi19 ? n55204 : n19317;
  assign n55206 = pi18 ? n32 : n55205;
  assign n55207 = pi17 ? n32 : n55206;
  assign n55208 = pi16 ? n32 : n55207;
  assign n55209 = pi19 ? n1969 : ~n589;
  assign n55210 = pi18 ? n32 : n55209;
  assign n55211 = pi17 ? n32 : n55210;
  assign n55212 = pi16 ? n32 : n55211;
  assign n55213 = pi15 ? n55208 : n55212;
  assign n55214 = pi14 ? n16452 : n55213;
  assign n55215 = pi21 ? n14399 : n10445;
  assign n55216 = pi20 ? n32 : n55215;
  assign n55217 = pi19 ? n55216 : n32;
  assign n55218 = pi18 ? n32 : n55217;
  assign n55219 = pi17 ? n32 : n55218;
  assign n55220 = pi16 ? n32 : n55219;
  assign n55221 = pi19 ? n30521 : n32;
  assign n55222 = pi18 ? n32 : n55221;
  assign n55223 = pi17 ? n32 : n55222;
  assign n55224 = pi16 ? n32 : n55223;
  assign n55225 = pi15 ? n55220 : n55224;
  assign n55226 = pi14 ? n55225 : n55160;
  assign n55227 = pi13 ? n55214 : n55226;
  assign n55228 = pi15 ? n21928 : n23340;
  assign n55229 = pi20 ? n32 : n19604;
  assign n55230 = pi19 ? n55229 : ~n617;
  assign n55231 = pi18 ? n32 : n55230;
  assign n55232 = pi17 ? n32 : n55231;
  assign n55233 = pi16 ? n32 : n55232;
  assign n55234 = pi19 ? n40454 : ~n617;
  assign n55235 = pi18 ? n32 : n55234;
  assign n55236 = pi17 ? n32 : n55235;
  assign n55237 = pi16 ? n32 : n55236;
  assign n55238 = pi15 ? n55233 : n55237;
  assign n55239 = pi14 ? n55228 : n55238;
  assign n55240 = pi19 ? n53174 : n32;
  assign n55241 = pi18 ? n32 : n55240;
  assign n55242 = pi17 ? n32 : n55241;
  assign n55243 = pi16 ? n32 : n55242;
  assign n55244 = pi15 ? n55243 : n15123;
  assign n55245 = pi14 ? n55244 : n648;
  assign n55246 = pi13 ? n55239 : n55245;
  assign n55247 = pi12 ? n55227 : n55246;
  assign n55248 = pi11 ? n55247 : n40402;
  assign n55249 = pi10 ? n55202 : n55248;
  assign n55250 = pi09 ? n17493 : n55249;
  assign n55251 = pi08 ? n55184 : n55250;
  assign n55252 = pi07 ? n55106 : n55251;
  assign n55253 = pi14 ? n40412 : n54939;
  assign n55254 = pi13 ? n32 : n55253;
  assign n55255 = pi12 ? n32 : n55254;
  assign n55256 = pi15 ? n16832 : n40660;
  assign n55257 = pi15 ? n54862 : n32;
  assign n55258 = pi14 ? n55256 : n55257;
  assign n55259 = pi18 ? n32 : n24054;
  assign n55260 = pi17 ? n32 : n55259;
  assign n55261 = pi16 ? n32 : n55260;
  assign n55262 = pi15 ? n23484 : n55261;
  assign n55263 = pi20 ? n321 : ~n7487;
  assign n55264 = pi19 ? n32 : ~n55263;
  assign n55265 = pi18 ? n32 : n55264;
  assign n55266 = pi17 ? n32 : n55265;
  assign n55267 = pi16 ? n32 : n55266;
  assign n55268 = pi20 ? n266 : ~n274;
  assign n55269 = pi19 ? n507 : ~n55268;
  assign n55270 = pi18 ? n32 : n55269;
  assign n55271 = pi17 ? n32 : n55270;
  assign n55272 = pi16 ? n32 : n55271;
  assign n55273 = pi15 ? n55267 : n55272;
  assign n55274 = pi14 ? n55262 : n55273;
  assign n55275 = pi13 ? n55258 : n55274;
  assign n55276 = pi20 ? n1319 : n243;
  assign n55277 = pi19 ? n519 : ~n55276;
  assign n55278 = pi18 ? n32 : n55277;
  assign n55279 = pi17 ? n32 : n55278;
  assign n55280 = pi16 ? n32 : n55279;
  assign n55281 = pi15 ? n24700 : n55280;
  assign n55282 = pi14 ? n15847 : n55281;
  assign n55283 = pi19 ? n519 : ~n6042;
  assign n55284 = pi18 ? n32 : n55283;
  assign n55285 = pi17 ? n32 : n55284;
  assign n55286 = pi16 ? n32 : n55285;
  assign n55287 = pi15 ? n15080 : n55286;
  assign n55288 = pi15 ? n37998 : n24874;
  assign n55289 = pi14 ? n55287 : n55288;
  assign n55290 = pi13 ? n55282 : n55289;
  assign n55291 = pi12 ? n55275 : n55290;
  assign n55292 = pi11 ? n55255 : n55291;
  assign n55293 = pi18 ? n32 : n21576;
  assign n55294 = pi17 ? n32 : n55293;
  assign n55295 = pi16 ? n32 : n55294;
  assign n55296 = pi15 ? n55295 : n50949;
  assign n55297 = pi18 ? n32 : n24306;
  assign n55298 = pi17 ? n32 : n55297;
  assign n55299 = pi16 ? n32 : n55298;
  assign n55300 = pi15 ? n26663 : n55299;
  assign n55301 = pi14 ? n55296 : n55300;
  assign n55302 = pi21 ? n32 : ~n9485;
  assign n55303 = pi20 ? n32 : n55302;
  assign n55304 = pi19 ? n55303 : ~n349;
  assign n55305 = pi18 ? n32 : n55304;
  assign n55306 = pi17 ? n32 : n55305;
  assign n55307 = pi16 ? n32 : n55306;
  assign n55308 = pi15 ? n55307 : n23443;
  assign n55309 = pi15 ? n25598 : n14790;
  assign n55310 = pi14 ? n55308 : n55309;
  assign n55311 = pi13 ? n55301 : n55310;
  assign n55312 = pi15 ? n27317 : n32;
  assign n55313 = pi14 ? n14975 : n55312;
  assign n55314 = pi13 ? n55313 : n40463;
  assign n55315 = pi12 ? n55311 : n55314;
  assign n55316 = pi11 ? n55315 : n32;
  assign n55317 = pi10 ? n55292 : n55316;
  assign n55318 = pi09 ? n17493 : n55317;
  assign n55319 = pi14 ? n17279 : n54939;
  assign n55320 = pi13 ? n32 : n55319;
  assign n55321 = pi12 ? n32 : n55320;
  assign n55322 = pi14 ? n55256 : n40562;
  assign n55323 = pi20 ? n1331 : ~n274;
  assign n55324 = pi19 ? n507 : ~n55323;
  assign n55325 = pi18 ? n32 : n55324;
  assign n55326 = pi17 ? n32 : n55325;
  assign n55327 = pi16 ? n32 : n55326;
  assign n55328 = pi15 ? n55267 : n55327;
  assign n55329 = pi14 ? n55262 : n55328;
  assign n55330 = pi13 ? n55322 : n55329;
  assign n55331 = pi20 ? n518 : n243;
  assign n55332 = pi19 ? n1840 : ~n55331;
  assign n55333 = pi18 ? n32 : n55332;
  assign n55334 = pi17 ? n32 : n55333;
  assign n55335 = pi16 ? n32 : n55334;
  assign n55336 = pi15 ? n24700 : n55335;
  assign n55337 = pi14 ? n15847 : n55336;
  assign n55338 = pi13 ? n55337 : n55289;
  assign n55339 = pi12 ? n55330 : n55338;
  assign n55340 = pi11 ? n55321 : n55339;
  assign n55341 = pi19 ? n519 : n247;
  assign n55342 = pi18 ? n32 : n55341;
  assign n55343 = pi17 ? n32 : n55342;
  assign n55344 = pi16 ? n32 : n55343;
  assign n55345 = pi15 ? n55295 : n55344;
  assign n55346 = pi19 ? n6398 : n1757;
  assign n55347 = pi18 ? n32 : n55346;
  assign n55348 = pi17 ? n32 : n55347;
  assign n55349 = pi16 ? n32 : n55348;
  assign n55350 = pi15 ? n26663 : n55349;
  assign n55351 = pi14 ? n55345 : n55350;
  assign n55352 = pi15 ? n40173 : n26663;
  assign n55353 = pi19 ? n1840 : ~n813;
  assign n55354 = pi18 ? n32 : n55353;
  assign n55355 = pi17 ? n32 : n55354;
  assign n55356 = pi16 ? n32 : n55355;
  assign n55357 = pi15 ? n55356 : n21928;
  assign n55358 = pi14 ? n55352 : n55357;
  assign n55359 = pi13 ? n55351 : n55358;
  assign n55360 = pi19 ? n15096 : n32;
  assign n55361 = pi18 ? n32 : n55360;
  assign n55362 = pi17 ? n32 : n55361;
  assign n55363 = pi16 ? n32 : n55362;
  assign n55364 = pi15 ? n55363 : n32;
  assign n55365 = pi15 ? n15119 : n15123;
  assign n55366 = pi14 ? n55364 : n55365;
  assign n55367 = pi13 ? n55366 : n32;
  assign n55368 = pi12 ? n55359 : n55367;
  assign n55369 = pi11 ? n55368 : n32;
  assign n55370 = pi10 ? n55340 : n55369;
  assign n55371 = pi09 ? n17493 : n55370;
  assign n55372 = pi08 ? n55318 : n55371;
  assign n55373 = pi14 ? n17279 : n40562;
  assign n55374 = pi13 ? n32 : n55373;
  assign n55375 = pi12 ? n32 : n55374;
  assign n55376 = pi15 ? n16392 : n40660;
  assign n55377 = pi14 ? n55376 : n25818;
  assign n55378 = pi19 ? n594 : ~n6298;
  assign n55379 = pi18 ? n32 : n55378;
  assign n55380 = pi17 ? n32 : n55379;
  assign n55381 = pi16 ? n32 : n55380;
  assign n55382 = pi15 ? n25888 : n55381;
  assign n55383 = pi15 ? n24247 : n14985;
  assign n55384 = pi14 ? n55382 : n55383;
  assign n55385 = pi13 ? n55377 : n55384;
  assign n55386 = pi14 ? n15847 : n40233;
  assign n55387 = pi19 ? n472 : ~n349;
  assign n55388 = pi18 ? n32 : n55387;
  assign n55389 = pi17 ? n32 : n55388;
  assign n55390 = pi16 ? n32 : n55389;
  assign n55391 = pi19 ? n472 : ~n4406;
  assign n55392 = pi18 ? n32 : n55391;
  assign n55393 = pi17 ? n32 : n55392;
  assign n55394 = pi16 ? n32 : n55393;
  assign n55395 = pi15 ? n55394 : n50949;
  assign n55396 = pi14 ? n55390 : n55395;
  assign n55397 = pi13 ? n55386 : n55396;
  assign n55398 = pi12 ? n55385 : n55397;
  assign n55399 = pi11 ? n55375 : n55398;
  assign n55400 = pi19 ? n507 : n3495;
  assign n55401 = pi18 ? n32 : n55400;
  assign n55402 = pi17 ? n32 : n55401;
  assign n55403 = pi16 ? n32 : n55402;
  assign n55404 = pi15 ? n37779 : n55403;
  assign n55405 = pi15 ? n32 : n15834;
  assign n55406 = pi14 ? n55404 : n55405;
  assign n55407 = pi19 ? n1785 : n1885;
  assign n55408 = pi18 ? n32 : n55407;
  assign n55409 = pi17 ? n32 : n55408;
  assign n55410 = pi16 ? n32 : n55409;
  assign n55411 = pi15 ? n55410 : n15263;
  assign n55412 = pi14 ? n55411 : n15127;
  assign n55413 = pi13 ? n55406 : n55412;
  assign n55414 = pi14 ? n22540 : n15267;
  assign n55415 = pi13 ? n55414 : n32;
  assign n55416 = pi12 ? n55413 : n55415;
  assign n55417 = pi11 ? n55416 : n32;
  assign n55418 = pi10 ? n55399 : n55417;
  assign n55419 = pi09 ? n17493 : n55418;
  assign n55420 = pi19 ? n2141 : ~n236;
  assign n55421 = pi18 ? n32 : n55420;
  assign n55422 = pi17 ? n32 : n55421;
  assign n55423 = pi16 ? n32 : n55422;
  assign n55424 = pi20 ? n7839 : ~n32;
  assign n55425 = pi19 ? n2141 : ~n55424;
  assign n55426 = pi18 ? n32 : n55425;
  assign n55427 = pi17 ? n32 : n55426;
  assign n55428 = pi16 ? n32 : n55427;
  assign n55429 = pi15 ? n55423 : n55428;
  assign n55430 = pi19 ? n32 : ~n3775;
  assign n55431 = pi18 ? n32 : n55430;
  assign n55432 = pi17 ? n32 : n55431;
  assign n55433 = pi16 ? n32 : n55432;
  assign n55434 = pi15 ? n24247 : n55433;
  assign n55435 = pi14 ? n55429 : n55434;
  assign n55436 = pi13 ? n55377 : n55435;
  assign n55437 = pi19 ? n594 : n247;
  assign n55438 = pi18 ? n32 : n55437;
  assign n55439 = pi17 ? n32 : n55438;
  assign n55440 = pi16 ? n32 : n55439;
  assign n55441 = pi15 ? n55295 : n55440;
  assign n55442 = pi14 ? n24247 : n55441;
  assign n55443 = pi13 ? n55386 : n55442;
  assign n55444 = pi12 ? n55436 : n55443;
  assign n55445 = pi11 ? n55375 : n55444;
  assign n55446 = pi19 ? n2141 : ~n4406;
  assign n55447 = pi18 ? n32 : n55446;
  assign n55448 = pi17 ? n32 : n55447;
  assign n55449 = pi16 ? n32 : n55448;
  assign n55450 = pi19 ? n2141 : n3495;
  assign n55451 = pi18 ? n32 : n55450;
  assign n55452 = pi17 ? n32 : n55451;
  assign n55453 = pi16 ? n32 : n55452;
  assign n55454 = pi15 ? n55449 : n55453;
  assign n55455 = pi15 ? n15263 : n15834;
  assign n55456 = pi14 ? n55454 : n55455;
  assign n55457 = pi15 ? n15834 : n32;
  assign n55458 = pi14 ? n55457 : n32;
  assign n55459 = pi13 ? n55456 : n55458;
  assign n55460 = pi12 ? n55459 : n32;
  assign n55461 = pi11 ? n55460 : n32;
  assign n55462 = pi10 ? n55445 : n55461;
  assign n55463 = pi09 ? n17493 : n55462;
  assign n55464 = pi08 ? n55419 : n55463;
  assign n55465 = pi07 ? n55372 : n55464;
  assign n55466 = pi06 ? n55252 : n55465;
  assign n55467 = pi15 ? n32 : n15927;
  assign n55468 = pi14 ? n17279 : n55467;
  assign n55469 = pi13 ? n32 : n55468;
  assign n55470 = pi12 ? n32 : n55469;
  assign n55471 = pi19 ? n32 : n23233;
  assign n55472 = pi18 ? n32 : n55471;
  assign n55473 = pi17 ? n32 : n55472;
  assign n55474 = pi16 ? n32 : n55473;
  assign n55475 = pi15 ? n16298 : n55474;
  assign n55476 = pi14 ? n15847 : n55475;
  assign n55477 = pi20 ? n357 : n6229;
  assign n55478 = pi19 ? n32 : n55477;
  assign n55479 = pi18 ? n32 : n55478;
  assign n55480 = pi17 ? n32 : n55479;
  assign n55481 = pi16 ? n32 : n55480;
  assign n55482 = pi15 ? n23250 : n55481;
  assign n55483 = pi19 ? n594 : n4342;
  assign n55484 = pi18 ? n32 : n55483;
  assign n55485 = pi17 ? n32 : n55484;
  assign n55486 = pi16 ? n32 : n55485;
  assign n55487 = pi15 ? n16392 : n55486;
  assign n55488 = pi14 ? n55482 : n55487;
  assign n55489 = pi13 ? n55476 : n55488;
  assign n55490 = pi15 ? n55486 : n16452;
  assign n55491 = pi19 ? n594 : ~n4406;
  assign n55492 = pi18 ? n32 : n55491;
  assign n55493 = pi17 ? n32 : n55492;
  assign n55494 = pi16 ? n32 : n55493;
  assign n55495 = pi15 ? n55494 : n15362;
  assign n55496 = pi14 ? n55490 : n55495;
  assign n55497 = pi15 ? n15362 : n15637;
  assign n55498 = pi19 ? n1574 : n247;
  assign n55499 = pi18 ? n32 : n55498;
  assign n55500 = pi17 ? n32 : n55499;
  assign n55501 = pi16 ? n32 : n55500;
  assign n55502 = pi15 ? n16606 : n55501;
  assign n55503 = pi14 ? n55497 : n55502;
  assign n55504 = pi13 ? n55496 : n55503;
  assign n55505 = pi12 ? n55489 : n55504;
  assign n55506 = pi11 ? n55470 : n55505;
  assign n55507 = pi19 ? n1574 : ~n589;
  assign n55508 = pi18 ? n32 : n55507;
  assign n55509 = pi17 ? n32 : n55508;
  assign n55510 = pi16 ? n32 : n55509;
  assign n55511 = pi19 ? n1574 : n9724;
  assign n55512 = pi18 ? n32 : n55511;
  assign n55513 = pi17 ? n32 : n55512;
  assign n55514 = pi16 ? n32 : n55513;
  assign n55515 = pi15 ? n55510 : n55514;
  assign n55516 = pi15 ? n32 : n22733;
  assign n55517 = pi14 ? n55515 : n55516;
  assign n55518 = pi15 ? n22733 : n22923;
  assign n55519 = pi14 ? n55518 : n22923;
  assign n55520 = pi13 ? n55517 : n55519;
  assign n55521 = pi12 ? n55520 : n32;
  assign n55522 = pi11 ? n55521 : n32;
  assign n55523 = pi10 ? n55506 : n55522;
  assign n55524 = pi09 ? n17493 : n55523;
  assign n55525 = pi15 ? n16485 : n15847;
  assign n55526 = pi20 ? n7839 : ~n141;
  assign n55527 = pi19 ? n32 : n55526;
  assign n55528 = pi18 ? n32 : n55527;
  assign n55529 = pi17 ? n32 : n55528;
  assign n55530 = pi16 ? n32 : n55529;
  assign n55531 = pi15 ? n55530 : n55474;
  assign n55532 = pi14 ? n55525 : n55531;
  assign n55533 = pi19 ? n32 : n49477;
  assign n55534 = pi18 ? n32 : n55533;
  assign n55535 = pi17 ? n32 : n55534;
  assign n55536 = pi16 ? n32 : n55535;
  assign n55537 = pi15 ? n55536 : n15847;
  assign n55538 = pi14 ? n23250 : n55537;
  assign n55539 = pi13 ? n55532 : n55538;
  assign n55540 = pi15 ? n55295 : n15507;
  assign n55541 = pi14 ? n39042 : n55540;
  assign n55542 = pi15 ? n15507 : n15501;
  assign n55543 = pi14 ? n55542 : n16452;
  assign n55544 = pi13 ? n55541 : n55543;
  assign n55545 = pi12 ? n55539 : n55544;
  assign n55546 = pi11 ? n55470 : n55545;
  assign n55547 = pi14 ? n24719 : n32;
  assign n55548 = pi15 ? n32 : n24274;
  assign n55549 = pi14 ? n55548 : n40595;
  assign n55550 = pi13 ? n55547 : n55549;
  assign n55551 = pi12 ? n55550 : n32;
  assign n55552 = pi11 ? n55551 : n32;
  assign n55553 = pi10 ? n55546 : n55552;
  assign n55554 = pi09 ? n17493 : n55553;
  assign n55555 = pi08 ? n55524 : n55554;
  assign n55556 = pi15 ? n32 : n16485;
  assign n55557 = pi14 ? n17279 : n55556;
  assign n55558 = pi13 ? n32 : n55557;
  assign n55559 = pi12 ? n32 : n55558;
  assign n55560 = pi21 ? n124 : ~n206;
  assign n55561 = pi20 ? n55560 : ~n141;
  assign n55562 = pi19 ? n32 : n55561;
  assign n55563 = pi18 ? n32 : n55562;
  assign n55564 = pi17 ? n32 : n55563;
  assign n55565 = pi16 ? n32 : n55564;
  assign n55566 = pi15 ? n37772 : n55565;
  assign n55567 = pi14 ? n55525 : n55566;
  assign n55568 = pi19 ? n32 : n12854;
  assign n55569 = pi18 ? n32 : n55568;
  assign n55570 = pi17 ? n32 : n55569;
  assign n55571 = pi16 ? n32 : n55570;
  assign n55572 = pi15 ? n15847 : n55571;
  assign n55573 = pi14 ? n23623 : n55572;
  assign n55574 = pi13 ? n55567 : n55573;
  assign n55575 = pi19 ? n32 : n44487;
  assign n55576 = pi18 ? n32 : n55575;
  assign n55577 = pi17 ? n32 : n55576;
  assign n55578 = pi16 ? n32 : n55577;
  assign n55579 = pi21 ? n10445 : ~n206;
  assign n55580 = pi20 ? n55579 : n32;
  assign n55581 = pi19 ? n32 : n55580;
  assign n55582 = pi18 ? n32 : n55581;
  assign n55583 = pi17 ? n32 : n55582;
  assign n55584 = pi16 ? n32 : n55583;
  assign n55585 = pi15 ? n55578 : n55584;
  assign n55586 = pi14 ? n55585 : n15834;
  assign n55587 = pi21 ? n51 : n174;
  assign n55588 = pi20 ? n55587 : n32;
  assign n55589 = pi19 ? n32 : n55588;
  assign n55590 = pi18 ? n32 : n55589;
  assign n55591 = pi17 ? n32 : n55590;
  assign n55592 = pi16 ? n32 : n55591;
  assign n55593 = pi15 ? n55592 : n16452;
  assign n55594 = pi21 ? n1009 : ~n206;
  assign n55595 = pi20 ? n55594 : n32;
  assign n55596 = pi19 ? n32 : n55595;
  assign n55597 = pi18 ? n32 : n55596;
  assign n55598 = pi17 ? n32 : n55597;
  assign n55599 = pi16 ? n32 : n55598;
  assign n55600 = pi15 ? n55599 : n24274;
  assign n55601 = pi14 ? n55593 : n55600;
  assign n55602 = pi13 ? n55586 : n55601;
  assign n55603 = pi12 ? n55574 : n55602;
  assign n55604 = pi11 ? n55559 : n55603;
  assign n55605 = pi21 ? n8275 : n32;
  assign n55606 = pi20 ? n55605 : n32;
  assign n55607 = pi19 ? n32 : n55606;
  assign n55608 = pi18 ? n32 : n55607;
  assign n55609 = pi17 ? n32 : n55608;
  assign n55610 = pi16 ? n32 : n55609;
  assign n55611 = pi15 ? n55610 : n15834;
  assign n55612 = pi14 ? n55611 : n16109;
  assign n55613 = pi13 ? n55612 : n32;
  assign n55614 = pi12 ? n55613 : n32;
  assign n55615 = pi11 ? n55614 : n32;
  assign n55616 = pi10 ? n55604 : n55615;
  assign n55617 = pi09 ? n17493 : n55616;
  assign n55618 = pi15 ? n25708 : n15847;
  assign n55619 = pi14 ? n55618 : n37772;
  assign n55620 = pi13 ? n55619 : n55573;
  assign n55621 = pi19 ? n32 : n9644;
  assign n55622 = pi18 ? n32 : n55621;
  assign n55623 = pi17 ? n32 : n55622;
  assign n55624 = pi16 ? n32 : n55623;
  assign n55625 = pi15 ? n55578 : n55624;
  assign n55626 = pi14 ? n55625 : n15834;
  assign n55627 = pi21 ? n16649 : n174;
  assign n55628 = pi20 ? n55627 : n32;
  assign n55629 = pi19 ? n32 : n55628;
  assign n55630 = pi18 ? n32 : n55629;
  assign n55631 = pi17 ? n32 : n55630;
  assign n55632 = pi16 ? n32 : n55631;
  assign n55633 = pi20 ? n54511 : n32;
  assign n55634 = pi19 ? n32 : n55633;
  assign n55635 = pi18 ? n32 : n55634;
  assign n55636 = pi17 ? n32 : n55635;
  assign n55637 = pi16 ? n32 : n55636;
  assign n55638 = pi15 ? n55632 : n55637;
  assign n55639 = pi21 ? n13784 : ~n206;
  assign n55640 = pi20 ? n55639 : n32;
  assign n55641 = pi19 ? n32 : n55640;
  assign n55642 = pi18 ? n32 : n55641;
  assign n55643 = pi17 ? n32 : n55642;
  assign n55644 = pi16 ? n32 : n55643;
  assign n55645 = pi15 ? n55644 : n32;
  assign n55646 = pi14 ? n55638 : n55645;
  assign n55647 = pi13 ? n55626 : n55646;
  assign n55648 = pi12 ? n55620 : n55647;
  assign n55649 = pi11 ? n55559 : n55648;
  assign n55650 = pi15 ? n16105 : n23741;
  assign n55651 = pi14 ? n24578 : n55650;
  assign n55652 = pi13 ? n55651 : n23327;
  assign n55653 = pi12 ? n55652 : n32;
  assign n55654 = pi11 ? n55653 : n32;
  assign n55655 = pi10 ? n55649 : n55654;
  assign n55656 = pi09 ? n17493 : n55655;
  assign n55657 = pi08 ? n55617 : n55656;
  assign n55658 = pi07 ? n55555 : n55657;
  assign n55659 = pi20 ? n501 : ~n141;
  assign n55660 = pi19 ? n32 : n55659;
  assign n55661 = pi18 ? n32 : n55660;
  assign n55662 = pi17 ? n32 : n55661;
  assign n55663 = pi16 ? n32 : n55662;
  assign n55664 = pi15 ? n15847 : n55663;
  assign n55665 = pi14 ? n17279 : n55664;
  assign n55666 = pi13 ? n32 : n55665;
  assign n55667 = pi12 ? n32 : n55666;
  assign n55668 = pi20 ? n653 : ~n321;
  assign n55669 = pi19 ? n32 : n55668;
  assign n55670 = pi18 ? n32 : n55669;
  assign n55671 = pi17 ? n32 : n55670;
  assign n55672 = pi16 ? n32 : n55671;
  assign n55673 = pi15 ? n55672 : n17188;
  assign n55674 = pi14 ? n55673 : n17188;
  assign n55675 = pi15 ? n16352 : n15695;
  assign n55676 = pi15 ? n15847 : n15695;
  assign n55677 = pi14 ? n55675 : n55676;
  assign n55678 = pi13 ? n55674 : n55677;
  assign n55679 = pi15 ? n15531 : n16319;
  assign n55680 = pi15 ? n16101 : n25211;
  assign n55681 = pi14 ? n55679 : n55680;
  assign n55682 = pi21 ? n16649 : ~n206;
  assign n55683 = pi20 ? n55682 : n32;
  assign n55684 = pi19 ? n32 : n55683;
  assign n55685 = pi18 ? n32 : n55684;
  assign n55686 = pi17 ? n32 : n55685;
  assign n55687 = pi16 ? n32 : n55686;
  assign n55688 = pi15 ? n55687 : n55637;
  assign n55689 = pi21 ? n48999 : ~n206;
  assign n55690 = pi20 ? n55689 : n32;
  assign n55691 = pi19 ? n32 : n55690;
  assign n55692 = pi18 ? n32 : n55691;
  assign n55693 = pi17 ? n32 : n55692;
  assign n55694 = pi16 ? n32 : n55693;
  assign n55695 = pi15 ? n55694 : n15700;
  assign n55696 = pi14 ? n55688 : n55695;
  assign n55697 = pi13 ? n55681 : n55696;
  assign n55698 = pi12 ? n55678 : n55697;
  assign n55699 = pi11 ? n55667 : n55698;
  assign n55700 = pi14 ? n24578 : n23421;
  assign n55701 = pi13 ? n55700 : n32;
  assign n55702 = pi12 ? n55701 : n32;
  assign n55703 = pi11 ? n55702 : n32;
  assign n55704 = pi10 ? n55699 : n55703;
  assign n55705 = pi09 ? n17493 : n55704;
  assign n55706 = pi14 ? n17279 : n16485;
  assign n55707 = pi13 ? n32 : n55706;
  assign n55708 = pi12 ? n32 : n55707;
  assign n55709 = pi15 ? n17363 : n17188;
  assign n55710 = pi14 ? n55709 : n17188;
  assign n55711 = pi20 ? n12244 : ~n749;
  assign n55712 = pi19 ? n32 : n55711;
  assign n55713 = pi18 ? n32 : n55712;
  assign n55714 = pi17 ? n32 : n55713;
  assign n55715 = pi16 ? n32 : n55714;
  assign n55716 = pi15 ? n55715 : n15695;
  assign n55717 = pi15 ? n15695 : n15863;
  assign n55718 = pi14 ? n55716 : n55717;
  assign n55719 = pi13 ? n55710 : n55718;
  assign n55720 = pi15 ? n40690 : n24874;
  assign n55721 = pi14 ? n55679 : n55720;
  assign n55722 = pi21 ? n51 : ~n206;
  assign n55723 = pi20 ? n55722 : n32;
  assign n55724 = pi19 ? n32 : n55723;
  assign n55725 = pi18 ? n32 : n55724;
  assign n55726 = pi17 ? n32 : n55725;
  assign n55727 = pi16 ? n32 : n55726;
  assign n55728 = pi15 ? n55727 : n16452;
  assign n55729 = pi15 ? n16298 : n15700;
  assign n55730 = pi14 ? n55728 : n55729;
  assign n55731 = pi13 ? n55721 : n55730;
  assign n55732 = pi12 ? n55719 : n55731;
  assign n55733 = pi11 ? n55708 : n55732;
  assign n55734 = pi10 ? n55733 : n40699;
  assign n55735 = pi09 ? n17493 : n55734;
  assign n55736 = pi08 ? n55705 : n55735;
  assign n55737 = pi14 ? n40663 : n16232;
  assign n55738 = pi13 ? n55710 : n55737;
  assign n55739 = pi15 ? n16298 : n16319;
  assign n55740 = pi14 ? n55739 : n38238;
  assign n55741 = pi14 ? n16452 : n40705;
  assign n55742 = pi13 ? n55740 : n55741;
  assign n55743 = pi12 ? n55738 : n55742;
  assign n55744 = pi11 ? n55708 : n55743;
  assign n55745 = pi10 ? n55744 : n40712;
  assign n55746 = pi09 ? n17493 : n55745;
  assign n55747 = pi15 ? n16485 : n16251;
  assign n55748 = pi14 ? n17279 : n55747;
  assign n55749 = pi13 ? n32 : n55748;
  assign n55750 = pi12 ? n32 : n55749;
  assign n55751 = pi20 ? n653 : n564;
  assign n55752 = pi19 ? n32 : n55751;
  assign n55753 = pi18 ? n32 : n55752;
  assign n55754 = pi17 ? n32 : n55753;
  assign n55755 = pi16 ? n32 : n55754;
  assign n55756 = pi15 ? n55755 : n17188;
  assign n55757 = pi14 ? n55756 : n17188;
  assign n55758 = pi13 ? n55757 : n40664;
  assign n55759 = pi15 ? n16293 : n23981;
  assign n55760 = pi15 ? n39569 : n16452;
  assign n55761 = pi14 ? n55759 : n55760;
  assign n55762 = pi13 ? n55761 : n40717;
  assign n55763 = pi12 ? n55758 : n55762;
  assign n55764 = pi11 ? n55750 : n55763;
  assign n55765 = pi10 ? n55764 : n32;
  assign n55766 = pi09 ? n17493 : n55765;
  assign n55767 = pi08 ? n55746 : n55766;
  assign n55768 = pi07 ? n55736 : n55767;
  assign n55769 = pi06 ? n55658 : n55768;
  assign n55770 = pi05 ? n55466 : n55769;
  assign n55771 = pi14 ? n17488 : n16392;
  assign n55772 = pi13 ? n32 : n55771;
  assign n55773 = pi12 ? n32 : n55772;
  assign n55774 = pi11 ? n32 : n55773;
  assign n55775 = pi10 ? n32 : n55774;
  assign n55776 = pi15 ? n17387 : n17188;
  assign n55777 = pi14 ? n55776 : n51504;
  assign n55778 = pi13 ? n32 : n55777;
  assign n55779 = pi12 ? n32 : n55778;
  assign n55780 = pi15 ? n17121 : n17188;
  assign n55781 = pi15 ? n17188 : n16629;
  assign n55782 = pi14 ? n55780 : n55781;
  assign n55783 = pi20 ? n321 : n274;
  assign n55784 = pi19 ? n32 : n55783;
  assign n55785 = pi18 ? n32 : n55784;
  assign n55786 = pi17 ? n32 : n55785;
  assign n55787 = pi16 ? n32 : n55786;
  assign n55788 = pi15 ? n55787 : n15847;
  assign n55789 = pi19 ? n32 : n6350;
  assign n55790 = pi18 ? n32 : n55789;
  assign n55791 = pi17 ? n32 : n55790;
  assign n55792 = pi16 ? n32 : n55791;
  assign n55793 = pi15 ? n15847 : n55792;
  assign n55794 = pi14 ? n55788 : n55793;
  assign n55795 = pi13 ? n55782 : n55794;
  assign n55796 = pi14 ? n16378 : n16515;
  assign n55797 = pi13 ? n55796 : n40740;
  assign n55798 = pi12 ? n55795 : n55797;
  assign n55799 = pi11 ? n55779 : n55798;
  assign n55800 = pi10 ? n55799 : n32;
  assign n55801 = pi09 ? n55775 : n55800;
  assign n55802 = pi15 ? n17367 : n17188;
  assign n55803 = pi14 ? n55802 : n55781;
  assign n55804 = pi20 ? n1839 : n274;
  assign n55805 = pi19 ? n32 : n55804;
  assign n55806 = pi18 ? n32 : n55805;
  assign n55807 = pi17 ? n32 : n55806;
  assign n55808 = pi16 ? n32 : n55807;
  assign n55809 = pi15 ? n55808 : n16333;
  assign n55810 = pi15 ? n16333 : n16392;
  assign n55811 = pi14 ? n55809 : n55810;
  assign n55812 = pi13 ? n55803 : n55811;
  assign n55813 = pi14 ? n32 : n16515;
  assign n55814 = pi13 ? n55813 : n40750;
  assign n55815 = pi12 ? n55812 : n55814;
  assign n55816 = pi11 ? n55779 : n55815;
  assign n55817 = pi10 ? n55816 : n32;
  assign n55818 = pi09 ? n55775 : n55817;
  assign n55819 = pi08 ? n55801 : n55818;
  assign n55820 = pi13 ? n32 : n40587;
  assign n55821 = pi12 ? n32 : n55820;
  assign n55822 = pi19 ? n32 : n31611;
  assign n55823 = pi18 ? n32 : n55822;
  assign n55824 = pi17 ? n32 : n55823;
  assign n55825 = pi16 ? n32 : n55824;
  assign n55826 = pi15 ? n55825 : n16546;
  assign n55827 = pi14 ? n17273 : n55826;
  assign n55828 = pi15 ? n16333 : n52322;
  assign n55829 = pi15 ? n52322 : n32;
  assign n55830 = pi14 ? n55828 : n55829;
  assign n55831 = pi13 ? n55827 : n55830;
  assign n55832 = pi13 ? n24564 : n32;
  assign n55833 = pi12 ? n55831 : n55832;
  assign n55834 = pi11 ? n55821 : n55833;
  assign n55835 = pi10 ? n55834 : n32;
  assign n55836 = pi09 ? n55775 : n55835;
  assign n55837 = pi14 ? n17273 : n16940;
  assign n55838 = pi13 ? n32 : n55837;
  assign n55839 = pi12 ? n32 : n55838;
  assign n55840 = pi15 ? n16546 : n16392;
  assign n55841 = pi14 ? n55840 : n40562;
  assign n55842 = pi13 ? n55827 : n55841;
  assign n55843 = pi12 ? n55842 : n55832;
  assign n55844 = pi11 ? n55839 : n55843;
  assign n55845 = pi10 ? n55844 : n32;
  assign n55846 = pi09 ? n55775 : n55845;
  assign n55847 = pi08 ? n55836 : n55846;
  assign n55848 = pi07 ? n55819 : n55847;
  assign n55849 = pi14 ? n17273 : n16392;
  assign n55850 = pi13 ? n32 : n55849;
  assign n55851 = pi12 ? n32 : n55850;
  assign n55852 = pi20 ? n175 : ~n141;
  assign n55853 = pi19 ? n32 : n55852;
  assign n55854 = pi18 ? n32 : n55853;
  assign n55855 = pi17 ? n32 : n55854;
  assign n55856 = pi16 ? n32 : n55855;
  assign n55857 = pi15 ? n16392 : n55856;
  assign n55858 = pi15 ? n55825 : n16606;
  assign n55859 = pi14 ? n55857 : n55858;
  assign n55860 = pi14 ? n55840 : n16392;
  assign n55861 = pi13 ? n55859 : n55860;
  assign n55862 = pi12 ? n55861 : n40774;
  assign n55863 = pi11 ? n55851 : n55862;
  assign n55864 = pi10 ? n55863 : n32;
  assign n55865 = pi09 ? n17493 : n55864;
  assign n55866 = pi15 ? n16392 : n39670;
  assign n55867 = pi20 ? n151 : ~n141;
  assign n55868 = pi19 ? n32 : n55867;
  assign n55869 = pi18 ? n32 : n55868;
  assign n55870 = pi17 ? n32 : n55869;
  assign n55871 = pi16 ? n32 : n55870;
  assign n55872 = pi15 ? n55871 : n24495;
  assign n55873 = pi14 ? n55866 : n55872;
  assign n55874 = pi13 ? n55873 : n16392;
  assign n55875 = pi12 ? n55874 : n40781;
  assign n55876 = pi11 ? n55851 : n55875;
  assign n55877 = pi10 ? n55876 : n32;
  assign n55878 = pi09 ? n17493 : n55877;
  assign n55879 = pi08 ? n55865 : n55878;
  assign n55880 = pi14 ? n32 : n25633;
  assign n55881 = pi13 ? n32 : n55880;
  assign n55882 = pi12 ? n32 : n55881;
  assign n55883 = pi14 ? n24496 : n55872;
  assign n55884 = pi13 ? n55883 : n40787;
  assign n55885 = pi12 ? n55884 : n32;
  assign n55886 = pi11 ? n55882 : n55885;
  assign n55887 = pi10 ? n55886 : n32;
  assign n55888 = pi09 ? n17493 : n55887;
  assign n55889 = pi13 ? n40855 : n40787;
  assign n55890 = pi12 ? n55889 : n32;
  assign n55891 = pi11 ? n55882 : n55890;
  assign n55892 = pi10 ? n55891 : n32;
  assign n55893 = pi09 ? n17493 : n55892;
  assign n55894 = pi08 ? n55888 : n55893;
  assign n55895 = pi07 ? n55879 : n55894;
  assign n55896 = pi06 ? n55848 : n55895;
  assign n55897 = pi15 ? n17036 : n16392;
  assign n55898 = pi14 ? n25492 : n55897;
  assign n55899 = pi13 ? n17269 : n55898;
  assign n55900 = pi12 ? n32 : n55899;
  assign n55901 = pi14 ? n36851 : n25959;
  assign n55902 = pi14 ? n17039 : n40797;
  assign n55903 = pi13 ? n55901 : n55902;
  assign n55904 = pi12 ? n55903 : n40802;
  assign n55905 = pi11 ? n55900 : n55904;
  assign n55906 = pi10 ? n55905 : n32;
  assign n55907 = pi09 ? n17493 : n55906;
  assign n55908 = pi15 ? n17036 : n16965;
  assign n55909 = pi14 ? n25492 : n55908;
  assign n55910 = pi13 ? n17269 : n55909;
  assign n55911 = pi12 ? n32 : n55910;
  assign n55912 = pi15 ? n17188 : n16965;
  assign n55913 = pi14 ? n17273 : n55912;
  assign n55914 = pi13 ? n55913 : n40809;
  assign n55915 = pi12 ? n55914 : n32;
  assign n55916 = pi11 ? n55911 : n55915;
  assign n55917 = pi10 ? n55916 : n32;
  assign n55918 = pi09 ? n17493 : n55917;
  assign n55919 = pi08 ? n55907 : n55918;
  assign n55920 = pi14 ? n25492 : n17070;
  assign n55921 = pi13 ? n17269 : n55920;
  assign n55922 = pi12 ? n32 : n55921;
  assign n55923 = pi14 ? n17273 : n27858;
  assign n55924 = pi13 ? n55923 : n40820;
  assign n55925 = pi12 ? n55924 : n32;
  assign n55926 = pi11 ? n55922 : n55925;
  assign n55927 = pi10 ? n55926 : n32;
  assign n55928 = pi09 ? n17493 : n55927;
  assign n55929 = pi15 ? n32 : n16919;
  assign n55930 = pi14 ? n32 : n55929;
  assign n55931 = pi14 ? n17090 : n17100;
  assign n55932 = pi13 ? n55930 : n55931;
  assign n55933 = pi12 ? n32 : n55932;
  assign n55934 = pi14 ? n17273 : n17036;
  assign n55935 = pi13 ? n55934 : n40820;
  assign n55936 = pi12 ? n55935 : n32;
  assign n55937 = pi11 ? n55933 : n55936;
  assign n55938 = pi10 ? n55937 : n32;
  assign n55939 = pi09 ? n17493 : n55938;
  assign n55940 = pi08 ? n55928 : n55939;
  assign n55941 = pi07 ? n55919 : n55940;
  assign n55942 = pi13 ? n32 : n51972;
  assign n55943 = pi15 ? n17090 : n17188;
  assign n55944 = pi14 ? n55943 : n17189;
  assign n55945 = pi13 ? n55930 : n55944;
  assign n55946 = pi12 ? n55942 : n55945;
  assign n55947 = pi14 ? n37568 : n17036;
  assign n55948 = pi13 ? n55947 : n40837;
  assign n55949 = pi12 ? n55948 : n32;
  assign n55950 = pi11 ? n55946 : n55949;
  assign n55951 = pi10 ? n55950 : n32;
  assign n55952 = pi09 ? n17493 : n55951;
  assign n55953 = pi14 ? n17188 : n32;
  assign n55954 = pi13 ? n17269 : n55953;
  assign n55955 = pi12 ? n55942 : n55954;
  assign n55956 = pi14 ? n25492 : n17133;
  assign n55957 = pi13 ? n55956 : n40848;
  assign n55958 = pi12 ? n55957 : n32;
  assign n55959 = pi11 ? n55955 : n55958;
  assign n55960 = pi10 ? n55959 : n32;
  assign n55961 = pi09 ? n17493 : n55960;
  assign n55962 = pi08 ? n55952 : n55961;
  assign n55963 = pi14 ? n32 : n17183;
  assign n55964 = pi13 ? n55963 : n55953;
  assign n55965 = pi12 ? n32 : n55964;
  assign n55966 = pi13 ? n55956 : n32;
  assign n55967 = pi12 ? n55966 : n32;
  assign n55968 = pi11 ? n55965 : n55967;
  assign n55969 = pi10 ? n55968 : n32;
  assign n55970 = pi09 ? n17493 : n55969;
  assign n55971 = pi13 ? n55963 : n17375;
  assign n55972 = pi12 ? n32 : n55971;
  assign n55973 = pi14 ? n17273 : n17100;
  assign n55974 = pi13 ? n55973 : n32;
  assign n55975 = pi12 ? n55974 : n32;
  assign n55976 = pi11 ? n55972 : n55975;
  assign n55977 = pi10 ? n55976 : n32;
  assign n55978 = pi09 ? n17493 : n55977;
  assign n55979 = pi08 ? n55970 : n55978;
  assign n55980 = pi07 ? n55962 : n55979;
  assign n55981 = pi06 ? n55941 : n55980;
  assign n55982 = pi05 ? n55896 : n55981;
  assign n55983 = pi04 ? n55770 : n55982;
  assign n55984 = pi03 ? n54938 : n55983;
  assign n55985 = pi13 ? n17313 : n32;
  assign n55986 = pi12 ? n32 : n55985;
  assign n55987 = pi11 ? n55986 : n40877;
  assign n55988 = pi10 ? n55987 : n32;
  assign n55989 = pi09 ? n17493 : n55988;
  assign n55990 = pi09 ? n17493 : n40884;
  assign n55991 = pi08 ? n55989 : n55990;
  assign n55992 = pi07 ? n55991 : n55990;
  assign n55993 = pi07 ? n55990 : n17568;
  assign n55994 = pi06 ? n55992 : n55993;
  assign n55995 = pi05 ? n55994 : n17568;
  assign n55996 = pi04 ? n55995 : n32;
  assign n55997 = pi07 ? n17595 : n17614;
  assign n55998 = pi06 ? n55997 : n17614;
  assign n55999 = pi05 ? n32 : n55998;
  assign n56000 = pi04 ? n32 : n55999;
  assign n56001 = pi03 ? n55996 : n56000;
  assign n56002 = pi02 ? n55984 : n56001;
  assign n56003 = pi07 ? n17614 : n17601;
  assign n56004 = pi06 ? n56003 : n17601;
  assign n56005 = pi06 ? n17601 : n32;
  assign n56006 = pi05 ? n56004 : n56005;
  assign n56007 = pi04 ? n56006 : n32;
  assign n56008 = pi03 ? n17614 : n56007;
  assign n56009 = pi02 ? n56008 : n32;
  assign n56010 = pi01 ? n56002 : n56009;
  assign n56011 = pi00 ? n52477 : n56010;
  assign n56012 = pi16 ? n1683 : ~n2144;
  assign n56013 = pi15 ? n32 : n56012;
  assign n56014 = pi16 ? n1834 : ~n1834;
  assign n56015 = pi16 ? n1581 : ~n1834;
  assign n56016 = pi15 ? n56014 : n56015;
  assign n56017 = pi14 ? n56013 : n56016;
  assign n56018 = pi16 ? n1581 : ~n1581;
  assign n56019 = pi16 ? n1594 : ~n1834;
  assign n56020 = pi15 ? n56018 : n56019;
  assign n56021 = pi14 ? n56020 : n56015;
  assign n56022 = pi13 ? n56017 : n56021;
  assign n56023 = pi12 ? n32 : n56022;
  assign n56024 = pi16 ? n1471 : ~n2144;
  assign n56025 = pi19 ? n266 : n18678;
  assign n56026 = pi18 ? n863 : ~n56025;
  assign n56027 = pi17 ? n32 : n56026;
  assign n56028 = pi17 ? n19904 : n1833;
  assign n56029 = pi16 ? n56027 : ~n56028;
  assign n56030 = pi15 ? n56024 : n56029;
  assign n56031 = pi14 ? n56030 : n28048;
  assign n56032 = pi14 ? n17638 : n18455;
  assign n56033 = pi13 ? n56031 : n56032;
  assign n56034 = pi18 ? n18331 : n18568;
  assign n56035 = pi17 ? n32 : n56034;
  assign n56036 = pi20 ? n17671 : n1324;
  assign n56037 = pi19 ? n18571 : ~n56036;
  assign n56038 = pi19 ? n41755 : n9641;
  assign n56039 = pi18 ? n56037 : ~n56038;
  assign n56040 = pi20 ? n1324 : n287;
  assign n56041 = pi21 ? n259 : ~n7107;
  assign n56042 = pi20 ? n18173 : n56041;
  assign n56043 = pi19 ? n56040 : ~n56042;
  assign n56044 = pi18 ? n56043 : n32;
  assign n56045 = pi17 ? n56039 : ~n56044;
  assign n56046 = pi16 ? n56035 : ~n56045;
  assign n56047 = pi16 ? n19234 : n17850;
  assign n56048 = pi15 ? n56046 : n56047;
  assign n56049 = pi15 ? n17851 : n40978;
  assign n56050 = pi14 ? n56048 : n56049;
  assign n56051 = pi13 ? n17684 : n56050;
  assign n56052 = pi12 ? n56033 : n56051;
  assign n56053 = pi11 ? n56023 : n56052;
  assign n56054 = pi20 ? n32 : n11574;
  assign n56055 = pi19 ? n9007 : n56054;
  assign n56056 = pi18 ? n56055 : ~n32;
  assign n56057 = pi17 ? n32 : n56056;
  assign n56058 = pi16 ? n1233 : ~n56057;
  assign n56059 = pi15 ? n17698 : n56058;
  assign n56060 = pi21 ? n405 : n242;
  assign n56061 = pi20 ? n32 : n56060;
  assign n56062 = pi19 ? n32 : n56061;
  assign n56063 = pi18 ? n56062 : ~n32;
  assign n56064 = pi17 ? n32 : n56063;
  assign n56065 = pi16 ? n1135 : ~n56064;
  assign n56066 = pi15 ? n29519 : n56065;
  assign n56067 = pi14 ? n56059 : n56066;
  assign n56068 = pi13 ? n41007 : n56067;
  assign n56069 = pi12 ? n41006 : n56068;
  assign n56070 = pi16 ? n1135 : ~n1705;
  assign n56071 = pi15 ? n56070 : n29875;
  assign n56072 = pi16 ? n1135 : ~n1843;
  assign n56073 = pi14 ? n56071 : n56072;
  assign n56074 = pi20 ? n220 : ~n2358;
  assign n56075 = pi20 ? n13171 : ~n9488;
  assign n56076 = pi19 ? n56074 : ~n56075;
  assign n56077 = pi18 ? n29658 : n56076;
  assign n56078 = pi17 ? n32 : n56077;
  assign n56079 = pi20 ? n18624 : ~n220;
  assign n56080 = pi19 ? n56079 : n32;
  assign n56081 = pi18 ? n56080 : n41030;
  assign n56082 = pi17 ? n56081 : n1322;
  assign n56083 = pi16 ? n56078 : ~n56082;
  assign n56084 = pi15 ? n29403 : n56083;
  assign n56085 = pi20 ? n220 : ~n1319;
  assign n56086 = pi19 ? n9037 : ~n56085;
  assign n56087 = pi18 ? n56086 : ~n32;
  assign n56088 = pi17 ? n28147 : n56087;
  assign n56089 = pi16 ? n28143 : ~n56088;
  assign n56090 = pi21 ? n309 : n242;
  assign n56091 = pi20 ? n266 : ~n56090;
  assign n56092 = pi19 ? n9037 : ~n56091;
  assign n56093 = pi18 ? n56092 : ~n32;
  assign n56094 = pi17 ? n28147 : n56093;
  assign n56095 = pi16 ? n28143 : ~n56094;
  assign n56096 = pi15 ? n56089 : n56095;
  assign n56097 = pi14 ? n56084 : n56096;
  assign n56098 = pi13 ? n56073 : n56097;
  assign n56099 = pi18 ? n46097 : n32;
  assign n56100 = pi17 ? n17768 : n56099;
  assign n56101 = pi16 ? n32 : n56100;
  assign n56102 = pi18 ? n728 : n237;
  assign n56103 = pi17 ? n32 : n56102;
  assign n56104 = pi19 ? n1757 : n267;
  assign n56105 = pi18 ? n56104 : n32;
  assign n56106 = pi17 ? n28194 : ~n56105;
  assign n56107 = pi16 ? n56103 : ~n56106;
  assign n56108 = pi15 ? n56101 : n56107;
  assign n56109 = pi14 ? n17765 : n56108;
  assign n56110 = pi13 ? n17748 : n56109;
  assign n56111 = pi12 ? n56098 : n56110;
  assign n56112 = pi11 ? n56069 : n56111;
  assign n56113 = pi10 ? n56053 : n56112;
  assign n56114 = pi09 ? n32 : n56113;
  assign n56115 = pi16 ? n1834 : ~n1581;
  assign n56116 = pi15 ? n32 : n56115;
  assign n56117 = pi15 ? n56015 : n56019;
  assign n56118 = pi14 ? n56116 : n56117;
  assign n56119 = pi16 ? n1594 : ~n1577;
  assign n56120 = pi15 ? n56018 : n56119;
  assign n56121 = pi16 ? n1581 : ~n18985;
  assign n56122 = pi16 ? n1581 : ~n1577;
  assign n56123 = pi15 ? n56121 : n56122;
  assign n56124 = pi14 ? n56120 : n56123;
  assign n56125 = pi13 ? n56118 : n56124;
  assign n56126 = pi12 ? n32 : n56125;
  assign n56127 = pi19 ? n32 : n14319;
  assign n56128 = pi18 ? n56127 : ~n32;
  assign n56129 = pi17 ? n32 : n56128;
  assign n56130 = pi16 ? n56129 : ~n1834;
  assign n56131 = pi17 ? n19904 : n1576;
  assign n56132 = pi16 ? n56027 : ~n56131;
  assign n56133 = pi15 ? n56130 : n56132;
  assign n56134 = pi14 ? n56133 : n28233;
  assign n56135 = pi15 ? n32 : n17825;
  assign n56136 = pi14 ? n32 : n56135;
  assign n56137 = pi13 ? n56134 : n56136;
  assign n56138 = pi15 ? n17800 : n17682;
  assign n56139 = pi14 ? n17794 : n56138;
  assign n56140 = pi18 ? n29364 : n18405;
  assign n56141 = pi17 ? n32 : n56140;
  assign n56142 = pi20 ? n18282 : n17669;
  assign n56143 = pi19 ? n18409 : ~n56142;
  assign n56144 = pi20 ? n17669 : ~n19731;
  assign n56145 = pi19 ? n56144 : n18073;
  assign n56146 = pi18 ? n56143 : ~n56145;
  assign n56147 = pi20 ? n17669 : n287;
  assign n56148 = pi20 ? n18832 : n2019;
  assign n56149 = pi19 ? n56147 : ~n56148;
  assign n56150 = pi18 ? n56149 : n32;
  assign n56151 = pi17 ? n56146 : ~n56150;
  assign n56152 = pi16 ? n56141 : ~n56151;
  assign n56153 = pi16 ? n19234 : n18162;
  assign n56154 = pi15 ? n56152 : n56153;
  assign n56155 = pi20 ? n32 : n13785;
  assign n56156 = pi19 ? n32 : n56155;
  assign n56157 = pi18 ? n56156 : n32;
  assign n56158 = pi17 ? n32 : n56157;
  assign n56159 = pi16 ? n32 : n56158;
  assign n56160 = pi15 ? n56159 : n41166;
  assign n56161 = pi14 ? n56154 : n56160;
  assign n56162 = pi13 ? n56139 : n56161;
  assign n56163 = pi12 ? n56137 : n56162;
  assign n56164 = pi11 ? n56126 : n56163;
  assign n56165 = pi15 ? n41179 : n17825;
  assign n56166 = pi14 ? n41175 : n56165;
  assign n56167 = pi13 ? n56166 : n41183;
  assign n56168 = pi20 ? n32 : n18256;
  assign n56169 = pi19 ? n9007 : n56168;
  assign n56170 = pi18 ? n56169 : ~n32;
  assign n56171 = pi17 ? n32 : n56170;
  assign n56172 = pi16 ? n1233 : ~n56171;
  assign n56173 = pi15 ? n17822 : n56172;
  assign n56174 = pi15 ? n29519 : n28947;
  assign n56175 = pi14 ? n56173 : n56174;
  assign n56176 = pi13 ? n41186 : n56175;
  assign n56177 = pi12 ? n56167 : n56176;
  assign n56178 = pi19 ? n32 : n56054;
  assign n56179 = pi18 ? n56178 : ~n32;
  assign n56180 = pi17 ? n32 : n56179;
  assign n56181 = pi16 ? n1135 : ~n56180;
  assign n56182 = pi15 ? n29676 : n56181;
  assign n56183 = pi16 ? n1233 : ~n1323;
  assign n56184 = pi15 ? n28947 : n56183;
  assign n56185 = pi14 ? n56182 : n56184;
  assign n56186 = pi16 ? n19652 : ~n1594;
  assign n56187 = pi19 ? n28130 : n17649;
  assign n56188 = pi18 ? n335 : n56187;
  assign n56189 = pi17 ? n32 : n56188;
  assign n56190 = pi20 ? n518 : n439;
  assign n56191 = pi19 ? n32 : n56190;
  assign n56192 = pi18 ? n56080 : n56191;
  assign n56193 = pi17 ? n56192 : n1593;
  assign n56194 = pi16 ? n56189 : ~n56193;
  assign n56195 = pi15 ? n56186 : n56194;
  assign n56196 = pi14 ? n56195 : n56096;
  assign n56197 = pi13 ? n56185 : n56196;
  assign n56198 = pi19 ? n1757 : n6057;
  assign n56199 = pi18 ? n56198 : n32;
  assign n56200 = pi17 ? n28194 : ~n56199;
  assign n56201 = pi16 ? n56103 : ~n56200;
  assign n56202 = pi15 ? n56101 : n56201;
  assign n56203 = pi14 ? n17765 : n56202;
  assign n56204 = pi13 ? n17748 : n56203;
  assign n56205 = pi12 ? n56197 : n56204;
  assign n56206 = pi11 ? n56177 : n56205;
  assign n56207 = pi10 ? n56164 : n56206;
  assign n56208 = pi09 ? n32 : n56207;
  assign n56209 = pi08 ? n56114 : n56208;
  assign n56210 = pi07 ? n32 : n56209;
  assign n56211 = pi06 ? n32 : n56210;
  assign n56212 = pi16 ? n1834 : ~n1683;
  assign n56213 = pi15 ? n32 : n56212;
  assign n56214 = pi16 ? n1581 : ~n1683;
  assign n56215 = pi14 ? n56213 : n56214;
  assign n56216 = pi15 ? n56019 : n18979;
  assign n56217 = pi15 ? n30304 : n43521;
  assign n56218 = pi14 ? n56216 : n56217;
  assign n56219 = pi13 ? n56215 : n56218;
  assign n56220 = pi12 ? n32 : n56219;
  assign n56221 = pi15 ? n43574 : n17885;
  assign n56222 = pi14 ? n56221 : n32;
  assign n56223 = pi13 ? n56222 : n17887;
  assign n56224 = pi20 ? n448 : n175;
  assign n56225 = pi19 ? n32 : n56224;
  assign n56226 = pi19 ? n29270 : n8622;
  assign n56227 = pi18 ? n56225 : n56226;
  assign n56228 = pi20 ? n339 : n310;
  assign n56229 = pi19 ? n56228 : ~n4670;
  assign n56230 = pi18 ? n56229 : n1676;
  assign n56231 = pi17 ? n56227 : ~n56230;
  assign n56232 = pi16 ? n41019 : n56231;
  assign n56233 = pi15 ? n56232 : n18972;
  assign n56234 = pi14 ? n17895 : n56233;
  assign n56235 = pi18 ? n28178 : ~n32;
  assign n56236 = pi17 ? n32 : n56235;
  assign n56237 = pi19 ? n32 : n29470;
  assign n56238 = pi18 ? n56237 : n29474;
  assign n56239 = pi20 ? n310 : ~n18415;
  assign n56240 = pi19 ? n56239 : ~n1324;
  assign n56241 = pi18 ? n56240 : n32;
  assign n56242 = pi17 ? n56238 : ~n56241;
  assign n56243 = pi16 ? n56236 : ~n56242;
  assign n56244 = pi19 ? n17652 : n30044;
  assign n56245 = pi18 ? n29658 : n56244;
  assign n56246 = pi17 ? n32 : n56245;
  assign n56247 = pi19 ? n36181 : ~n6822;
  assign n56248 = pi20 ? n333 : ~n9194;
  assign n56249 = pi19 ? n56248 : n17652;
  assign n56250 = pi18 ? n56247 : ~n56249;
  assign n56251 = pi19 ? n17670 : ~n31309;
  assign n56252 = pi18 ? n56251 : n32;
  assign n56253 = pi17 ? n56250 : ~n56252;
  assign n56254 = pi16 ? n56246 : ~n56253;
  assign n56255 = pi15 ? n56243 : n56254;
  assign n56256 = pi14 ? n56255 : n41350;
  assign n56257 = pi13 ? n56234 : n56256;
  assign n56258 = pi12 ? n56223 : n56257;
  assign n56259 = pi11 ? n56220 : n56258;
  assign n56260 = pi14 ? n17903 : n41552;
  assign n56261 = pi13 ? n41378 : n56260;
  assign n56262 = pi20 ? n18253 : n18281;
  assign n56263 = pi19 ? n28081 : ~n56262;
  assign n56264 = pi18 ? n312 : ~n56263;
  assign n56265 = pi17 ? n32 : n56264;
  assign n56266 = pi20 ? n12884 : n309;
  assign n56267 = pi19 ? n35635 : ~n56266;
  assign n56268 = pi20 ? n287 : n13171;
  assign n56269 = pi20 ? n17669 : n17652;
  assign n56270 = pi19 ? n56268 : ~n56269;
  assign n56271 = pi18 ? n56267 : n56270;
  assign n56272 = pi20 ? n333 : ~n314;
  assign n56273 = pi20 ? n1817 : n22910;
  assign n56274 = pi19 ? n56272 : n56273;
  assign n56275 = pi18 ? n56274 : ~n32;
  assign n56276 = pi17 ? n56271 : ~n56275;
  assign n56277 = pi16 ? n56265 : n56276;
  assign n56278 = pi20 ? n32 : n22910;
  assign n56279 = pi19 ? n32 : n56278;
  assign n56280 = pi18 ? n56279 : ~n32;
  assign n56281 = pi17 ? n32 : n56280;
  assign n56282 = pi16 ? n1135 : ~n56281;
  assign n56283 = pi15 ? n56277 : n56282;
  assign n56284 = pi15 ? n29676 : n41405;
  assign n56285 = pi14 ? n56283 : n56284;
  assign n56286 = pi13 ? n41387 : n56285;
  assign n56287 = pi12 ? n56261 : n56286;
  assign n56288 = pi17 ? n32 : n30233;
  assign n56289 = pi16 ? n1214 : ~n56288;
  assign n56290 = pi15 ? n29875 : n56289;
  assign n56291 = pi20 ? n32 : n18610;
  assign n56292 = pi19 ? n32 : n56291;
  assign n56293 = pi18 ? n56292 : ~n32;
  assign n56294 = pi17 ? n32 : n56293;
  assign n56295 = pi16 ? n1214 : ~n56294;
  assign n56296 = pi15 ? n56295 : n42685;
  assign n56297 = pi14 ? n56290 : n56296;
  assign n56298 = pi19 ? n343 : ~n507;
  assign n56299 = pi18 ? n56298 : n32;
  assign n56300 = pi17 ? n28422 : n56299;
  assign n56301 = pi16 ? n19804 : n56300;
  assign n56302 = pi15 ? n30025 : n56301;
  assign n56303 = pi19 ? n208 : ~n22558;
  assign n56304 = pi18 ? n56303 : n32;
  assign n56305 = pi17 ? n28428 : n56304;
  assign n56306 = pi16 ? n32 : n56305;
  assign n56307 = pi15 ? n56306 : n17937;
  assign n56308 = pi14 ? n56302 : n56307;
  assign n56309 = pi13 ? n56297 : n56308;
  assign n56310 = pi17 ? n28450 : n17979;
  assign n56311 = pi16 ? n32 : n56310;
  assign n56312 = pi19 ? n28456 : ~n17982;
  assign n56313 = pi18 ? n56312 : ~n32;
  assign n56314 = pi17 ? n32 : n56313;
  assign n56315 = pi16 ? n1233 : ~n56314;
  assign n56316 = pi15 ? n56311 : n56315;
  assign n56317 = pi14 ? n17973 : n56316;
  assign n56318 = pi13 ? n17960 : n56317;
  assign n56319 = pi12 ? n56309 : n56318;
  assign n56320 = pi11 ? n56287 : n56319;
  assign n56321 = pi10 ? n56259 : n56320;
  assign n56322 = pi09 ? n32 : n56321;
  assign n56323 = pi15 ? n32 : n56214;
  assign n56324 = pi16 ? n1594 : ~n1683;
  assign n56325 = pi15 ? n56324 : n56214;
  assign n56326 = pi14 ? n56323 : n56325;
  assign n56327 = pi18 ? n936 : n1676;
  assign n56328 = pi17 ? n32 : n56327;
  assign n56329 = pi16 ? n1594 : ~n56328;
  assign n56330 = pi16 ? n1233 : ~n1678;
  assign n56331 = pi15 ? n56329 : n56330;
  assign n56332 = pi16 ? n29318 : ~n1678;
  assign n56333 = pi15 ? n41479 : n56332;
  assign n56334 = pi14 ? n56331 : n56333;
  assign n56335 = pi13 ? n56326 : n56334;
  assign n56336 = pi12 ? n32 : n56335;
  assign n56337 = pi15 ? n56330 : n17894;
  assign n56338 = pi14 ? n56337 : n18008;
  assign n56339 = pi13 ? n56338 : n18003;
  assign n56340 = pi19 ? n32 : n28483;
  assign n56341 = pi18 ? n56340 : n56226;
  assign n56342 = pi18 ? n56229 : ~n32;
  assign n56343 = pi17 ? n56341 : ~n56342;
  assign n56344 = pi16 ? n41019 : n56343;
  assign n56345 = pi15 ? n56344 : n32;
  assign n56346 = pi14 ? n29508 : n56345;
  assign n56347 = pi18 ? n56240 : ~n618;
  assign n56348 = pi17 ? n56238 : ~n56347;
  assign n56349 = pi16 ? n56236 : ~n56348;
  assign n56350 = pi19 ? n17670 : ~n17652;
  assign n56351 = pi18 ? n56350 : ~n618;
  assign n56352 = pi17 ? n56250 : ~n56351;
  assign n56353 = pi16 ? n56246 : ~n56352;
  assign n56354 = pi15 ? n56349 : n56353;
  assign n56355 = pi14 ? n56354 : n41531;
  assign n56356 = pi13 ? n56346 : n56355;
  assign n56357 = pi12 ? n56339 : n56356;
  assign n56358 = pi11 ? n56336 : n56357;
  assign n56359 = pi18 ? n41548 : ~n1676;
  assign n56360 = pi17 ? n3282 : n56359;
  assign n56361 = pi16 ? n32 : n56360;
  assign n56362 = pi15 ? n32 : n56361;
  assign n56363 = pi14 ? n17891 : n56362;
  assign n56364 = pi13 ? n41547 : n56363;
  assign n56365 = pi21 ? n140 : n313;
  assign n56366 = pi20 ? n32 : n56365;
  assign n56367 = pi19 ? n32 : n56366;
  assign n56368 = pi19 ? n43407 : ~n41294;
  assign n56369 = pi18 ? n56367 : ~n56368;
  assign n56370 = pi17 ? n32 : n56369;
  assign n56371 = pi20 ? n18415 : ~n18762;
  assign n56372 = pi19 ? n56371 : ~n49221;
  assign n56373 = pi20 ? n17665 : ~n20396;
  assign n56374 = pi20 ? n3523 : n6822;
  assign n56375 = pi19 ? n56373 : n56374;
  assign n56376 = pi18 ? n56372 : ~n56375;
  assign n56377 = pi20 ? n1817 : n1385;
  assign n56378 = pi19 ? n56272 : n56377;
  assign n56379 = pi18 ? n56378 : ~n32;
  assign n56380 = pi17 ? n56376 : ~n56379;
  assign n56381 = pi16 ? n56370 : n56380;
  assign n56382 = pi18 ? n17912 : ~n32;
  assign n56383 = pi17 ? n32 : n56382;
  assign n56384 = pi16 ? n1233 : ~n56383;
  assign n56385 = pi15 ? n56381 : n56384;
  assign n56386 = pi20 ? n32 : ~n2077;
  assign n56387 = pi19 ? n32 : n56386;
  assign n56388 = pi18 ? n56387 : ~n32;
  assign n56389 = pi17 ? n32 : n56388;
  assign n56390 = pi16 ? n1135 : ~n56389;
  assign n56391 = pi15 ? n29676 : n56390;
  assign n56392 = pi14 ? n56385 : n56391;
  assign n56393 = pi13 ? n41555 : n56392;
  assign n56394 = pi12 ? n56364 : n56393;
  assign n56395 = pi21 ? n206 : ~n2076;
  assign n56396 = pi20 ? n32 : n56395;
  assign n56397 = pi19 ? n32 : n56396;
  assign n56398 = pi18 ? n56397 : ~n32;
  assign n56399 = pi17 ? n32 : n56398;
  assign n56400 = pi16 ? n1233 : ~n56399;
  assign n56401 = pi16 ? n19652 : ~n56288;
  assign n56402 = pi15 ? n56400 : n56401;
  assign n56403 = pi14 ? n56402 : n56296;
  assign n56404 = pi15 ? n28947 : n56301;
  assign n56405 = pi19 ? n208 : ~n1508;
  assign n56406 = pi18 ? n56405 : n32;
  assign n56407 = pi17 ? n28428 : n56406;
  assign n56408 = pi16 ? n32 : n56407;
  assign n56409 = pi15 ? n56408 : n17937;
  assign n56410 = pi14 ? n56404 : n56409;
  assign n56411 = pi13 ? n56403 : n56410;
  assign n56412 = pi19 ? n594 : n13632;
  assign n56413 = pi18 ? n56412 : n32;
  assign n56414 = pi17 ? n32 : n56413;
  assign n56415 = pi16 ? n32 : n56414;
  assign n56416 = pi15 ? n17945 : n56415;
  assign n56417 = pi19 ? n32 : n18041;
  assign n56418 = pi18 ? n56417 : n32;
  assign n56419 = pi17 ? n32 : n56418;
  assign n56420 = pi16 ? n32 : n56419;
  assign n56421 = pi19 ? n322 : n28408;
  assign n56422 = pi18 ? n56421 : n32;
  assign n56423 = pi17 ? n32 : n56422;
  assign n56424 = pi16 ? n32 : n56423;
  assign n56425 = pi15 ? n56420 : n56424;
  assign n56426 = pi14 ? n56416 : n56425;
  assign n56427 = pi19 ? n4126 : n36073;
  assign n56428 = pi18 ? n56427 : n32;
  assign n56429 = pi17 ? n18395 : n56428;
  assign n56430 = pi16 ? n32 : n56429;
  assign n56431 = pi21 ? n10182 : ~n173;
  assign n56432 = pi20 ? n32 : n56431;
  assign n56433 = pi19 ? n32 : n56432;
  assign n56434 = pi18 ? n56433 : n28557;
  assign n56435 = pi17 ? n32 : n56434;
  assign n56436 = pi19 ? n28565 : n17982;
  assign n56437 = pi18 ? n56436 : n32;
  assign n56438 = pi17 ? n28564 : ~n56437;
  assign n56439 = pi16 ? n56435 : ~n56438;
  assign n56440 = pi15 ? n56430 : n56439;
  assign n56441 = pi14 ? n18053 : n56440;
  assign n56442 = pi13 ? n56426 : n56441;
  assign n56443 = pi12 ? n56411 : n56442;
  assign n56444 = pi11 ? n56394 : n56443;
  assign n56445 = pi10 ? n56358 : n56444;
  assign n56446 = pi09 ? n32 : n56445;
  assign n56447 = pi08 ? n56322 : n56446;
  assign n56448 = pi20 ? n18129 : ~n18415;
  assign n56449 = pi19 ? n56448 : ~n30044;
  assign n56450 = pi18 ? n32 : n56449;
  assign n56451 = pi17 ? n32 : n56450;
  assign n56452 = pi19 ? n36181 : ~n47881;
  assign n56453 = pi20 ? n1331 : ~n2358;
  assign n56454 = pi19 ? n23180 : n56453;
  assign n56455 = pi18 ? n56452 : n56454;
  assign n56456 = pi19 ? n6683 : ~n19596;
  assign n56457 = pi18 ? n56456 : ~n32;
  assign n56458 = pi17 ? n56455 : ~n56457;
  assign n56459 = pi16 ? n56451 : n56458;
  assign n56460 = pi16 ? n1581 : ~n3356;
  assign n56461 = pi15 ? n56459 : n56460;
  assign n56462 = pi16 ? n1594 : ~n3356;
  assign n56463 = pi15 ? n56462 : n56460;
  assign n56464 = pi14 ? n56461 : n56463;
  assign n56465 = pi20 ? n2358 : ~n206;
  assign n56466 = pi19 ? n56465 : n29023;
  assign n56467 = pi18 ? n29021 : n56466;
  assign n56468 = pi19 ? n1757 : ~n28686;
  assign n56469 = pi18 ? n56468 : ~n32;
  assign n56470 = pi17 ? n56467 : ~n56469;
  assign n56471 = pi16 ? n29019 : n56470;
  assign n56472 = pi15 ? n18979 : n56471;
  assign n56473 = pi14 ? n19349 : n56472;
  assign n56474 = pi13 ? n56464 : n56473;
  assign n56475 = pi12 ? n32 : n56474;
  assign n56476 = pi16 ? n1705 : ~n3356;
  assign n56477 = pi15 ? n56476 : n18008;
  assign n56478 = pi14 ? n56477 : n18080;
  assign n56479 = pi14 ? n17997 : n18092;
  assign n56480 = pi13 ? n56478 : n56479;
  assign n56481 = pi20 ? n321 : ~n18762;
  assign n56482 = pi19 ? n56481 : ~n428;
  assign n56483 = pi18 ? n56482 : ~n18076;
  assign n56484 = pi17 ? n41654 : ~n56483;
  assign n56485 = pi16 ? n41651 : n56484;
  assign n56486 = pi15 ? n18137 : n56485;
  assign n56487 = pi14 ? n18121 : n56486;
  assign n56488 = pi19 ? n4670 : n342;
  assign n56489 = pi18 ? n32 : n56488;
  assign n56490 = pi18 ? n18397 : ~n32;
  assign n56491 = pi17 ? n56489 : n56490;
  assign n56492 = pi16 ? n1214 : ~n56491;
  assign n56493 = pi18 ? n36402 : ~n3350;
  assign n56494 = pi17 ? n41668 : ~n56493;
  assign n56495 = pi16 ? n41666 : ~n56494;
  assign n56496 = pi15 ? n56492 : n56495;
  assign n56497 = pi14 ? n56496 : n41682;
  assign n56498 = pi13 ? n56487 : n56497;
  assign n56499 = pi12 ? n56480 : n56498;
  assign n56500 = pi11 ? n56475 : n56499;
  assign n56501 = pi15 ? n41862 : n28620;
  assign n56502 = pi14 ? n41859 : n56501;
  assign n56503 = pi15 ? n28627 : n17891;
  assign n56504 = pi14 ? n17891 : n56503;
  assign n56505 = pi13 ? n56502 : n56504;
  assign n56506 = pi15 ? n32 : n17894;
  assign n56507 = pi14 ? n56506 : n32;
  assign n56508 = pi16 ? n1233 : ~n28804;
  assign n56509 = pi17 ? n32 : n44150;
  assign n56510 = pi16 ? n1233 : ~n56509;
  assign n56511 = pi15 ? n56508 : n56510;
  assign n56512 = pi15 ? n42857 : n29240;
  assign n56513 = pi14 ? n56511 : n56512;
  assign n56514 = pi13 ? n56507 : n56513;
  assign n56515 = pi12 ? n56505 : n56514;
  assign n56516 = pi20 ? n32 : n7108;
  assign n56517 = pi19 ? n32 : n56516;
  assign n56518 = pi18 ? n56517 : ~n32;
  assign n56519 = pi17 ? n32 : n56518;
  assign n56520 = pi16 ? n1233 : ~n56519;
  assign n56521 = pi15 ? n42685 : n56520;
  assign n56522 = pi16 ? n1233 : ~n56288;
  assign n56523 = pi19 ? n32 : n54022;
  assign n56524 = pi18 ? n56523 : ~n32;
  assign n56525 = pi17 ? n32 : n56524;
  assign n56526 = pi16 ? n1233 : ~n56525;
  assign n56527 = pi15 ? n56522 : n56526;
  assign n56528 = pi14 ? n56521 : n56527;
  assign n56529 = pi20 ? n32 : n18624;
  assign n56530 = pi19 ? n32 : n56529;
  assign n56531 = pi20 ? n18832 : n314;
  assign n56532 = pi19 ? n41868 : ~n56531;
  assign n56533 = pi18 ? n56530 : ~n56532;
  assign n56534 = pi17 ? n32 : n56533;
  assign n56535 = pi20 ? n18415 : ~n405;
  assign n56536 = pi20 ? n174 : n333;
  assign n56537 = pi19 ? n56535 : ~n56536;
  assign n56538 = pi20 ? n20944 : ~n333;
  assign n56539 = pi19 ? n56538 : ~n28081;
  assign n56540 = pi18 ? n56537 : n56539;
  assign n56541 = pi20 ? n174 : n9863;
  assign n56542 = pi21 ? n309 : n1939;
  assign n56543 = pi20 ? n32 : n56542;
  assign n56544 = pi19 ? n56541 : n56543;
  assign n56545 = pi18 ? n56544 : ~n32;
  assign n56546 = pi17 ? n56540 : ~n56545;
  assign n56547 = pi16 ? n56534 : n56546;
  assign n56548 = pi19 ? n208 : ~n56291;
  assign n56549 = pi18 ? n56548 : n32;
  assign n56550 = pi17 ? n32 : n56549;
  assign n56551 = pi16 ? n32 : n56550;
  assign n56552 = pi15 ? n56547 : n56551;
  assign n56553 = pi15 ? n18859 : n17846;
  assign n56554 = pi14 ? n56552 : n56553;
  assign n56555 = pi13 ? n56528 : n56554;
  assign n56556 = pi19 ? n33683 : n17766;
  assign n56557 = pi18 ? n1395 : ~n56556;
  assign n56558 = pi17 ? n32 : n56557;
  assign n56559 = pi17 ? n32 : n18206;
  assign n56560 = pi16 ? n56558 : ~n56559;
  assign n56561 = pi15 ? n18196 : n56560;
  assign n56562 = pi18 ? n1613 : n32;
  assign n56563 = pi17 ? n32 : n56562;
  assign n56564 = pi16 ? n56563 : n18216;
  assign n56565 = pi18 ? n23194 : n28682;
  assign n56566 = pi17 ? n32 : n56565;
  assign n56567 = pi18 ? n37675 : ~n32;
  assign n56568 = pi17 ? n28688 : n56567;
  assign n56569 = pi16 ? n56566 : ~n56568;
  assign n56570 = pi15 ? n56564 : n56569;
  assign n56571 = pi14 ? n56561 : n56570;
  assign n56572 = pi13 ? n18192 : n56571;
  assign n56573 = pi12 ? n56555 : n56572;
  assign n56574 = pi11 ? n56515 : n56573;
  assign n56575 = pi10 ? n56500 : n56574;
  assign n56576 = pi09 ? n32 : n56575;
  assign n56577 = pi20 ? n18408 : ~n6822;
  assign n56578 = pi20 ? n9641 : n6085;
  assign n56579 = pi19 ? n56577 : ~n56578;
  assign n56580 = pi18 ? n858 : n56579;
  assign n56581 = pi17 ? n32 : n56580;
  assign n56582 = pi20 ? n448 : ~n18253;
  assign n56583 = pi20 ? n6822 : ~n9488;
  assign n56584 = pi19 ? n56582 : n56583;
  assign n56585 = pi20 ? n29452 : n9194;
  assign n56586 = pi20 ? n9488 : ~n17669;
  assign n56587 = pi19 ? n56585 : n56586;
  assign n56588 = pi18 ? n56584 : ~n56587;
  assign n56589 = pi20 ? n17669 : ~n18073;
  assign n56590 = pi19 ? n56589 : ~n44185;
  assign n56591 = pi18 ? n56590 : ~n32;
  assign n56592 = pi17 ? n56588 : n56591;
  assign n56593 = pi16 ? n56581 : ~n56592;
  assign n56594 = pi16 ? n1594 : ~n3352;
  assign n56595 = pi15 ? n56593 : n56594;
  assign n56596 = pi16 ? n1581 : ~n3352;
  assign n56597 = pi15 ? n43933 : n56596;
  assign n56598 = pi14 ? n56595 : n56597;
  assign n56599 = pi18 ? n32 : ~n18076;
  assign n56600 = pi17 ? n32 : n56599;
  assign n56601 = pi16 ? n1233 : ~n56600;
  assign n56602 = pi20 ? n820 : ~n11107;
  assign n56603 = pi19 ? n56602 : n28850;
  assign n56604 = pi18 ? n28848 : n56603;
  assign n56605 = pi19 ? n5614 : ~n28854;
  assign n56606 = pi18 ? n56605 : ~n359;
  assign n56607 = pi17 ? n56604 : ~n56606;
  assign n56608 = pi16 ? n28845 : n56607;
  assign n56609 = pi15 ? n56601 : n56608;
  assign n56610 = pi14 ? n44289 : n56609;
  assign n56611 = pi13 ? n56598 : n56610;
  assign n56612 = pi12 ? n32 : n56611;
  assign n56613 = pi16 ? n1705 : ~n3352;
  assign n56614 = pi15 ? n56613 : n19172;
  assign n56615 = pi18 ? n18075 : n359;
  assign n56616 = pi17 ? n18072 : n56615;
  assign n56617 = pi16 ? n32 : n56616;
  assign n56618 = pi15 ? n56617 : n32;
  assign n56619 = pi14 ? n56614 : n56618;
  assign n56620 = pi14 ? n18143 : n18238;
  assign n56621 = pi13 ? n56619 : n56620;
  assign n56622 = pi18 ? n56482 : ~n359;
  assign n56623 = pi17 ? n41654 : ~n56622;
  assign n56624 = pi16 ? n41651 : n56623;
  assign n56625 = pi15 ? n18289 : n56624;
  assign n56626 = pi14 ? n18273 : n56625;
  assign n56627 = pi18 ? n209 : ~n9170;
  assign n56628 = pi17 ? n32 : n56627;
  assign n56629 = pi16 ? n56628 : ~n56491;
  assign n56630 = pi18 ? n36402 : ~n237;
  assign n56631 = pi17 ? n41668 : ~n56630;
  assign n56632 = pi16 ? n41666 : ~n56631;
  assign n56633 = pi15 ? n56629 : n56632;
  assign n56634 = pi14 ? n56633 : n41851;
  assign n56635 = pi13 ? n56626 : n56634;
  assign n56636 = pi12 ? n56621 : n56635;
  assign n56637 = pi11 ? n56612 : n56636;
  assign n56638 = pi18 ? n41366 : n3350;
  assign n56639 = pi17 ? n41365 : ~n56638;
  assign n56640 = pi16 ? n32 : n56639;
  assign n56641 = pi15 ? n41693 : n56640;
  assign n56642 = pi18 ? n41695 : n3350;
  assign n56643 = pi17 ? n8193 : ~n56642;
  assign n56644 = pi16 ? n32 : n56643;
  assign n56645 = pi15 ? n56644 : n28727;
  assign n56646 = pi14 ? n56641 : n56645;
  assign n56647 = pi15 ? n28732 : n18439;
  assign n56648 = pi14 ? n18439 : n56647;
  assign n56649 = pi13 ? n56646 : n56648;
  assign n56650 = pi18 ? n222 : n1676;
  assign n56651 = pi17 ? n32 : n56650;
  assign n56652 = pi16 ? n1135 : ~n56651;
  assign n56653 = pi18 ? n19350 : n1676;
  assign n56654 = pi17 ? n32 : n56653;
  assign n56655 = pi16 ? n1233 : ~n56654;
  assign n56656 = pi15 ? n56652 : n56655;
  assign n56657 = pi16 ? n1214 : ~n43707;
  assign n56658 = pi15 ? n56186 : n56657;
  assign n56659 = pi14 ? n56656 : n56658;
  assign n56660 = pi13 ? n32 : n56659;
  assign n56661 = pi12 ? n56649 : n56660;
  assign n56662 = pi18 ? n17819 : ~n32;
  assign n56663 = pi17 ? n32 : n56662;
  assign n56664 = pi16 ? n1233 : ~n56663;
  assign n56665 = pi16 ? n1135 : ~n56519;
  assign n56666 = pi15 ? n56664 : n56665;
  assign n56667 = pi17 ? n28638 : n30233;
  assign n56668 = pi16 ? n1135 : ~n56667;
  assign n56669 = pi16 ? n1135 : ~n2144;
  assign n56670 = pi15 ? n56668 : n56669;
  assign n56671 = pi14 ? n56666 : n56670;
  assign n56672 = pi20 ? n9491 : n18415;
  assign n56673 = pi19 ? n41868 : ~n56672;
  assign n56674 = pi18 ? n29681 : ~n56673;
  assign n56675 = pi17 ? n32 : n56674;
  assign n56676 = pi19 ? n41878 : ~n1612;
  assign n56677 = pi18 ? n56676 : n32;
  assign n56678 = pi17 ? n41877 : n56677;
  assign n56679 = pi16 ? n56675 : n56678;
  assign n56680 = pi15 ? n56679 : n28766;
  assign n56681 = pi19 ? n28781 : ~n2141;
  assign n56682 = pi18 ? n56681 : n32;
  assign n56683 = pi17 ? n28780 : n56682;
  assign n56684 = pi16 ? n28773 : n56683;
  assign n56685 = pi15 ? n56684 : n17846;
  assign n56686 = pi14 ? n56680 : n56685;
  assign n56687 = pi13 ? n56671 : n56686;
  assign n56688 = pi18 ? n209 : ~n56556;
  assign n56689 = pi17 ? n32 : n56688;
  assign n56690 = pi16 ? n56689 : ~n56559;
  assign n56691 = pi15 ? n18355 : n56690;
  assign n56692 = pi18 ? n12172 : n32;
  assign n56693 = pi17 ? n32 : n56692;
  assign n56694 = pi16 ? n56693 : n18216;
  assign n56695 = pi20 ? n32 : n55594;
  assign n56696 = pi19 ? n32 : n56695;
  assign n56697 = pi18 ? n56696 : n28682;
  assign n56698 = pi17 ? n32 : n56697;
  assign n56699 = pi19 ? n22185 : ~n1818;
  assign n56700 = pi18 ? n56699 : ~n32;
  assign n56701 = pi17 ? n28688 : n56700;
  assign n56702 = pi16 ? n56698 : ~n56701;
  assign n56703 = pi15 ? n56694 : n56702;
  assign n56704 = pi14 ? n56691 : n56703;
  assign n56705 = pi13 ? n18351 : n56704;
  assign n56706 = pi12 ? n56687 : n56705;
  assign n56707 = pi11 ? n56661 : n56706;
  assign n56708 = pi10 ? n56637 : n56707;
  assign n56709 = pi09 ? n32 : n56708;
  assign n56710 = pi08 ? n56576 : n56709;
  assign n56711 = pi07 ? n56447 : n56710;
  assign n56712 = pi18 ? n863 : ~n21194;
  assign n56713 = pi17 ? n32 : n56712;
  assign n56714 = pi18 ? n28827 : n237;
  assign n56715 = pi17 ? n28825 : n56714;
  assign n56716 = pi16 ? n56713 : ~n56715;
  assign n56717 = pi16 ? n1594 : ~n1944;
  assign n56718 = pi15 ? n56716 : n56717;
  assign n56719 = pi14 ? n56718 : n19831;
  assign n56720 = pi18 ? n5657 : n9012;
  assign n56721 = pi19 ? n267 : ~n207;
  assign n56722 = pi18 ? n56721 : n1942;
  assign n56723 = pi17 ? n56720 : n56722;
  assign n56724 = pi16 ? n1214 : ~n56723;
  assign n56725 = pi15 ? n19711 : n56724;
  assign n56726 = pi17 ? n16982 : ~n42286;
  assign n56727 = pi16 ? n29318 : ~n56726;
  assign n56728 = pi15 ? n43787 : n56727;
  assign n56729 = pi14 ? n56725 : n56728;
  assign n56730 = pi13 ? n56719 : n56729;
  assign n56731 = pi12 ? n32 : n56730;
  assign n56732 = pi21 ? n8275 : ~n174;
  assign n56733 = pi20 ? n32 : n56732;
  assign n56734 = pi19 ? n32 : n56733;
  assign n56735 = pi18 ? n56734 : ~n28478;
  assign n56736 = pi17 ? n32 : n56735;
  assign n56737 = pi19 ? n28483 : n41508;
  assign n56738 = pi18 ? n28482 : n56737;
  assign n56739 = pi18 ? n43087 : ~n237;
  assign n56740 = pi17 ? n56738 : ~n56739;
  assign n56741 = pi16 ? n56736 : ~n56740;
  assign n56742 = pi15 ? n56741 : n28858;
  assign n56743 = pi20 ? n18253 : ~n6822;
  assign n56744 = pi19 ? n448 : ~n56743;
  assign n56745 = pi18 ? n858 : n56744;
  assign n56746 = pi17 ? n32 : n56745;
  assign n56747 = pi19 ? n56578 : n18783;
  assign n56748 = pi19 ? n56224 : n30571;
  assign n56749 = pi18 ? n56747 : n56748;
  assign n56750 = pi18 ? n42004 : n54;
  assign n56751 = pi17 ? n56749 : n56750;
  assign n56752 = pi16 ? n56746 : n56751;
  assign n56753 = pi15 ? n56752 : n32;
  assign n56754 = pi14 ? n56742 : n56753;
  assign n56755 = pi15 ? n19172 : n18381;
  assign n56756 = pi14 ? n32 : n56755;
  assign n56757 = pi13 ? n56754 : n56756;
  assign n56758 = pi15 ? n18420 : n19166;
  assign n56759 = pi14 ? n18401 : n56758;
  assign n56760 = pi18 ? n6059 : n38;
  assign n56761 = pi17 ? n18929 : n56760;
  assign n56762 = pi16 ? n32 : n56761;
  assign n56763 = pi19 ? n49001 : ~n32;
  assign n56764 = pi18 ? n42037 : ~n56763;
  assign n56765 = pi17 ? n42045 : ~n56764;
  assign n56766 = pi16 ? n42044 : ~n56765;
  assign n56767 = pi15 ? n56762 : n56766;
  assign n56768 = pi21 ? n7410 : ~n32;
  assign n56769 = pi20 ? n56768 : ~n32;
  assign n56770 = pi19 ? n56769 : ~n32;
  assign n56771 = pi18 ? n32 : n56770;
  assign n56772 = pi17 ? n42056 : ~n56771;
  assign n56773 = pi16 ? n32 : n56772;
  assign n56774 = pi15 ? n42053 : n56773;
  assign n56775 = pi14 ? n56767 : n56774;
  assign n56776 = pi13 ? n56759 : n56775;
  assign n56777 = pi12 ? n56757 : n56776;
  assign n56778 = pi11 ? n56731 : n56777;
  assign n56779 = pi18 ? n248 : n56770;
  assign n56780 = pi17 ? n42067 : ~n56779;
  assign n56781 = pi16 ? n32 : n56780;
  assign n56782 = pi15 ? n56781 : n42217;
  assign n56783 = pi18 ? n42081 : n3350;
  assign n56784 = pi17 ? n17119 : ~n56783;
  assign n56785 = pi16 ? n32 : n56784;
  assign n56786 = pi15 ? n56785 : n18008;
  assign n56787 = pi14 ? n56782 : n56786;
  assign n56788 = pi13 ? n56787 : n28932;
  assign n56789 = pi15 ? n17891 : n18008;
  assign n56790 = pi17 ? n32 : n28407;
  assign n56791 = pi16 ? n32 : n56790;
  assign n56792 = pi15 ? n32 : n56791;
  assign n56793 = pi14 ? n56789 : n56792;
  assign n56794 = pi18 ? n940 : n1676;
  assign n56795 = pi17 ? n32 : n56794;
  assign n56796 = pi16 ? n1135 : ~n56795;
  assign n56797 = pi18 ? n209 : n1676;
  assign n56798 = pi17 ? n32 : n56797;
  assign n56799 = pi16 ? n1233 : ~n56798;
  assign n56800 = pi15 ? n56796 : n56799;
  assign n56801 = pi15 ? n29519 : n30025;
  assign n56802 = pi14 ? n56800 : n56801;
  assign n56803 = pi13 ? n56793 : n56802;
  assign n56804 = pi12 ? n56788 : n56803;
  assign n56805 = pi16 ? n1233 : ~n43707;
  assign n56806 = pi17 ? n32 : n4520;
  assign n56807 = pi16 ? n1233 : ~n56806;
  assign n56808 = pi15 ? n56805 : n56807;
  assign n56809 = pi16 ? n41062 : ~n1471;
  assign n56810 = pi19 ? n18084 : n28578;
  assign n56811 = pi18 ? n41200 : ~n56810;
  assign n56812 = pi17 ? n32 : n56811;
  assign n56813 = pi19 ? n45789 : ~n32;
  assign n56814 = pi19 ? n6398 : ~n48495;
  assign n56815 = pi18 ? n56813 : ~n56814;
  assign n56816 = pi19 ? n50852 : ~n594;
  assign n56817 = pi18 ? n56816 : n32;
  assign n56818 = pi17 ? n56815 : n56817;
  assign n56819 = pi16 ? n56812 : n56818;
  assign n56820 = pi15 ? n56809 : n56819;
  assign n56821 = pi14 ? n56808 : n56820;
  assign n56822 = pi19 ? n32 : ~n24763;
  assign n56823 = pi18 ? n56822 : ~n32;
  assign n56824 = pi17 ? n32 : n56823;
  assign n56825 = pi16 ? n28949 : ~n56824;
  assign n56826 = pi15 ? n43526 : n56825;
  assign n56827 = pi14 ? n56826 : n18461;
  assign n56828 = pi13 ? n56821 : n56827;
  assign n56829 = pi19 ? n18496 : n342;
  assign n56830 = pi18 ? n222 : ~n56829;
  assign n56831 = pi17 ? n32 : n56830;
  assign n56832 = pi16 ? n56831 : ~n18508;
  assign n56833 = pi15 ? n18495 : n56832;
  assign n56834 = pi18 ? n1012 : n5657;
  assign n56835 = pi17 ? n32 : n56834;
  assign n56836 = pi16 ? n56835 : n28275;
  assign n56837 = pi15 ? n1015 : n56836;
  assign n56838 = pi14 ? n56833 : n56837;
  assign n56839 = pi13 ? n18486 : n56838;
  assign n56840 = pi12 ? n56828 : n56839;
  assign n56841 = pi11 ? n56804 : n56840;
  assign n56842 = pi10 ? n56778 : n56841;
  assign n56843 = pi09 ? n32 : n56842;
  assign n56844 = pi15 ? n56716 : n32185;
  assign n56845 = pi14 ? n56844 : n32185;
  assign n56846 = pi18 ? n56721 : n814;
  assign n56847 = pi17 ? n56720 : n56846;
  assign n56848 = pi16 ? n1214 : ~n56847;
  assign n56849 = pi15 ? n19711 : n56848;
  assign n56850 = pi18 ? n18520 : ~n237;
  assign n56851 = pi17 ? n18518 : ~n56850;
  assign n56852 = pi16 ? n1135 : ~n56851;
  assign n56853 = pi15 ? n56852 : n29135;
  assign n56854 = pi14 ? n56849 : n56853;
  assign n56855 = pi13 ? n56845 : n56854;
  assign n56856 = pi12 ? n32 : n56855;
  assign n56857 = pi18 ? n30697 : n41286;
  assign n56858 = pi17 ? n32 : n56857;
  assign n56859 = pi19 ? n7480 : ~n32;
  assign n56860 = pi18 ? n30335 : ~n56859;
  assign n56861 = pi17 ? n30333 : ~n56860;
  assign n56862 = pi16 ? n56858 : ~n56861;
  assign n56863 = pi18 ? n29026 : ~n18521;
  assign n56864 = pi17 ? n29025 : ~n56863;
  assign n56865 = pi16 ? n29019 : n56864;
  assign n56866 = pi15 ? n56862 : n56865;
  assign n56867 = pi19 ? n357 : n32344;
  assign n56868 = pi18 ? n32 : n56867;
  assign n56869 = pi17 ? n32 : n56868;
  assign n56870 = pi19 ? n4491 : n357;
  assign n56871 = pi18 ? n56870 : n358;
  assign n56872 = pi17 ? n56871 : n18533;
  assign n56873 = pi16 ? n56869 : n56872;
  assign n56874 = pi15 ? n56873 : n57;
  assign n56875 = pi14 ? n56866 : n56874;
  assign n56876 = pi15 ? n19172 : n18545;
  assign n56877 = pi14 ? n29050 : n56876;
  assign n56878 = pi13 ? n56875 : n56877;
  assign n56879 = pi15 ? n18582 : n19166;
  assign n56880 = pi14 ? n18565 : n56879;
  assign n56881 = pi16 ? n32 : n42498;
  assign n56882 = pi18 ? n42037 : ~n1942;
  assign n56883 = pi17 ? n42045 : ~n56882;
  assign n56884 = pi16 ? n42193 : ~n56883;
  assign n56885 = pi15 ? n56881 : n56884;
  assign n56886 = pi14 ? n56885 : n42205;
  assign n56887 = pi13 ? n56880 : n56886;
  assign n56888 = pi12 ? n56878 : n56887;
  assign n56889 = pi11 ? n56856 : n56888;
  assign n56890 = pi18 ? n42076 : n237;
  assign n56891 = pi17 ? n42073 : ~n56890;
  assign n56892 = pi16 ? n32 : n56891;
  assign n56893 = pi15 ? n42214 : n56892;
  assign n56894 = pi18 ? n42081 : n237;
  assign n56895 = pi17 ? n17119 : ~n56894;
  assign n56896 = pi16 ? n32 : n56895;
  assign n56897 = pi15 ? n56896 : n18008;
  assign n56898 = pi14 ? n56893 : n56897;
  assign n56899 = pi15 ? n17903 : n18142;
  assign n56900 = pi14 ? n29079 : n56899;
  assign n56901 = pi13 ? n56898 : n56900;
  assign n56902 = pi15 ? n17903 : n18008;
  assign n56903 = pi14 ? n56902 : n56792;
  assign n56904 = pi18 ? n940 : n618;
  assign n56905 = pi17 ? n32 : n56904;
  assign n56906 = pi16 ? n1233 : ~n56905;
  assign n56907 = pi18 ? n209 : n618;
  assign n56908 = pi17 ? n32 : n56907;
  assign n56909 = pi16 ? n1135 : ~n56908;
  assign n56910 = pi15 ? n56906 : n56909;
  assign n56911 = pi18 ? n863 : n1676;
  assign n56912 = pi17 ? n32 : n56911;
  assign n56913 = pi16 ? n1135 : ~n56912;
  assign n56914 = pi15 ? n56796 : n56913;
  assign n56915 = pi14 ? n56910 : n56914;
  assign n56916 = pi13 ? n56903 : n56915;
  assign n56917 = pi12 ? n56901 : n56916;
  assign n56918 = pi16 ? n1135 : ~n56806;
  assign n56919 = pi15 ? n43708 : n56918;
  assign n56920 = pi16 ? n41208 : ~n1471;
  assign n56921 = pi18 ? n341 : ~n9578;
  assign n56922 = pi17 ? n32 : n56921;
  assign n56923 = pi16 ? n56922 : ~n1834;
  assign n56924 = pi15 ? n56920 : n56923;
  assign n56925 = pi14 ? n56919 : n56924;
  assign n56926 = pi13 ? n56925 : n56827;
  assign n56927 = pi16 ? n1014 : n17855;
  assign n56928 = pi16 ? n56835 : n17706;
  assign n56929 = pi15 ? n56927 : n56928;
  assign n56930 = pi14 ? n56833 : n56929;
  assign n56931 = pi13 ? n18635 : n56930;
  assign n56932 = pi12 ? n56926 : n56931;
  assign n56933 = pi11 ? n56917 : n56932;
  assign n56934 = pi10 ? n56889 : n56933;
  assign n56935 = pi09 ? n32 : n56934;
  assign n56936 = pi08 ? n56843 : n56935;
  assign n56937 = pi19 ? n18129 : ~n18778;
  assign n56938 = pi18 ? n863 : ~n56937;
  assign n56939 = pi17 ? n32 : n56938;
  assign n56940 = pi19 ? n18782 : n358;
  assign n56941 = pi18 ? n56940 : n32;
  assign n56942 = pi18 ? n28876 : n1813;
  assign n56943 = pi17 ? n56941 : n56942;
  assign n56944 = pi16 ? n56939 : ~n56943;
  assign n56945 = pi15 ? n56944 : n18798;
  assign n56946 = pi15 ? n44993 : n32185;
  assign n56947 = pi14 ? n56945 : n56946;
  assign n56948 = pi16 ? n1233 : ~n42601;
  assign n56949 = pi15 ? n56948 : n44537;
  assign n56950 = pi18 ? n18647 : n237;
  assign n56951 = pi17 ? n18646 : n56950;
  assign n56952 = pi16 ? n1233 : ~n56951;
  assign n56953 = pi16 ? n29318 : ~n1815;
  assign n56954 = pi15 ? n56952 : n56953;
  assign n56955 = pi14 ? n56949 : n56954;
  assign n56956 = pi13 ? n56947 : n56955;
  assign n56957 = pi12 ? n32 : n56956;
  assign n56958 = pi18 ? n6145 : n1813;
  assign n56959 = pi17 ? n13946 : n56958;
  assign n56960 = pi16 ? n1471 : ~n56959;
  assign n56961 = pi15 ? n45734 : n56960;
  assign n56962 = pi14 ? n56961 : n18663;
  assign n56963 = pi18 ? n18668 : ~n814;
  assign n56964 = pi17 ? n18667 : n56963;
  assign n56965 = pi16 ? n32 : n56964;
  assign n56966 = pi15 ? n56965 : n18672;
  assign n56967 = pi14 ? n32 : n56966;
  assign n56968 = pi13 ? n56962 : n56967;
  assign n56969 = pi14 ? n18683 : n19333;
  assign n56970 = pi18 ? n42297 : n814;
  assign n56971 = pi17 ? n42294 : ~n56970;
  assign n56972 = pi16 ? n32 : n56971;
  assign n56973 = pi15 ? n42288 : n56972;
  assign n56974 = pi19 ? n10447 : ~n32;
  assign n56975 = pi18 ? n42310 : n56974;
  assign n56976 = pi17 ? n17346 : ~n56975;
  assign n56977 = pi16 ? n32 : n56976;
  assign n56978 = pi15 ? n42309 : n56977;
  assign n56979 = pi14 ? n56973 : n56978;
  assign n56980 = pi13 ? n56969 : n56979;
  assign n56981 = pi12 ? n56968 : n56980;
  assign n56982 = pi11 ? n56957 : n56981;
  assign n56983 = pi18 ? n42319 : n56974;
  assign n56984 = pi17 ? n23052 : ~n56983;
  assign n56985 = pi16 ? n32 : n56984;
  assign n56986 = pi18 ? n13182 : n237;
  assign n56987 = pi17 ? n23052 : ~n56986;
  assign n56988 = pi16 ? n32 : n56987;
  assign n56989 = pi15 ? n56985 : n56988;
  assign n56990 = pi15 ? n42428 : n18142;
  assign n56991 = pi14 ? n56989 : n56990;
  assign n56992 = pi15 ? n18439 : n18142;
  assign n56993 = pi14 ? n18594 : n56992;
  assign n56994 = pi13 ? n56991 : n56993;
  assign n56995 = pi15 ? n17637 : n29780;
  assign n56996 = pi14 ? n17885 : n56995;
  assign n56997 = pi16 ? n1135 : ~n56905;
  assign n56998 = pi15 ? n56997 : n56909;
  assign n56999 = pi15 ? n29676 : n28947;
  assign n57000 = pi14 ? n56998 : n56999;
  assign n57001 = pi13 ? n56996 : n57000;
  assign n57002 = pi12 ? n56994 : n57001;
  assign n57003 = pi20 ? n32 : n18245;
  assign n57004 = pi19 ? n32 : n57003;
  assign n57005 = pi20 ? n6050 : ~n9488;
  assign n57006 = pi19 ? n47656 : ~n57005;
  assign n57007 = pi18 ? n57004 : ~n57006;
  assign n57008 = pi17 ? n32 : n57007;
  assign n57009 = pi19 ? n29918 : n17974;
  assign n57010 = pi19 ? n2250 : n275;
  assign n57011 = pi18 ? n57009 : n57010;
  assign n57012 = pi19 ? n1818 : n322;
  assign n57013 = pi18 ? n57012 : n1676;
  assign n57014 = pi17 ? n57011 : n57013;
  assign n57015 = pi16 ? n57008 : ~n57014;
  assign n57016 = pi18 ? n4519 : n1676;
  assign n57017 = pi17 ? n32 : n57016;
  assign n57018 = pi16 ? n1233 : ~n57017;
  assign n57019 = pi15 ? n57015 : n57018;
  assign n57020 = pi15 ? n43577 : n43574;
  assign n57021 = pi14 ? n57019 : n57020;
  assign n57022 = pi15 ? n41122 : n17915;
  assign n57023 = pi14 ? n57022 : n18707;
  assign n57024 = pi13 ? n57021 : n57023;
  assign n57025 = pi20 ? n785 : n1324;
  assign n57026 = pi19 ? n44193 : ~n57025;
  assign n57027 = pi18 ? n47982 : n57026;
  assign n57028 = pi17 ? n32 : n57027;
  assign n57029 = pi20 ? n32 : ~n2385;
  assign n57030 = pi19 ? n29297 : ~n57029;
  assign n57031 = pi18 ? n57030 : ~n32;
  assign n57032 = pi17 ? n29296 : n57031;
  assign n57033 = pi16 ? n57028 : ~n57032;
  assign n57034 = pi15 ? n18740 : n57033;
  assign n57035 = pi18 ? n1012 : n20164;
  assign n57036 = pi17 ? n32 : n57035;
  assign n57037 = pi16 ? n57036 : n17855;
  assign n57038 = pi15 ? n1015 : n57037;
  assign n57039 = pi14 ? n57034 : n57038;
  assign n57040 = pi13 ? n18736 : n57039;
  assign n57041 = pi12 ? n57024 : n57040;
  assign n57042 = pi11 ? n57002 : n57041;
  assign n57043 = pi10 ? n56982 : n57042;
  assign n57044 = pi09 ? n32 : n57043;
  assign n57045 = pi15 ? n29601 : n29729;
  assign n57046 = pi15 ? n44993 : n20034;
  assign n57047 = pi14 ? n57045 : n57046;
  assign n57048 = pi17 ? n32 : n2314;
  assign n57049 = pi16 ? n1135 : ~n57048;
  assign n57050 = pi18 ? n341 : n18753;
  assign n57051 = pi17 ? n32 : n57050;
  assign n57052 = pi18 ? n18764 : ~n30435;
  assign n57053 = pi17 ? n18760 : ~n57052;
  assign n57054 = pi16 ? n57051 : ~n57053;
  assign n57055 = pi15 ? n57049 : n57054;
  assign n57056 = pi19 ? n41311 : n1464;
  assign n57057 = pi18 ? n6071 : n57056;
  assign n57058 = pi19 ? n6171 : n274;
  assign n57059 = pi18 ? n57058 : n814;
  assign n57060 = pi17 ? n57057 : n57059;
  assign n57061 = pi16 ? n1135 : ~n57060;
  assign n57062 = pi16 ? n29318 : ~n1808;
  assign n57063 = pi15 ? n57061 : n57062;
  assign n57064 = pi14 ? n57055 : n57063;
  assign n57065 = pi13 ? n57047 : n57064;
  assign n57066 = pi12 ? n42387 : n57065;
  assign n57067 = pi15 ? n57062 : n29328;
  assign n57068 = pi14 ? n57067 : n18663;
  assign n57069 = pi18 ? n18790 : ~n814;
  assign n57070 = pi17 ? n18788 : n57069;
  assign n57071 = pi16 ? n18781 : n57070;
  assign n57072 = pi15 ? n57071 : n18794;
  assign n57073 = pi14 ? n32 : n57072;
  assign n57074 = pi13 ? n57068 : n57073;
  assign n57075 = pi14 ? n18800 : n19333;
  assign n57076 = pi17 ? n42411 : ~n56970;
  assign n57077 = pi16 ? n32 : n57076;
  assign n57078 = pi15 ? n42408 : n57077;
  assign n57079 = pi14 ? n57078 : n42421;
  assign n57080 = pi13 ? n57075 : n57079;
  assign n57081 = pi12 ? n57074 : n57080;
  assign n57082 = pi11 ? n57066 : n57081;
  assign n57083 = pi18 ? n13182 : n1942;
  assign n57084 = pi17 ? n23052 : ~n57083;
  assign n57085 = pi16 ? n32 : n57084;
  assign n57086 = pi15 ? n42322 : n57085;
  assign n57087 = pi14 ? n57086 : n42429;
  assign n57088 = pi15 ? n18439 : n18294;
  assign n57089 = pi14 ? n18814 : n57088;
  assign n57090 = pi13 ? n57087 : n57089;
  assign n57091 = pi15 ? n17637 : n29875;
  assign n57092 = pi14 ? n17885 : n57091;
  assign n57093 = pi18 ? n940 : ~n18076;
  assign n57094 = pi17 ? n32 : n57093;
  assign n57095 = pi16 ? n1233 : ~n57094;
  assign n57096 = pi15 ? n57095 : n29875;
  assign n57097 = pi15 ? n56906 : n28947;
  assign n57098 = pi14 ? n57096 : n57097;
  assign n57099 = pi13 ? n57092 : n57098;
  assign n57100 = pi12 ? n57090 : n57099;
  assign n57101 = pi17 ? n32 : n57013;
  assign n57102 = pi16 ? n1135 : ~n57101;
  assign n57103 = pi16 ? n1135 : ~n56383;
  assign n57104 = pi15 ? n57102 : n57103;
  assign n57105 = pi14 ? n57104 : n43574;
  assign n57106 = pi15 ? n41122 : n17825;
  assign n57107 = pi14 ? n57106 : n18853;
  assign n57108 = pi13 ? n57105 : n57107;
  assign n57109 = pi20 ? n5854 : ~n9491;
  assign n57110 = pi19 ? n57109 : ~n57025;
  assign n57111 = pi18 ? n47982 : n57110;
  assign n57112 = pi17 ? n32 : n57111;
  assign n57113 = pi20 ? n5854 : ~n831;
  assign n57114 = pi20 ? n32 : ~n9361;
  assign n57115 = pi19 ? n57113 : ~n57114;
  assign n57116 = pi18 ? n57115 : ~n32;
  assign n57117 = pi17 ? n29396 : n57116;
  assign n57118 = pi16 ? n57112 : ~n57117;
  assign n57119 = pi15 ? n18859 : n57118;
  assign n57120 = pi19 ? n32 : n472;
  assign n57121 = pi18 ? n57120 : n32;
  assign n57122 = pi17 ? n32 : n57121;
  assign n57123 = pi16 ? n1014 : n57122;
  assign n57124 = pi15 ? n57123 : n57037;
  assign n57125 = pi14 ? n57119 : n57124;
  assign n57126 = pi13 ? n18736 : n57125;
  assign n57127 = pi12 ? n57108 : n57126;
  assign n57128 = pi11 ? n57100 : n57127;
  assign n57129 = pi10 ? n57082 : n57128;
  assign n57130 = pi09 ? n32 : n57129;
  assign n57131 = pi08 ? n57044 : n57130;
  assign n57132 = pi07 ? n56936 : n57131;
  assign n57133 = pi06 ? n56711 : n57132;
  assign n57134 = pi05 ? n56211 : n57133;
  assign n57135 = pi04 ? n32 : n57134;
  assign n57136 = pi14 ? n34363 : n32;
  assign n57137 = pi20 ? n1611 : n1331;
  assign n57138 = pi19 ? n28370 : n57137;
  assign n57139 = pi18 ? n863 : n57138;
  assign n57140 = pi17 ? n32 : n57139;
  assign n57141 = pi19 ? n18106 : ~n24055;
  assign n57142 = pi19 ? n23346 : ~n35996;
  assign n57143 = pi18 ? n57141 : n57142;
  assign n57144 = pi19 ? n29270 : n47731;
  assign n57145 = pi18 ? n57144 : n350;
  assign n57146 = pi17 ? n57143 : n57145;
  assign n57147 = pi16 ? n57140 : ~n57146;
  assign n57148 = pi15 ? n32 : n57147;
  assign n57149 = pi14 ? n18906 : n57148;
  assign n57150 = pi13 ? n57136 : n57149;
  assign n57151 = pi14 ? n29601 : n44537;
  assign n57152 = pi20 ? n16168 : ~n32;
  assign n57153 = pi19 ? n57152 : ~n32;
  assign n57154 = pi18 ? n32 : n57153;
  assign n57155 = pi17 ? n32 : n57154;
  assign n57156 = pi16 ? n1233 : ~n57155;
  assign n57157 = pi18 ? n366 : n18882;
  assign n57158 = pi17 ? n32 : n57157;
  assign n57159 = pi16 ? n57158 : n32;
  assign n57160 = pi15 ? n57156 : n57159;
  assign n57161 = pi15 ? n32185 : n29845;
  assign n57162 = pi14 ? n57160 : n57161;
  assign n57163 = pi13 ? n57151 : n57162;
  assign n57164 = pi12 ? n57150 : n57163;
  assign n57165 = pi15 ? n29845 : n19531;
  assign n57166 = pi14 ? n57165 : n18906;
  assign n57167 = pi18 ? n18920 : ~n822;
  assign n57168 = pi17 ? n18917 : ~n57167;
  assign n57169 = pi16 ? n18913 : ~n57168;
  assign n57170 = pi15 ? n57169 : n18932;
  assign n57171 = pi14 ? n19333 : n57170;
  assign n57172 = pi13 ? n57166 : n57171;
  assign n57173 = pi18 ? n9012 : n1813;
  assign n57174 = pi17 ? n1124 : n57173;
  assign n57175 = pi16 ? n18938 : ~n57174;
  assign n57176 = pi18 ? n42514 : ~n237;
  assign n57177 = pi17 ? n42513 : n57176;
  assign n57178 = pi16 ? n32 : n57177;
  assign n57179 = pi15 ? n57175 : n57178;
  assign n57180 = pi20 ? n785 : n357;
  assign n57181 = pi19 ? n57180 : n29473;
  assign n57182 = pi18 ? n17058 : ~n57181;
  assign n57183 = pi18 ? n29478 : n32;
  assign n57184 = pi17 ? n57182 : n57183;
  assign n57185 = pi16 ? n32 : n57184;
  assign n57186 = pi15 ? n57185 : n18531;
  assign n57187 = pi14 ? n57179 : n57186;
  assign n57188 = pi18 ? n42536 : n20023;
  assign n57189 = pi17 ? n32 : ~n57188;
  assign n57190 = pi16 ? n32 : n57189;
  assign n57191 = pi15 ? n42534 : n57190;
  assign n57192 = pi15 ? n19536 : n19459;
  assign n57193 = pi14 ? n57191 : n57192;
  assign n57194 = pi13 ? n57187 : n57193;
  assign n57195 = pi12 ? n57172 : n57194;
  assign n57196 = pi11 ? n57164 : n57195;
  assign n57197 = pi14 ? n42654 : n29499;
  assign n57198 = pi14 ? n29504 : n30211;
  assign n57199 = pi13 ? n57197 : n57198;
  assign n57200 = pi19 ? n322 : ~n32090;
  assign n57201 = pi18 ? n57200 : n618;
  assign n57202 = pi17 ? n32 : n57201;
  assign n57203 = pi16 ? n1214 : ~n57202;
  assign n57204 = pi18 ? n863 : n3350;
  assign n57205 = pi17 ? n32 : n57204;
  assign n57206 = pi16 ? n1135 : ~n57205;
  assign n57207 = pi15 ? n57203 : n57206;
  assign n57208 = pi14 ? n32 : n57207;
  assign n57209 = pi16 ? n1135 : ~n57094;
  assign n57210 = pi15 ? n57209 : n29676;
  assign n57211 = pi18 ? n43221 : ~n28876;
  assign n57212 = pi17 ? n32 : n57211;
  assign n57213 = pi19 ? n4491 : n43029;
  assign n57214 = pi18 ? n57213 : n19232;
  assign n57215 = pi17 ? n57214 : n3380;
  assign n57216 = pi16 ? n57212 : ~n57215;
  assign n57217 = pi16 ? n1233 : ~n41489;
  assign n57218 = pi15 ? n57216 : n57217;
  assign n57219 = pi14 ? n57210 : n57218;
  assign n57220 = pi13 ? n57208 : n57219;
  assign n57221 = pi12 ? n57199 : n57220;
  assign n57222 = pi18 ? n940 : ~n17994;
  assign n57223 = pi17 ? n32 : n57222;
  assign n57224 = pi16 ? n1233 : ~n57223;
  assign n57225 = pi15 ? n57224 : n56330;
  assign n57226 = pi18 ? n323 : n32;
  assign n57227 = pi17 ? n32 : n57226;
  assign n57228 = pi16 ? n32 : n57227;
  assign n57229 = pi15 ? n19100 : n57228;
  assign n57230 = pi14 ? n57225 : n57229;
  assign n57231 = pi18 ? n42558 : n32;
  assign n57232 = pi17 ? n32 : n57231;
  assign n57233 = pi16 ? n32 : n57232;
  assign n57234 = pi15 ? n57233 : n18977;
  assign n57235 = pi16 ? n18981 : ~n1577;
  assign n57236 = pi15 ? n18979 : n57235;
  assign n57237 = pi14 ? n57234 : n57236;
  assign n57238 = pi13 ? n57230 : n57237;
  assign n57239 = pi16 ? n18991 : ~n1577;
  assign n57240 = pi15 ? n57239 : n18995;
  assign n57241 = pi14 ? n57240 : n19005;
  assign n57242 = pi20 ? n266 : n11107;
  assign n57243 = pi19 ? n507 : n57242;
  assign n57244 = pi18 ? n57243 : ~n32;
  assign n57245 = pi17 ? n32 : n57244;
  assign n57246 = pi16 ? n1135 : ~n57245;
  assign n57247 = pi15 ? n57246 : n33585;
  assign n57248 = pi18 ? n127 : n16449;
  assign n57249 = pi17 ? n32 : n57248;
  assign n57250 = pi16 ? n57249 : n17850;
  assign n57251 = pi18 ? n4127 : ~n32;
  assign n57252 = pi17 ? n32 : n57251;
  assign n57253 = pi16 ? n1233 : ~n57252;
  assign n57254 = pi15 ? n57250 : n57253;
  assign n57255 = pi14 ? n57247 : n57254;
  assign n57256 = pi13 ? n57241 : n57255;
  assign n57257 = pi12 ? n57238 : n57256;
  assign n57258 = pi11 ? n57221 : n57257;
  assign n57259 = pi10 ? n57196 : n57258;
  assign n57260 = pi09 ? n32 : n57259;
  assign n57261 = pi15 ? n18904 : n19628;
  assign n57262 = pi14 ? n57261 : n32;
  assign n57263 = pi20 ? n820 : n18245;
  assign n57264 = pi19 ? n57263 : ~n41325;
  assign n57265 = pi18 ? n1862 : n57264;
  assign n57266 = pi17 ? n32 : n57265;
  assign n57267 = pi20 ? n18129 : ~n18173;
  assign n57268 = pi20 ? n339 : n18245;
  assign n57269 = pi19 ? n57267 : ~n57268;
  assign n57270 = pi20 ? n18245 : ~n428;
  assign n57271 = pi19 ? n43838 : ~n57270;
  assign n57272 = pi18 ? n57269 : n57271;
  assign n57273 = pi18 ? n42564 : n3336;
  assign n57274 = pi17 ? n57272 : n57273;
  assign n57275 = pi16 ? n57266 : ~n57274;
  assign n57276 = pi15 ? n32 : n57275;
  assign n57277 = pi14 ? n18906 : n57276;
  assign n57278 = pi13 ? n57262 : n57277;
  assign n57279 = pi16 ? n1135 : ~n3338;
  assign n57280 = pi14 ? n57279 : n30941;
  assign n57281 = pi17 ? n32 : n43016;
  assign n57282 = pi16 ? n1135 : ~n57281;
  assign n57283 = pi18 ? n341 : n18882;
  assign n57284 = pi17 ? n32 : n57283;
  assign n57285 = pi16 ? n57284 : n32;
  assign n57286 = pi15 ? n57282 : n57285;
  assign n57287 = pi15 ? n29601 : n29845;
  assign n57288 = pi14 ? n57286 : n57287;
  assign n57289 = pi13 ? n57280 : n57288;
  assign n57290 = pi12 ? n57278 : n57289;
  assign n57291 = pi21 ? n9326 : n32;
  assign n57292 = pi20 ? n57291 : n32;
  assign n57293 = pi19 ? n57292 : n32;
  assign n57294 = pi18 ? n32 : n57293;
  assign n57295 = pi17 ? n32 : n57294;
  assign n57296 = pi16 ? n32 : n57295;
  assign n57297 = pi15 ? n29845 : n57296;
  assign n57298 = pi14 ? n57297 : n19032;
  assign n57299 = pi15 ? n18661 : n18805;
  assign n57300 = pi16 ? n19037 : ~n57168;
  assign n57301 = pi15 ? n57300 : n19041;
  assign n57302 = pi14 ? n57299 : n57301;
  assign n57303 = pi13 ? n57298 : n57302;
  assign n57304 = pi16 ? n19048 : ~n57174;
  assign n57305 = pi15 ? n57304 : n57178;
  assign n57306 = pi18 ? n17118 : ~n57181;
  assign n57307 = pi17 ? n57306 : n57183;
  assign n57308 = pi16 ? n32 : n57307;
  assign n57309 = pi15 ? n57308 : n18531;
  assign n57310 = pi14 ? n57305 : n57309;
  assign n57311 = pi18 ? n42641 : n20023;
  assign n57312 = pi17 ? n32 : ~n57311;
  assign n57313 = pi16 ? n32 : n57312;
  assign n57314 = pi15 ? n42639 : n57313;
  assign n57315 = pi15 ? n18814 : n19459;
  assign n57316 = pi14 ? n57314 : n57315;
  assign n57317 = pi13 ? n57310 : n57316;
  assign n57318 = pi12 ? n57303 : n57317;
  assign n57319 = pi11 ? n57290 : n57318;
  assign n57320 = pi18 ? n11884 : n814;
  assign n57321 = pi17 ? n32 : ~n57320;
  assign n57322 = pi16 ? n32 : n57321;
  assign n57323 = pi18 ? n936 : ~n814;
  assign n57324 = pi17 ? n32 : n57323;
  assign n57325 = pi16 ? n32 : n57324;
  assign n57326 = pi15 ? n57322 : n57325;
  assign n57327 = pi14 ? n57326 : n29647;
  assign n57328 = pi18 ? n32 : ~n56974;
  assign n57329 = pi17 ? n32 : n57328;
  assign n57330 = pi16 ? n32 : n57329;
  assign n57331 = pi15 ? n32 : n57330;
  assign n57332 = pi14 ? n29652 : n57331;
  assign n57333 = pi13 ? n57327 : n57332;
  assign n57334 = pi18 ? n57200 : ~n32;
  assign n57335 = pi17 ? n32 : n57334;
  assign n57336 = pi16 ? n1214 : ~n57335;
  assign n57337 = pi19 ? n40268 : ~n32;
  assign n57338 = pi18 ? n863 : n57337;
  assign n57339 = pi17 ? n32 : n57338;
  assign n57340 = pi16 ? n1233 : ~n57339;
  assign n57341 = pi15 ? n57336 : n57340;
  assign n57342 = pi14 ? n17997 : n57341;
  assign n57343 = pi18 ? n940 : ~n359;
  assign n57344 = pi17 ? n32 : n57343;
  assign n57345 = pi16 ? n1233 : ~n57344;
  assign n57346 = pi18 ? n751 : ~n18076;
  assign n57347 = pi17 ? n32 : n57346;
  assign n57348 = pi16 ? n1233 : ~n57347;
  assign n57349 = pi15 ? n57345 : n57348;
  assign n57350 = pi16 ? n1135 : ~n41489;
  assign n57351 = pi15 ? n57095 : n57350;
  assign n57352 = pi14 ? n57349 : n57351;
  assign n57353 = pi13 ? n57342 : n57352;
  assign n57354 = pi12 ? n57333 : n57353;
  assign n57355 = pi16 ? n1135 : ~n1678;
  assign n57356 = pi15 ? n56997 : n57355;
  assign n57357 = pi15 ? n18979 : n57228;
  assign n57358 = pi14 ? n57356 : n57357;
  assign n57359 = pi15 ? n57233 : n19098;
  assign n57360 = pi15 ? n19100 : n57235;
  assign n57361 = pi14 ? n57359 : n57360;
  assign n57362 = pi13 ? n57358 : n57361;
  assign n57363 = pi16 ? n18991 : ~n1834;
  assign n57364 = pi15 ? n57363 : n18995;
  assign n57365 = pi14 ? n57364 : n19005;
  assign n57366 = pi20 ? n274 : n11107;
  assign n57367 = pi19 ? n507 : n57366;
  assign n57368 = pi18 ? n57367 : ~n32;
  assign n57369 = pi17 ? n32 : n57368;
  assign n57370 = pi16 ? n1135 : ~n57369;
  assign n57371 = pi18 ? n10058 : ~n32;
  assign n57372 = pi17 ? n32 : n57371;
  assign n57373 = pi16 ? n1135 : ~n57372;
  assign n57374 = pi15 ? n57370 : n57373;
  assign n57375 = pi14 ? n57374 : n57254;
  assign n57376 = pi13 ? n57365 : n57375;
  assign n57377 = pi12 ? n57362 : n57376;
  assign n57378 = pi11 ? n57354 : n57377;
  assign n57379 = pi10 ? n57319 : n57378;
  assign n57380 = pi09 ? n32 : n57379;
  assign n57381 = pi08 ? n57260 : n57380;
  assign n57382 = pi15 ? n19235 : n19628;
  assign n57383 = pi14 ? n57382 : n32;
  assign n57384 = pi15 ? n32 : n32806;
  assign n57385 = pi14 ? n20746 : n57384;
  assign n57386 = pi13 ? n57383 : n57385;
  assign n57387 = pi15 ? n29601 : n32806;
  assign n57388 = pi14 ? n32806 : n57387;
  assign n57389 = pi19 ? n7014 : ~n32;
  assign n57390 = pi18 ? n32 : n57389;
  assign n57391 = pi17 ? n32 : n57390;
  assign n57392 = pi16 ? n1233 : ~n57391;
  assign n57393 = pi15 ? n57392 : n31146;
  assign n57394 = pi16 ? n1471 : ~n2540;
  assign n57395 = pi15 ? n29601 : n57394;
  assign n57396 = pi14 ? n57393 : n57395;
  assign n57397 = pi13 ? n57388 : n57396;
  assign n57398 = pi12 ? n57386 : n57397;
  assign n57399 = pi20 ? n9488 : n29452;
  assign n57400 = pi19 ? n29458 : n57399;
  assign n57401 = pi20 ? n1324 : n6822;
  assign n57402 = pi20 ? n29452 : ~n17669;
  assign n57403 = pi19 ? n57401 : ~n57402;
  assign n57404 = pi18 ? n57400 : ~n57403;
  assign n57405 = pi19 ? n19134 : ~n18281;
  assign n57406 = pi18 ? n57405 : ~n19121;
  assign n57407 = pi17 ? n57404 : ~n57406;
  assign n57408 = pi16 ? n29738 : n57407;
  assign n57409 = pi15 ? n57408 : n19145;
  assign n57410 = pi14 ? n57409 : n19147;
  assign n57411 = pi13 ? n57410 : n19157;
  assign n57412 = pi17 ? n42761 : ~n2325;
  assign n57413 = pi16 ? n32 : n57412;
  assign n57414 = pi18 ? n42768 : n237;
  assign n57415 = pi17 ? n42765 : ~n57414;
  assign n57416 = pi16 ? n32 : n57415;
  assign n57417 = pi15 ? n57413 : n57416;
  assign n57418 = pi19 ? n857 : n448;
  assign n57419 = pi18 ? n32 : n57418;
  assign n57420 = pi20 ? n17671 : n342;
  assign n57421 = pi19 ? n28338 : n57420;
  assign n57422 = pi18 ? n57421 : n6867;
  assign n57423 = pi17 ? n57419 : n57422;
  assign n57424 = pi16 ? n32 : n57423;
  assign n57425 = pi15 ? n57424 : n19628;
  assign n57426 = pi14 ? n57417 : n57425;
  assign n57427 = pi18 ? n2387 : ~n350;
  assign n57428 = pi17 ? n32 : n57427;
  assign n57429 = pi16 ? n32 : n57428;
  assign n57430 = pi15 ? n42785 : n57429;
  assign n57431 = pi18 ? n2387 : ~n20023;
  assign n57432 = pi17 ? n32 : n57431;
  assign n57433 = pi16 ? n32 : n57432;
  assign n57434 = pi18 ? n42799 : ~n20023;
  assign n57435 = pi17 ? n42798 : n57434;
  assign n57436 = pi16 ? n42795 : n57435;
  assign n57437 = pi15 ? n57433 : n57436;
  assign n57438 = pi14 ? n57430 : n57437;
  assign n57439 = pi13 ? n57426 : n57438;
  assign n57440 = pi12 ? n57411 : n57439;
  assign n57441 = pi11 ? n57398 : n57440;
  assign n57442 = pi15 ? n19073 : n19166;
  assign n57443 = pi14 ? n42946 : n57442;
  assign n57444 = pi15 ? n18814 : n19166;
  assign n57445 = pi14 ? n57444 : n58;
  assign n57446 = pi13 ? n57443 : n57445;
  assign n57447 = pi18 ? n17848 : ~n32;
  assign n57448 = pi17 ? n32 : n57447;
  assign n57449 = pi16 ? n1135 : ~n57448;
  assign n57450 = pi16 ? n1135 : ~n28030;
  assign n57451 = pi15 ? n57449 : n57450;
  assign n57452 = pi14 ? n28612 : n57451;
  assign n57453 = pi18 ? n940 : ~n38;
  assign n57454 = pi17 ? n32 : n57453;
  assign n57455 = pi16 ? n1135 : ~n57454;
  assign n57456 = pi15 ? n57455 : n29676;
  assign n57457 = pi16 ? n19200 : ~n1471;
  assign n57458 = pi18 ? n863 : ~n18076;
  assign n57459 = pi17 ? n32 : n57458;
  assign n57460 = pi16 ? n1135 : ~n57459;
  assign n57461 = pi15 ? n57457 : n57460;
  assign n57462 = pi14 ? n57456 : n57461;
  assign n57463 = pi13 ? n57452 : n57462;
  assign n57464 = pi12 ? n57446 : n57463;
  assign n57465 = pi16 ? n1233 : ~n57459;
  assign n57466 = pi15 ? n57465 : n43933;
  assign n57467 = pi18 ? n702 : ~n1676;
  assign n57468 = pi17 ? n32 : n57467;
  assign n57469 = pi16 ? n32 : n57468;
  assign n57470 = pi15 ? n56330 : n57469;
  assign n57471 = pi14 ? n57466 : n57470;
  assign n57472 = pi13 ? n57471 : n19207;
  assign n57473 = pi20 ? n287 : ~n1076;
  assign n57474 = pi19 ? n18728 : ~n57473;
  assign n57475 = pi18 ? n4380 : n57474;
  assign n57476 = pi17 ? n32 : n57475;
  assign n57477 = pi20 ? n342 : n4279;
  assign n57478 = pi20 ? n5854 : ~n405;
  assign n57479 = pi19 ? n57477 : n57478;
  assign n57480 = pi20 ? n6621 : ~n310;
  assign n57481 = pi19 ? n32509 : ~n57480;
  assign n57482 = pi18 ? n57479 : ~n57481;
  assign n57483 = pi20 ? n309 : n101;
  assign n57484 = pi19 ? n29682 : n57483;
  assign n57485 = pi18 ? n57484 : ~n32;
  assign n57486 = pi17 ? n57482 : ~n57485;
  assign n57487 = pi16 ? n57476 : n57486;
  assign n57488 = pi15 ? n19217 : n57487;
  assign n57489 = pi14 ? n19214 : n57488;
  assign n57490 = pi22 ? n173 : n65;
  assign n57491 = pi21 ? n206 : ~n57490;
  assign n57492 = pi20 ? n32 : n57491;
  assign n57493 = pi19 ? n32 : n57492;
  assign n57494 = pi18 ? n57493 : ~n32;
  assign n57495 = pi17 ? n32 : n57494;
  assign n57496 = pi16 ? n42855 : ~n57495;
  assign n57497 = pi15 ? n57496 : n43373;
  assign n57498 = pi18 ? n1012 : n16234;
  assign n57499 = pi17 ? n32 : n57498;
  assign n57500 = pi16 ? n57499 : n17836;
  assign n57501 = pi16 ? n1233 : ~n2144;
  assign n57502 = pi15 ? n57500 : n57501;
  assign n57503 = pi14 ? n57497 : n57502;
  assign n57504 = pi13 ? n57489 : n57503;
  assign n57505 = pi12 ? n57472 : n57504;
  assign n57506 = pi11 ? n57464 : n57505;
  assign n57507 = pi10 ? n57441 : n57506;
  assign n57508 = pi09 ? n32 : n57507;
  assign n57509 = pi15 ? n32 : n31854;
  assign n57510 = pi14 ? n20746 : n57509;
  assign n57511 = pi13 ? n57383 : n57510;
  assign n57512 = pi15 ? n30941 : n31854;
  assign n57513 = pi14 ? n45477 : n57512;
  assign n57514 = pi18 ? n32 : n289;
  assign n57515 = pi17 ? n32 : n57514;
  assign n57516 = pi16 ? n1135 : ~n57515;
  assign n57517 = pi15 ? n57516 : n31146;
  assign n57518 = pi15 ? n57279 : n57394;
  assign n57519 = pi14 ? n57517 : n57518;
  assign n57520 = pi13 ? n57513 : n57519;
  assign n57521 = pi12 ? n57511 : n57520;
  assign n57522 = pi20 ? n18129 : n266;
  assign n57523 = pi19 ? n29618 : n57522;
  assign n57524 = pi20 ? n2358 : n18415;
  assign n57525 = pi19 ? n57524 : ~n28152;
  assign n57526 = pi18 ? n57523 : ~n57525;
  assign n57527 = pi19 ? n19249 : ~n17665;
  assign n57528 = pi18 ? n57527 : ~n19137;
  assign n57529 = pi17 ? n57526 : ~n57528;
  assign n57530 = pi16 ? n29851 : n57529;
  assign n57531 = pi15 ? n57530 : n19145;
  assign n57532 = pi14 ? n57531 : n19147;
  assign n57533 = pi13 ? n57532 : n19157;
  assign n57534 = pi17 ? n42919 : ~n2325;
  assign n57535 = pi16 ? n32 : n57534;
  assign n57536 = pi15 ? n57535 : n57416;
  assign n57537 = pi15 ? n17903 : n19628;
  assign n57538 = pi14 ? n57536 : n57537;
  assign n57539 = pi15 ? n42930 : n57429;
  assign n57540 = pi14 ? n57539 : n42938;
  assign n57541 = pi13 ? n57538 : n57540;
  assign n57542 = pi12 ? n57533 : n57541;
  assign n57543 = pi11 ? n57521 : n57542;
  assign n57544 = pi18 ? n23504 : n1813;
  assign n57545 = pi17 ? n42812 : n57544;
  assign n57546 = pi16 ? n42810 : ~n57545;
  assign n57547 = pi15 ? n57546 : n19706;
  assign n57548 = pi14 ? n57547 : n29869;
  assign n57549 = pi14 ? n29871 : n19333;
  assign n57550 = pi13 ? n57548 : n57549;
  assign n57551 = pi18 ? n32 : ~n54;
  assign n57552 = pi17 ? n32 : n57551;
  assign n57553 = pi16 ? n1135 : ~n57552;
  assign n57554 = pi18 ? n863 : n1942;
  assign n57555 = pi17 ? n32 : n57554;
  assign n57556 = pi16 ? n1135 : ~n57555;
  assign n57557 = pi15 ? n57553 : n57556;
  assign n57558 = pi14 ? n32 : n57557;
  assign n57559 = pi15 ? n29676 : n57345;
  assign n57560 = pi16 ? n19200 : ~n57344;
  assign n57561 = pi15 ? n57560 : n57460;
  assign n57562 = pi14 ? n57559 : n57561;
  assign n57563 = pi13 ? n57558 : n57562;
  assign n57564 = pi12 ? n57550 : n57563;
  assign n57565 = pi15 ? n57460 : n19349;
  assign n57566 = pi15 ? n57355 : n29902;
  assign n57567 = pi14 ? n57565 : n57566;
  assign n57568 = pi13 ? n57567 : n19290;
  assign n57569 = pi19 ? n29682 : n28565;
  assign n57570 = pi18 ? n57569 : ~n32;
  assign n57571 = pi17 ? n57482 : ~n57570;
  assign n57572 = pi16 ? n57476 : n57571;
  assign n57573 = pi15 ? n19217 : n57572;
  assign n57574 = pi14 ? n19214 : n57573;
  assign n57575 = pi21 ? n206 : ~n14158;
  assign n57576 = pi20 ? n32 : n57575;
  assign n57577 = pi19 ? n32 : n57576;
  assign n57578 = pi18 ? n57577 : ~n32;
  assign n57579 = pi17 ? n32 : n57578;
  assign n57580 = pi16 ? n42855 : ~n57579;
  assign n57581 = pi20 ? n32 : ~n67;
  assign n57582 = pi19 ? n32 : n57581;
  assign n57583 = pi18 ? n57582 : ~n32;
  assign n57584 = pi17 ? n32 : n57583;
  assign n57585 = pi16 ? n1214 : ~n57584;
  assign n57586 = pi15 ? n57580 : n57585;
  assign n57587 = pi14 ? n57586 : n57502;
  assign n57588 = pi13 ? n57574 : n57587;
  assign n57589 = pi12 ? n57568 : n57588;
  assign n57590 = pi11 ? n57564 : n57589;
  assign n57591 = pi10 ? n57543 : n57590;
  assign n57592 = pi09 ? n32 : n57591;
  assign n57593 = pi08 ? n57508 : n57592;
  assign n57594 = pi07 ? n57381 : n57593;
  assign n57595 = pi14 ? n19621 : n32;
  assign n57596 = pi16 ? n1233 : ~n2540;
  assign n57597 = pi15 ? n29601 : n57596;
  assign n57598 = pi14 ? n42986 : n57597;
  assign n57599 = pi13 ? n57595 : n57598;
  assign n57600 = pi15 ? n57596 : n29601;
  assign n57601 = pi15 ? n31146 : n31856;
  assign n57602 = pi14 ? n57600 : n57601;
  assign n57603 = pi15 ? n31854 : n31146;
  assign n57604 = pi19 ? n311 : ~n358;
  assign n57605 = pi18 ? n32 : n57604;
  assign n57606 = pi17 ? n32 : n57605;
  assign n57607 = pi16 ? n57606 : ~n2320;
  assign n57608 = pi15 ? n29729 : n57607;
  assign n57609 = pi14 ? n57603 : n57608;
  assign n57610 = pi13 ? n57602 : n57609;
  assign n57611 = pi12 ? n57599 : n57610;
  assign n57612 = pi15 ? n165 : n19531;
  assign n57613 = pi19 ? n32 : n17652;
  assign n57614 = pi18 ? n32 : n57613;
  assign n57615 = pi19 ? n29290 : ~n17652;
  assign n57616 = pi18 ? n57615 : ~n237;
  assign n57617 = pi17 ? n57614 : n57616;
  assign n57618 = pi16 ? n32 : n57617;
  assign n57619 = pi15 ? n18657 : n57618;
  assign n57620 = pi14 ? n57612 : n57619;
  assign n57621 = pi13 ? n19327 : n57620;
  assign n57622 = pi17 ? n2750 : ~n2325;
  assign n57623 = pi16 ? n32 : n57622;
  assign n57624 = pi15 ? n57623 : n32;
  assign n57625 = pi14 ? n57624 : n19691;
  assign n57626 = pi18 ? n32 : ~n43015;
  assign n57627 = pi17 ? n32 : n57626;
  assign n57628 = pi16 ? n32 : n57627;
  assign n57629 = pi15 ? n19264 : n57628;
  assign n57630 = pi14 ? n57629 : n19628;
  assign n57631 = pi13 ? n57625 : n57630;
  assign n57632 = pi12 ? n57621 : n57631;
  assign n57633 = pi11 ? n57611 : n57632;
  assign n57634 = pi18 ? n33807 : ~n20023;
  assign n57635 = pi17 ? n43031 : n57634;
  assign n57636 = pi16 ? n32 : n57635;
  assign n57637 = pi15 ? n57636 : n18661;
  assign n57638 = pi14 ? n57637 : n19334;
  assign n57639 = pi15 ? n19172 : n18535;
  assign n57640 = pi14 ? n18536 : n57639;
  assign n57641 = pi13 ? n57638 : n57640;
  assign n57642 = pi16 ? n1471 : ~n4729;
  assign n57643 = pi17 ? n32 : n4381;
  assign n57644 = pi16 ? n1214 : ~n57643;
  assign n57645 = pi15 ? n57642 : n57644;
  assign n57646 = pi16 ? n1233 : ~n57552;
  assign n57647 = pi14 ? n57645 : n57646;
  assign n57648 = pi15 ? n28947 : n31707;
  assign n57649 = pi14 ? n56174 : n57648;
  assign n57650 = pi13 ? n57647 : n57649;
  assign n57651 = pi12 ? n57641 : n57650;
  assign n57652 = pi15 ? n31707 : n44289;
  assign n57653 = pi18 ? n702 : ~n618;
  assign n57654 = pi17 ? n32 : n57653;
  assign n57655 = pi16 ? n32 : n57654;
  assign n57656 = pi18 ? n36761 : ~n618;
  assign n57657 = pi17 ? n32 : n57656;
  assign n57658 = pi16 ? n32 : n57657;
  assign n57659 = pi15 ? n57655 : n57658;
  assign n57660 = pi14 ? n57652 : n57659;
  assign n57661 = pi13 ? n57660 : n19355;
  assign n57662 = pi18 ? n917 : ~n32;
  assign n57663 = pi17 ? n32 : n57662;
  assign n57664 = pi16 ? n1214 : ~n57663;
  assign n57665 = pi15 ? n18309 : n57664;
  assign n57666 = pi14 ? n19362 : n57665;
  assign n57667 = pi22 ? n32 : ~n33;
  assign n57668 = pi21 ? n32 : ~n57667;
  assign n57669 = pi20 ? n32 : n57668;
  assign n57670 = pi19 ? n32 : n57669;
  assign n57671 = pi18 ? n57670 : ~n32;
  assign n57672 = pi17 ? n32 : n57671;
  assign n57673 = pi16 ? n43068 : ~n57672;
  assign n57674 = pi15 ? n57673 : n28992;
  assign n57675 = pi20 ? n32 : n13674;
  assign n57676 = pi19 ? n32 : n57675;
  assign n57677 = pi18 ? n57676 : ~n32;
  assign n57678 = pi17 ? n32 : n57677;
  assign n57679 = pi16 ? n1233 : ~n57678;
  assign n57680 = pi15 ? n57679 : n43529;
  assign n57681 = pi14 ? n57674 : n57680;
  assign n57682 = pi13 ? n57666 : n57681;
  assign n57683 = pi12 ? n57661 : n57682;
  assign n57684 = pi11 ? n57651 : n57683;
  assign n57685 = pi10 ? n57633 : n57684;
  assign n57686 = pi09 ? n32 : n57685;
  assign n57687 = pi16 ? n1135 : ~n2320;
  assign n57688 = pi15 ? n30941 : n57687;
  assign n57689 = pi14 ? n19326 : n57688;
  assign n57690 = pi13 ? n57595 : n57689;
  assign n57691 = pi15 ? n57687 : n31854;
  assign n57692 = pi16 ? n1214 : ~n2320;
  assign n57693 = pi15 ? n31146 : n57692;
  assign n57694 = pi14 ? n57691 : n57693;
  assign n57695 = pi16 ? n1233 : ~n2320;
  assign n57696 = pi15 ? n57695 : n31146;
  assign n57697 = pi14 ? n57696 : n57608;
  assign n57698 = pi13 ? n57694 : n57697;
  assign n57699 = pi12 ? n57690 : n57698;
  assign n57700 = pi15 ? n19235 : n165;
  assign n57701 = pi14 ? n19325 : n57700;
  assign n57702 = pi13 ? n57701 : n57620;
  assign n57703 = pi15 ? n19628 : n19694;
  assign n57704 = pi14 ? n57703 : n19264;
  assign n57705 = pi13 ? n57625 : n57704;
  assign n57706 = pi12 ? n57702 : n57705;
  assign n57707 = pi11 ? n57699 : n57706;
  assign n57708 = pi17 ? n18560 : n20095;
  assign n57709 = pi16 ? n32 : n57708;
  assign n57710 = pi15 ? n57709 : n18657;
  assign n57711 = pi14 ? n57710 : n19399;
  assign n57712 = pi15 ? n19172 : n18531;
  assign n57713 = pi14 ? n43103 : n57712;
  assign n57714 = pi13 ? n57711 : n57713;
  assign n57715 = pi18 ? n32 : ~n18802;
  assign n57716 = pi17 ? n32 : n57715;
  assign n57717 = pi16 ? n1135 : ~n57716;
  assign n57718 = pi17 ? n32 : n43909;
  assign n57719 = pi16 ? n1135 : ~n57718;
  assign n57720 = pi15 ? n57717 : n57719;
  assign n57721 = pi14 ? n57645 : n57720;
  assign n57722 = pi18 ? n863 : ~n54;
  assign n57723 = pi17 ? n32 : n57722;
  assign n57724 = pi16 ? n1233 : ~n57723;
  assign n57725 = pi15 ? n29676 : n57724;
  assign n57726 = pi15 ? n57724 : n31707;
  assign n57727 = pi14 ? n57725 : n57726;
  assign n57728 = pi13 ? n57721 : n57727;
  assign n57729 = pi12 ? n57714 : n57728;
  assign n57730 = pi15 ? n31707 : n19476;
  assign n57731 = pi14 ? n57730 : n57659;
  assign n57732 = pi16 ? n19352 : ~n1683;
  assign n57733 = pi15 ? n19349 : n57732;
  assign n57734 = pi14 ? n19348 : n57733;
  assign n57735 = pi13 ? n57731 : n57734;
  assign n57736 = pi16 ? n19358 : ~n1683;
  assign n57737 = pi15 ? n57736 : n19361;
  assign n57738 = pi19 ? n32 : n30659;
  assign n57739 = pi18 ? n57738 : ~n32;
  assign n57740 = pi17 ? n32 : n57739;
  assign n57741 = pi16 ? n19652 : ~n57740;
  assign n57742 = pi15 ? n18309 : n57741;
  assign n57743 = pi14 ? n57737 : n57742;
  assign n57744 = pi16 ? n43068 : ~n56806;
  assign n57745 = pi16 ? n1214 : ~n56281;
  assign n57746 = pi15 ? n57744 : n57745;
  assign n57747 = pi14 ? n57746 : n43529;
  assign n57748 = pi13 ? n57743 : n57747;
  assign n57749 = pi12 ? n57735 : n57748;
  assign n57750 = pi11 ? n57729 : n57749;
  assign n57751 = pi10 ? n57707 : n57750;
  assign n57752 = pi09 ? n32 : n57751;
  assign n57753 = pi08 ? n57686 : n57752;
  assign n57754 = pi14 ? n30520 : n32;
  assign n57755 = pi15 ? n57596 : n57695;
  assign n57756 = pi14 ? n19447 : n57755;
  assign n57757 = pi13 ? n57754 : n57756;
  assign n57758 = pi15 ? n57692 : n31856;
  assign n57759 = pi15 ? n31854 : n57692;
  assign n57760 = pi14 ? n57758 : n57759;
  assign n57761 = pi14 ? n57758 : n19435;
  assign n57762 = pi13 ? n57760 : n57761;
  assign n57763 = pi12 ? n57757 : n57762;
  assign n57764 = pi18 ? n56721 : ~n237;
  assign n57765 = pi17 ? n35241 : n57764;
  assign n57766 = pi16 ? n32 : n57765;
  assign n57767 = pi15 ? n32 : n57766;
  assign n57768 = pi14 ? n32 : n57767;
  assign n57769 = pi13 ? n19448 : n57768;
  assign n57770 = pi17 ? n3067 : ~n2136;
  assign n57771 = pi16 ? n32 : n57770;
  assign n57772 = pi15 ? n57771 : n18657;
  assign n57773 = pi19 ? n8064 : n32;
  assign n57774 = pi18 ? n32 : n57773;
  assign n57775 = pi17 ? n32 : n57774;
  assign n57776 = pi16 ? n32 : n57775;
  assign n57777 = pi15 ? n19235 : n57776;
  assign n57778 = pi14 ? n57772 : n57777;
  assign n57779 = pi21 ? n405 : n124;
  assign n57780 = pi20 ? n57779 : n32;
  assign n57781 = pi19 ? n57780 : n32;
  assign n57782 = pi18 ? n32 : n57781;
  assign n57783 = pi17 ? n32 : n57782;
  assign n57784 = pi16 ? n32 : n57783;
  assign n57785 = pi15 ? n19531 : n57784;
  assign n57786 = pi21 ? n7107 : ~n140;
  assign n57787 = pi20 ? n57786 : n32;
  assign n57788 = pi19 ? n57787 : n32;
  assign n57789 = pi18 ? n32 : n57788;
  assign n57790 = pi17 ? n32 : n57789;
  assign n57791 = pi16 ? n32 : n57790;
  assign n57792 = pi21 ? n100 : n140;
  assign n57793 = pi20 ? n57792 : ~n32;
  assign n57794 = pi19 ? n57793 : ~n32;
  assign n57795 = pi18 ? n32 : ~n57794;
  assign n57796 = pi17 ? n32 : n57795;
  assign n57797 = pi16 ? n32 : n57796;
  assign n57798 = pi15 ? n57791 : n57797;
  assign n57799 = pi14 ? n57785 : n57798;
  assign n57800 = pi13 ? n57778 : n57799;
  assign n57801 = pi12 ? n57769 : n57800;
  assign n57802 = pi11 ? n57763 : n57801;
  assign n57803 = pi20 ? n9618 : ~n32;
  assign n57804 = pi19 ? n57803 : ~n32;
  assign n57805 = pi18 ? n32 : ~n57804;
  assign n57806 = pi17 ? n32 : n57805;
  assign n57807 = pi16 ? n32 : n57806;
  assign n57808 = pi15 ? n57807 : n57296;
  assign n57809 = pi14 ? n57808 : n18531;
  assign n57810 = pi15 ? n32 : n30096;
  assign n57811 = pi14 ? n20583 : n57810;
  assign n57812 = pi13 ? n57809 : n57811;
  assign n57813 = pi17 ? n32 : n49539;
  assign n57814 = pi16 ? n1471 : ~n57813;
  assign n57815 = pi15 ? n57814 : n57449;
  assign n57816 = pi16 ? n1233 : ~n57718;
  assign n57817 = pi15 ? n19100 : n57816;
  assign n57818 = pi14 ? n57815 : n57817;
  assign n57819 = pi18 ? n940 : ~n18802;
  assign n57820 = pi17 ? n32 : n57819;
  assign n57821 = pi16 ? n1233 : ~n57820;
  assign n57822 = pi15 ? n57821 : n28947;
  assign n57823 = pi15 ? n28947 : n57556;
  assign n57824 = pi14 ? n57822 : n57823;
  assign n57825 = pi13 ? n57818 : n57824;
  assign n57826 = pi12 ? n57812 : n57825;
  assign n57827 = pi15 ? n57556 : n43787;
  assign n57828 = pi18 ? n702 : ~n3350;
  assign n57829 = pi17 ? n32 : n57828;
  assign n57830 = pi16 ? n32 : n57829;
  assign n57831 = pi15 ? n57830 : n18594;
  assign n57832 = pi14 ? n57827 : n57831;
  assign n57833 = pi13 ? n57832 : n19482;
  assign n57834 = pi20 ? n220 : ~n274;
  assign n57835 = pi19 ? n32 : ~n57834;
  assign n57836 = pi18 ? n32 : n57835;
  assign n57837 = pi17 ? n32 : n57836;
  assign n57838 = pi20 ? n5854 : n246;
  assign n57839 = pi19 ? n57838 : ~n11899;
  assign n57840 = pi20 ? n309 : ~n206;
  assign n57841 = pi20 ? n5854 : ~n287;
  assign n57842 = pi19 ? n57840 : ~n57841;
  assign n57843 = pi18 ? n57839 : ~n57842;
  assign n57844 = pi20 ? n175 : ~n287;
  assign n57845 = pi19 ? n57844 : n2033;
  assign n57846 = pi18 ? n57845 : ~n618;
  assign n57847 = pi17 ? n57843 : n57846;
  assign n57848 = pi16 ? n57837 : n57847;
  assign n57849 = pi18 ? n28178 : n1676;
  assign n57850 = pi17 ? n32 : n57849;
  assign n57851 = pi16 ? n1214 : ~n57850;
  assign n57852 = pi15 ? n57848 : n57851;
  assign n57853 = pi14 ? n19489 : n57852;
  assign n57854 = pi16 ? n1046 : ~n57643;
  assign n57855 = pi16 ? n1135 : ~n18985;
  assign n57856 = pi15 ? n57854 : n57855;
  assign n57857 = pi16 ? n1233 : ~n18985;
  assign n57858 = pi15 ? n57857 : n43529;
  assign n57859 = pi14 ? n57856 : n57858;
  assign n57860 = pi13 ? n57853 : n57859;
  assign n57861 = pi12 ? n57833 : n57860;
  assign n57862 = pi11 ? n57826 : n57861;
  assign n57863 = pi10 ? n57802 : n57862;
  assign n57864 = pi09 ? n32 : n57863;
  assign n57865 = pi14 ? n30520 : n92;
  assign n57866 = pi15 ? n31854 : n32021;
  assign n57867 = pi14 ? n19447 : n57866;
  assign n57868 = pi13 ? n57865 : n57867;
  assign n57869 = pi15 ? n32153 : n31856;
  assign n57870 = pi15 ? n57596 : n32153;
  assign n57871 = pi14 ? n57869 : n57870;
  assign n57872 = pi14 ? n57869 : n19510;
  assign n57873 = pi13 ? n57871 : n57872;
  assign n57874 = pi12 ? n57868 : n57873;
  assign n57875 = pi14 ? n19520 : n19621;
  assign n57876 = pi13 ? n57875 : n57768;
  assign n57877 = pi15 ? n57771 : n32;
  assign n57878 = pi15 ? n30155 : n19814;
  assign n57879 = pi14 ? n57877 : n57878;
  assign n57880 = pi15 ? n19531 : n18904;
  assign n57881 = pi15 ? n19531 : n20089;
  assign n57882 = pi14 ? n57880 : n57881;
  assign n57883 = pi13 ? n57879 : n57882;
  assign n57884 = pi12 ? n57876 : n57883;
  assign n57885 = pi11 ? n57874 : n57884;
  assign n57886 = pi18 ? n32 : ~n20194;
  assign n57887 = pi17 ? n32 : n57886;
  assign n57888 = pi16 ? n32 : n57887;
  assign n57889 = pi15 ? n57888 : n19691;
  assign n57890 = pi14 ? n57889 : n43338;
  assign n57891 = pi18 ? n32 : n2662;
  assign n57892 = pi17 ? n32 : n57891;
  assign n57893 = pi16 ? n32 : n57892;
  assign n57894 = pi15 ? n32 : n57893;
  assign n57895 = pi14 ? n32 : n57894;
  assign n57896 = pi13 ? n57890 : n57895;
  assign n57897 = pi15 ? n57814 : n18979;
  assign n57898 = pi18 ? n32 : ~n18658;
  assign n57899 = pi17 ? n32 : n57898;
  assign n57900 = pi16 ? n1135 : ~n57899;
  assign n57901 = pi18 ? n32 : ~n18521;
  assign n57902 = pi17 ? n32 : n57901;
  assign n57903 = pi16 ? n1135 : ~n57902;
  assign n57904 = pi15 ? n57900 : n57903;
  assign n57905 = pi14 ? n57897 : n57904;
  assign n57906 = pi18 ? n863 : ~n18532;
  assign n57907 = pi17 ? n32 : n57906;
  assign n57908 = pi16 ? n1233 : ~n57907;
  assign n57909 = pi15 ? n29676 : n57908;
  assign n57910 = pi15 ? n57908 : n57556;
  assign n57911 = pi14 ? n57909 : n57910;
  assign n57912 = pi13 ? n57905 : n57911;
  assign n57913 = pi12 ? n57896 : n57912;
  assign n57914 = pi15 ? n57556 : n31707;
  assign n57915 = pi14 ? n57914 : n57831;
  assign n57916 = pi13 ? n57915 : n19565;
  assign n57917 = pi20 ? n7839 : ~n274;
  assign n57918 = pi19 ? n1817 : ~n57917;
  assign n57919 = pi18 ? n1819 : n57918;
  assign n57920 = pi17 ? n32 : n57919;
  assign n57921 = pi20 ? n354 : ~n9491;
  assign n57922 = pi19 ? n57838 : ~n57921;
  assign n57923 = pi20 ? n309 : n12884;
  assign n57924 = pi20 ? n21111 : ~n206;
  assign n57925 = pi19 ? n57923 : ~n57924;
  assign n57926 = pi18 ? n57922 : ~n57925;
  assign n57927 = pi20 ? n18415 : n206;
  assign n57928 = pi20 ? n18415 : n266;
  assign n57929 = pi19 ? n57927 : n57928;
  assign n57930 = pi18 ? n57929 : n618;
  assign n57931 = pi17 ? n57926 : ~n57930;
  assign n57932 = pi16 ? n57920 : n57931;
  assign n57933 = pi18 ? n4127 : n1676;
  assign n57934 = pi17 ? n32 : n57933;
  assign n57935 = pi16 ? n1214 : ~n57934;
  assign n57936 = pi15 ? n57932 : n57935;
  assign n57937 = pi14 ? n19489 : n57936;
  assign n57938 = pi18 ? n4380 : n1676;
  assign n57939 = pi17 ? n32 : n57938;
  assign n57940 = pi16 ? n1046 : ~n57939;
  assign n57941 = pi21 ? n32 : n6898;
  assign n57942 = pi20 ? n32 : n57941;
  assign n57943 = pi19 ? n32 : n57942;
  assign n57944 = pi18 ? n57943 : ~n32;
  assign n57945 = pi17 ? n32 : n57944;
  assign n57946 = pi16 ? n1135 : ~n57945;
  assign n57947 = pi15 ? n57940 : n57946;
  assign n57948 = pi14 ? n57947 : n57858;
  assign n57949 = pi13 ? n57937 : n57948;
  assign n57950 = pi12 ? n57916 : n57949;
  assign n57951 = pi11 ? n57913 : n57950;
  assign n57952 = pi10 ? n57885 : n57951;
  assign n57953 = pi09 ? n32 : n57952;
  assign n57954 = pi08 ? n57864 : n57953;
  assign n57955 = pi07 ? n57753 : n57954;
  assign n57956 = pi06 ? n57594 : n57955;
  assign n57957 = pi15 ? n19868 : n32;
  assign n57958 = pi14 ? n57957 : n19925;
  assign n57959 = pi18 ? n858 : ~n56244;
  assign n57960 = pi17 ? n32 : n57959;
  assign n57961 = pi20 ? n6050 : n17652;
  assign n57962 = pi19 ? n36181 : ~n57961;
  assign n57963 = pi20 ? n17652 : n29457;
  assign n57964 = pi20 ? n17652 : ~n6621;
  assign n57965 = pi19 ? n57963 : n57964;
  assign n57966 = pi18 ? n57962 : ~n57965;
  assign n57967 = pi19 ? n57480 : n2180;
  assign n57968 = pi18 ? n57967 : n18532;
  assign n57969 = pi17 ? n57966 : n57968;
  assign n57970 = pi16 ? n57960 : n57969;
  assign n57971 = pi15 ? n19503 : n57970;
  assign n57972 = pi15 ? n31856 : n32153;
  assign n57973 = pi14 ? n57971 : n57972;
  assign n57974 = pi13 ? n57958 : n57973;
  assign n57975 = pi15 ? n32021 : n57692;
  assign n57976 = pi14 ? n57975 : n57972;
  assign n57977 = pi15 ? n32153 : n31854;
  assign n57978 = pi14 ? n57977 : n19592;
  assign n57979 = pi13 ? n57976 : n57978;
  assign n57980 = pi12 ? n57974 : n57979;
  assign n57981 = pi14 ? n19235 : n34363;
  assign n57982 = pi13 ? n19619 : n57981;
  assign n57983 = pi18 ? n35798 : n350;
  assign n57984 = pi17 ? n32 : ~n57983;
  assign n57985 = pi16 ? n32 : n57984;
  assign n57986 = pi15 ? n57985 : n19936;
  assign n57987 = pi14 ? n57986 : n19936;
  assign n57988 = pi18 ? n32 : n19121;
  assign n57989 = pi17 ? n32 : n57988;
  assign n57990 = pi16 ? n32 : n57989;
  assign n57991 = pi17 ? n43341 : n19812;
  assign n57992 = pi16 ? n32 : n57991;
  assign n57993 = pi15 ? n57990 : n57992;
  assign n57994 = pi14 ? n43338 : n57993;
  assign n57995 = pi13 ? n57987 : n57994;
  assign n57996 = pi12 ? n57982 : n57995;
  assign n57997 = pi11 ? n57980 : n57996;
  assign n57998 = pi18 ? n17848 : n19688;
  assign n57999 = pi17 ? n32 : n57998;
  assign n58000 = pi16 ? n32 : n57999;
  assign n58001 = pi15 ? n19691 : n58000;
  assign n58002 = pi14 ? n58001 : n30209;
  assign n58003 = pi15 ? n32 : n20282;
  assign n58004 = pi14 ? n32 : n58003;
  assign n58005 = pi13 ? n58002 : n58004;
  assign n58006 = pi16 ? n1471 : ~n1683;
  assign n58007 = pi15 ? n58006 : n19100;
  assign n58008 = pi18 ? n209 : ~n18658;
  assign n58009 = pi17 ? n32 : n58008;
  assign n58010 = pi16 ? n1233 : ~n58009;
  assign n58011 = pi15 ? n19100 : n58010;
  assign n58012 = pi14 ? n58007 : n58011;
  assign n58013 = pi18 ? n684 : ~n18658;
  assign n58014 = pi17 ? n32 : n58013;
  assign n58015 = pi16 ? n1233 : ~n58014;
  assign n58016 = pi15 ? n58015 : n28947;
  assign n58017 = pi14 ? n58016 : n20034;
  assign n58018 = pi13 ? n58012 : n58017;
  assign n58019 = pi12 ? n58005 : n58018;
  assign n58020 = pi19 ? n18261 : n29682;
  assign n58021 = pi18 ? n42108 : n58020;
  assign n58022 = pi17 ? n32 : n58021;
  assign n58023 = pi20 ? n2180 : n5854;
  assign n58024 = pi19 ? n1076 : n58023;
  assign n58025 = pi18 ? n58024 : ~n43356;
  assign n58026 = pi18 ? n43360 : ~n1942;
  assign n58027 = pi17 ? n58025 : ~n58026;
  assign n58028 = pi16 ? n58022 : ~n58027;
  assign n58029 = pi15 ? n19831 : n58028;
  assign n58030 = pi14 ? n58029 : n30956;
  assign n58031 = pi13 ? n58030 : n19659;
  assign n58032 = pi18 ? n4343 : n32;
  assign n58033 = pi17 ? n58032 : n18437;
  assign n58034 = pi16 ? n32 : n58033;
  assign n58035 = pi17 ? n1219 : ~n18324;
  assign n58036 = pi16 ? n32 : ~n58035;
  assign n58037 = pi15 ? n58034 : n58036;
  assign n58038 = pi14 ? n19667 : n58037;
  assign n58039 = pi18 ? n1592 : n1676;
  assign n58040 = pi17 ? n2005 : ~n58039;
  assign n58041 = pi16 ? n1471 : n58040;
  assign n58042 = pi16 ? n1214 : ~n57448;
  assign n58043 = pi15 ? n58041 : n58042;
  assign n58044 = pi15 ? n19100 : n43577;
  assign n58045 = pi14 ? n58043 : n58044;
  assign n58046 = pi13 ? n58038 : n58045;
  assign n58047 = pi12 ? n58031 : n58046;
  assign n58048 = pi11 ? n58019 : n58047;
  assign n58049 = pi10 ? n57997 : n58048;
  assign n58050 = pi09 ? n32 : n58049;
  assign n58051 = pi20 ? n333 : n6822;
  assign n58052 = pi19 ? n58051 : n56578;
  assign n58053 = pi18 ? n1862 : ~n58052;
  assign n58054 = pi17 ? n32 : n58053;
  assign n58055 = pi20 ? n310 : n6822;
  assign n58056 = pi19 ? n56582 : n58055;
  assign n58057 = pi20 ? n6822 : n310;
  assign n58058 = pi20 ? n6822 : ~n395;
  assign n58059 = pi19 ? n58057 : n58058;
  assign n58060 = pi18 ? n58056 : n58059;
  assign n58061 = pi20 ? n18173 : ~n310;
  assign n58062 = pi19 ? n58061 : n501;
  assign n58063 = pi21 ? n174 : n85;
  assign n58064 = pi20 ? n58063 : n32;
  assign n58065 = pi19 ? n58064 : n32;
  assign n58066 = pi18 ? n58062 : n58065;
  assign n58067 = pi17 ? n58060 : ~n58066;
  assign n58068 = pi16 ? n58054 : ~n58067;
  assign n58069 = pi15 ? n156 : n58068;
  assign n58070 = pi16 ? n1214 : ~n2306;
  assign n58071 = pi15 ? n31856 : n58070;
  assign n58072 = pi14 ? n58069 : n58071;
  assign n58073 = pi13 ? n57958 : n58072;
  assign n58074 = pi16 ? n1233 : ~n2306;
  assign n58075 = pi15 ? n58074 : n32153;
  assign n58076 = pi21 ? n32 : n48999;
  assign n58077 = pi20 ? n58076 : ~n32;
  assign n58078 = pi19 ? n58077 : ~n32;
  assign n58079 = pi18 ? n32 : n58078;
  assign n58080 = pi17 ? n32 : n58079;
  assign n58081 = pi16 ? n1214 : ~n58080;
  assign n58082 = pi15 ? n32153 : n58081;
  assign n58083 = pi14 ? n58075 : n58082;
  assign n58084 = pi15 ? n58070 : n45572;
  assign n58085 = pi17 ? n19579 : ~n1933;
  assign n58086 = pi16 ? n32 : n58085;
  assign n58087 = pi15 ? n58086 : n19591;
  assign n58088 = pi14 ? n58084 : n58087;
  assign n58089 = pi13 ? n58083 : n58088;
  assign n58090 = pi12 ? n58073 : n58089;
  assign n58091 = pi14 ? n19617 : n19758;
  assign n58092 = pi18 ? n32 : ~n20345;
  assign n58093 = pi17 ? n32 : n58092;
  assign n58094 = pi16 ? n32 : n58093;
  assign n58095 = pi15 ? n91 : n58094;
  assign n58096 = pi14 ? n19235 : n58095;
  assign n58097 = pi13 ? n58091 : n58096;
  assign n58098 = pi15 ? n57985 : n19814;
  assign n58099 = pi14 ? n58098 : n43419;
  assign n58100 = pi17 ? n43423 : n19934;
  assign n58101 = pi16 ? n32 : n58100;
  assign n58102 = pi15 ? n30199 : n58101;
  assign n58103 = pi14 ? n43421 : n58102;
  assign n58104 = pi13 ? n58099 : n58103;
  assign n58105 = pi12 ? n58097 : n58104;
  assign n58106 = pi11 ? n58090 : n58105;
  assign n58107 = pi15 ? n19814 : n43498;
  assign n58108 = pi14 ? n58107 : n30263;
  assign n58109 = pi14 ? n32 : n19763;
  assign n58110 = pi13 ? n58108 : n58109;
  assign n58111 = pi15 ? n58006 : n18979;
  assign n58112 = pi18 ? n32 : ~n6867;
  assign n58113 = pi17 ? n32 : n58112;
  assign n58114 = pi16 ? n1135 : ~n58113;
  assign n58115 = pi16 ? n1135 : ~n46460;
  assign n58116 = pi15 ? n58114 : n58115;
  assign n58117 = pi14 ? n58111 : n58116;
  assign n58118 = pi16 ? n1135 : ~n58014;
  assign n58119 = pi18 ? n863 : ~n18658;
  assign n58120 = pi17 ? n32 : n58119;
  assign n58121 = pi16 ? n1135 : ~n58120;
  assign n58122 = pi15 ? n58118 : n58121;
  assign n58123 = pi15 ? n20034 : n32185;
  assign n58124 = pi14 ? n58122 : n58123;
  assign n58125 = pi13 ? n58117 : n58124;
  assign n58126 = pi12 ? n58110 : n58125;
  assign n58127 = pi19 ? n18762 : n43437;
  assign n58128 = pi18 ? n46574 : n58127;
  assign n58129 = pi17 ? n32 : n58128;
  assign n58130 = pi20 ? n501 : ~n18762;
  assign n58131 = pi19 ? n43441 : n58130;
  assign n58132 = pi18 ? n58131 : ~n43444;
  assign n58133 = pi18 ? n43447 : ~n1942;
  assign n58134 = pi17 ? n58132 : ~n58133;
  assign n58135 = pi16 ? n58129 : ~n58134;
  assign n58136 = pi15 ? n43787 : n58135;
  assign n58137 = pi14 ? n58136 : n30956;
  assign n58138 = pi17 ? n19655 : n2123;
  assign n58139 = pi16 ? n1214 : ~n58138;
  assign n58140 = pi15 ? n19711 : n58139;
  assign n58141 = pi14 ? n19650 : n58140;
  assign n58142 = pi13 ? n58137 : n58141;
  assign n58143 = pi18 ? n4380 : ~n618;
  assign n58144 = pi17 ? n1219 : ~n58143;
  assign n58145 = pi16 ? n32 : ~n58144;
  assign n58146 = pi15 ? n58034 : n58145;
  assign n58147 = pi14 ? n19667 : n58146;
  assign n58148 = pi18 ? n1592 : n618;
  assign n58149 = pi17 ? n2005 : ~n58148;
  assign n58150 = pi16 ? n1471 : n58149;
  assign n58151 = pi15 ? n58150 : n58042;
  assign n58152 = pi14 ? n58151 : n58044;
  assign n58153 = pi13 ? n58147 : n58152;
  assign n58154 = pi12 ? n58142 : n58153;
  assign n58155 = pi11 ? n58126 : n58154;
  assign n58156 = pi10 ? n58106 : n58155;
  assign n58157 = pi09 ? n32 : n58156;
  assign n58158 = pi08 ? n58050 : n58157;
  assign n58159 = pi14 ? n32 : n181;
  assign n58160 = pi13 ? n32 : n58159;
  assign n58161 = pi12 ? n32 : n58160;
  assign n58162 = pi11 ? n32 : n58161;
  assign n58163 = pi10 ? n32 : n58162;
  assign n58164 = pi15 ? n20531 : n32;
  assign n58165 = pi14 ? n58164 : n19869;
  assign n58166 = pi16 ? n1705 : ~n1934;
  assign n58167 = pi15 ? n116 : n58166;
  assign n58168 = pi19 ? n18330 : n28481;
  assign n58169 = pi18 ? n341 : ~n58168;
  assign n58170 = pi17 ? n32 : n58169;
  assign n58171 = pi20 ? n18337 : n29457;
  assign n58172 = pi19 ? n41134 : n58171;
  assign n58173 = pi21 ? n173 : ~n313;
  assign n58174 = pi20 ? n29457 : ~n58173;
  assign n58175 = pi19 ? n58174 : n11107;
  assign n58176 = pi18 ? n58172 : n58175;
  assign n58177 = pi20 ? n18624 : ~n18073;
  assign n58178 = pi20 ? n28553 : n18415;
  assign n58179 = pi19 ? n58177 : ~n58178;
  assign n58180 = pi19 ? n13172 : n32;
  assign n58181 = pi18 ? n58179 : ~n58180;
  assign n58182 = pi17 ? n58176 : n58181;
  assign n58183 = pi16 ? n58170 : ~n58182;
  assign n58184 = pi15 ? n58183 : n58070;
  assign n58185 = pi14 ? n58167 : n58184;
  assign n58186 = pi13 ? n58165 : n58185;
  assign n58187 = pi15 ? n58070 : n32153;
  assign n58188 = pi20 ? n18610 : ~n32;
  assign n58189 = pi19 ? n58188 : ~n32;
  assign n58190 = pi18 ? n32 : n58189;
  assign n58191 = pi17 ? n32 : n58190;
  assign n58192 = pi16 ? n1135 : ~n58191;
  assign n58193 = pi15 ? n32153 : n58192;
  assign n58194 = pi14 ? n58187 : n58193;
  assign n58195 = pi15 ? n34377 : n19503;
  assign n58196 = pi14 ? n58195 : n19744;
  assign n58197 = pi13 ? n58194 : n58196;
  assign n58198 = pi12 ? n58186 : n58197;
  assign n58199 = pi13 ? n19756 : n42477;
  assign n58200 = pi18 ? n17848 : n4689;
  assign n58201 = pi17 ? n32 : n58200;
  assign n58202 = pi16 ? n32 : n58201;
  assign n58203 = pi15 ? n58202 : n19942;
  assign n58204 = pi19 ? n25151 : n32;
  assign n58205 = pi18 ? n17848 : n58204;
  assign n58206 = pi17 ? n32 : n58205;
  assign n58207 = pi16 ? n32 : n58206;
  assign n58208 = pi18 ? n32 : n58204;
  assign n58209 = pi17 ? n32 : n58208;
  assign n58210 = pi16 ? n32 : n58209;
  assign n58211 = pi15 ? n58207 : n58210;
  assign n58212 = pi14 ? n58203 : n58211;
  assign n58213 = pi13 ? n43495 : n58212;
  assign n58214 = pi12 ? n58199 : n58213;
  assign n58215 = pi11 ? n58198 : n58214;
  assign n58216 = pi14 ? n30368 : n30300;
  assign n58217 = pi13 ? n58216 : n167;
  assign n58218 = pi15 ? n42182 : n18979;
  assign n58219 = pi16 ? n1135 : ~n47718;
  assign n58220 = pi15 ? n30941 : n58219;
  assign n58221 = pi14 ? n58218 : n58220;
  assign n58222 = pi15 ? n33708 : n19100;
  assign n58223 = pi14 ? n58222 : n20104;
  assign n58224 = pi13 ? n58221 : n58223;
  assign n58225 = pi12 ? n58217 : n58224;
  assign n58226 = pi15 ? n20034 : n19264;
  assign n58227 = pi14 ? n58226 : n19166;
  assign n58228 = pi13 ? n58227 : n19783;
  assign n58229 = pi15 ? n19787 : n18297;
  assign n58230 = pi16 ? n129 : n42353;
  assign n58231 = pi17 ? n1219 : ~n29201;
  assign n58232 = pi16 ? n465 : ~n58231;
  assign n58233 = pi15 ? n58230 : n58232;
  assign n58234 = pi14 ? n58229 : n58233;
  assign n58235 = pi17 ? n1227 : ~n2123;
  assign n58236 = pi16 ? n20208 : n58235;
  assign n58237 = pi16 ? n1135 : ~n56328;
  assign n58238 = pi15 ? n58236 : n58237;
  assign n58239 = pi15 ? n43529 : n18979;
  assign n58240 = pi14 ? n58238 : n58239;
  assign n58241 = pi13 ? n58234 : n58240;
  assign n58242 = pi12 ? n58228 : n58241;
  assign n58243 = pi11 ? n58225 : n58242;
  assign n58244 = pi10 ? n58215 : n58243;
  assign n58245 = pi09 ? n58163 : n58244;
  assign n58246 = pi19 ? n32 : n20937;
  assign n58247 = pi18 ? n58246 : n28484;
  assign n58248 = pi19 ? n18789 : n3495;
  assign n58249 = pi18 ? n58248 : n430;
  assign n58250 = pi17 ? n58247 : n58249;
  assign n58251 = pi16 ? n1233 : ~n58250;
  assign n58252 = pi15 ? n58251 : n45969;
  assign n58253 = pi14 ? n58167 : n58252;
  assign n58254 = pi13 ? n58165 : n58253;
  assign n58255 = pi15 ? n32153 : n57596;
  assign n58256 = pi14 ? n45969 : n58255;
  assign n58257 = pi15 ? n46354 : n20315;
  assign n58258 = pi14 ? n58257 : n19744;
  assign n58259 = pi13 ? n58256 : n58258;
  assign n58260 = pi12 ? n58254 : n58259;
  assign n58261 = pi15 ? n19753 : n32;
  assign n58262 = pi14 ? n58261 : n19755;
  assign n58263 = pi13 ? n58262 : n42477;
  assign n58264 = pi18 ? n32 : n6315;
  assign n58265 = pi17 ? n32 : n58264;
  assign n58266 = pi16 ? n32 : n58265;
  assign n58267 = pi15 ? n30207 : n58266;
  assign n58268 = pi14 ? n58203 : n58267;
  assign n58269 = pi13 ? n43556 : n58268;
  assign n58270 = pi12 ? n58263 : n58269;
  assign n58271 = pi11 ? n58260 : n58270;
  assign n58272 = pi18 ? n30295 : n19933;
  assign n58273 = pi17 ? n32 : n58272;
  assign n58274 = pi16 ? n32 : n58273;
  assign n58275 = pi15 ? n19936 : n58274;
  assign n58276 = pi14 ? n58275 : n30369;
  assign n58277 = pi13 ? n58276 : n21122;
  assign n58278 = pi15 ? n42182 : n19100;
  assign n58279 = pi18 ? n209 : ~n19688;
  assign n58280 = pi17 ? n32 : n58279;
  assign n58281 = pi16 ? n1233 : ~n58280;
  assign n58282 = pi15 ? n32806 : n58281;
  assign n58283 = pi14 ? n58278 : n58282;
  assign n58284 = pi18 ? n684 : ~n6867;
  assign n58285 = pi17 ? n32 : n58284;
  assign n58286 = pi16 ? n1233 : ~n58285;
  assign n58287 = pi15 ? n58286 : n58114;
  assign n58288 = pi15 ? n20104 : n44537;
  assign n58289 = pi14 ? n58287 : n58288;
  assign n58290 = pi13 ? n58283 : n58289;
  assign n58291 = pi12 ? n58277 : n58290;
  assign n58292 = pi15 ? n32185 : n19264;
  assign n58293 = pi14 ? n58292 : n19166;
  assign n58294 = pi13 ? n58293 : n19834;
  assign n58295 = pi16 ? n32 : n51150;
  assign n58296 = pi15 ? n19787 : n58295;
  assign n58297 = pi17 ? n18718 : n18140;
  assign n58298 = pi16 ? n32 : n58297;
  assign n58299 = pi18 ? n56517 : n18076;
  assign n58300 = pi17 ? n1219 : ~n58299;
  assign n58301 = pi16 ? n465 : ~n58300;
  assign n58302 = pi15 ? n58298 : n58301;
  assign n58303 = pi14 ? n58296 : n58302;
  assign n58304 = pi18 ? n1575 : n1676;
  assign n58305 = pi17 ? n32 : n58304;
  assign n58306 = pi16 ? n1233 : ~n58305;
  assign n58307 = pi15 ? n58236 : n58306;
  assign n58308 = pi15 ? n43577 : n18979;
  assign n58309 = pi14 ? n58307 : n58308;
  assign n58310 = pi13 ? n58303 : n58309;
  assign n58311 = pi12 ? n58294 : n58310;
  assign n58312 = pi11 ? n58291 : n58311;
  assign n58313 = pi10 ? n58271 : n58312;
  assign n58314 = pi09 ? n58163 : n58313;
  assign n58315 = pi08 ? n58245 : n58314;
  assign n58316 = pi07 ? n58158 : n58315;
  assign n58317 = pi14 ? n20139 : n32;
  assign n58318 = pi16 ? n1705 : ~n2530;
  assign n58319 = pi15 ? n180 : n58318;
  assign n58320 = pi15 ? n58318 : n45969;
  assign n58321 = pi14 ? n58319 : n58320;
  assign n58322 = pi13 ? n58317 : n58321;
  assign n58323 = pi15 ? n45969 : n31828;
  assign n58324 = pi15 ? n32153 : n32021;
  assign n58325 = pi14 ? n58323 : n58324;
  assign n58326 = pi15 ? n46354 : n180;
  assign n58327 = pi14 ? n58326 : n19857;
  assign n58328 = pi13 ? n58325 : n58327;
  assign n58329 = pi12 ? n58322 : n58328;
  assign n58330 = pi18 ? n9012 : n32;
  assign n58331 = pi17 ? n32 : n58330;
  assign n58332 = pi16 ? n32 : n58331;
  assign n58333 = pi20 ? n18415 : ~n9488;
  assign n58334 = pi19 ? n58333 : ~n44753;
  assign n58335 = pi18 ? n58334 : ~n43643;
  assign n58336 = pi17 ? n43655 : n58335;
  assign n58337 = pi16 ? n32 : n58336;
  assign n58338 = pi15 ? n58332 : n58337;
  assign n58339 = pi14 ? n32 : n58338;
  assign n58340 = pi13 ? n19863 : n58339;
  assign n58341 = pi21 ? n206 : ~n48999;
  assign n58342 = pi20 ? n58341 : n32;
  assign n58343 = pi19 ? n58342 : n32;
  assign n58344 = pi18 ? n43677 : n58343;
  assign n58345 = pi17 ? n32 : n58344;
  assign n58346 = pi16 ? n32 : n58345;
  assign n58347 = pi15 ? n58346 : n43684;
  assign n58348 = pi20 ? n8661 : n32;
  assign n58349 = pi19 ? n58348 : n32;
  assign n58350 = pi18 ? n32 : n58349;
  assign n58351 = pi17 ? n32 : n58350;
  assign n58352 = pi16 ? n32 : n58351;
  assign n58353 = pi15 ? n58352 : n19942;
  assign n58354 = pi14 ? n58347 : n58353;
  assign n58355 = pi13 ? n43676 : n58354;
  assign n58356 = pi12 ? n58340 : n58355;
  assign n58357 = pi11 ? n58329 : n58356;
  assign n58358 = pi15 ? n30534 : n30431;
  assign n58359 = pi14 ? n58358 : n30439;
  assign n58360 = pi15 ? n32 : n20646;
  assign n58361 = pi14 ? n32 : n58360;
  assign n58362 = pi13 ? n58359 : n58361;
  assign n58363 = pi18 ? n4380 : n57389;
  assign n58364 = pi17 ? n32 : n58363;
  assign n58365 = pi16 ? n1135 : ~n58364;
  assign n58366 = pi17 ? n19886 : n1978;
  assign n58367 = pi16 ? n1135 : ~n58366;
  assign n58368 = pi15 ? n58365 : n58367;
  assign n58369 = pi14 ? n31707 : n58368;
  assign n58370 = pi15 ? n19100 : n29601;
  assign n58371 = pi15 ? n30941 : n20104;
  assign n58372 = pi14 ? n58370 : n58371;
  assign n58373 = pi13 ? n58369 : n58372;
  assign n58374 = pi12 ? n58362 : n58373;
  assign n58375 = pi18 ? n936 : ~n1813;
  assign n58376 = pi17 ? n32 : n58375;
  assign n58377 = pi16 ? n32 : n58376;
  assign n58378 = pi15 ? n58377 : n19706;
  assign n58379 = pi14 ? n58378 : n19902;
  assign n58380 = pi13 ? n58379 : n19911;
  assign n58381 = pi15 ? n18688 : n41;
  assign n58382 = pi15 ? n18008 : n57460;
  assign n58383 = pi14 ? n58381 : n58382;
  assign n58384 = pi18 ? n858 : n618;
  assign n58385 = pi17 ? n30475 : n58384;
  assign n58386 = pi16 ? n1135 : ~n58385;
  assign n58387 = pi15 ? n58386 : n19100;
  assign n58388 = pi15 ? n19100 : n57355;
  assign n58389 = pi14 ? n58387 : n58388;
  assign n58390 = pi13 ? n58383 : n58389;
  assign n58391 = pi12 ? n58380 : n58390;
  assign n58392 = pi11 ? n58374 : n58391;
  assign n58393 = pi10 ? n58357 : n58392;
  assign n58394 = pi09 ? n32 : n58393;
  assign n58395 = pi16 ? n1705 : ~n2300;
  assign n58396 = pi16 ? n1214 : ~n2300;
  assign n58397 = pi15 ? n58395 : n58396;
  assign n58398 = pi14 ? n58319 : n58397;
  assign n58399 = pi13 ? n58317 : n58398;
  assign n58400 = pi16 ? n1233 : ~n2300;
  assign n58401 = pi15 ? n58396 : n58400;
  assign n58402 = pi14 ? n58401 : n58324;
  assign n58403 = pi15 ? n58400 : n13392;
  assign n58404 = pi14 ? n58403 : n19857;
  assign n58405 = pi13 ? n58402 : n58404;
  assign n58406 = pi12 ? n58399 : n58405;
  assign n58407 = pi15 ? n19856 : n32;
  assign n58408 = pi14 ? n58407 : n20140;
  assign n58409 = pi13 ? n58408 : n58339;
  assign n58410 = pi15 ? n43764 : n19531;
  assign n58411 = pi14 ? n58410 : n43773;
  assign n58412 = pi18 ? n43677 : n20249;
  assign n58413 = pi17 ? n32 : n58412;
  assign n58414 = pi16 ? n32 : n58413;
  assign n58415 = pi15 ? n58414 : n43684;
  assign n58416 = pi15 ? n19384 : n20258;
  assign n58417 = pi14 ? n58415 : n58416;
  assign n58418 = pi13 ? n58411 : n58417;
  assign n58419 = pi12 ? n58409 : n58418;
  assign n58420 = pi11 ? n58406 : n58419;
  assign n58421 = pi18 ? n21255 : n4689;
  assign n58422 = pi17 ? n32 : n58421;
  assign n58423 = pi16 ? n32 : n58422;
  assign n58424 = pi15 ? n58423 : n30537;
  assign n58425 = pi14 ? n58424 : n30544;
  assign n58426 = pi15 ? n32 : n19996;
  assign n58427 = pi14 ? n32 : n58426;
  assign n58428 = pi13 ? n58425 : n58427;
  assign n58429 = pi16 ? n1233 : ~n57515;
  assign n58430 = pi15 ? n43787 : n58429;
  assign n58431 = pi18 ? n4380 : n289;
  assign n58432 = pi17 ? n32 : n58431;
  assign n58433 = pi16 ? n1233 : ~n58432;
  assign n58434 = pi18 ? n496 : ~n162;
  assign n58435 = pi17 ? n19886 : n58434;
  assign n58436 = pi16 ? n1233 : ~n58435;
  assign n58437 = pi15 ? n58433 : n58436;
  assign n58438 = pi14 ? n58430 : n58437;
  assign n58439 = pi18 ? n32 : ~n162;
  assign n58440 = pi17 ? n32 : n58439;
  assign n58441 = pi16 ? n1135 : ~n58440;
  assign n58442 = pi15 ? n58441 : n30941;
  assign n58443 = pi15 ? n30941 : n44537;
  assign n58444 = pi14 ? n58442 : n58443;
  assign n58445 = pi13 ? n58438 : n58444;
  assign n58446 = pi12 ? n58428 : n58445;
  assign n58447 = pi15 ? n18428 : n32;
  assign n58448 = pi15 ? n19172 : n28947;
  assign n58449 = pi14 ? n58447 : n58448;
  assign n58450 = pi18 ? n858 : n3350;
  assign n58451 = pi17 ? n30475 : n58450;
  assign n58452 = pi16 ? n1135 : ~n58451;
  assign n58453 = pi15 ? n58452 : n19100;
  assign n58454 = pi15 ? n19100 : n19349;
  assign n58455 = pi14 ? n58453 : n58454;
  assign n58456 = pi13 ? n58449 : n58455;
  assign n58457 = pi12 ? n19954 : n58456;
  assign n58458 = pi11 ? n58446 : n58457;
  assign n58459 = pi10 ? n58420 : n58458;
  assign n58460 = pi09 ? n32 : n58459;
  assign n58461 = pi08 ? n58394 : n58460;
  assign n58462 = pi17 ? n20834 : n2410;
  assign n58463 = pi16 ? n1135 : ~n58462;
  assign n58464 = pi15 ? n58318 : n58463;
  assign n58465 = pi14 ? n58397 : n58464;
  assign n58466 = pi13 ? n30921 : n58465;
  assign n58467 = pi18 ? n32 : n30575;
  assign n58468 = pi17 ? n32 : n58467;
  assign n58469 = pi16 ? n1214 : ~n58468;
  assign n58470 = pi16 ? n1135 : ~n58468;
  assign n58471 = pi15 ? n58469 : n58470;
  assign n58472 = pi15 ? n31828 : n58070;
  assign n58473 = pi14 ? n58471 : n58472;
  assign n58474 = pi20 ? n18129 : ~n314;
  assign n58475 = pi20 ? n18173 : n18408;
  assign n58476 = pi19 ? n58474 : ~n58475;
  assign n58477 = pi18 ? n356 : ~n58476;
  assign n58478 = pi17 ? n32 : n58477;
  assign n58479 = pi19 ? n18782 : n6085;
  assign n58480 = pi20 ? n17665 : n6085;
  assign n58481 = pi19 ? n58480 : n9488;
  assign n58482 = pi18 ? n58479 : n58481;
  assign n58483 = pi19 ? n28749 : n6822;
  assign n58484 = pi21 ? n313 : ~n100;
  assign n58485 = pi20 ? n58484 : n32;
  assign n58486 = pi19 ? n58485 : n32;
  assign n58487 = pi18 ? n58483 : ~n58486;
  assign n58488 = pi17 ? n58482 : n58487;
  assign n58489 = pi16 ? n58478 : ~n58488;
  assign n58490 = pi15 ? n58489 : n32;
  assign n58491 = pi14 ? n58490 : n19972;
  assign n58492 = pi13 ? n58473 : n58491;
  assign n58493 = pi12 ? n58466 : n58492;
  assign n58494 = pi19 ? n44078 : ~n33544;
  assign n58495 = pi18 ? n58494 : ~n32;
  assign n58496 = pi17 ? n32 : ~n58495;
  assign n58497 = pi16 ? n32 : n58496;
  assign n58498 = pi15 ? n32 : n58497;
  assign n58499 = pi19 ? n28685 : ~n342;
  assign n58500 = pi18 ? n58499 : ~n177;
  assign n58501 = pi17 ? n32 : ~n58500;
  assign n58502 = pi16 ? n32 : n58501;
  assign n58503 = pi19 ? n9644 : n32;
  assign n58504 = pi18 ? n43872 : n58503;
  assign n58505 = pi17 ? n3282 : n58504;
  assign n58506 = pi16 ? n32 : n58505;
  assign n58507 = pi15 ? n58502 : n58506;
  assign n58508 = pi14 ? n58498 : n58507;
  assign n58509 = pi13 ? n19978 : n58508;
  assign n58510 = pi18 ? n43677 : n20320;
  assign n58511 = pi17 ? n32 : n58510;
  assign n58512 = pi16 ? n32 : n58511;
  assign n58513 = pi15 ? n58512 : n43889;
  assign n58514 = pi14 ? n43885 : n58513;
  assign n58515 = pi18 ? n43892 : n20320;
  assign n58516 = pi17 ? n32 : n58515;
  assign n58517 = pi16 ? n32 : n58516;
  assign n58518 = pi19 ? n7230 : ~n32;
  assign n58519 = pi18 ? n43896 : ~n58518;
  assign n58520 = pi17 ? n32 : n58519;
  assign n58521 = pi16 ? n32 : n58520;
  assign n58522 = pi15 ? n58517 : n58521;
  assign n58523 = pi18 ? n858 : n113;
  assign n58524 = pi17 ? n32 : n58523;
  assign n58525 = pi16 ? n32 : n58524;
  assign n58526 = pi18 ? n30607 : ~n344;
  assign n58527 = pi17 ? n32 : n58526;
  assign n58528 = pi16 ? n32 : n58527;
  assign n58529 = pi15 ? n58525 : n58528;
  assign n58530 = pi14 ? n58522 : n58529;
  assign n58531 = pi13 ? n58514 : n58530;
  assign n58532 = pi12 ? n58509 : n58531;
  assign n58533 = pi11 ? n58493 : n58532;
  assign n58534 = pi15 ? n30723 : n30537;
  assign n58535 = pi14 ? n58534 : n32;
  assign n58536 = pi13 ? n58535 : n93;
  assign n58537 = pi18 ? n17118 : n237;
  assign n58538 = pi17 ? n32 : n58537;
  assign n58539 = pi16 ? n1135 : ~n58538;
  assign n58540 = pi18 ? n17118 : n289;
  assign n58541 = pi17 ? n32 : n58540;
  assign n58542 = pi16 ? n1135 : ~n58541;
  assign n58543 = pi15 ? n58539 : n58542;
  assign n58544 = pi18 ? n20007 : n289;
  assign n58545 = pi17 ? n32 : n58544;
  assign n58546 = pi16 ? n1135 : ~n58545;
  assign n58547 = pi17 ? n20011 : n1978;
  assign n58548 = pi16 ? n1135 : ~n58547;
  assign n58549 = pi15 ? n58546 : n58548;
  assign n58550 = pi14 ? n58543 : n58549;
  assign n58551 = pi16 ? n1233 : ~n58440;
  assign n58552 = pi15 ? n58551 : n32806;
  assign n58553 = pi14 ? n58552 : n30941;
  assign n58554 = pi13 ? n58550 : n58553;
  assign n58555 = pi12 ? n58536 : n58554;
  assign n58556 = pi17 ? n20021 : n19396;
  assign n58557 = pi16 ? n32 : n58556;
  assign n58558 = pi15 ? n58557 : n20028;
  assign n58559 = pi14 ? n19628 : n58558;
  assign n58560 = pi13 ? n58559 : n20038;
  assign n58561 = pi15 ? n41 : n43925;
  assign n58562 = pi14 ? n57 : n58561;
  assign n58563 = pi18 ? n936 : n237;
  assign n58564 = pi17 ? n32752 : n58563;
  assign n58565 = pi16 ? n1214 : ~n58564;
  assign n58566 = pi15 ? n58565 : n43933;
  assign n58567 = pi17 ? n32 : n58450;
  assign n58568 = pi16 ? n1233 : ~n58567;
  assign n58569 = pi15 ? n58568 : n19476;
  assign n58570 = pi14 ? n58566 : n58569;
  assign n58571 = pi13 ? n58562 : n58570;
  assign n58572 = pi12 ? n58560 : n58571;
  assign n58573 = pi11 ? n58555 : n58572;
  assign n58574 = pi10 ? n58533 : n58573;
  assign n58575 = pi09 ? n32 : n58574;
  assign n58576 = pi16 ? n1705 : ~n3625;
  assign n58577 = pi17 ? n20834 : n2531;
  assign n58578 = pi16 ? n1233 : ~n58577;
  assign n58579 = pi15 ? n58576 : n58578;
  assign n58580 = pi14 ? n58397 : n58579;
  assign n58581 = pi13 ? n30921 : n58580;
  assign n58582 = pi17 ? n32 : n3333;
  assign n58583 = pi16 ? n1214 : ~n58582;
  assign n58584 = pi16 ? n1135 : ~n58582;
  assign n58585 = pi15 ? n58583 : n58584;
  assign n58586 = pi20 ? n2077 : ~n32;
  assign n58587 = pi19 ? n58586 : ~n32;
  assign n58588 = pi18 ? n32 : n58587;
  assign n58589 = pi17 ? n32 : n58588;
  assign n58590 = pi16 ? n1214 : ~n58589;
  assign n58591 = pi15 ? n58400 : n58590;
  assign n58592 = pi14 ? n58585 : n58591;
  assign n58593 = pi20 ? n17671 : n18282;
  assign n58594 = pi19 ? n58593 : n58480;
  assign n58595 = pi18 ? n29658 : n58594;
  assign n58596 = pi17 ? n32 : n58595;
  assign n58597 = pi19 ? n41134 : ~n41240;
  assign n58598 = pi20 ? n3523 : ~n18408;
  assign n58599 = pi19 ? n58598 : n28750;
  assign n58600 = pi18 ? n58597 : n58599;
  assign n58601 = pi20 ? n175 : n18129;
  assign n58602 = pi19 ? n9536 : ~n58601;
  assign n58603 = pi20 ? n17669 : n32;
  assign n58604 = pi19 ? n58603 : n32;
  assign n58605 = pi18 ? n58602 : ~n58604;
  assign n58606 = pi17 ? n58600 : ~n58605;
  assign n58607 = pi16 ? n58596 : n58606;
  assign n58608 = pi15 ? n58607 : n32;
  assign n58609 = pi14 ? n58608 : n20048;
  assign n58610 = pi13 ? n58592 : n58609;
  assign n58611 = pi12 ? n58581 : n58610;
  assign n58612 = pi18 ? n43976 : ~n43756;
  assign n58613 = pi17 ? n36054 : n58612;
  assign n58614 = pi16 ? n32 : n58613;
  assign n58615 = pi15 ? n58502 : n58614;
  assign n58616 = pi14 ? n58498 : n58615;
  assign n58617 = pi13 ? n20054 : n58616;
  assign n58618 = pi15 ? n58512 : n43985;
  assign n58619 = pi14 ? n43885 : n58618;
  assign n58620 = pi15 ? n58517 : n43899;
  assign n58621 = pi18 ? n30607 : ~n2304;
  assign n58622 = pi17 ? n32 : n58621;
  assign n58623 = pi16 ? n32 : n58622;
  assign n58624 = pi15 ? n17637 : n58623;
  assign n58625 = pi14 ? n58620 : n58624;
  assign n58626 = pi13 ? n58619 : n58625;
  assign n58627 = pi12 ? n58617 : n58626;
  assign n58628 = pi11 ? n58611 : n58627;
  assign n58629 = pi18 ? n30616 : n20249;
  assign n58630 = pi17 ? n32 : n58629;
  assign n58631 = pi16 ? n32 : n58630;
  assign n58632 = pi15 ? n58631 : n30726;
  assign n58633 = pi14 ? n58632 : n32;
  assign n58634 = pi14 ? n32 : n19504;
  assign n58635 = pi13 ? n58633 : n58634;
  assign n58636 = pi16 ? n1233 : ~n58538;
  assign n58637 = pi18 ? n17118 : n20267;
  assign n58638 = pi17 ? n32 : n58637;
  assign n58639 = pi16 ? n1233 : ~n58638;
  assign n58640 = pi15 ? n58636 : n58639;
  assign n58641 = pi18 ? n20007 : n20267;
  assign n58642 = pi17 ? n32 : n58641;
  assign n58643 = pi16 ? n1233 : ~n58642;
  assign n58644 = pi18 ? n496 : ~n19232;
  assign n58645 = pi17 ? n20011 : n58644;
  assign n58646 = pi16 ? n1233 : ~n58645;
  assign n58647 = pi15 ? n58643 : n58646;
  assign n58648 = pi14 ? n58640 : n58647;
  assign n58649 = pi18 ? n32 : ~n19232;
  assign n58650 = pi17 ? n32 : n58649;
  assign n58651 = pi16 ? n1135 : ~n58650;
  assign n58652 = pi15 ? n58651 : n57279;
  assign n58653 = pi14 ? n58652 : n57279;
  assign n58654 = pi13 ? n58648 : n58653;
  assign n58655 = pi12 ? n58635 : n58654;
  assign n58656 = pi17 ? n20021 : n18487;
  assign n58657 = pi16 ? n32 : n58656;
  assign n58658 = pi15 ? n58657 : n20099;
  assign n58659 = pi14 ? n19694 : n58658;
  assign n58660 = pi13 ? n58659 : n20108;
  assign n58661 = pi15 ? n18688 : n44005;
  assign n58662 = pi14 ? n20110 : n58661;
  assign n58663 = pi13 ? n58662 : n58570;
  assign n58664 = pi12 ? n58660 : n58663;
  assign n58665 = pi11 ? n58655 : n58664;
  assign n58666 = pi10 ? n58628 : n58665;
  assign n58667 = pi09 ? n32 : n58666;
  assign n58668 = pi08 ? n58575 : n58667;
  assign n58669 = pi07 ? n58461 : n58668;
  assign n58670 = pi06 ? n58316 : n58669;
  assign n58671 = pi05 ? n57956 : n58670;
  assign n58672 = pi18 ? n32 : ~n3786;
  assign n58673 = pi17 ? n32 : n58672;
  assign n58674 = pi16 ? n32 : n58673;
  assign n58675 = pi15 ? n58674 : n12788;
  assign n58676 = pi18 ? n36162 : n32413;
  assign n58677 = pi17 ? n1480 : ~n58676;
  assign n58678 = pi16 ? n32 : n58677;
  assign n58679 = pi15 ? n58678 : n29729;
  assign n58680 = pi14 ? n58675 : n58679;
  assign n58681 = pi15 ? n58576 : n47261;
  assign n58682 = pi20 ? n6621 : n1331;
  assign n58683 = pi19 ? n58682 : ~n207;
  assign n58684 = pi18 ? n48399 : n58683;
  assign n58685 = pi20 ? n1817 : n518;
  assign n58686 = pi20 ? n7839 : n246;
  assign n58687 = pi19 ? n58685 : ~n58686;
  assign n58688 = pi18 ? n58687 : n532;
  assign n58689 = pi17 ? n58684 : ~n58688;
  assign n58690 = pi16 ? n41019 : n58689;
  assign n58691 = pi19 ? n16304 : n5614;
  assign n58692 = pi18 ? n58691 : n423;
  assign n58693 = pi17 ? n18655 : n58692;
  assign n58694 = pi16 ? n1135 : ~n58693;
  assign n58695 = pi15 ? n58690 : n58694;
  assign n58696 = pi14 ? n58681 : n58695;
  assign n58697 = pi13 ? n58680 : n58696;
  assign n58698 = pi17 ? n32 : n24786;
  assign n58699 = pi16 ? n1135 : ~n58698;
  assign n58700 = pi15 ? n58699 : n58583;
  assign n58701 = pi18 ? n341 : ~n9012;
  assign n58702 = pi17 ? n32 : n58701;
  assign n58703 = pi16 ? n58702 : ~n2530;
  assign n58704 = pi19 ? n28578 : n32;
  assign n58705 = pi18 ? n366 : ~n58704;
  assign n58706 = pi17 ? n32 : n58705;
  assign n58707 = pi16 ? n58706 : ~n3625;
  assign n58708 = pi15 ? n58703 : n58707;
  assign n58709 = pi14 ? n58700 : n58708;
  assign n58710 = pi14 ? n20127 : n20779;
  assign n58711 = pi13 ? n58709 : n58710;
  assign n58712 = pi12 ? n58697 : n58711;
  assign n58713 = pi14 ? n20126 : n20053;
  assign n58714 = pi20 ? n3523 : n3843;
  assign n58715 = pi20 ? n3843 : ~n9491;
  assign n58716 = pi19 ? n58714 : n58715;
  assign n58717 = pi18 ? n58716 : n2662;
  assign n58718 = pi17 ? n3282 : n58717;
  assign n58719 = pi16 ? n32 : n58718;
  assign n58720 = pi18 ? n30779 : n34724;
  assign n58721 = pi17 ? n2954 : ~n58720;
  assign n58722 = pi16 ? n32 : n58721;
  assign n58723 = pi15 ? n58719 : n58722;
  assign n58724 = pi17 ? n32 : n33156;
  assign n58725 = pi16 ? n32 : n58724;
  assign n58726 = pi15 ? n58725 : n44224;
  assign n58727 = pi14 ? n58723 : n58726;
  assign n58728 = pi13 ? n58713 : n58727;
  assign n58729 = pi21 ? n405 : ~n9326;
  assign n58730 = pi20 ? n58729 : n32;
  assign n58731 = pi19 ? n58730 : n32;
  assign n58732 = pi18 ? n44105 : n58731;
  assign n58733 = pi17 ? n16450 : n58732;
  assign n58734 = pi16 ? n32 : n58733;
  assign n58735 = pi20 ? n406 : ~n32;
  assign n58736 = pi19 ? n58735 : ~n32;
  assign n58737 = pi18 ? n44110 : ~n58736;
  assign n58738 = pi17 ? n16317 : n58737;
  assign n58739 = pi16 ? n32 : n58738;
  assign n58740 = pi15 ? n58734 : n58739;
  assign n58741 = pi18 ? n4127 : n20320;
  assign n58742 = pi17 ? n32 : n58741;
  assign n58743 = pi16 ? n32 : n58742;
  assign n58744 = pi15 ? n58743 : n30929;
  assign n58745 = pi14 ? n58740 : n58744;
  assign n58746 = pi13 ? n44104 : n58745;
  assign n58747 = pi12 ? n58728 : n58746;
  assign n58748 = pi11 ? n58712 : n58747;
  assign n58749 = pi16 ? n1471 : ~n1471;
  assign n58750 = pi19 ? n9101 : ~n32;
  assign n58751 = pi18 ? n32 : n58750;
  assign n58752 = pi17 ? n32 : n58751;
  assign n58753 = pi16 ? n1135 : ~n58752;
  assign n58754 = pi15 ? n58749 : n58753;
  assign n58755 = pi14 ? n32 : n58754;
  assign n58756 = pi13 ? n44256 : n58755;
  assign n58757 = pi21 ? n206 : ~n85;
  assign n58758 = pi20 ? n58757 : ~n32;
  assign n58759 = pi19 ? n58758 : ~n32;
  assign n58760 = pi18 ? n4380 : n58759;
  assign n58761 = pi17 ? n16103 : n58760;
  assign n58762 = pi16 ? n1135 : ~n58761;
  assign n58763 = pi15 ? n31253 : n58762;
  assign n58764 = pi18 ? n4380 : n20345;
  assign n58765 = pi17 ? n32 : n58764;
  assign n58766 = pi16 ? n1135 : ~n58765;
  assign n58767 = pi18 ? n20166 : ~n6059;
  assign n58768 = pi17 ? n20165 : n58767;
  assign n58769 = pi16 ? n1135 : ~n58768;
  assign n58770 = pi15 ? n58766 : n58769;
  assign n58771 = pi14 ? n58763 : n58770;
  assign n58772 = pi18 ? n32 : n53735;
  assign n58773 = pi17 ? n32 : n58772;
  assign n58774 = pi16 ? n19652 : ~n58773;
  assign n58775 = pi18 ? n37939 : ~n6303;
  assign n58776 = pi17 ? n32 : n58775;
  assign n58777 = pi20 ? n820 : n7939;
  assign n58778 = pi20 ? n18540 : n354;
  assign n58779 = pi19 ? n58777 : n58778;
  assign n58780 = pi18 ? n58779 : ~n44136;
  assign n58781 = pi18 ? n44140 : ~n1548;
  assign n58782 = pi17 ? n58780 : n58781;
  assign n58783 = pi16 ? n58776 : n58782;
  assign n58784 = pi15 ? n58774 : n58783;
  assign n58785 = pi14 ? n57596 : n58784;
  assign n58786 = pi13 ? n58771 : n58785;
  assign n58787 = pi12 ? n58756 : n58786;
  assign n58788 = pi15 ? n20212 : n18661;
  assign n58789 = pi14 ? n20206 : n58788;
  assign n58790 = pi13 ? n20199 : n58789;
  assign n58791 = pi16 ? n270 : n18660;
  assign n58792 = pi17 ? n30877 : n18533;
  assign n58793 = pi16 ? n270 : n58792;
  assign n58794 = pi15 ? n58791 : n58793;
  assign n58795 = pi17 ? n1542 : n44925;
  assign n58796 = pi16 ? n1214 : ~n58795;
  assign n58797 = pi15 ? n58796 : n19711;
  assign n58798 = pi14 ? n58794 : n58797;
  assign n58799 = pi18 ? n936 : n56974;
  assign n58800 = pi17 ? n32 : n58799;
  assign n58801 = pi16 ? n1214 : ~n58800;
  assign n58802 = pi15 ? n58801 : n43933;
  assign n58803 = pi16 ? n1233 : ~n41825;
  assign n58804 = pi18 ? n209 : ~n46569;
  assign n58805 = pi17 ? n32 : n58804;
  assign n58806 = pi18 ? n20020 : n32;
  assign n58807 = pi17 ? n58806 : n2325;
  assign n58808 = pi16 ? n58805 : ~n58807;
  assign n58809 = pi15 ? n58803 : n58808;
  assign n58810 = pi14 ? n58802 : n58809;
  assign n58811 = pi13 ? n58798 : n58810;
  assign n58812 = pi12 ? n58790 : n58811;
  assign n58813 = pi11 ? n58787 : n58812;
  assign n58814 = pi10 ? n58748 : n58813;
  assign n58815 = pi09 ? n32 : n58814;
  assign n58816 = pi19 ? n41493 : ~n18778;
  assign n58817 = pi18 ? n41321 : ~n58816;
  assign n58818 = pi17 ? n32 : n58817;
  assign n58819 = pi19 ? n58480 : n18129;
  assign n58820 = pi18 ? n58479 : n58819;
  assign n58821 = pi19 ? n29002 : n17671;
  assign n58822 = pi18 ? n58821 : n3786;
  assign n58823 = pi17 ? n58820 : n58822;
  assign n58824 = pi16 ? n58818 : ~n58823;
  assign n58825 = pi20 ? n175 : n141;
  assign n58826 = pi19 ? n58825 : ~n32;
  assign n58827 = pi18 ? n24064 : n58826;
  assign n58828 = pi17 ? n19529 : n58827;
  assign n58829 = pi16 ? n1135 : ~n58828;
  assign n58830 = pi15 ? n58824 : n58829;
  assign n58831 = pi14 ? n47339 : n58830;
  assign n58832 = pi13 ? n58680 : n58831;
  assign n58833 = pi18 ? n32 : n20680;
  assign n58834 = pi17 ? n32 : n58833;
  assign n58835 = pi16 ? n1233 : ~n58834;
  assign n58836 = pi15 ? n58835 : n58583;
  assign n58837 = pi16 ? n1233 : ~n3788;
  assign n58838 = pi15 ? n58703 : n58837;
  assign n58839 = pi14 ? n58836 : n58838;
  assign n58840 = pi15 ? n19972 : n20779;
  assign n58841 = pi14 ? n30915 : n58840;
  assign n58842 = pi13 ? n58839 : n58841;
  assign n58843 = pi12 ? n58832 : n58842;
  assign n58844 = pi13 ? n20228 : n58727;
  assign n58845 = pi18 ? n4127 : n13086;
  assign n58846 = pi17 ? n32 : n58845;
  assign n58847 = pi16 ? n32 : n58846;
  assign n58848 = pi18 ? n7038 : ~n430;
  assign n58849 = pi17 ? n32 : n58848;
  assign n58850 = pi16 ? n32 : n58849;
  assign n58851 = pi15 ? n58847 : n58850;
  assign n58852 = pi14 ? n44243 : n58851;
  assign n58853 = pi13 ? n44235 : n58852;
  assign n58854 = pi12 ? n58844 : n58853;
  assign n58855 = pi11 ? n58843 : n58854;
  assign n58856 = pi19 ? n11575 : ~n32;
  assign n58857 = pi18 ? n32 : n58856;
  assign n58858 = pi17 ? n32 : n58857;
  assign n58859 = pi16 ? n1233 : ~n58858;
  assign n58860 = pi15 ? n58749 : n58859;
  assign n58861 = pi14 ? n32 : n58860;
  assign n58862 = pi13 ? n44256 : n58861;
  assign n58863 = pi16 ? n1233 : ~n31252;
  assign n58864 = pi18 ? n4380 : n58750;
  assign n58865 = pi17 ? n16103 : n58864;
  assign n58866 = pi16 ? n1233 : ~n58865;
  assign n58867 = pi15 ? n58863 : n58866;
  assign n58868 = pi18 ? n4380 : n1078;
  assign n58869 = pi17 ? n32 : n58868;
  assign n58870 = pi16 ? n1233 : ~n58869;
  assign n58871 = pi18 ? n20166 : ~n58204;
  assign n58872 = pi17 ? n20165 : n58871;
  assign n58873 = pi16 ? n1233 : ~n58872;
  assign n58874 = pi15 ? n58870 : n58873;
  assign n58875 = pi14 ? n58867 : n58874;
  assign n58876 = pi18 ? n1592 : ~n5854;
  assign n58877 = pi17 ? n32 : n58876;
  assign n58878 = pi19 ? n31675 : n44318;
  assign n58879 = pi20 ? n1817 : n4279;
  assign n58880 = pi19 ? n58879 : n44265;
  assign n58881 = pi18 ? n58878 : ~n58880;
  assign n58882 = pi18 ? n44270 : ~n1548;
  assign n58883 = pi17 ? n58881 : n58882;
  assign n58884 = pi16 ? n58877 : n58883;
  assign n58885 = pi15 ? n31856 : n58884;
  assign n58886 = pi14 ? n57691 : n58885;
  assign n58887 = pi13 ? n58875 : n58886;
  assign n58888 = pi12 ? n58862 : n58887;
  assign n58889 = pi15 ? n20212 : n18657;
  assign n58890 = pi14 ? n20278 : n58889;
  assign n58891 = pi13 ? n20199 : n58890;
  assign n58892 = pi16 ? n270 : n19530;
  assign n58893 = pi17 ? n30877 : n18803;
  assign n58894 = pi16 ? n270 : n58893;
  assign n58895 = pi15 ? n58892 : n58894;
  assign n58896 = pi17 ? n1542 : n3100;
  assign n58897 = pi16 ? n1214 : ~n58896;
  assign n58898 = pi18 ? n32 : n31156;
  assign n58899 = pi17 ? n32 : n58898;
  assign n58900 = pi16 ? n1214 : ~n58899;
  assign n58901 = pi15 ? n58897 : n58900;
  assign n58902 = pi14 ? n58895 : n58901;
  assign n58903 = pi17 ? n32 : n3367;
  assign n58904 = pi16 ? n1214 : ~n58903;
  assign n58905 = pi15 ? n58904 : n43933;
  assign n58906 = pi14 ? n58905 : n58809;
  assign n58907 = pi13 ? n58902 : n58906;
  assign n58908 = pi12 ? n58891 : n58907;
  assign n58909 = pi11 ? n58888 : n58908;
  assign n58910 = pi10 ? n58855 : n58909;
  assign n58911 = pi09 ? n32 : n58910;
  assign n58912 = pi08 ? n58815 : n58911;
  assign n58913 = pi15 ? n23561 : n12788;
  assign n58914 = pi18 ? n36162 : n1601;
  assign n58915 = pi17 ? n1480 : ~n58914;
  assign n58916 = pi16 ? n32 : n58915;
  assign n58917 = pi15 ? n58916 : n31146;
  assign n58918 = pi14 ? n58913 : n58917;
  assign n58919 = pi19 ? n32 : ~n18266;
  assign n58920 = pi20 ? n19731 : ~n18253;
  assign n58921 = pi19 ? n58920 : ~n7939;
  assign n58922 = pi18 ? n58919 : n58921;
  assign n58923 = pi20 ? n18415 : n6822;
  assign n58924 = pi19 ? n58923 : ~n1368;
  assign n58925 = pi20 ? n18129 : n141;
  assign n58926 = pi19 ? n58925 : ~n32;
  assign n58927 = pi18 ? n58924 : n58926;
  assign n58928 = pi17 ? n58922 : ~n58927;
  assign n58929 = pi16 ? n41651 : n58928;
  assign n58930 = pi15 ? n58929 : n46774;
  assign n58931 = pi18 ? n32 : n23312;
  assign n58932 = pi17 ? n32 : n58931;
  assign n58933 = pi16 ? n1214 : ~n58932;
  assign n58934 = pi15 ? n35359 : n58933;
  assign n58935 = pi14 ? n58930 : n58934;
  assign n58936 = pi13 ? n58918 : n58935;
  assign n58937 = pi16 ? n1135 : ~n58834;
  assign n58938 = pi15 ? n58937 : n35359;
  assign n58939 = pi18 ? n209 : ~n36678;
  assign n58940 = pi17 ? n32 : n58939;
  assign n58941 = pi16 ? n58940 : ~n3625;
  assign n58942 = pi20 ? n32 : n18281;
  assign n58943 = pi19 ? n32 : n58942;
  assign n58944 = pi19 ? n6074 : n18832;
  assign n58945 = pi18 ? n58943 : n58944;
  assign n58946 = pi17 ? n32 : n58945;
  assign n58947 = pi17 ? n19432 : n58931;
  assign n58948 = pi16 ? n58946 : ~n58947;
  assign n58949 = pi15 ? n58941 : n58948;
  assign n58950 = pi14 ? n58938 : n58949;
  assign n58951 = pi14 ? n30915 : n20302;
  assign n58952 = pi13 ? n58950 : n58951;
  assign n58953 = pi12 ? n58936 : n58952;
  assign n58954 = pi19 ? n221 : n266;
  assign n58955 = pi18 ? n58954 : ~n237;
  assign n58956 = pi17 ? n32 : n58955;
  assign n58957 = pi16 ? n32 : n58956;
  assign n58958 = pi15 ? n32 : n58957;
  assign n58959 = pi14 ? n58958 : n44355;
  assign n58960 = pi13 ? n20307 : n58959;
  assign n58961 = pi15 ? n44360 : n44500;
  assign n58962 = pi14 ? n58961 : n44378;
  assign n58963 = pi15 ? n33618 : n44511;
  assign n58964 = pi18 ? n863 : n13389;
  assign n58965 = pi17 ? n32 : n58964;
  assign n58966 = pi16 ? n32 : n58965;
  assign n58967 = pi15 ? n58966 : n31014;
  assign n58968 = pi14 ? n58963 : n58967;
  assign n58969 = pi13 ? n58962 : n58968;
  assign n58970 = pi12 ? n58960 : n58969;
  assign n58971 = pi11 ? n58953 : n58970;
  assign n58972 = pi18 ? n17848 : n44957;
  assign n58973 = pi17 ? n32 : n58972;
  assign n58974 = pi16 ? n1135 : ~n58973;
  assign n58975 = pi15 ? n58749 : n58974;
  assign n58976 = pi14 ? n32 : n58975;
  assign n58977 = pi13 ? n44393 : n58976;
  assign n58978 = pi18 ? n4380 : n1548;
  assign n58979 = pi17 ? n32 : n58978;
  assign n58980 = pi16 ? n1135 : ~n58979;
  assign n58981 = pi18 ? n4380 : n58189;
  assign n58982 = pi17 ? n32 : n58981;
  assign n58983 = pi16 ? n1135 : ~n58982;
  assign n58984 = pi15 ? n58980 : n58983;
  assign n58985 = pi18 ? n4380 : n2304;
  assign n58986 = pi17 ? n32 : n58985;
  assign n58987 = pi16 ? n1135 : ~n58986;
  assign n58988 = pi15 ? n58987 : n32021;
  assign n58989 = pi14 ? n58984 : n58988;
  assign n58990 = pi15 ? n45572 : n57695;
  assign n58991 = pi18 ? n30848 : ~n44398;
  assign n58992 = pi18 ? n44400 : ~n2318;
  assign n58993 = pi17 ? n58991 : n58992;
  assign n58994 = pi16 ? n30847 : n58993;
  assign n58995 = pi15 ? n45573 : n58994;
  assign n58996 = pi14 ? n58990 : n58995;
  assign n58997 = pi13 ? n58989 : n58996;
  assign n58998 = pi12 ? n58977 : n58997;
  assign n58999 = pi17 ? n58806 : n18655;
  assign n59000 = pi16 ? n270 : n58999;
  assign n59001 = pi17 ? n30877 : n18659;
  assign n59002 = pi16 ? n919 : n59001;
  assign n59003 = pi15 ? n59000 : n59002;
  assign n59004 = pi14 ? n59003 : n44439;
  assign n59005 = pi17 ? n29699 : n2136;
  assign n59006 = pi16 ? n19652 : ~n59005;
  assign n59007 = pi15 ? n59006 : n43787;
  assign n59008 = pi14 ? n59007 : n19778;
  assign n59009 = pi13 ? n59004 : n59008;
  assign n59010 = pi12 ? n20408 : n59009;
  assign n59011 = pi11 ? n58998 : n59010;
  assign n59012 = pi10 ? n58971 : n59011;
  assign n59013 = pi09 ? n32 : n59012;
  assign n59014 = pi20 ? n18173 : ~n3523;
  assign n59015 = pi19 ? n32 : ~n59014;
  assign n59016 = pi19 ? n19087 : n246;
  assign n59017 = pi18 ? n59015 : n59016;
  assign n59018 = pi20 ? n339 : n18415;
  assign n59019 = pi19 ? n59018 : ~n175;
  assign n59020 = pi20 ? n6621 : n141;
  assign n59021 = pi19 ? n59020 : ~n32;
  assign n59022 = pi18 ? n59019 : n59021;
  assign n59023 = pi17 ? n59017 : ~n59022;
  assign n59024 = pi16 ? n19804 : n59023;
  assign n59025 = pi15 ? n59024 : n46774;
  assign n59026 = pi16 ? n1214 : ~n35367;
  assign n59027 = pi15 ? n46441 : n59026;
  assign n59028 = pi14 ? n59025 : n59027;
  assign n59029 = pi13 ? n58918 : n59028;
  assign n59030 = pi18 ? n32 : n54689;
  assign n59031 = pi17 ? n32 : n59030;
  assign n59032 = pi16 ? n1135 : ~n59031;
  assign n59033 = pi15 ? n59032 : n35162;
  assign n59034 = pi18 ? n209 : ~n34189;
  assign n59035 = pi17 ? n32 : n59034;
  assign n59036 = pi16 ? n59035 : ~n3625;
  assign n59037 = pi20 ? n9488 : ~n6303;
  assign n59038 = pi19 ? n59037 : ~n32;
  assign n59039 = pi18 ? n59038 : ~n32;
  assign n59040 = pi20 ? n1611 : n339;
  assign n59041 = pi19 ? n59040 : ~n32;
  assign n59042 = pi18 ? n32 : n59041;
  assign n59043 = pi17 ? n59039 : ~n59042;
  assign n59044 = pi16 ? n42505 : n59043;
  assign n59045 = pi15 ? n59036 : n59044;
  assign n59046 = pi14 ? n59033 : n59045;
  assign n59047 = pi14 ? n20302 : n13952;
  assign n59048 = pi13 ? n59046 : n59047;
  assign n59049 = pi12 ? n59029 : n59048;
  assign n59050 = pi15 ? n44877 : n31135;
  assign n59051 = pi14 ? n44512 : n59050;
  assign n59052 = pi13 ? n44508 : n59051;
  assign n59053 = pi12 ? n58960 : n59052;
  assign n59054 = pi11 ? n59049 : n59053;
  assign n59055 = pi21 ? n206 : n7478;
  assign n59056 = pi20 ? n59055 : ~n32;
  assign n59057 = pi19 ? n59056 : ~n32;
  assign n59058 = pi18 ? n17848 : n59057;
  assign n59059 = pi17 ? n32 : n59058;
  assign n59060 = pi16 ? n1233 : ~n59059;
  assign n59061 = pi15 ? n58749 : n59060;
  assign n59062 = pi14 ? n32 : n59061;
  assign n59063 = pi13 ? n43242 : n59062;
  assign n59064 = pi16 ? n1233 : ~n58979;
  assign n59065 = pi18 ? n4380 : n1266;
  assign n59066 = pi17 ? n32 : n59065;
  assign n59067 = pi16 ? n1233 : ~n59066;
  assign n59068 = pi15 ? n59064 : n59067;
  assign n59069 = pi18 ? n4380 : n430;
  assign n59070 = pi17 ? n32 : n59069;
  assign n59071 = pi16 ? n1233 : ~n59070;
  assign n59072 = pi15 ? n59071 : n45572;
  assign n59073 = pi14 ? n59068 : n59072;
  assign n59074 = pi17 ? n32 : n3093;
  assign n59075 = pi16 ? n1135 : ~n59074;
  assign n59076 = pi15 ? n59075 : n58994;
  assign n59077 = pi14 ? n32021 : n59076;
  assign n59078 = pi13 ? n59073 : n59077;
  assign n59079 = pi12 ? n59063 : n59078;
  assign n59080 = pi17 ? n16103 : n57988;
  assign n59081 = pi16 ? n32 : n59080;
  assign n59082 = pi15 ? n59081 : n20364;
  assign n59083 = pi14 ? n59082 : n20378;
  assign n59084 = pi18 ? n20459 : n162;
  assign n59085 = pi17 ? n20457 : n59084;
  assign n59086 = pi16 ? n32 : n59085;
  assign n59087 = pi15 ? n59086 : n18904;
  assign n59088 = pi14 ? n20390 : n59087;
  assign n59089 = pi13 ? n59083 : n59088;
  assign n59090 = pi17 ? n30877 : n32;
  assign n59091 = pi16 ? n919 : n59090;
  assign n59092 = pi15 ? n59000 : n59091;
  assign n59093 = pi17 ? n29699 : n42600;
  assign n59094 = pi16 ? n1214 : ~n59093;
  assign n59095 = pi15 ? n20104 : n59094;
  assign n59096 = pi14 ? n59092 : n59095;
  assign n59097 = pi16 ? n1214 : ~n59005;
  assign n59098 = pi15 ? n59097 : n43787;
  assign n59099 = pi15 ? n19778 : n19831;
  assign n59100 = pi14 ? n59098 : n59099;
  assign n59101 = pi13 ? n59096 : n59100;
  assign n59102 = pi12 ? n59089 : n59101;
  assign n59103 = pi11 ? n59079 : n59102;
  assign n59104 = pi10 ? n59054 : n59103;
  assign n59105 = pi09 ? n32 : n59104;
  assign n59106 = pi08 ? n59013 : n59105;
  assign n59107 = pi07 ? n58912 : n59106;
  assign n59108 = pi15 ? n23614 : n23561;
  assign n59109 = pi19 ? n54302 : n32;
  assign n59110 = pi18 ? n9012 : n59109;
  assign n59111 = pi17 ? n19803 : n59110;
  assign n59112 = pi16 ? n32 : n59111;
  assign n59113 = pi19 ? n3692 : n507;
  assign n59114 = pi18 ? n10078 : n59113;
  assign n59115 = pi19 ? n1490 : ~n44694;
  assign n59116 = pi18 ? n59115 : n532;
  assign n59117 = pi17 ? n59114 : ~n59116;
  assign n59118 = pi16 ? n32 : n59117;
  assign n59119 = pi15 ? n59112 : n59118;
  assign n59120 = pi14 ? n59108 : n59119;
  assign n59121 = pi19 ? n9589 : n32;
  assign n59122 = pi18 ? n30968 : n59121;
  assign n59123 = pi17 ? n32 : n59122;
  assign n59124 = pi16 ? n32 : n59123;
  assign n59125 = pi15 ? n59124 : n32;
  assign n59126 = pi18 ? n32 : ~n1601;
  assign n59127 = pi17 ? n32 : n59126;
  assign n59128 = pi16 ? n32 : n59127;
  assign n59129 = pi14 ? n59125 : n59128;
  assign n59130 = pi13 ? n59120 : n59129;
  assign n59131 = pi16 ? n1471 : ~n2654;
  assign n59132 = pi15 ? n59131 : n47261;
  assign n59133 = pi15 ? n35162 : n13952;
  assign n59134 = pi14 ? n59132 : n59133;
  assign n59135 = pi15 ? n13952 : n20477;
  assign n59136 = pi14 ? n59135 : n20477;
  assign n59137 = pi13 ? n59134 : n59136;
  assign n59138 = pi12 ? n59130 : n59137;
  assign n59139 = pi14 ? n20487 : n147;
  assign n59140 = pi18 ? n28876 : n18532;
  assign n59141 = pi17 ? n32 : n59140;
  assign n59142 = pi16 ? n32 : n59141;
  assign n59143 = pi19 ? n507 : n1076;
  assign n59144 = pi19 ? n43838 : n32;
  assign n59145 = pi18 ? n59143 : n59144;
  assign n59146 = pi17 ? n32 : n59145;
  assign n59147 = pi16 ? n32 : n59146;
  assign n59148 = pi15 ? n59142 : n59147;
  assign n59149 = pi18 ? n44615 : n31186;
  assign n59150 = pi17 ? n32 : n59149;
  assign n59151 = pi16 ? n32 : n59150;
  assign n59152 = pi15 ? n59151 : n44621;
  assign n59153 = pi14 ? n59148 : n59152;
  assign n59154 = pi13 ? n59139 : n59153;
  assign n59155 = pi18 ? n880 : ~n20680;
  assign n59156 = pi17 ? n32 : n59155;
  assign n59157 = pi16 ? n32 : n59156;
  assign n59158 = pi15 ? n33135 : n59157;
  assign n59159 = pi14 ? n59158 : n44634;
  assign n59160 = pi20 ? n18624 : ~n141;
  assign n59161 = pi19 ? n59160 : n32;
  assign n59162 = pi18 ? n463 : n59161;
  assign n59163 = pi17 ? n32 : n59162;
  assign n59164 = pi16 ? n32 : n59163;
  assign n59165 = pi15 ? n59164 : n20048;
  assign n59166 = pi15 ? n31343 : n31229;
  assign n59167 = pi14 ? n59165 : n59166;
  assign n59168 = pi13 ? n59159 : n59167;
  assign n59169 = pi12 ? n59154 : n59168;
  assign n59170 = pi11 ? n59138 : n59169;
  assign n59171 = pi18 ? n268 : ~n18532;
  assign n59172 = pi17 ? n32 : n59171;
  assign n59173 = pi16 ? n1135 : ~n59172;
  assign n59174 = pi21 ? n32 : ~n6898;
  assign n59175 = pi20 ? n59174 : n32;
  assign n59176 = pi19 ? n59175 : n32;
  assign n59177 = pi18 ? n751 : ~n59176;
  assign n59178 = pi17 ? n32 : n59177;
  assign n59179 = pi16 ? n1135 : ~n59178;
  assign n59180 = pi15 ? n59173 : n59179;
  assign n59181 = pi14 ? n32 : n59180;
  assign n59182 = pi13 ? n32 : n59181;
  assign n59183 = pi16 ? n1135 : ~n36009;
  assign n59184 = pi18 ? n32 : n34724;
  assign n59185 = pi17 ? n32 : n59184;
  assign n59186 = pi16 ? n1135 : ~n59185;
  assign n59187 = pi15 ? n59183 : n59186;
  assign n59188 = pi18 ? n940 : n34724;
  assign n59189 = pi17 ? n32 : n59188;
  assign n59190 = pi16 ? n1135 : ~n59189;
  assign n59191 = pi15 ? n59190 : n34377;
  assign n59192 = pi14 ? n59187 : n59191;
  assign n59193 = pi18 ? n31071 : ~n344;
  assign n59194 = pi17 ? n31260 : n59193;
  assign n59195 = pi16 ? n919 : n59194;
  assign n59196 = pi15 ? n59195 : n20550;
  assign n59197 = pi14 ? n32021 : n59196;
  assign n59198 = pi13 ? n59192 : n59197;
  assign n59199 = pi12 ? n59182 : n59198;
  assign n59200 = pi15 ? n32 : n19030;
  assign n59201 = pi14 ? n20578 : n59200;
  assign n59202 = pi13 ? n20574 : n59201;
  assign n59203 = pi18 ? n16847 : ~n19020;
  assign n59204 = pi17 ? n33128 : n59203;
  assign n59205 = pi16 ? n3283 : ~n59204;
  assign n59206 = pi15 ? n59205 : n44681;
  assign n59207 = pi14 ? n59206 : n44692;
  assign n59208 = pi17 ? n44699 : n42600;
  assign n59209 = pi16 ? n44697 : ~n59208;
  assign n59210 = pi15 ? n59209 : n43787;
  assign n59211 = pi17 ? n29510 : n2136;
  assign n59212 = pi16 ? n1233 : ~n59211;
  assign n59213 = pi15 ? n32185 : n59212;
  assign n59214 = pi14 ? n59210 : n59213;
  assign n59215 = pi13 ? n59207 : n59214;
  assign n59216 = pi12 ? n59202 : n59215;
  assign n59217 = pi11 ? n59199 : n59216;
  assign n59218 = pi10 ? n59170 : n59217;
  assign n59219 = pi09 ? n32 : n59218;
  assign n59220 = pi18 ? n32 : n59121;
  assign n59221 = pi17 ? n32 : n59220;
  assign n59222 = pi16 ? n32 : n59221;
  assign n59223 = pi15 ? n59222 : n32;
  assign n59224 = pi19 ? n8247 : ~n32;
  assign n59225 = pi18 ? n32 : ~n59224;
  assign n59226 = pi17 ? n32 : n59225;
  assign n59227 = pi16 ? n32 : n59226;
  assign n59228 = pi14 ? n59223 : n59227;
  assign n59229 = pi13 ? n59120 : n59228;
  assign n59230 = pi16 ? n1471 : ~n2426;
  assign n59231 = pi16 ? n19652 : ~n2654;
  assign n59232 = pi15 ? n59230 : n59231;
  assign n59233 = pi15 ? n46655 : n486;
  assign n59234 = pi14 ? n59232 : n59233;
  assign n59235 = pi13 ? n59234 : n20477;
  assign n59236 = pi12 ? n59229 : n59235;
  assign n59237 = pi20 ? n4279 : ~n339;
  assign n59238 = pi19 ? n59237 : n32;
  assign n59239 = pi18 ? n59143 : n59238;
  assign n59240 = pi17 ? n32 : n59239;
  assign n59241 = pi16 ? n32 : n59240;
  assign n59242 = pi15 ? n59142 : n59241;
  assign n59243 = pi14 ? n59242 : n44785;
  assign n59244 = pi13 ? n20592 : n59243;
  assign n59245 = pi18 ? n880 : ~n54689;
  assign n59246 = pi17 ? n32 : n59245;
  assign n59247 = pi16 ? n32 : n59246;
  assign n59248 = pi15 ? n11429 : n59247;
  assign n59249 = pi14 ? n59248 : n44796;
  assign n59250 = pi15 ? n59222 : n13684;
  assign n59251 = pi20 ? n2385 : ~n141;
  assign n59252 = pi19 ? n59251 : n32;
  assign n59253 = pi18 ? n268 : n59252;
  assign n59254 = pi17 ? n32 : n59253;
  assign n59255 = pi16 ? n32 : n59254;
  assign n59256 = pi15 ? n59255 : n31346;
  assign n59257 = pi14 ? n59250 : n59256;
  assign n59258 = pi13 ? n59249 : n59257;
  assign n59259 = pi12 ? n59244 : n59258;
  assign n59260 = pi11 ? n59236 : n59259;
  assign n59261 = pi18 ? n268 : n30435;
  assign n59262 = pi17 ? n32 : n59261;
  assign n59263 = pi16 ? n1135 : ~n59262;
  assign n59264 = pi19 ? n21588 : n32;
  assign n59265 = pi18 ? n751 : ~n59264;
  assign n59266 = pi17 ? n32 : n59265;
  assign n59267 = pi16 ? n1135 : ~n59266;
  assign n59268 = pi15 ? n59263 : n59267;
  assign n59269 = pi14 ? n32 : n59268;
  assign n59270 = pi13 ? n32 : n59269;
  assign n59271 = pi20 ? n33737 : n32;
  assign n59272 = pi19 ? n59271 : n32;
  assign n59273 = pi18 ? n32 : ~n59272;
  assign n59274 = pi17 ? n32 : n59273;
  assign n59275 = pi16 ? n1135 : ~n59274;
  assign n59276 = pi19 ? n12008 : ~n32;
  assign n59277 = pi18 ? n32 : n59276;
  assign n59278 = pi17 ? n32 : n59277;
  assign n59279 = pi16 ? n1135 : ~n59278;
  assign n59280 = pi15 ? n59275 : n59279;
  assign n59281 = pi15 ? n59190 : n58074;
  assign n59282 = pi14 ? n59280 : n59281;
  assign n59283 = pi14 ? n58074 : n59196;
  assign n59284 = pi13 ? n59282 : n59283;
  assign n59285 = pi12 ? n59270 : n59284;
  assign n59286 = pi17 ? n20566 : n31051;
  assign n59287 = pi16 ? n1471 : ~n59286;
  assign n59288 = pi17 ? n20570 : n2537;
  assign n59289 = pi16 ? n1471 : ~n59288;
  assign n59290 = pi15 ? n59287 : n59289;
  assign n59291 = pi14 ? n20564 : n59290;
  assign n59292 = pi15 ? n19235 : n20646;
  assign n59293 = pi14 ? n20578 : n59292;
  assign n59294 = pi13 ? n59291 : n59293;
  assign n59295 = pi18 ? n16847 : ~n162;
  assign n59296 = pi17 ? n33128 : n59295;
  assign n59297 = pi16 ? n3283 : ~n59296;
  assign n59298 = pi15 ? n59297 : n44812;
  assign n59299 = pi18 ? n44683 : n350;
  assign n59300 = pi17 ? n2736 : ~n59299;
  assign n59301 = pi16 ? n32 : n59300;
  assign n59302 = pi17 ? n21288 : n1807;
  assign n59303 = pi16 ? n44689 : ~n59302;
  assign n59304 = pi15 ? n59301 : n59303;
  assign n59305 = pi14 ? n59298 : n59304;
  assign n59306 = pi16 ? n1135 : ~n59211;
  assign n59307 = pi15 ? n32185 : n59306;
  assign n59308 = pi14 ? n59210 : n59307;
  assign n59309 = pi13 ? n59305 : n59308;
  assign n59310 = pi12 ? n59294 : n59309;
  assign n59311 = pi11 ? n59285 : n59310;
  assign n59312 = pi10 ? n59260 : n59311;
  assign n59313 = pi09 ? n32 : n59312;
  assign n59314 = pi08 ? n59219 : n59313;
  assign n59315 = pi15 ? n12784 : n12788;
  assign n59316 = pi19 ? n57522 : ~n29614;
  assign n59317 = pi18 ? n28053 : n59316;
  assign n59318 = pi17 ? n32 : n59317;
  assign n59319 = pi20 ? n1324 : n18762;
  assign n59320 = pi19 ? n29618 : ~n59319;
  assign n59321 = pi20 ? n357 : n17652;
  assign n59322 = pi19 ? n59321 : n12884;
  assign n59323 = pi18 ? n59320 : ~n59322;
  assign n59324 = pi20 ? n2358 : n321;
  assign n59325 = pi19 ? n247 : ~n59324;
  assign n59326 = pi18 ? n59325 : ~n13070;
  assign n59327 = pi17 ? n59323 : ~n59326;
  assign n59328 = pi16 ? n59318 : n59327;
  assign n59329 = pi20 ? n175 : n9488;
  assign n59330 = pi19 ? n32 : n59329;
  assign n59331 = pi18 ? n32 : n59330;
  assign n59332 = pi17 ? n32 : n59331;
  assign n59333 = pi20 ? n4279 : n2180;
  assign n59334 = pi19 ? n18778 : ~n59333;
  assign n59335 = pi20 ? n18282 : n2180;
  assign n59336 = pi19 ? n18924 : n59335;
  assign n59337 = pi18 ? n59334 : ~n59336;
  assign n59338 = pi20 ? n17652 : ~n9491;
  assign n59339 = pi19 ? n59338 : ~n43833;
  assign n59340 = pi19 ? n15051 : ~n32;
  assign n59341 = pi18 ? n59339 : ~n59340;
  assign n59342 = pi17 ? n59337 : ~n59341;
  assign n59343 = pi16 ? n59332 : ~n59342;
  assign n59344 = pi15 ? n59328 : n59343;
  assign n59345 = pi14 ? n59315 : n59344;
  assign n59346 = pi19 ? n12680 : ~n32;
  assign n59347 = pi18 ? n32 : ~n59346;
  assign n59348 = pi17 ? n32 : n59347;
  assign n59349 = pi16 ? n32 : n59348;
  assign n59350 = pi14 ? n20591 : n59349;
  assign n59351 = pi13 ? n59345 : n59350;
  assign n59352 = pi15 ? n59230 : n46991;
  assign n59353 = pi15 ? n46991 : n32;
  assign n59354 = pi14 ? n59352 : n59353;
  assign n59355 = pi15 ? n20477 : n20660;
  assign n59356 = pi14 ? n59355 : n20660;
  assign n59357 = pi13 ? n59354 : n59356;
  assign n59358 = pi12 ? n59351 : n59357;
  assign n59359 = pi15 ? n32 : n21755;
  assign n59360 = pi14 ? n59359 : n44865;
  assign n59361 = pi13 ? n20666 : n59360;
  assign n59362 = pi18 ? n863 : n21724;
  assign n59363 = pi17 ? n32 : n59362;
  assign n59364 = pi16 ? n32 : n59363;
  assign n59365 = pi15 ? n20982 : n59364;
  assign n59366 = pi14 ? n44874 : n59365;
  assign n59367 = pi20 ? n8644 : ~n243;
  assign n59368 = pi19 ? n59367 : n32;
  assign n59369 = pi18 ? n268 : n59368;
  assign n59370 = pi17 ? n32 : n59369;
  assign n59371 = pi16 ? n32 : n59370;
  assign n59372 = pi15 ? n59371 : n31511;
  assign n59373 = pi15 ? n20862 : n146;
  assign n59374 = pi14 ? n59372 : n59373;
  assign n59375 = pi13 ? n59366 : n59374;
  assign n59376 = pi12 ? n59361 : n59375;
  assign n59377 = pi11 ? n59358 : n59376;
  assign n59378 = pi18 ? n940 : ~n4671;
  assign n59379 = pi17 ? n32 : n59378;
  assign n59380 = pi16 ? n1233 : ~n59379;
  assign n59381 = pi15 ? n29601 : n59380;
  assign n59382 = pi14 ? n19504 : n59381;
  assign n59383 = pi13 ? n22048 : n59382;
  assign n59384 = pi18 ? n4380 : ~n6059;
  assign n59385 = pi17 ? n32 : n59384;
  assign n59386 = pi16 ? n1233 : ~n59385;
  assign n59387 = pi21 ? n206 : n13585;
  assign n59388 = pi20 ? n59387 : ~n32;
  assign n59389 = pi19 ? n59388 : ~n32;
  assign n59390 = pi18 ? n940 : n59389;
  assign n59391 = pi17 ? n32 : n59390;
  assign n59392 = pi16 ? n1233 : ~n59391;
  assign n59393 = pi15 ? n59386 : n59392;
  assign n59394 = pi16 ? n1135 : ~n2300;
  assign n59395 = pi15 ? n59394 : n34377;
  assign n59396 = pi14 ? n59393 : n59395;
  assign n59397 = pi18 ? n31071 : ~n2304;
  assign n59398 = pi17 ? n31260 : n59397;
  assign n59399 = pi16 ? n919 : n59398;
  assign n59400 = pi15 ? n59399 : n20720;
  assign n59401 = pi14 ? n34377 : n59400;
  assign n59402 = pi13 ? n59396 : n59401;
  assign n59403 = pi12 ? n59383 : n59402;
  assign n59404 = pi15 ? n20740 : n91;
  assign n59405 = pi14 ? n59404 : n19235;
  assign n59406 = pi13 ? n20742 : n59405;
  assign n59407 = pi17 ? n36949 : ~n59295;
  assign n59408 = pi16 ? n32 : n59407;
  assign n59409 = pi15 ? n59408 : n44913;
  assign n59410 = pi14 ? n59409 : n44923;
  assign n59411 = pi18 ? n32 : ~n19654;
  assign n59412 = pi17 ? n31659 : n59411;
  assign n59413 = pi16 ? n3438 : ~n59412;
  assign n59414 = pi16 ? n1233 : ~n44928;
  assign n59415 = pi15 ? n59413 : n59414;
  assign n59416 = pi18 ? n32 : n56859;
  assign n59417 = pi17 ? n32 : n59416;
  assign n59418 = pi16 ? n1233 : ~n59417;
  assign n59419 = pi20 ? n32 : n52168;
  assign n59420 = pi19 ? n32 : n59419;
  assign n59421 = pi19 ? n31482 : n33524;
  assign n59422 = pi18 ? n59420 : ~n59421;
  assign n59423 = pi17 ? n32 : n59422;
  assign n59424 = pi20 ? n820 : ~n342;
  assign n59425 = pi20 ? n6050 : n974;
  assign n59426 = pi19 ? n59424 : n59425;
  assign n59427 = pi18 ? n59426 : ~n32;
  assign n59428 = pi17 ? n59427 : ~n42600;
  assign n59429 = pi16 ? n59423 : n59428;
  assign n59430 = pi15 ? n59418 : n59429;
  assign n59431 = pi14 ? n59415 : n59430;
  assign n59432 = pi13 ? n59410 : n59431;
  assign n59433 = pi12 ? n59406 : n59432;
  assign n59434 = pi11 ? n59403 : n59433;
  assign n59435 = pi10 ? n59377 : n59434;
  assign n59436 = pi09 ? n32 : n59435;
  assign n59437 = pi19 ? n57399 : ~n29453;
  assign n59438 = pi18 ? n41285 : n59437;
  assign n59439 = pi17 ? n32 : n59438;
  assign n59440 = pi20 ? n974 : n428;
  assign n59441 = pi19 ? n29458 : ~n59440;
  assign n59442 = pi19 ? n29657 : n246;
  assign n59443 = pi18 ? n59441 : ~n59442;
  assign n59444 = pi20 ? n314 : n501;
  assign n59445 = pi19 ? n9169 : ~n59444;
  assign n59446 = pi18 ? n59445 : ~n13070;
  assign n59447 = pi17 ? n59443 : ~n59446;
  assign n59448 = pi16 ? n59439 : n59447;
  assign n59449 = pi18 ? n32 : n58246;
  assign n59450 = pi17 ? n32 : n59449;
  assign n59451 = pi20 ? n342 : n1076;
  assign n59452 = pi19 ? n18571 : ~n59451;
  assign n59453 = pi20 ? n18282 : n32;
  assign n59454 = pi19 ? n59453 : n19596;
  assign n59455 = pi18 ? n59452 : ~n59454;
  assign n59456 = pi20 ? n9491 : n18173;
  assign n59457 = pi19 ? n59338 : ~n59456;
  assign n59458 = pi20 ? n1324 : n243;
  assign n59459 = pi19 ? n59458 : ~n32;
  assign n59460 = pi18 ? n59457 : ~n59459;
  assign n59461 = pi17 ? n59455 : ~n59460;
  assign n59462 = pi16 ? n59450 : ~n59461;
  assign n59463 = pi15 ? n59448 : n59462;
  assign n59464 = pi14 ? n59315 : n59463;
  assign n59465 = pi19 ? n34295 : ~n32;
  assign n59466 = pi18 ? n32 : ~n59465;
  assign n59467 = pi17 ? n32 : n59466;
  assign n59468 = pi16 ? n32 : n59467;
  assign n59469 = pi14 ? n20591 : n59468;
  assign n59470 = pi13 ? n59464 : n59469;
  assign n59471 = pi16 ? n29327 : ~n2120;
  assign n59472 = pi15 ? n59471 : n36601;
  assign n59473 = pi15 ? n47256 : n32;
  assign n59474 = pi14 ? n59472 : n59473;
  assign n59475 = pi15 ? n20660 : n20756;
  assign n59476 = pi14 ? n59475 : n20758;
  assign n59477 = pi13 ? n59474 : n59476;
  assign n59478 = pi12 ? n59470 : n59477;
  assign n59479 = pi18 ? n32 : n31593;
  assign n59480 = pi17 ? n32 : n59479;
  assign n59481 = pi16 ? n32 : n59480;
  assign n59482 = pi15 ? n59371 : n59481;
  assign n59483 = pi14 ? n59482 : n31516;
  assign n59484 = pi13 ? n44969 : n59483;
  assign n59485 = pi12 ? n59361 : n59484;
  assign n59486 = pi11 ? n59478 : n59485;
  assign n59487 = pi18 ? n940 : ~n20671;
  assign n59488 = pi17 ? n32 : n59487;
  assign n59489 = pi16 ? n1135 : ~n59488;
  assign n59490 = pi15 ? n30941 : n59489;
  assign n59491 = pi14 ? n19504 : n59490;
  assign n59492 = pi13 ? n32 : n59491;
  assign n59493 = pi20 ? n11107 : n32;
  assign n59494 = pi19 ? n59493 : n32;
  assign n59495 = pi18 ? n4380 : ~n59494;
  assign n59496 = pi17 ? n32 : n59495;
  assign n59497 = pi16 ? n1135 : ~n59496;
  assign n59498 = pi20 ? n18624 : ~n32;
  assign n59499 = pi19 ? n59498 : ~n32;
  assign n59500 = pi18 ? n940 : n59499;
  assign n59501 = pi17 ? n32 : n59500;
  assign n59502 = pi16 ? n1135 : ~n59501;
  assign n59503 = pi15 ? n59497 : n59502;
  assign n59504 = pi15 ? n59394 : n31828;
  assign n59505 = pi14 ? n59503 : n59504;
  assign n59506 = pi16 ? n568 : n59194;
  assign n59507 = pi15 ? n59506 : n20720;
  assign n59508 = pi14 ? n46354 : n59507;
  assign n59509 = pi13 ? n59505 : n59508;
  assign n59510 = pi12 ? n59492 : n59509;
  assign n59511 = pi18 ? n20725 : n344;
  assign n59512 = pi17 ? n2733 : ~n59511;
  assign n59513 = pi16 ? n32 : n59512;
  assign n59514 = pi15 ? n59513 : n20733;
  assign n59515 = pi14 ? n59514 : n20741;
  assign n59516 = pi15 ? n20740 : n19503;
  assign n59517 = pi14 ? n59516 : n19621;
  assign n59518 = pi13 ? n59515 : n59517;
  assign n59519 = pi17 ? n44679 : ~n3337;
  assign n59520 = pi16 ? n32 : n59519;
  assign n59521 = pi15 ? n59408 : n59520;
  assign n59522 = pi14 ? n59521 : n44923;
  assign n59523 = pi17 ? n31659 : n1807;
  assign n59524 = pi16 ? n3438 : ~n59523;
  assign n59525 = pi15 ? n59524 : n32185;
  assign n59526 = pi20 ? n18261 : n1611;
  assign n59527 = pi19 ? n59526 : n29033;
  assign n59528 = pi18 ? n19082 : n59527;
  assign n59529 = pi17 ? n32 : n59528;
  assign n59530 = pi20 ? n2358 : ~n1076;
  assign n59531 = pi19 ? n59530 : n42075;
  assign n59532 = pi18 ? n59531 : ~n18532;
  assign n59533 = pi17 ? n59532 : ~n42600;
  assign n59534 = pi16 ? n59529 : n59533;
  assign n59535 = pi15 ? n59418 : n59534;
  assign n59536 = pi14 ? n59525 : n59535;
  assign n59537 = pi13 ? n59522 : n59536;
  assign n59538 = pi12 ? n59518 : n59537;
  assign n59539 = pi11 ? n59510 : n59538;
  assign n59540 = pi10 ? n59486 : n59539;
  assign n59541 = pi09 ? n32 : n59540;
  assign n59542 = pi08 ? n59436 : n59541;
  assign n59543 = pi07 ? n59314 : n59542;
  assign n59544 = pi06 ? n59107 : n59543;
  assign n59545 = pi15 ? n21232 : n32;
  assign n59546 = pi17 ? n32 : n5077;
  assign n59547 = pi18 ? n6118 : n32381;
  assign n59548 = pi17 ? n32 : n59547;
  assign n59549 = pi16 ? n59546 : ~n59548;
  assign n59550 = pi15 ? n59549 : n45947;
  assign n59551 = pi14 ? n59545 : n59550;
  assign n59552 = pi18 ? n32 : ~n34229;
  assign n59553 = pi17 ? n32 : n59552;
  assign n59554 = pi16 ? n32 : n59553;
  assign n59555 = pi15 ? n32 : n59554;
  assign n59556 = pi16 ? n1471 : ~n2415;
  assign n59557 = pi15 ? n59556 : n47471;
  assign n59558 = pi14 ? n59555 : n59557;
  assign n59559 = pi13 ? n59551 : n59558;
  assign n59560 = pi16 ? n1233 : ~n2415;
  assign n59561 = pi15 ? n47256 : n59560;
  assign n59562 = pi14 ? n59561 : n20838;
  assign n59563 = pi15 ? n13948 : n20836;
  assign n59564 = pi14 ? n59563 : n20838;
  assign n59565 = pi13 ? n59562 : n59564;
  assign n59566 = pi12 ? n59559 : n59565;
  assign n59567 = pi19 ? n507 : n28076;
  assign n59568 = pi18 ? n59567 : ~n822;
  assign n59569 = pi17 ? n32 : n59568;
  assign n59570 = pi16 ? n32 : n59569;
  assign n59571 = pi15 ? n59570 : n33101;
  assign n59572 = pi14 ? n59571 : n45050;
  assign n59573 = pi13 ? n20842 : n59572;
  assign n59574 = pi18 ? n4127 : n31785;
  assign n59575 = pi17 ? n32 : n59574;
  assign n59576 = pi16 ? n32 : n59575;
  assign n59577 = pi15 ? n19972 : n59576;
  assign n59578 = pi14 ? n45056 : n59577;
  assign n59579 = pi15 ? n21153 : n45060;
  assign n59580 = pi14 ? n59579 : n20416;
  assign n59581 = pi13 ? n59578 : n59580;
  assign n59582 = pi12 ? n59573 : n59581;
  assign n59583 = pi11 ? n59566 : n59582;
  assign n59584 = pi18 ? n880 : n32413;
  assign n59585 = pi17 ? n32 : n59584;
  assign n59586 = pi16 ? n1471 : ~n59585;
  assign n59587 = pi18 ? n4380 : n32413;
  assign n59588 = pi17 ? n32 : n59587;
  assign n59589 = pi16 ? n1214 : ~n59588;
  assign n59590 = pi15 ? n59586 : n59589;
  assign n59591 = pi18 ? n940 : ~n143;
  assign n59592 = pi17 ? n32 : n59591;
  assign n59593 = pi16 ? n1233 : ~n59592;
  assign n59594 = pi15 ? n31526 : n59593;
  assign n59595 = pi14 ? n59590 : n59594;
  assign n59596 = pi13 ? n44299 : n59595;
  assign n59597 = pi18 ? n32 : n31102;
  assign n59598 = pi17 ? n32 : n59597;
  assign n59599 = pi16 ? n1233 : ~n59598;
  assign n59600 = pi15 ? n42961 : n59599;
  assign n59601 = pi16 ? n19652 : ~n3625;
  assign n59602 = pi15 ? n59601 : n31828;
  assign n59603 = pi14 ? n59600 : n59602;
  assign n59604 = pi18 ? n341 : ~n31643;
  assign n59605 = pi17 ? n32 : n59604;
  assign n59606 = pi18 ? n31650 : n430;
  assign n59607 = pi17 ? n31649 : ~n59606;
  assign n59608 = pi16 ? n59605 : n59607;
  assign n59609 = pi15 ? n31828 : n59608;
  assign n59610 = pi14 ? n59609 : n20905;
  assign n59611 = pi13 ? n59603 : n59610;
  assign n59612 = pi12 ? n59596 : n59611;
  assign n59613 = pi15 ? n20949 : n19503;
  assign n59614 = pi18 ? n6145 : n20267;
  assign n59615 = pi17 ? n32 : n59614;
  assign n59616 = pi16 ? n1683 : ~n59615;
  assign n59617 = pi15 ? n20955 : n59616;
  assign n59618 = pi14 ? n59613 : n59617;
  assign n59619 = pi13 ? n20932 : n59618;
  assign n59620 = pi15 ? n31862 : n31695;
  assign n59621 = pi14 ? n59620 : n45118;
  assign n59622 = pi18 ? n268 : n33017;
  assign n59623 = pi17 ? n32 : n59622;
  assign n59624 = pi19 ? n349 : ~n221;
  assign n59625 = pi18 ? n59624 : ~n32;
  assign n59626 = pi17 ? n59625 : ~n43016;
  assign n59627 = pi16 ? n59623 : n59626;
  assign n59628 = pi15 ? n59627 : n32185;
  assign n59629 = pi17 ? n20165 : n1807;
  assign n59630 = pi16 ? n1233 : ~n59629;
  assign n59631 = pi18 ? n32 : ~n20172;
  assign n59632 = pi17 ? n32 : n59631;
  assign n59633 = pi16 ? n59632 : ~n57048;
  assign n59634 = pi15 ? n59630 : n59633;
  assign n59635 = pi14 ? n59628 : n59634;
  assign n59636 = pi13 ? n59621 : n59635;
  assign n59637 = pi12 ? n59619 : n59636;
  assign n59638 = pi11 ? n59612 : n59637;
  assign n59639 = pi10 ? n59583 : n59638;
  assign n59640 = pi09 ? n32 : n59639;
  assign n59641 = pi13 ? n32 : n49586;
  assign n59642 = pi12 ? n32 : n59641;
  assign n59643 = pi11 ? n32 : n59642;
  assign n59644 = pi10 ? n32 : n59643;
  assign n59645 = pi18 ? n6145 : n32381;
  assign n59646 = pi17 ? n32 : n59645;
  assign n59647 = pi16 ? n59546 : ~n59646;
  assign n59648 = pi15 ? n59647 : n45947;
  assign n59649 = pi14 ? n21558 : n59648;
  assign n59650 = pi18 ? n32 : ~n53436;
  assign n59651 = pi17 ? n32 : n59650;
  assign n59652 = pi16 ? n32 : n59651;
  assign n59653 = pi15 ? n32 : n59652;
  assign n59654 = pi16 ? n1471 : ~n2409;
  assign n59655 = pi15 ? n59654 : n47471;
  assign n59656 = pi14 ? n59653 : n59655;
  assign n59657 = pi13 ? n59649 : n59656;
  assign n59658 = pi15 ? n47256 : n34146;
  assign n59659 = pi14 ? n59658 : n20969;
  assign n59660 = pi14 ? n59563 : n20969;
  assign n59661 = pi13 ? n59659 : n59660;
  assign n59662 = pi12 ? n59657 : n59661;
  assign n59663 = pi13 ? n20838 : n59572;
  assign n59664 = pi15 ? n12095 : n45060;
  assign n59665 = pi14 ? n59664 : n20416;
  assign n59666 = pi13 ? n59578 : n59665;
  assign n59667 = pi12 ? n59663 : n59666;
  assign n59668 = pi11 ? n59662 : n59667;
  assign n59669 = pi17 ? n32 : n33884;
  assign n59670 = pi16 ? n1471 : ~n59669;
  assign n59671 = pi16 ? n1214 : ~n31442;
  assign n59672 = pi15 ? n59670 : n59671;
  assign n59673 = pi18 ? n940 : ~n13949;
  assign n59674 = pi17 ? n32 : n59673;
  assign n59675 = pi16 ? n1135 : ~n59674;
  assign n59676 = pi15 ? n31443 : n59675;
  assign n59677 = pi14 ? n59672 : n59676;
  assign n59678 = pi13 ? n32 : n59677;
  assign n59679 = pi18 ? n880 : ~n143;
  assign n59680 = pi17 ? n32 : n59679;
  assign n59681 = pi16 ? n1135 : ~n59680;
  assign n59682 = pi15 ? n59681 : n35162;
  assign n59683 = pi15 ? n58396 : n59394;
  assign n59684 = pi14 ? n59682 : n59683;
  assign n59685 = pi13 ? n59684 : n59610;
  assign n59686 = pi12 ? n59678 : n59685;
  assign n59687 = pi15 ? n21017 : n19503;
  assign n59688 = pi15 ? n91 : n59616;
  assign n59689 = pi14 ? n59687 : n59688;
  assign n59690 = pi13 ? n20932 : n59689;
  assign n59691 = pi17 ? n3067 : ~n1807;
  assign n59692 = pi16 ? n32 : n59691;
  assign n59693 = pi15 ? n31862 : n59692;
  assign n59694 = pi14 ? n59693 : n45174;
  assign n59695 = pi16 ? n1135 : ~n59629;
  assign n59696 = pi16 ? n59632 : ~n2326;
  assign n59697 = pi15 ? n59695 : n59696;
  assign n59698 = pi14 ? n59628 : n59697;
  assign n59699 = pi13 ? n59694 : n59698;
  assign n59700 = pi12 ? n59690 : n59699;
  assign n59701 = pi11 ? n59686 : n59700;
  assign n59702 = pi10 ? n59668 : n59701;
  assign n59703 = pi09 ? n59644 : n59702;
  assign n59704 = pi08 ? n59640 : n59703;
  assign n59705 = pi14 ? n32 : n21326;
  assign n59706 = pi13 ? n32 : n59705;
  assign n59707 = pi12 ? n32 : n59706;
  assign n59708 = pi11 ? n32 : n59707;
  assign n59709 = pi10 ? n32 : n59708;
  assign n59710 = pi18 ? n32 : n22159;
  assign n59711 = pi17 ? n32 : n59710;
  assign n59712 = pi16 ? n1934 : ~n59711;
  assign n59713 = pi15 ? n59712 : n20831;
  assign n59714 = pi14 ? n21553 : n59713;
  assign n59715 = pi16 ? n1214 : ~n2409;
  assign n59716 = pi15 ? n59654 : n59715;
  assign n59717 = pi14 ? n59653 : n59716;
  assign n59718 = pi13 ? n59714 : n59717;
  assign n59719 = pi14 ? n36601 : n20836;
  assign n59720 = pi15 ? n13948 : n21033;
  assign n59721 = pi14 ? n59720 : n21035;
  assign n59722 = pi13 ? n59719 : n59721;
  assign n59723 = pi12 ? n59718 : n59722;
  assign n59724 = pi13 ? n32 : n45225;
  assign n59725 = pi20 ? n8644 : ~n1940;
  assign n59726 = pi19 ? n59725 : n32;
  assign n59727 = pi18 ? n268 : n59726;
  assign n59728 = pi17 ? n32 : n59727;
  assign n59729 = pi16 ? n32 : n59728;
  assign n59730 = pi20 ? n206 : ~n10446;
  assign n59731 = pi19 ? n59730 : n32;
  assign n59732 = pi18 ? n684 : n59731;
  assign n59733 = pi17 ? n32 : n59732;
  assign n59734 = pi16 ? n32 : n59733;
  assign n59735 = pi15 ? n59729 : n59734;
  assign n59736 = pi14 ? n45233 : n59735;
  assign n59737 = pi15 ? n12095 : n45239;
  assign n59738 = pi14 ? n59737 : n486;
  assign n59739 = pi13 ? n59736 : n59738;
  assign n59740 = pi12 ? n59724 : n59739;
  assign n59741 = pi11 ? n59723 : n59740;
  assign n59742 = pi15 ? n59670 : n31443;
  assign n59743 = pi14 ? n59742 : n59676;
  assign n59744 = pi13 ? n32 : n59743;
  assign n59745 = pi18 ? n21066 : ~n13377;
  assign n59746 = pi17 ? n32 : n59745;
  assign n59747 = pi16 ? n1135 : ~n59746;
  assign n59748 = pi15 ? n59747 : n46774;
  assign n59749 = pi15 ? n59601 : n58400;
  assign n59750 = pi14 ? n59748 : n59749;
  assign n59751 = pi15 ? n58400 : n21079;
  assign n59752 = pi14 ? n59751 : n21088;
  assign n59753 = pi13 ? n59750 : n59752;
  assign n59754 = pi12 ? n59744 : n59753;
  assign n59755 = pi18 ? n6145 : n20345;
  assign n59756 = pi17 ? n32 : n59755;
  assign n59757 = pi16 ? n1683 : ~n59756;
  assign n59758 = pi15 ? n19503 : n59757;
  assign n59759 = pi14 ? n43466 : n59758;
  assign n59760 = pi13 ? n21119 : n59759;
  assign n59761 = pi19 ? n358 : n6303;
  assign n59762 = pi18 ? n17927 : ~n59761;
  assign n59763 = pi17 ? n32 : n59762;
  assign n59764 = pi17 ? n19432 : n31057;
  assign n59765 = pi16 ? n59763 : ~n59764;
  assign n59766 = pi15 ? n59765 : n32185;
  assign n59767 = pi20 ? n2358 : n18762;
  assign n59768 = pi19 ? n59767 : n18540;
  assign n59769 = pi18 ? n341 : n59768;
  assign n59770 = pi17 ? n32 : n59769;
  assign n59771 = pi20 ? n18540 : n266;
  assign n59772 = pi19 ? n59771 : ~n45863;
  assign n59773 = pi20 ? n5854 : ~n18129;
  assign n59774 = pi19 ? n59773 : ~n349;
  assign n59775 = pi18 ? n59772 : ~n59774;
  assign n59776 = pi17 ? n59775 : ~n57390;
  assign n59777 = pi16 ? n59770 : n59776;
  assign n59778 = pi15 ? n59777 : n31687;
  assign n59779 = pi14 ? n59766 : n59778;
  assign n59780 = pi13 ? n45291 : n59779;
  assign n59781 = pi12 ? n59760 : n59780;
  assign n59782 = pi11 ? n59754 : n59781;
  assign n59783 = pi10 ? n59741 : n59782;
  assign n59784 = pi09 ? n59709 : n59783;
  assign n59785 = pi14 ? n32 : n14613;
  assign n59786 = pi13 ? n32 : n59785;
  assign n59787 = pi12 ? n32 : n59786;
  assign n59788 = pi11 ? n32 : n59787;
  assign n59789 = pi10 ? n32 : n59788;
  assign n59790 = pi15 ? n59712 : n20836;
  assign n59791 = pi14 ? n21553 : n59790;
  assign n59792 = pi20 ? n321 : n1475;
  assign n59793 = pi19 ? n59792 : ~n32;
  assign n59794 = pi18 ? n32 : ~n59793;
  assign n59795 = pi17 ? n32 : n59794;
  assign n59796 = pi16 ? n32 : n59795;
  assign n59797 = pi15 ? n32 : n59796;
  assign n59798 = pi16 ? n1471 : ~n2293;
  assign n59799 = pi16 ? n1214 : ~n2293;
  assign n59800 = pi15 ? n59798 : n59799;
  assign n59801 = pi14 ? n59797 : n59800;
  assign n59802 = pi13 ? n59791 : n59801;
  assign n59803 = pi14 ? n34146 : n21326;
  assign n59804 = pi15 ? n13943 : n21033;
  assign n59805 = pi14 ? n59804 : n21035;
  assign n59806 = pi13 ? n59803 : n59805;
  assign n59807 = pi12 ? n59802 : n59806;
  assign n59808 = pi15 ? n21141 : n20831;
  assign n59809 = pi14 ? n20969 : n59808;
  assign n59810 = pi18 ? n4428 : ~n605;
  assign n59811 = pi17 ? n32 : n59810;
  assign n59812 = pi16 ? n32 : n59811;
  assign n59813 = pi15 ? n45216 : n59812;
  assign n59814 = pi15 ? n45049 : n22036;
  assign n59815 = pi14 ? n59813 : n59814;
  assign n59816 = pi13 ? n59809 : n59815;
  assign n59817 = pi15 ? n31788 : n59734;
  assign n59818 = pi14 ? n45339 : n59817;
  assign n59819 = pi15 ? n12091 : n45345;
  assign n59820 = pi14 ? n59819 : n32;
  assign n59821 = pi13 ? n59818 : n59820;
  assign n59822 = pi12 ? n59816 : n59821;
  assign n59823 = pi11 ? n59807 : n59822;
  assign n59824 = pi15 ? n59670 : n31526;
  assign n59825 = pi18 ? n940 : ~n20474;
  assign n59826 = pi17 ? n32 : n59825;
  assign n59827 = pi16 ? n1233 : ~n59826;
  assign n59828 = pi15 ? n31526 : n59827;
  assign n59829 = pi14 ? n59824 : n59828;
  assign n59830 = pi13 ? n32 : n59829;
  assign n59831 = pi20 ? n1385 : ~n339;
  assign n59832 = pi19 ? n59831 : n32;
  assign n59833 = pi18 ? n21066 : ~n59832;
  assign n59834 = pi17 ? n32 : n59833;
  assign n59835 = pi16 ? n1233 : ~n59834;
  assign n59836 = pi15 ? n59835 : n46774;
  assign n59837 = pi14 ? n59836 : n47262;
  assign n59838 = pi15 ? n59394 : n21079;
  assign n59839 = pi14 ? n59838 : n21190;
  assign n59840 = pi13 ? n59837 : n59839;
  assign n59841 = pi12 ? n59830 : n59840;
  assign n59842 = pi15 ? n180 : n20538;
  assign n59843 = pi18 ? n6118 : n20345;
  assign n59844 = pi17 ? n32 : n59843;
  assign n59845 = pi16 ? n1683 : ~n59844;
  assign n59846 = pi15 ? n19503 : n59845;
  assign n59847 = pi14 ? n59842 : n59846;
  assign n59848 = pi13 ? n21203 : n59847;
  assign n59849 = pi17 ? n31691 : ~n2319;
  assign n59850 = pi16 ? n32 : n59849;
  assign n59851 = pi15 ? n59850 : n31864;
  assign n59852 = pi14 ? n59851 : n45367;
  assign n59853 = pi16 ? n1135 : ~n31058;
  assign n59854 = pi16 ? n1233 : ~n57281;
  assign n59855 = pi15 ? n59853 : n59854;
  assign n59856 = pi19 ? n22038 : n11107;
  assign n59857 = pi18 ? n341 : n59856;
  assign n59858 = pi17 ? n32 : n59857;
  assign n59859 = pi20 ? n11107 : n266;
  assign n59860 = pi20 ? n207 : n501;
  assign n59861 = pi19 ? n59859 : ~n59860;
  assign n59862 = pi20 ? n18261 : n32;
  assign n59863 = pi19 ? n59862 : n349;
  assign n59864 = pi18 ? n59861 : n59863;
  assign n59865 = pi17 ? n59864 : ~n57390;
  assign n59866 = pi16 ? n59858 : n59865;
  assign n59867 = pi15 ? n59866 : n31687;
  assign n59868 = pi14 ? n59855 : n59867;
  assign n59869 = pi13 ? n59852 : n59868;
  assign n59870 = pi12 ? n59848 : n59869;
  assign n59871 = pi11 ? n59841 : n59870;
  assign n59872 = pi10 ? n59823 : n59871;
  assign n59873 = pi09 ? n59789 : n59872;
  assign n59874 = pi08 ? n59784 : n59873;
  assign n59875 = pi07 ? n59704 : n59874;
  assign n59876 = pi14 ? n32 : n658;
  assign n59877 = pi13 ? n32 : n59876;
  assign n59878 = pi12 ? n32 : n59877;
  assign n59879 = pi11 ? n32 : n59878;
  assign n59880 = pi10 ? n32 : n59879;
  assign n59881 = pi15 ? n14613 : n59654;
  assign n59882 = pi19 ? n57844 : n3495;
  assign n59883 = pi20 ? n18834 : n7487;
  assign n59884 = pi19 ? n59883 : n32;
  assign n59885 = pi18 ? n59882 : n59884;
  assign n59886 = pi17 ? n19529 : n59885;
  assign n59887 = pi16 ? n32 : n59886;
  assign n59888 = pi20 ? n207 : ~n7487;
  assign n59889 = pi19 ? n59888 : ~n32;
  assign n59890 = pi18 ? n32 : ~n59889;
  assign n59891 = pi17 ? n32 : n59890;
  assign n59892 = pi16 ? n32 : n59891;
  assign n59893 = pi15 ? n59887 : n59892;
  assign n59894 = pi14 ? n59881 : n59893;
  assign n59895 = pi20 ? n207 : ~n439;
  assign n59896 = pi19 ? n59895 : ~n32;
  assign n59897 = pi18 ? n32 : ~n59896;
  assign n59898 = pi17 ? n32 : n59897;
  assign n59899 = pi16 ? n32 : n59898;
  assign n59900 = pi15 ? n59899 : n47471;
  assign n59901 = pi16 ? n1233 : ~n2293;
  assign n59902 = pi15 ? n59799 : n59901;
  assign n59903 = pi14 ? n59900 : n59902;
  assign n59904 = pi13 ? n59894 : n59903;
  assign n59905 = pi15 ? n34044 : n32;
  assign n59906 = pi14 ? n59905 : n21326;
  assign n59907 = pi15 ? n13943 : n14397;
  assign n59908 = pi14 ? n59907 : n21217;
  assign n59909 = pi13 ? n59906 : n59908;
  assign n59910 = pi12 ? n59904 : n59909;
  assign n59911 = pi19 ? n32 : n17669;
  assign n59912 = pi18 ? n59911 : n19194;
  assign n59913 = pi17 ? n32 : n59912;
  assign n59914 = pi16 ? n32 : n59913;
  assign n59915 = pi15 ? n59914 : n22167;
  assign n59916 = pi14 ? n32 : n59915;
  assign n59917 = pi13 ? n59916 : n45441;
  assign n59918 = pi18 ? n8819 : ~n605;
  assign n59919 = pi17 ? n32 : n59918;
  assign n59920 = pi16 ? n32 : n59919;
  assign n59921 = pi15 ? n59920 : n32;
  assign n59922 = pi20 ? n32 : n52880;
  assign n59923 = pi19 ? n59922 : ~n32;
  assign n59924 = pi18 ? n880 : ~n59923;
  assign n59925 = pi17 ? n32 : n59924;
  assign n59926 = pi16 ? n32 : n59925;
  assign n59927 = pi15 ? n32219 : n59926;
  assign n59928 = pi14 ? n59921 : n59927;
  assign n59929 = pi15 ? n45812 : n13948;
  assign n59930 = pi14 ? n59929 : n21558;
  assign n59931 = pi13 ? n59928 : n59930;
  assign n59932 = pi12 ? n59917 : n59931;
  assign n59933 = pi11 ? n59910 : n59932;
  assign n59934 = pi14 ? n32 : n31120;
  assign n59935 = pi15 ? n31146 : n30941;
  assign n59936 = pi20 ? n266 : n481;
  assign n59937 = pi19 ? n59936 : n32;
  assign n59938 = pi18 ? n21255 : ~n59937;
  assign n59939 = pi17 ? n32 : n59938;
  assign n59940 = pi16 ? n1135 : ~n59939;
  assign n59941 = pi15 ? n30941 : n59940;
  assign n59942 = pi14 ? n59935 : n59941;
  assign n59943 = pi13 ? n59934 : n59942;
  assign n59944 = pi18 ? n32 : n1349;
  assign n59945 = pi17 ? n32 : n59944;
  assign n59946 = pi16 ? n1135 : ~n59945;
  assign n59947 = pi15 ? n46774 : n35359;
  assign n59948 = pi14 ? n59946 : n59947;
  assign n59949 = pi15 ? n35359 : n21268;
  assign n59950 = pi14 ? n59949 : n21278;
  assign n59951 = pi13 ? n59948 : n59950;
  assign n59952 = pi12 ? n59943 : n59951;
  assign n59953 = pi15 ? n21302 : n180;
  assign n59954 = pi14 ? n21291 : n59953;
  assign n59955 = pi18 ? n268 : n32061;
  assign n59956 = pi17 ? n32 : n59955;
  assign n59957 = pi17 ? n19170 : n20313;
  assign n59958 = pi16 ? n59956 : n59957;
  assign n59959 = pi15 ? n180 : n59958;
  assign n59960 = pi18 ? n32 : n32061;
  assign n59961 = pi17 ? n32 : n59960;
  assign n59962 = pi19 ? n17766 : ~n18502;
  assign n59963 = pi18 ? n59962 : ~n58856;
  assign n59964 = pi17 ? n19170 : n59963;
  assign n59965 = pi16 ? n59961 : n59964;
  assign n59966 = pi16 ? n45482 : ~n1934;
  assign n59967 = pi15 ? n59965 : n59966;
  assign n59968 = pi14 ? n59959 : n59967;
  assign n59969 = pi13 ? n59954 : n59968;
  assign n59970 = pi21 ? n405 : ~n85;
  assign n59971 = pi20 ? n59970 : ~n32;
  assign n59972 = pi19 ? n59971 : ~n32;
  assign n59973 = pi18 ? n32 : n59972;
  assign n59974 = pi17 ? n32 : n59973;
  assign n59975 = pi16 ? n1233 : ~n59974;
  assign n59976 = pi17 ? n45514 : n57514;
  assign n59977 = pi16 ? n1233 : ~n59976;
  assign n59978 = pi15 ? n59975 : n59977;
  assign n59979 = pi17 ? n45518 : ~n2537;
  assign n59980 = pi16 ? n32 : n59979;
  assign n59981 = pi17 ? n18017 : n3337;
  assign n59982 = pi16 ? n45587 : ~n59981;
  assign n59983 = pi15 ? n59980 : n59982;
  assign n59984 = pi14 ? n59978 : n59983;
  assign n59985 = pi13 ? n45512 : n59984;
  assign n59986 = pi12 ? n59969 : n59985;
  assign n59987 = pi11 ? n59952 : n59986;
  assign n59988 = pi10 ? n59933 : n59987;
  assign n59989 = pi09 ? n59880 : n59988;
  assign n59990 = pi14 ? n32 : n21319;
  assign n59991 = pi13 ? n32 : n59990;
  assign n59992 = pi12 ? n32 : n59991;
  assign n59993 = pi11 ? n32 : n59992;
  assign n59994 = pi10 ? n32 : n59993;
  assign n59995 = pi16 ? n1471 : ~n3769;
  assign n59996 = pi15 ? n32 : n59995;
  assign n59997 = pi14 ? n59996 : n59893;
  assign n59998 = pi17 ? n32 : n2868;
  assign n59999 = pi16 ? n1214 : ~n59998;
  assign n60000 = pi15 ? n59899 : n59999;
  assign n60001 = pi15 ? n48747 : n47710;
  assign n60002 = pi14 ? n60000 : n60001;
  assign n60003 = pi13 ? n59997 : n60002;
  assign n60004 = pi15 ? n34044 : n21319;
  assign n60005 = pi14 ? n60004 : n32128;
  assign n60006 = pi13 ? n60005 : n59908;
  assign n60007 = pi12 ? n60003 : n60006;
  assign n60008 = pi20 ? n310 : ~n11048;
  assign n60009 = pi19 ? n60008 : n32;
  assign n60010 = pi18 ? n50152 : n60009;
  assign n60011 = pi17 ? n32 : n60010;
  assign n60012 = pi16 ? n32 : n60011;
  assign n60013 = pi15 ? n60012 : n22167;
  assign n60014 = pi14 ? n21326 : n60013;
  assign n60015 = pi13 ? n60014 : n45441;
  assign n60016 = pi14 ? n59921 : n32219;
  assign n60017 = pi19 ? n39001 : n32;
  assign n60018 = pi18 ? n863 : n60017;
  assign n60019 = pi17 ? n32 : n60018;
  assign n60020 = pi16 ? n32 : n60019;
  assign n60021 = pi15 ? n60020 : n13952;
  assign n60022 = pi14 ? n60021 : n21558;
  assign n60023 = pi13 ? n60016 : n60022;
  assign n60024 = pi12 ? n60015 : n60023;
  assign n60025 = pi11 ? n60007 : n60024;
  assign n60026 = pi15 ? n31146 : n29601;
  assign n60027 = pi18 ? n21255 : ~n21330;
  assign n60028 = pi17 ? n32 : n60027;
  assign n60029 = pi16 ? n1233 : ~n60028;
  assign n60030 = pi15 ? n29601 : n60029;
  assign n60031 = pi14 ? n60026 : n60030;
  assign n60032 = pi13 ? n59934 : n60031;
  assign n60033 = pi16 ? n1233 : ~n2426;
  assign n60034 = pi15 ? n60033 : n46655;
  assign n60035 = pi14 ? n60034 : n46774;
  assign n60036 = pi15 ? n35162 : n21268;
  assign n60037 = pi14 ? n60036 : n21278;
  assign n60038 = pi13 ? n60035 : n60037;
  assign n60039 = pi12 ? n60032 : n60038;
  assign n60040 = pi18 ? n21299 : n20525;
  assign n60041 = pi17 ? n21298 : ~n60040;
  assign n60042 = pi16 ? n21294 : n60041;
  assign n60043 = pi15 ? n60042 : n13392;
  assign n60044 = pi14 ? n21366 : n60043;
  assign n60045 = pi17 ? n19170 : n178;
  assign n60046 = pi16 ? n59956 : n60045;
  assign n60047 = pi15 ? n20136 : n60046;
  assign n60048 = pi20 ? n16008 : ~n32;
  assign n60049 = pi19 ? n60048 : ~n32;
  assign n60050 = pi18 ? n59962 : ~n60049;
  assign n60051 = pi17 ? n19170 : n60050;
  assign n60052 = pi16 ? n59961 : n60051;
  assign n60053 = pi15 ? n60052 : n59966;
  assign n60054 = pi14 ? n60047 : n60053;
  assign n60055 = pi13 ? n60044 : n60054;
  assign n60056 = pi17 ? n45490 : ~n1933;
  assign n60057 = pi16 ? n23483 : n60056;
  assign n60058 = pi15 ? n60057 : n45497;
  assign n60059 = pi14 ? n60058 : n45581;
  assign n60060 = pi19 ? n6652 : ~n32;
  assign n60061 = pi18 ? n32 : n60060;
  assign n60062 = pi17 ? n45514 : n60061;
  assign n60063 = pi16 ? n1233 : ~n60062;
  assign n60064 = pi15 ? n59975 : n60063;
  assign n60065 = pi14 ? n60064 : n59983;
  assign n60066 = pi13 ? n60059 : n60065;
  assign n60067 = pi12 ? n60055 : n60066;
  assign n60068 = pi11 ? n60039 : n60067;
  assign n60069 = pi10 ? n60025 : n60068;
  assign n60070 = pi09 ? n59994 : n60069;
  assign n60071 = pi08 ? n59989 : n60070;
  assign n60072 = pi15 ? n21464 : n21389;
  assign n60073 = pi14 ? n32 : n60072;
  assign n60074 = pi13 ? n32 : n60073;
  assign n60075 = pi12 ? n32 : n60074;
  assign n60076 = pi11 ? n32 : n60075;
  assign n60077 = pi10 ? n32 : n60076;
  assign n60078 = pi20 ? n32 : n9667;
  assign n60079 = pi19 ? n60078 : ~n32;
  assign n60080 = pi18 ? n32 : n60079;
  assign n60081 = pi17 ? n32 : n60080;
  assign n60082 = pi16 ? n31442 : ~n60081;
  assign n60083 = pi15 ? n32 : n60082;
  assign n60084 = pi19 ? n32 : n35481;
  assign n60085 = pi18 ? n32 : n60084;
  assign n60086 = pi17 ? n32 : n60085;
  assign n60087 = pi20 ? n428 : n11107;
  assign n60088 = pi19 ? n36181 : ~n60087;
  assign n60089 = pi20 ? n5854 : n17652;
  assign n60090 = pi19 ? n6314 : n60089;
  assign n60091 = pi18 ? n60088 : ~n60090;
  assign n60092 = pi20 ? n310 : ~n501;
  assign n60093 = pi19 ? n60092 : ~n17652;
  assign n60094 = pi18 ? n60093 : ~n41055;
  assign n60095 = pi17 ? n60091 : ~n60094;
  assign n60096 = pi16 ? n60086 : ~n60095;
  assign n60097 = pi15 ? n14397 : n60096;
  assign n60098 = pi14 ? n60083 : n60097;
  assign n60099 = pi15 ? n32692 : n59999;
  assign n60100 = pi14 ? n60099 : n47710;
  assign n60101 = pi13 ? n60098 : n60100;
  assign n60102 = pi15 ? n34146 : n21319;
  assign n60103 = pi14 ? n60102 : n32128;
  assign n60104 = pi15 ? n13943 : n21389;
  assign n60105 = pi14 ? n60104 : n21391;
  assign n60106 = pi13 ? n60103 : n60105;
  assign n60107 = pi12 ? n60101 : n60106;
  assign n60108 = pi15 ? n11654 : n45640;
  assign n60109 = pi14 ? n32 : n60108;
  assign n60110 = pi13 ? n60109 : n45648;
  assign n60111 = pi18 ? n880 : ~n32919;
  assign n60112 = pi17 ? n32 : n60111;
  assign n60113 = pi16 ? n32 : n60112;
  assign n60114 = pi15 ? n34679 : n60113;
  assign n60115 = pi14 ? n45653 : n60114;
  assign n60116 = pi15 ? n60020 : n20831;
  assign n60117 = pi14 ? n60116 : n59545;
  assign n60118 = pi13 ? n60115 : n60117;
  assign n60119 = pi12 ? n60110 : n60118;
  assign n60120 = pi11 ? n60107 : n60119;
  assign n60121 = pi18 ? n16316 : n350;
  assign n60122 = pi17 ? n32 : n60121;
  assign n60123 = pi16 ? n1135 : ~n60122;
  assign n60124 = pi20 ? n2385 : ~n357;
  assign n60125 = pi19 ? n60124 : ~n32;
  assign n60126 = pi18 ? n21414 : n60125;
  assign n60127 = pi17 ? n32 : n60126;
  assign n60128 = pi16 ? n1135 : ~n60127;
  assign n60129 = pi15 ? n60123 : n60128;
  assign n60130 = pi14 ? n30941 : n60129;
  assign n60131 = pi13 ? n32 : n60130;
  assign n60132 = pi15 ? n46774 : n58837;
  assign n60133 = pi14 ? n46991 : n60132;
  assign n60134 = pi19 ? n30699 : n43441;
  assign n60135 = pi18 ? n28748 : ~n60134;
  assign n60136 = pi17 ? n32 : n60135;
  assign n60137 = pi19 ? n2180 : n18133;
  assign n60138 = pi19 ? n6050 : n30984;
  assign n60139 = pi18 ? n60137 : ~n60138;
  assign n60140 = pi18 ? n45670 : ~n44610;
  assign n60141 = pi17 ? n60139 : n60140;
  assign n60142 = pi16 ? n60136 : ~n60141;
  assign n60143 = pi15 ? n60142 : n21431;
  assign n60144 = pi14 ? n60143 : n21439;
  assign n60145 = pi13 ? n60133 : n60144;
  assign n60146 = pi12 ? n60131 : n60145;
  assign n60147 = pi15 ? n180 : n19969;
  assign n60148 = pi14 ? n21450 : n60147;
  assign n60149 = pi19 ? n207 : n8818;
  assign n60150 = pi18 ? n60149 : ~n20020;
  assign n60151 = pi18 ? n237 : ~n177;
  assign n60152 = pi17 ? n60150 : ~n60151;
  assign n60153 = pi16 ? n45692 : n60152;
  assign n60154 = pi15 ? n19969 : n60153;
  assign n60155 = pi17 ? n13946 : n2410;
  assign n60156 = pi16 ? n45699 : ~n60155;
  assign n60157 = pi15 ? n60156 : n45707;
  assign n60158 = pi14 ? n60154 : n60157;
  assign n60159 = pi13 ? n60148 : n60158;
  assign n60160 = pi18 ? n366 : ~n32337;
  assign n60161 = pi17 ? n32 : n60160;
  assign n60162 = pi20 ? n749 : n339;
  assign n60163 = pi19 ? n19596 : ~n60162;
  assign n60164 = pi19 ? n18200 : ~n8818;
  assign n60165 = pi18 ? n60163 : n60164;
  assign n60166 = pi18 ? n45747 : ~n20355;
  assign n60167 = pi17 ? n60165 : n60166;
  assign n60168 = pi16 ? n60161 : ~n60167;
  assign n60169 = pi15 ? n45572 : n60168;
  assign n60170 = pi20 ? n56060 : ~n32;
  assign n60171 = pi19 ? n60170 : ~n32;
  assign n60172 = pi18 ? n32 : n60171;
  assign n60173 = pi17 ? n45752 : ~n60172;
  assign n60174 = pi16 ? n32 : n60173;
  assign n60175 = pi18 ? n32 : n45755;
  assign n60176 = pi17 ? n32 : n60175;
  assign n60177 = pi16 ? n60176 : ~n45525;
  assign n60178 = pi15 ? n60174 : n60177;
  assign n60179 = pi14 ? n60169 : n60178;
  assign n60180 = pi13 ? n45733 : n60179;
  assign n60181 = pi12 ? n60159 : n60180;
  assign n60182 = pi11 ? n60146 : n60181;
  assign n60183 = pi10 ? n60120 : n60182;
  assign n60184 = pi09 ? n60077 : n60183;
  assign n60185 = pi18 ? n32 : n54044;
  assign n60186 = pi17 ? n32 : n60185;
  assign n60187 = pi16 ? n1214 : ~n60186;
  assign n60188 = pi15 ? n32692 : n60187;
  assign n60189 = pi16 ? n1135 : ~n2756;
  assign n60190 = pi16 ? n1233 : ~n3769;
  assign n60191 = pi15 ? n60189 : n60190;
  assign n60192 = pi14 ? n60188 : n60191;
  assign n60193 = pi13 ? n60098 : n60192;
  assign n60194 = pi15 ? n60190 : n21464;
  assign n60195 = pi14 ? n60194 : n21467;
  assign n60196 = pi15 ? n14156 : n21464;
  assign n60197 = pi14 ? n60196 : n21391;
  assign n60198 = pi13 ? n60195 : n60197;
  assign n60199 = pi12 ? n60193 : n60198;
  assign n60200 = pi14 ? n32128 : n60108;
  assign n60201 = pi13 ? n60200 : n45801;
  assign n60202 = pi21 ? n11402 : ~n32;
  assign n60203 = pi20 ? n32 : n60202;
  assign n60204 = pi19 ? n60203 : ~n32;
  assign n60205 = pi18 ? n880 : ~n60204;
  assign n60206 = pi17 ? n32 : n60205;
  assign n60207 = pi16 ? n32 : n60206;
  assign n60208 = pi15 ? n32219 : n60207;
  assign n60209 = pi14 ? n45806 : n60208;
  assign n60210 = pi20 ? n266 : n7487;
  assign n60211 = pi19 ? n60210 : n32;
  assign n60212 = pi18 ? n863 : n60211;
  assign n60213 = pi17 ? n32 : n60212;
  assign n60214 = pi16 ? n32 : n60213;
  assign n60215 = pi15 ? n60214 : n32;
  assign n60216 = pi14 ? n60215 : n21558;
  assign n60217 = pi13 ? n60209 : n60216;
  assign n60218 = pi12 ? n60201 : n60217;
  assign n60219 = pi11 ? n60199 : n60218;
  assign n60220 = pi20 ? n321 : ~n52;
  assign n60221 = pi19 ? n60220 : ~n32;
  assign n60222 = pi18 ? n16316 : n60221;
  assign n60223 = pi17 ? n32 : n60222;
  assign n60224 = pi16 ? n1233 : ~n60223;
  assign n60225 = pi20 ? n2385 : n1940;
  assign n60226 = pi19 ? n60225 : ~n32;
  assign n60227 = pi18 ? n21414 : n60226;
  assign n60228 = pi17 ? n32 : n60227;
  assign n60229 = pi16 ? n1233 : ~n60228;
  assign n60230 = pi15 ? n60224 : n60229;
  assign n60231 = pi14 ? n29601 : n60230;
  assign n60232 = pi13 ? n32 : n60231;
  assign n60233 = pi18 ? n1395 : ~n32247;
  assign n60234 = pi17 ? n32 : n60233;
  assign n60235 = pi19 ? n175 : n32;
  assign n60236 = pi20 ? n32 : ~n18415;
  assign n60237 = pi19 ? n32 : n60236;
  assign n60238 = pi18 ? n60235 : n60237;
  assign n60239 = pi18 ? n359 : n2424;
  assign n60240 = pi17 ? n60238 : n60239;
  assign n60241 = pi16 ? n60234 : ~n60240;
  assign n60242 = pi15 ? n60033 : n60241;
  assign n60243 = pi14 ? n60242 : n46655;
  assign n60244 = pi20 ? n448 : ~n501;
  assign n60245 = pi20 ? n501 : ~n448;
  assign n60246 = pi19 ? n60244 : ~n60245;
  assign n60247 = pi18 ? n1613 : n60246;
  assign n60248 = pi17 ? n32 : n60247;
  assign n60249 = pi19 ? n448 : n45824;
  assign n60250 = pi20 ? n310 : n1331;
  assign n60251 = pi19 ? n45826 : n60250;
  assign n60252 = pi18 ? n60249 : n60251;
  assign n60253 = pi18 ? n45832 : n13080;
  assign n60254 = pi17 ? n60252 : n60253;
  assign n60255 = pi16 ? n60248 : n60254;
  assign n60256 = pi15 ? n60255 : n21268;
  assign n60257 = pi15 ? n21273 : n21438;
  assign n60258 = pi14 ? n60256 : n60257;
  assign n60259 = pi13 ? n60243 : n60258;
  assign n60260 = pi12 ? n60232 : n60259;
  assign n60261 = pi18 ? n21443 : ~n532;
  assign n60262 = pi17 ? n32 : n60261;
  assign n60263 = pi16 ? n32 : n60262;
  assign n60264 = pi15 ? n60263 : n21449;
  assign n60265 = pi20 ? n13674 : n32;
  assign n60266 = pi19 ? n60265 : n32;
  assign n60267 = pi18 ? n32 : n60266;
  assign n60268 = pi17 ? n32 : n60267;
  assign n60269 = pi16 ? n32 : n60268;
  assign n60270 = pi15 ? n180 : n60269;
  assign n60271 = pi14 ? n60264 : n60270;
  assign n60272 = pi18 ? n237 : ~n69;
  assign n60273 = pi17 ? n60150 : ~n60272;
  assign n60274 = pi16 ? n45692 : n60273;
  assign n60275 = pi15 ? n20048 : n60274;
  assign n60276 = pi16 ? n45849 : ~n60155;
  assign n60277 = pi17 ? n45705 : ~n2305;
  assign n60278 = pi16 ? n45704 : n60277;
  assign n60279 = pi15 ? n60276 : n60278;
  assign n60280 = pi14 ? n60275 : n60279;
  assign n60281 = pi13 ? n60271 : n60280;
  assign n60282 = pi17 ? n45712 : ~n2305;
  assign n60283 = pi16 ? n32 : n60282;
  assign n60284 = pi15 ? n60283 : n45855;
  assign n60285 = pi14 ? n60284 : n45732;
  assign n60286 = pi18 ? n1190 : ~n32337;
  assign n60287 = pi17 ? n32 : n60286;
  assign n60288 = pi20 ? n749 : n314;
  assign n60289 = pi19 ? n19596 : ~n60288;
  assign n60290 = pi19 ? n32443 : ~n8818;
  assign n60291 = pi18 ? n60289 : n60290;
  assign n60292 = pi17 ? n60291 : n60166;
  assign n60293 = pi16 ? n60287 : ~n60292;
  assign n60294 = pi15 ? n45572 : n60293;
  assign n60295 = pi14 ? n60294 : n60178;
  assign n60296 = pi13 ? n60285 : n60295;
  assign n60297 = pi12 ? n60281 : n60296;
  assign n60298 = pi11 ? n60260 : n60297;
  assign n60299 = pi10 ? n60219 : n60298;
  assign n60300 = pi09 ? n60077 : n60299;
  assign n60301 = pi08 ? n60184 : n60300;
  assign n60302 = pi07 ? n60071 : n60301;
  assign n60303 = pi06 ? n59875 : n60302;
  assign n60304 = pi05 ? n59544 : n60303;
  assign n60305 = pi04 ? n58671 : n60304;
  assign n60306 = pi03 ? n57135 : n60305;
  assign n60307 = pi14 ? n32 : n21543;
  assign n60308 = pi13 ? n32 : n60307;
  assign n60309 = pi12 ? n32 : n60308;
  assign n60310 = pi11 ? n32 : n60309;
  assign n60311 = pi10 ? n32 : n60310;
  assign n60312 = pi19 ? n30040 : ~n30044;
  assign n60313 = pi18 ? n18908 : n60312;
  assign n60314 = pi17 ? n32 : n60313;
  assign n60315 = pi20 ? n310 : ~n18408;
  assign n60316 = pi19 ? n60315 : n17652;
  assign n60317 = pi18 ? n56247 : ~n60316;
  assign n60318 = pi20 ? n310 : ~n17652;
  assign n60319 = pi19 ? n60318 : ~n17652;
  assign n60320 = pi20 ? n18624 : ~n207;
  assign n60321 = pi19 ? n60320 : n32;
  assign n60322 = pi18 ? n60319 : ~n60321;
  assign n60323 = pi17 ? n60317 : ~n60322;
  assign n60324 = pi16 ? n60314 : n60323;
  assign n60325 = pi20 ? n6085 : ~n2180;
  assign n60326 = pi19 ? n60325 : ~n30040;
  assign n60327 = pi18 ? n4380 : n60326;
  assign n60328 = pi17 ? n32 : n60327;
  assign n60329 = pi19 ? n30044 : ~n501;
  assign n60330 = pi20 ? n5854 : ~n1331;
  assign n60331 = pi19 ? n60330 : n2180;
  assign n60332 = pi18 ? n60329 : ~n60331;
  assign n60333 = pi19 ? n29294 : ~n17669;
  assign n60334 = pi20 ? n310 : ~n10889;
  assign n60335 = pi19 ? n60334 : n32;
  assign n60336 = pi18 ? n60333 : ~n60335;
  assign n60337 = pi17 ? n60332 : ~n60336;
  assign n60338 = pi16 ? n60328 : n60337;
  assign n60339 = pi15 ? n60324 : n60338;
  assign n60340 = pi20 ? n3523 : n17671;
  assign n60341 = pi19 ? n60340 : n28481;
  assign n60342 = pi18 ? n32 : n60341;
  assign n60343 = pi17 ? n32 : n60342;
  assign n60344 = pi19 ? n41134 : n267;
  assign n60345 = pi19 ? n6314 : n274;
  assign n60346 = pi18 ? n60344 : n60345;
  assign n60347 = pi19 ? n22591 : n18129;
  assign n60348 = pi20 ? n12884 : n7388;
  assign n60349 = pi19 ? n60348 : n32;
  assign n60350 = pi18 ? n60347 : n60349;
  assign n60351 = pi17 ? n60346 : n60350;
  assign n60352 = pi16 ? n60343 : n60351;
  assign n60353 = pi15 ? n60352 : n21695;
  assign n60354 = pi14 ? n60339 : n60353;
  assign n60355 = pi19 ? n41233 : ~n502;
  assign n60356 = pi18 ? n312 : ~n60355;
  assign n60357 = pi17 ? n32 : n60356;
  assign n60358 = pi16 ? n60357 : ~n3769;
  assign n60359 = pi18 ? n936 : n350;
  assign n60360 = pi17 ? n32 : n60359;
  assign n60361 = pi16 ? n60360 : ~n3769;
  assign n60362 = pi15 ? n60358 : n60361;
  assign n60363 = pi17 ? n45886 : ~n21799;
  assign n60364 = pi16 ? n1135 : ~n60363;
  assign n60365 = pi17 ? n45886 : ~n14154;
  assign n60366 = pi16 ? n1135 : ~n60365;
  assign n60367 = pi15 ? n60364 : n60366;
  assign n60368 = pi14 ? n60362 : n60367;
  assign n60369 = pi13 ? n60354 : n60368;
  assign n60370 = pi18 ? n18402 : n45896;
  assign n60371 = pi17 ? n32 : n60370;
  assign n60372 = pi17 ? n45900 : n32;
  assign n60373 = pi16 ? n60371 : n60372;
  assign n60374 = pi15 ? n60373 : n21464;
  assign n60375 = pi14 ? n60374 : n21467;
  assign n60376 = pi13 ? n60375 : n21544;
  assign n60377 = pi12 ? n60369 : n60376;
  assign n60378 = pi18 ? n268 : ~n24344;
  assign n60379 = pi17 ? n32 : n60378;
  assign n60380 = pi16 ? n32 : n60379;
  assign n60381 = pi15 ? n32 : n60380;
  assign n60382 = pi14 ? n60381 : n45937;
  assign n60383 = pi13 ? n60382 : n45943;
  assign n60384 = pi20 ? n206 : ~n501;
  assign n60385 = pi19 ? n60384 : n32;
  assign n60386 = pi18 ? n863 : n60385;
  assign n60387 = pi17 ? n32 : n60386;
  assign n60388 = pi16 ? n32 : n60387;
  assign n60389 = pi15 ? n33020 : n60388;
  assign n60390 = pi14 ? n45948 : n60389;
  assign n60391 = pi14 ? n23063 : n22692;
  assign n60392 = pi13 ? n60390 : n60391;
  assign n60393 = pi12 ? n60383 : n60392;
  assign n60394 = pi11 ? n60377 : n60393;
  assign n60395 = pi14 ? n20844 : n20831;
  assign n60396 = pi20 ? n342 : ~n52;
  assign n60397 = pi19 ? n60396 : ~n32;
  assign n60398 = pi18 ? n32 : n60397;
  assign n60399 = pi17 ? n32 : n60398;
  assign n60400 = pi16 ? n1135 : ~n60399;
  assign n60401 = pi15 ? n60400 : n30941;
  assign n60402 = pi16 ? n1135 : ~n2415;
  assign n60403 = pi15 ? n31828 : n60402;
  assign n60404 = pi14 ? n60401 : n60403;
  assign n60405 = pi13 ? n60395 : n60404;
  assign n60406 = pi18 ? n42797 : n22705;
  assign n60407 = pi17 ? n32 : n60406;
  assign n60408 = pi16 ? n1135 : ~n60407;
  assign n60409 = pi15 ? n46441 : n60408;
  assign n60410 = pi14 ? n47256 : n60409;
  assign n60411 = pi13 ? n60410 : n21605;
  assign n60412 = pi12 ? n60405 : n60411;
  assign n60413 = pi15 ? n19805 : n19972;
  assign n60414 = pi14 ? n13375 : n60413;
  assign n60415 = pi18 ? n38127 : ~n4671;
  assign n60416 = pi17 ? n32 : n60415;
  assign n60417 = pi16 ? n1135 : ~n60416;
  assign n60418 = pi18 ? n6581 : n34724;
  assign n60419 = pi17 ? n32 : n60418;
  assign n60420 = pi16 ? n1214 : ~n60419;
  assign n60421 = pi15 ? n60417 : n60420;
  assign n60422 = pi15 ? n31828 : n45972;
  assign n60423 = pi14 ? n60421 : n60422;
  assign n60424 = pi13 ? n60414 : n60423;
  assign n60425 = pi18 ? n366 : ~n20164;
  assign n60426 = pi17 ? n32 : n60425;
  assign n60427 = pi19 ? n18678 : ~n4391;
  assign n60428 = pi18 ? n15241 : n60427;
  assign n60429 = pi17 ? n60428 : n2305;
  assign n60430 = pi16 ? n60426 : ~n60429;
  assign n60431 = pi18 ? n566 : n268;
  assign n60432 = pi17 ? n32 : n60431;
  assign n60433 = pi19 ? n20555 : ~n321;
  assign n60434 = pi18 ? n25760 : ~n60433;
  assign n60435 = pi17 ? n60434 : ~n1933;
  assign n60436 = pi16 ? n60432 : n60435;
  assign n60437 = pi15 ? n60430 : n60436;
  assign n60438 = pi19 ? n221 : n207;
  assign n60439 = pi18 ? n46003 : n60438;
  assign n60440 = pi21 ? n174 : ~n85;
  assign n60441 = pi20 ? n60440 : ~n32;
  assign n60442 = pi19 ? n60441 : ~n32;
  assign n60443 = pi18 ? n32 : n60442;
  assign n60444 = pi17 ? n60439 : ~n60443;
  assign n60445 = pi16 ? n46205 : n60444;
  assign n60446 = pi16 ? n15402 : n46012;
  assign n60447 = pi15 ? n60445 : n60446;
  assign n60448 = pi14 ? n60437 : n60447;
  assign n60449 = pi13 ? n45989 : n60448;
  assign n60450 = pi12 ? n60424 : n60449;
  assign n60451 = pi11 ? n60412 : n60450;
  assign n60452 = pi10 ? n60394 : n60451;
  assign n60453 = pi09 ? n60311 : n60452;
  assign n60454 = pi14 ? n32 : n21858;
  assign n60455 = pi13 ? n32 : n60454;
  assign n60456 = pi12 ? n32 : n60455;
  assign n60457 = pi11 ? n32 : n60456;
  assign n60458 = pi10 ? n32 : n60457;
  assign n60459 = pi19 ? n56743 : ~n56578;
  assign n60460 = pi18 ? n29364 : n60459;
  assign n60461 = pi17 ? n32 : n60460;
  assign n60462 = pi19 ? n56582 : n31723;
  assign n60463 = pi20 ? n310 : ~n18173;
  assign n60464 = pi19 ? n60463 : n333;
  assign n60465 = pi18 ? n60462 : n60464;
  assign n60466 = pi20 ? n3843 : ~n17652;
  assign n60467 = pi19 ? n60466 : n9488;
  assign n60468 = pi20 ? n17665 : n207;
  assign n60469 = pi19 ? n60468 : ~n32;
  assign n60470 = pi18 ? n60467 : n60469;
  assign n60471 = pi17 ? n60465 : n60470;
  assign n60472 = pi16 ? n60461 : ~n60471;
  assign n60473 = pi21 ? n7659 : ~n405;
  assign n60474 = pi20 ? n32 : n60473;
  assign n60475 = pi19 ? n32 : n60474;
  assign n60476 = pi20 ? n18282 : n1368;
  assign n60477 = pi19 ? n60476 : n42118;
  assign n60478 = pi18 ? n60475 : ~n60477;
  assign n60479 = pi17 ? n32 : n60478;
  assign n60480 = pi19 ? n30044 : ~n2180;
  assign n60481 = pi20 ? n5854 : n18253;
  assign n60482 = pi19 ? n60481 : n2180;
  assign n60483 = pi18 ? n60480 : ~n60482;
  assign n60484 = pi20 ? n5854 : ~n3695;
  assign n60485 = pi19 ? n60484 : ~n17669;
  assign n60486 = pi20 ? n310 : ~n53551;
  assign n60487 = pi19 ? n60486 : n32;
  assign n60488 = pi18 ? n60485 : ~n60487;
  assign n60489 = pi17 ? n60483 : ~n60488;
  assign n60490 = pi16 ? n60479 : n60489;
  assign n60491 = pi15 ? n60472 : n60490;
  assign n60492 = pi20 ? n1324 : n18253;
  assign n60493 = pi19 ? n60492 : n18409;
  assign n60494 = pi18 ? n32 : n60493;
  assign n60495 = pi17 ? n32 : n60494;
  assign n60496 = pi20 ? n18282 : n18540;
  assign n60497 = pi19 ? n28058 : ~n60496;
  assign n60498 = pi20 ? n354 : n18282;
  assign n60499 = pi19 ? n60498 : n18281;
  assign n60500 = pi18 ? n60497 : ~n60499;
  assign n60501 = pi20 ? n17652 : ~n1076;
  assign n60502 = pi19 ? n60501 : ~n18073;
  assign n60503 = pi20 ? n174 : ~n29949;
  assign n60504 = pi19 ? n60503 : ~n32;
  assign n60505 = pi18 ? n60502 : ~n60504;
  assign n60506 = pi17 ? n60500 : ~n60505;
  assign n60507 = pi16 ? n60495 : ~n60506;
  assign n60508 = pi18 ? n1370 : n359;
  assign n60509 = pi17 ? n32 : n60508;
  assign n60510 = pi16 ? n60509 : n21694;
  assign n60511 = pi15 ? n60507 : n60510;
  assign n60512 = pi14 ? n60491 : n60511;
  assign n60513 = pi19 ? n28823 : ~n315;
  assign n60514 = pi18 ? n41321 : ~n60513;
  assign n60515 = pi17 ? n32 : n60514;
  assign n60516 = pi16 ? n60515 : ~n3769;
  assign n60517 = pi18 ? n47993 : n30435;
  assign n60518 = pi17 ? n32 : n60517;
  assign n60519 = pi16 ? n60518 : ~n2518;
  assign n60520 = pi15 ? n60516 : n60519;
  assign n60521 = pi17 ? n45886 : ~n14150;
  assign n60522 = pi16 ? n1233 : ~n60521;
  assign n60523 = pi16 ? n1233 : ~n60363;
  assign n60524 = pi15 ? n60522 : n60523;
  assign n60525 = pi14 ? n60520 : n60524;
  assign n60526 = pi13 ? n60512 : n60525;
  assign n60527 = pi20 ? n974 : n1817;
  assign n60528 = pi19 ? n60527 : n56578;
  assign n60529 = pi18 ? n2197 : n60528;
  assign n60530 = pi17 ? n32 : n60529;
  assign n60531 = pi17 ? n42369 : n32;
  assign n60532 = pi16 ? n60530 : n60531;
  assign n60533 = pi15 ? n60532 : n387;
  assign n60534 = pi14 ? n60533 : n388;
  assign n60535 = pi13 ? n60534 : n32669;
  assign n60536 = pi12 ? n60526 : n60535;
  assign n60537 = pi20 ? n220 : ~n7388;
  assign n60538 = pi19 ? n60537 : ~n32;
  assign n60539 = pi18 ? n268 : ~n60538;
  assign n60540 = pi17 ? n32 : n60539;
  assign n60541 = pi16 ? n32 : n60540;
  assign n60542 = pi15 ? n21464 : n60541;
  assign n60543 = pi14 ? n60542 : n45937;
  assign n60544 = pi13 ? n60543 : n45943;
  assign n60545 = pi15 ? n32613 : n33020;
  assign n60546 = pi14 ? n45948 : n60545;
  assign n60547 = pi15 ? n21319 : n20836;
  assign n60548 = pi14 ? n60547 : n20969;
  assign n60549 = pi13 ? n60546 : n60548;
  assign n60550 = pi12 ? n60544 : n60549;
  assign n60551 = pi11 ? n60536 : n60550;
  assign n60552 = pi14 ? n20844 : n32;
  assign n60553 = pi15 ? n32021 : n30941;
  assign n60554 = pi19 ? n7604 : ~n32;
  assign n60555 = pi18 ? n32 : n60554;
  assign n60556 = pi17 ? n32 : n60555;
  assign n60557 = pi16 ? n1135 : ~n60556;
  assign n60558 = pi15 ? n60557 : n34146;
  assign n60559 = pi14 ? n60553 : n60558;
  assign n60560 = pi13 ? n60552 : n60559;
  assign n60561 = pi18 ? n42797 : n21257;
  assign n60562 = pi17 ? n32 : n60561;
  assign n60563 = pi16 ? n1135 : ~n60562;
  assign n60564 = pi15 ? n46991 : n60563;
  assign n60565 = pi14 ? n47256 : n60564;
  assign n60566 = pi13 ? n60565 : n21666;
  assign n60567 = pi12 ? n60560 : n60566;
  assign n60568 = pi15 ? n19805 : n20779;
  assign n60569 = pi14 ? n13375 : n60568;
  assign n60570 = pi18 ? n38127 : ~n20671;
  assign n60571 = pi17 ? n32 : n60570;
  assign n60572 = pi16 ? n1135 : ~n60571;
  assign n60573 = pi18 ? n6581 : n59276;
  assign n60574 = pi17 ? n32 : n60573;
  assign n60575 = pi16 ? n1214 : ~n60574;
  assign n60576 = pi15 ? n60572 : n60575;
  assign n60577 = pi15 ? n59394 : n46172;
  assign n60578 = pi14 ? n60576 : n60577;
  assign n60579 = pi13 ? n60569 : n60578;
  assign n60580 = pi17 ? n60439 : ~n3345;
  assign n60581 = pi16 ? n46205 : n60580;
  assign n60582 = pi17 ? n46011 : ~n45483;
  assign n60583 = pi16 ? n15402 : n60582;
  assign n60584 = pi15 ? n60581 : n60583;
  assign n60585 = pi14 ? n60437 : n60584;
  assign n60586 = pi13 ? n46068 : n60585;
  assign n60587 = pi12 ? n60579 : n60586;
  assign n60588 = pi11 ? n60567 : n60587;
  assign n60589 = pi10 ? n60551 : n60588;
  assign n60590 = pi09 ? n60458 : n60589;
  assign n60591 = pi08 ? n60453 : n60590;
  assign n60592 = pi15 ? n21786 : n21686;
  assign n60593 = pi14 ? n32 : n60592;
  assign n60594 = pi13 ? n32 : n60593;
  assign n60595 = pi12 ? n32 : n60594;
  assign n60596 = pi11 ? n32 : n60595;
  assign n60597 = pi10 ? n32 : n60596;
  assign n60598 = pi20 ? n9491 : ~n6822;
  assign n60599 = pi19 ? n43597 : n60598;
  assign n60600 = pi18 ? n32 : n60599;
  assign n60601 = pi17 ? n32 : n60600;
  assign n60602 = pi19 ? n56578 : n2019;
  assign n60603 = pi20 ? n1611 : n2019;
  assign n60604 = pi19 ? n60603 : ~n501;
  assign n60605 = pi18 ? n60602 : n60604;
  assign n60606 = pi20 ? n18762 : n974;
  assign n60607 = pi20 ? n974 : n1324;
  assign n60608 = pi19 ? n60606 : n60607;
  assign n60609 = pi20 ? n3843 : ~n266;
  assign n60610 = pi19 ? n60609 : ~n32;
  assign n60611 = pi18 ? n60608 : n60610;
  assign n60612 = pi17 ? n60605 : n60611;
  assign n60613 = pi16 ? n60601 : ~n60612;
  assign n60614 = pi19 ? n28161 : n1757;
  assign n60615 = pi18 ? n1139 : n60614;
  assign n60616 = pi17 ? n32 : n60615;
  assign n60617 = pi19 ? n4670 : ~n207;
  assign n60618 = pi18 ? n32 : n60617;
  assign n60619 = pi20 ? n32 : ~n58757;
  assign n60620 = pi19 ? n60619 : n32;
  assign n60621 = pi18 ? n4380 : n60620;
  assign n60622 = pi17 ? n60618 : n60621;
  assign n60623 = pi16 ? n60616 : n60622;
  assign n60624 = pi15 ? n60613 : n60623;
  assign n60625 = pi20 ? n175 : ~n18834;
  assign n60626 = pi20 ? n2019 : ~n18282;
  assign n60627 = pi19 ? n60625 : ~n60626;
  assign n60628 = pi18 ? n32 : n60627;
  assign n60629 = pi17 ? n32 : n60628;
  assign n60630 = pi20 ? n29457 : ~n29452;
  assign n60631 = pi20 ? n9641 : n18073;
  assign n60632 = pi19 ? n60630 : n60631;
  assign n60633 = pi20 ? n17669 : n9641;
  assign n60634 = pi19 ? n60633 : n406;
  assign n60635 = pi18 ? n60632 : n60634;
  assign n60636 = pi20 ? n1324 : n310;
  assign n60637 = pi19 ? n60636 : n18624;
  assign n60638 = pi20 ? n21111 : ~n1377;
  assign n60639 = pi19 ? n60638 : n32;
  assign n60640 = pi18 ? n60637 : ~n60639;
  assign n60641 = pi17 ? n60635 : n60640;
  assign n60642 = pi16 ? n60629 : ~n60641;
  assign n60643 = pi15 ? n60642 : n22381;
  assign n60644 = pi14 ? n60624 : n60643;
  assign n60645 = pi16 ? n2137 : ~n3769;
  assign n60646 = pi16 ? n1808 : ~n2518;
  assign n60647 = pi15 ? n60645 : n60646;
  assign n60648 = pi20 ? n17652 : n18282;
  assign n60649 = pi19 ? n60648 : n18782;
  assign n60650 = pi18 ? n29658 : n60649;
  assign n60651 = pi17 ? n32 : n60650;
  assign n60652 = pi20 ? n9194 : ~n321;
  assign n60653 = pi19 ? n60652 : n32;
  assign n60654 = pi18 ? n60653 : ~n350;
  assign n60655 = pi17 ? n60654 : n14150;
  assign n60656 = pi16 ? n60651 : n60655;
  assign n60657 = pi19 ? n9491 : ~n41340;
  assign n60658 = pi18 ? n42434 : n60657;
  assign n60659 = pi17 ? n32 : n60658;
  assign n60660 = pi19 ? n8562 : ~n32;
  assign n60661 = pi18 ? n60660 : n1353;
  assign n60662 = pi17 ? n60661 : ~n14154;
  assign n60663 = pi16 ? n60659 : ~n60662;
  assign n60664 = pi15 ? n60656 : n60663;
  assign n60665 = pi14 ? n60647 : n60664;
  assign n60666 = pi13 ? n60644 : n60665;
  assign n60667 = pi14 ? n21681 : n23466;
  assign n60668 = pi13 ? n60667 : n21688;
  assign n60669 = pi12 ? n60666 : n60668;
  assign n60670 = pi18 ? n356 : ~n23543;
  assign n60671 = pi17 ? n32 : n60670;
  assign n60672 = pi16 ? n32 : n60671;
  assign n60673 = pi15 ? n32 : n60672;
  assign n60674 = pi14 ? n60673 : n12079;
  assign n60675 = pi13 ? n60674 : n46147;
  assign n60676 = pi15 ? n21346 : n24213;
  assign n60677 = pi15 ? n46262 : n13948;
  assign n60678 = pi14 ? n60676 : n60677;
  assign n60679 = pi15 ? n14397 : n14613;
  assign n60680 = pi14 ? n60679 : n21035;
  assign n60681 = pi13 ? n60678 : n60680;
  assign n60682 = pi12 ? n60675 : n60681;
  assign n60683 = pi11 ? n60669 : n60682;
  assign n60684 = pi20 ? n2358 : ~n175;
  assign n60685 = pi19 ? n1165 : ~n60684;
  assign n60686 = pi18 ? n60685 : ~n31385;
  assign n60687 = pi17 ? n32 : n60686;
  assign n60688 = pi16 ? n32 : n60687;
  assign n60689 = pi15 ? n32717 : n60688;
  assign n60690 = pi14 ? n32 : n60689;
  assign n60691 = pi18 ? n16603 : n350;
  assign n60692 = pi17 ? n32 : n60691;
  assign n60693 = pi16 ? n1233 : ~n60692;
  assign n60694 = pi15 ? n46354 : n60693;
  assign n60695 = pi14 ? n60694 : n34044;
  assign n60696 = pi13 ? n60690 : n60695;
  assign n60697 = pi16 ? n129 : n21729;
  assign n60698 = pi15 ? n60033 : n60697;
  assign n60699 = pi14 ? n36601 : n60698;
  assign n60700 = pi13 ? n60699 : n21757;
  assign n60701 = pi12 ? n60696 : n60700;
  assign n60702 = pi15 ? n21762 : n32730;
  assign n60703 = pi15 ? n19805 : n13684;
  assign n60704 = pi14 ? n60702 : n60703;
  assign n60705 = pi18 ? n496 : ~n13681;
  assign n60706 = pi17 ? n32 : n60705;
  assign n60707 = pi16 ? n19652 : ~n60706;
  assign n60708 = pi15 ? n60707 : n58396;
  assign n60709 = pi14 ? n60708 : n60577;
  assign n60710 = pi13 ? n60704 : n60709;
  assign n60711 = pi17 ? n18487 : n59184;
  assign n60712 = pi16 ? n1471 : ~n60711;
  assign n60713 = pi15 ? n46188 : n60712;
  assign n60714 = pi14 ? n46183 : n60713;
  assign n60715 = pi19 ? n29705 : ~n39206;
  assign n60716 = pi18 ? n366 : ~n60715;
  assign n60717 = pi17 ? n32 : n60716;
  assign n60718 = pi19 ? n28686 : n34188;
  assign n60719 = pi19 ? n39206 : ~n4391;
  assign n60720 = pi18 ? n60718 : ~n60719;
  assign n60721 = pi17 ? n60720 : ~n2410;
  assign n60722 = pi16 ? n60717 : n60721;
  assign n60723 = pi19 ? n20555 : ~n31490;
  assign n60724 = pi18 ? n39110 : ~n60723;
  assign n60725 = pi17 ? n60724 : ~n1933;
  assign n60726 = pi16 ? n60432 : n60725;
  assign n60727 = pi15 ? n60722 : n60726;
  assign n60728 = pi19 ? n8631 : ~n32;
  assign n60729 = pi18 ? n32 : n60728;
  assign n60730 = pi17 ? n46210 : ~n60729;
  assign n60731 = pi16 ? n46205 : n60730;
  assign n60732 = pi15 ? n60731 : n91;
  assign n60733 = pi14 ? n60727 : n60732;
  assign n60734 = pi13 ? n60714 : n60733;
  assign n60735 = pi12 ? n60710 : n60734;
  assign n60736 = pi11 ? n60701 : n60735;
  assign n60737 = pi10 ? n60683 : n60736;
  assign n60738 = pi09 ? n60597 : n60737;
  assign n60739 = pi19 ? n43597 : n30040;
  assign n60740 = pi18 ? n32 : n60739;
  assign n60741 = pi17 ? n32 : n60740;
  assign n60742 = pi19 ? n30044 : ~n4279;
  assign n60743 = pi20 ? n5854 : n4279;
  assign n60744 = pi19 ? n60743 : n2180;
  assign n60745 = pi18 ? n60742 : ~n60744;
  assign n60746 = pi20 ? n5854 : ~n2358;
  assign n60747 = pi19 ? n60746 : ~n17669;
  assign n60748 = pi18 ? n60747 : ~n31972;
  assign n60749 = pi17 ? n60745 : ~n60748;
  assign n60750 = pi16 ? n60741 : ~n60749;
  assign n60751 = pi18 ? n1862 : n28164;
  assign n60752 = pi17 ? n32 : n60751;
  assign n60753 = pi16 ? n60752 : n60622;
  assign n60754 = pi15 ? n60750 : n60753;
  assign n60755 = pi20 ? n4279 : n1817;
  assign n60756 = pi19 ? n37233 : n60755;
  assign n60757 = pi18 ? n32 : n60756;
  assign n60758 = pi17 ? n32 : n60757;
  assign n60759 = pi19 ? n9197 : n9491;
  assign n60760 = pi19 ? n18410 : n7939;
  assign n60761 = pi18 ? n60759 : n60760;
  assign n60762 = pi20 ? n17669 : n29457;
  assign n60763 = pi19 ? n60762 : n287;
  assign n60764 = pi20 ? n5854 : ~n1377;
  assign n60765 = pi19 ? n60764 : n32;
  assign n60766 = pi18 ? n60763 : ~n60765;
  assign n60767 = pi17 ? n60761 : n60766;
  assign n60768 = pi16 ? n60758 : ~n60767;
  assign n60769 = pi15 ? n60768 : n21319;
  assign n60770 = pi14 ? n60754 : n60769;
  assign n60771 = pi16 ? n2137 : ~n2756;
  assign n60772 = pi16 ? n1808 : ~n2749;
  assign n60773 = pi15 ? n60771 : n60772;
  assign n60774 = pi17 ? n60654 : n22467;
  assign n60775 = pi16 ? n60651 : n60774;
  assign n60776 = pi17 ? n60661 : ~n14150;
  assign n60777 = pi16 ? n60659 : ~n60776;
  assign n60778 = pi15 ? n60775 : n60777;
  assign n60779 = pi14 ? n60773 : n60778;
  assign n60780 = pi13 ? n60770 : n60779;
  assign n60781 = pi14 ? n21787 : n21790;
  assign n60782 = pi15 ? n21543 : n21786;
  assign n60783 = pi14 ? n60782 : n21790;
  assign n60784 = pi13 ? n60781 : n60783;
  assign n60785 = pi12 ? n60780 : n60784;
  assign n60786 = pi19 ? n58685 : ~n32;
  assign n60787 = pi18 ? n341 : ~n60786;
  assign n60788 = pi17 ? n32 : n60787;
  assign n60789 = pi16 ? n32 : n60788;
  assign n60790 = pi15 ? n32 : n60789;
  assign n60791 = pi15 ? n12079 : n32468;
  assign n60792 = pi14 ? n60790 : n60791;
  assign n60793 = pi15 ? n32828 : n46138;
  assign n60794 = pi14 ? n60793 : n46255;
  assign n60795 = pi13 ? n60792 : n60794;
  assign n60796 = pi18 ? n32 : n22779;
  assign n60797 = pi17 ? n32 : n60796;
  assign n60798 = pi16 ? n32 : n60797;
  assign n60799 = pi15 ? n21346 : n60798;
  assign n60800 = pi14 ? n46263 : n60799;
  assign n60801 = pi15 ? n21695 : n32;
  assign n60802 = pi14 ? n60801 : n20836;
  assign n60803 = pi13 ? n60800 : n60802;
  assign n60804 = pi12 ? n60795 : n60803;
  assign n60805 = pi11 ? n60785 : n60804;
  assign n60806 = pi19 ? n32847 : ~n28965;
  assign n60807 = pi18 ? n60806 : ~n3508;
  assign n60808 = pi17 ? n32 : n60807;
  assign n60809 = pi16 ? n32 : n60808;
  assign n60810 = pi15 ? n32846 : n60809;
  assign n60811 = pi14 ? n32 : n60810;
  assign n60812 = pi16 ? n1135 : ~n60692;
  assign n60813 = pi15 ? n31828 : n60812;
  assign n60814 = pi16 ? n1135 : ~n2293;
  assign n60815 = pi14 ? n60813 : n60814;
  assign n60816 = pi13 ? n60811 : n60815;
  assign n60817 = pi15 ? n47256 : n21830;
  assign n60818 = pi14 ? n60402 : n60817;
  assign n60819 = pi13 ? n60818 : n21757;
  assign n60820 = pi12 ? n60816 : n60819;
  assign n60821 = pi18 ? n32 : n31396;
  assign n60822 = pi17 ? n32 : n60821;
  assign n60823 = pi16 ? n32 : n60822;
  assign n60824 = pi15 ? n21762 : n60823;
  assign n60825 = pi15 ? n32730 : n20301;
  assign n60826 = pi14 ? n60824 : n60825;
  assign n60827 = pi16 ? n1214 : ~n60706;
  assign n60828 = pi15 ? n60827 : n47261;
  assign n60829 = pi14 ? n60828 : n60577;
  assign n60830 = pi13 ? n60826 : n60829;
  assign n60831 = pi17 ? n60724 : ~n2305;
  assign n60832 = pi16 ? n60432 : n60831;
  assign n60833 = pi15 ? n60722 : n60832;
  assign n60834 = pi18 ? n32 : n19606;
  assign n60835 = pi17 ? n46210 : ~n60834;
  assign n60836 = pi16 ? n46205 : n60835;
  assign n60837 = pi15 ? n60836 : n19503;
  assign n60838 = pi14 ? n60833 : n60837;
  assign n60839 = pi13 ? n60714 : n60838;
  assign n60840 = pi12 ? n60830 : n60839;
  assign n60841 = pi11 ? n60820 : n60840;
  assign n60842 = pi10 ? n60805 : n60841;
  assign n60843 = pi09 ? n60597 : n60842;
  assign n60844 = pi08 ? n60738 : n60843;
  assign n60845 = pi07 ? n60591 : n60844;
  assign n60846 = pi20 ? n175 : ~n1611;
  assign n60847 = pi19 ? n60846 : n32;
  assign n60848 = pi18 ? n32 : n60847;
  assign n60849 = pi17 ? n32 : n60848;
  assign n60850 = pi16 ? n32 : n60849;
  assign n60851 = pi15 ? n21853 : n60850;
  assign n60852 = pi14 ? n32 : n60851;
  assign n60853 = pi13 ? n32 : n60852;
  assign n60854 = pi12 ? n32 : n60853;
  assign n60855 = pi11 ? n32 : n60854;
  assign n60856 = pi10 ? n32 : n60855;
  assign n60857 = pi15 ? n34852 : n14389;
  assign n60858 = pi14 ? n60857 : n23609;
  assign n60859 = pi16 ? n1683 : ~n2518;
  assign n60860 = pi16 ? n31442 : ~n2749;
  assign n60861 = pi15 ? n60859 : n60860;
  assign n60862 = pi19 ? n28786 : n5371;
  assign n60863 = pi18 ? n32 : ~n60862;
  assign n60864 = pi17 ? n32 : n60863;
  assign n60865 = pi17 ? n19907 : n21684;
  assign n60866 = pi16 ? n60864 : n60865;
  assign n60867 = pi15 ? n60866 : n32;
  assign n60868 = pi14 ? n60861 : n60867;
  assign n60869 = pi13 ? n60858 : n60868;
  assign n60870 = pi13 ? n60781 : n21855;
  assign n60871 = pi12 ? n60869 : n60870;
  assign n60872 = pi18 ? n209 : ~n323;
  assign n60873 = pi17 ? n32 : n60872;
  assign n60874 = pi16 ? n32 : n60873;
  assign n60875 = pi15 ? n60874 : n12289;
  assign n60876 = pi14 ? n60875 : n46327;
  assign n60877 = pi13 ? n60876 : n46333;
  assign n60878 = pi15 ? n54379 : n21543;
  assign n60879 = pi14 ? n32899 : n60878;
  assign n60880 = pi14 ? n21697 : n40399;
  assign n60881 = pi13 ? n60879 : n60880;
  assign n60882 = pi12 ? n60877 : n60881;
  assign n60883 = pi11 ? n60871 : n60882;
  assign n60884 = pi14 ? n31978 : n32923;
  assign n60885 = pi18 ? n15844 : n532;
  assign n60886 = pi17 ? n32 : n60885;
  assign n60887 = pi16 ? n1233 : ~n60886;
  assign n60888 = pi18 ? n16316 : n418;
  assign n60889 = pi17 ? n32 : n60888;
  assign n60890 = pi16 ? n1233 : ~n60889;
  assign n60891 = pi15 ? n60887 : n60890;
  assign n60892 = pi14 ? n60891 : n59901;
  assign n60893 = pi13 ? n60884 : n60892;
  assign n60894 = pi18 ? n29802 : ~n605;
  assign n60895 = pi17 ? n32 : n60894;
  assign n60896 = pi16 ? n568 : n60895;
  assign n60897 = pi15 ? n60896 : n21891;
  assign n60898 = pi14 ? n59560 : n60897;
  assign n60899 = pi13 ? n60898 : n21905;
  assign n60900 = pi12 ? n60893 : n60899;
  assign n60901 = pi15 ? n20048 : n23708;
  assign n60902 = pi19 ? n5855 : n1076;
  assign n60903 = pi18 ? n41883 : n60902;
  assign n60904 = pi17 ? n32 : n60903;
  assign n60905 = pi19 ? n22698 : ~n22701;
  assign n60906 = pi18 ? n43622 : n60905;
  assign n60907 = pi18 ? n32372 : ~n13949;
  assign n60908 = pi17 ? n60906 : ~n60907;
  assign n60909 = pi16 ? n60904 : n60908;
  assign n60910 = pi15 ? n13952 : n60909;
  assign n60911 = pi14 ? n60901 : n60910;
  assign n60912 = pi18 ? n6071 : n3786;
  assign n60913 = pi17 ? n32 : n60912;
  assign n60914 = pi16 ? n46369 : ~n60913;
  assign n60915 = pi16 ? n46373 : ~n3625;
  assign n60916 = pi15 ? n60914 : n60915;
  assign n60917 = pi14 ? n60916 : n46380;
  assign n60918 = pi13 ? n60911 : n60917;
  assign n60919 = pi17 ? n46393 : n58467;
  assign n60920 = pi16 ? n46390 : ~n60919;
  assign n60921 = pi15 ? n32980 : n60920;
  assign n60922 = pi14 ? n46387 : n60921;
  assign n60923 = pi18 ? n366 : ~n6581;
  assign n60924 = pi17 ? n32 : n60923;
  assign n60925 = pi20 ? n12062 : ~n32;
  assign n60926 = pi19 ? n60925 : ~n32;
  assign n60927 = pi18 ? n32 : n60926;
  assign n60928 = pi17 ? n46401 : n60927;
  assign n60929 = pi16 ? n60924 : ~n60928;
  assign n60930 = pi18 ? n566 : n4965;
  assign n60931 = pi17 ? n32 : n60930;
  assign n60932 = pi21 ? n206 : n10445;
  assign n60933 = pi20 ? n60932 : ~n32;
  assign n60934 = pi19 ? n60933 : ~n32;
  assign n60935 = pi18 ? n940 : n60934;
  assign n60936 = pi17 ? n46405 : ~n60935;
  assign n60937 = pi16 ? n60931 : n60936;
  assign n60938 = pi15 ? n60929 : n60937;
  assign n60939 = pi15 ? n20538 : n19503;
  assign n60940 = pi14 ? n60938 : n60939;
  assign n60941 = pi13 ? n60922 : n60940;
  assign n60942 = pi12 ? n60918 : n60941;
  assign n60943 = pi11 ? n60900 : n60942;
  assign n60944 = pi10 ? n60883 : n60943;
  assign n60945 = pi09 ? n60856 : n60944;
  assign n60946 = pi20 ? n175 : ~n342;
  assign n60947 = pi19 ? n60946 : n32;
  assign n60948 = pi18 ? n32 : n60947;
  assign n60949 = pi17 ? n32 : n60948;
  assign n60950 = pi16 ? n32 : n60949;
  assign n60951 = pi15 ? n21853 : n60950;
  assign n60952 = pi14 ? n32 : n60951;
  assign n60953 = pi13 ? n32 : n60952;
  assign n60954 = pi12 ? n32 : n60953;
  assign n60955 = pi11 ? n32 : n60954;
  assign n60956 = pi10 ? n32 : n60955;
  assign n60957 = pi16 ? n1683 : ~n2749;
  assign n60958 = pi16 ? n31442 : ~n2513;
  assign n60959 = pi15 ? n60957 : n60958;
  assign n60960 = pi17 ? n19907 : n20021;
  assign n60961 = pi16 ? n60864 : n60960;
  assign n60962 = pi15 ? n60961 : n32;
  assign n60963 = pi14 ? n60959 : n60962;
  assign n60964 = pi13 ? n60858 : n60963;
  assign n60965 = pi14 ? n21929 : n22133;
  assign n60966 = pi13 ? n60965 : n21932;
  assign n60967 = pi12 ? n60964 : n60966;
  assign n60968 = pi15 ? n60874 : n32885;
  assign n60969 = pi14 ? n60968 : n46327;
  assign n60970 = pi13 ? n60969 : n46333;
  assign n60971 = pi19 ? n17194 : n32;
  assign n60972 = pi18 ? n32 : n60971;
  assign n60973 = pi17 ? n32 : n60972;
  assign n60974 = pi16 ? n32 : n60973;
  assign n60975 = pi15 ? n60974 : n32;
  assign n60976 = pi14 ? n33021 : n60975;
  assign n60977 = pi14 ? n21697 : n32;
  assign n60978 = pi13 ? n60976 : n60977;
  assign n60979 = pi12 ? n60970 : n60978;
  assign n60980 = pi11 ? n60967 : n60979;
  assign n60981 = pi14 ? n31978 : n33033;
  assign n60982 = pi16 ? n1135 : ~n60886;
  assign n60983 = pi19 ? n42337 : ~n32;
  assign n60984 = pi18 ? n16316 : n60983;
  assign n60985 = pi17 ? n32 : n60984;
  assign n60986 = pi16 ? n1135 : ~n60985;
  assign n60987 = pi15 ? n60982 : n60986;
  assign n60988 = pi15 ? n47710 : n60814;
  assign n60989 = pi14 ? n60987 : n60988;
  assign n60990 = pi13 ? n60981 : n60989;
  assign n60991 = pi15 ? n34146 : n60402;
  assign n60992 = pi16 ? n919 : n60895;
  assign n60993 = pi15 ? n60992 : n21891;
  assign n60994 = pi14 ? n60991 : n60993;
  assign n60995 = pi13 ? n60994 : n21905;
  assign n60996 = pi12 ? n60990 : n60995;
  assign n60997 = pi15 ? n20301 : n23780;
  assign n60998 = pi18 ? n32372 : ~n20474;
  assign n60999 = pi17 ? n60906 : ~n60998;
  assign n61000 = pi16 ? n60904 : n60999;
  assign n61001 = pi15 ? n486 : n61000;
  assign n61002 = pi14 ? n60997 : n61001;
  assign n61003 = pi18 ? n6071 : n39007;
  assign n61004 = pi17 ? n32 : n61003;
  assign n61005 = pi16 ? n46460 : ~n61004;
  assign n61006 = pi16 ? n46463 : ~n3788;
  assign n61007 = pi15 ? n61005 : n61006;
  assign n61008 = pi15 ? n46559 : n44087;
  assign n61009 = pi14 ? n61007 : n61008;
  assign n61010 = pi13 ? n61002 : n61009;
  assign n61011 = pi17 ? n46401 : n2299;
  assign n61012 = pi16 ? n60924 : ~n61011;
  assign n61013 = pi21 ? n206 : n7659;
  assign n61014 = pi20 ? n61013 : ~n32;
  assign n61015 = pi19 ? n61014 : ~n32;
  assign n61016 = pi18 ? n940 : n61015;
  assign n61017 = pi17 ? n46405 : ~n61016;
  assign n61018 = pi16 ? n60931 : n61017;
  assign n61019 = pi15 ? n61012 : n61018;
  assign n61020 = pi15 ? n180 : n19874;
  assign n61021 = pi14 ? n61019 : n61020;
  assign n61022 = pi13 ? n46474 : n61021;
  assign n61023 = pi12 ? n61010 : n61022;
  assign n61024 = pi11 ? n60996 : n61023;
  assign n61025 = pi10 ? n60980 : n61024;
  assign n61026 = pi09 ? n60956 : n61025;
  assign n61027 = pi08 ? n60945 : n61026;
  assign n61028 = pi19 ? n30349 : n507;
  assign n61029 = pi20 ? n339 : ~n2140;
  assign n61030 = pi19 ? n61029 : n32;
  assign n61031 = pi18 ? n61028 : n61030;
  assign n61032 = pi17 ? n32 : n61031;
  assign n61033 = pi16 ? n32 : n61032;
  assign n61034 = pi15 ? n14790 : n61033;
  assign n61035 = pi14 ? n32 : n61034;
  assign n61036 = pi13 ? n32 : n61035;
  assign n61037 = pi12 ? n32 : n61036;
  assign n61038 = pi11 ? n32 : n61037;
  assign n61039 = pi10 ? n32 : n61038;
  assign n61040 = pi20 ? n4279 : n266;
  assign n61041 = pi19 ? n61040 : n32;
  assign n61042 = pi18 ? n32 : n61041;
  assign n61043 = pi17 ? n32 : n61042;
  assign n61044 = pi16 ? n32 : n61043;
  assign n61045 = pi15 ? n61044 : n22958;
  assign n61046 = pi14 ? n61045 : n22133;
  assign n61047 = pi16 ? n59546 : ~n2513;
  assign n61048 = pi15 ? n60957 : n61047;
  assign n61049 = pi18 ? n4380 : ~n17118;
  assign n61050 = pi17 ? n32 : n61049;
  assign n61051 = pi17 ? n36647 : ~n20021;
  assign n61052 = pi16 ? n61050 : ~n61051;
  assign n61053 = pi15 ? n61052 : n32;
  assign n61054 = pi14 ? n61048 : n61053;
  assign n61055 = pi13 ? n61046 : n61054;
  assign n61056 = pi14 ? n32 : n476;
  assign n61057 = pi14 ? n21790 : n48800;
  assign n61058 = pi13 ? n61056 : n61057;
  assign n61059 = pi12 ? n61055 : n61058;
  assign n61060 = pi14 ? n33088 : n21790;
  assign n61061 = pi14 ? n22009 : n21322;
  assign n61062 = pi13 ? n61060 : n61061;
  assign n61063 = pi12 ? n46522 : n61062;
  assign n61064 = pi11 ? n61059 : n61063;
  assign n61065 = pi14 ? n32 : n33102;
  assign n61066 = pi18 ? n32 : n2360;
  assign n61067 = pi17 ? n32 : n61066;
  assign n61068 = pi16 ? n1233 : ~n61067;
  assign n61069 = pi15 ? n60887 : n61068;
  assign n61070 = pi15 ? n60190 : n59901;
  assign n61071 = pi14 ? n61069 : n61070;
  assign n61072 = pi13 ? n61065 : n61071;
  assign n61073 = pi15 ? n34044 : n59560;
  assign n61074 = pi18 ? n29802 : ~n32381;
  assign n61075 = pi17 ? n32 : n61074;
  assign n61076 = pi16 ? n568 : n61075;
  assign n61077 = pi15 ? n61076 : n22028;
  assign n61078 = pi14 ? n61073 : n61077;
  assign n61079 = pi18 ? n22039 : n21229;
  assign n61080 = pi17 ? n32 : n61079;
  assign n61081 = pi16 ? n32 : n61080;
  assign n61082 = pi15 ? n22036 : n61081;
  assign n61083 = pi14 ? n22037 : n61082;
  assign n61084 = pi13 ? n61078 : n61083;
  assign n61085 = pi12 ? n61072 : n61084;
  assign n61086 = pi17 ? n46549 : n32743;
  assign n61087 = pi16 ? n46546 : ~n61086;
  assign n61088 = pi15 ? n486 : n61087;
  assign n61089 = pi14 ? n55021 : n61088;
  assign n61090 = pi15 ? n46774 : n46556;
  assign n61091 = pi14 ? n61090 : n46563;
  assign n61092 = pi13 ? n61089 : n61091;
  assign n61093 = pi17 ? n19170 : n46560;
  assign n61094 = pi16 ? n32 : n61093;
  assign n61095 = pi15 ? n61094 : n46584;
  assign n61096 = pi14 ? n46573 : n61095;
  assign n61097 = pi17 ? n46401 : n58467;
  assign n61098 = pi16 ? n60924 : ~n61097;
  assign n61099 = pi18 ? n30458 : n4965;
  assign n61100 = pi17 ? n32 : n61099;
  assign n61101 = pi20 ? n1368 : n32;
  assign n61102 = pi19 ? n61101 : n32;
  assign n61103 = pi18 ? n1592 : ~n61102;
  assign n61104 = pi17 ? n46591 : n61103;
  assign n61105 = pi16 ? n61100 : ~n61104;
  assign n61106 = pi15 ? n61098 : n61105;
  assign n61107 = pi16 ? n129 : n18561;
  assign n61108 = pi15 ? n116 : n61107;
  assign n61109 = pi14 ? n61106 : n61108;
  assign n61110 = pi13 ? n61096 : n61109;
  assign n61111 = pi12 ? n61092 : n61110;
  assign n61112 = pi11 ? n61085 : n61111;
  assign n61113 = pi10 ? n61064 : n61112;
  assign n61114 = pi09 ? n61039 : n61113;
  assign n61115 = pi15 ? n21853 : n61033;
  assign n61116 = pi14 ? n32 : n61115;
  assign n61117 = pi13 ? n32 : n61116;
  assign n61118 = pi12 ? n32 : n61117;
  assign n61119 = pi11 ? n32 : n61118;
  assign n61120 = pi10 ? n32 : n61119;
  assign n61121 = pi14 ? n61045 : n476;
  assign n61122 = pi16 ? n1683 : ~n2629;
  assign n61123 = pi16 ? n59546 : ~n2629;
  assign n61124 = pi15 ? n61122 : n61123;
  assign n61125 = pi14 ? n61124 : n61053;
  assign n61126 = pi13 ? n61121 : n61125;
  assign n61127 = pi15 ? n21928 : n648;
  assign n61128 = pi15 ? n648 : n21853;
  assign n61129 = pi14 ? n61127 : n61128;
  assign n61130 = pi13 ? n47691 : n61129;
  assign n61131 = pi12 ? n61126 : n61130;
  assign n61132 = pi15 ? n12518 : n12515;
  assign n61133 = pi14 ? n61132 : n46514;
  assign n61134 = pi15 ? n46331 : n13920;
  assign n61135 = pi14 ? n61134 : n46520;
  assign n61136 = pi13 ? n61133 : n61135;
  assign n61137 = pi15 ? n13920 : n22006;
  assign n61138 = pi14 ? n61137 : n21790;
  assign n61139 = pi14 ? n23466 : n21322;
  assign n61140 = pi13 ? n61138 : n61139;
  assign n61141 = pi12 ? n61136 : n61140;
  assign n61142 = pi11 ? n61131 : n61141;
  assign n61143 = pi20 ? n32 : n6886;
  assign n61144 = pi19 ? n61143 : ~n32;
  assign n61145 = pi18 ? n32 : n61144;
  assign n61146 = pi17 ? n32 : n61145;
  assign n61147 = pi16 ? n1135 : ~n61146;
  assign n61148 = pi15 ? n60982 : n61147;
  assign n61149 = pi15 ? n60189 : n47710;
  assign n61150 = pi14 ? n61148 : n61149;
  assign n61151 = pi13 ? n61065 : n61150;
  assign n61152 = pi15 ? n60814 : n34146;
  assign n61153 = pi18 ? n29802 : ~n532;
  assign n61154 = pi17 ? n32 : n61153;
  assign n61155 = pi16 ? n919 : n61154;
  assign n61156 = pi15 ? n61155 : n22100;
  assign n61157 = pi14 ? n61152 : n61156;
  assign n61158 = pi18 ? n22107 : n20753;
  assign n61159 = pi17 ? n32 : n61158;
  assign n61160 = pi16 ? n32 : n61159;
  assign n61161 = pi15 ? n22036 : n61160;
  assign n61162 = pi14 ? n22105 : n61161;
  assign n61163 = pi13 ? n61157 : n61162;
  assign n61164 = pi12 ? n61151 : n61163;
  assign n61165 = pi15 ? n13952 : n21232;
  assign n61166 = pi18 ? n323 : ~n483;
  assign n61167 = pi17 ? n46549 : n61166;
  assign n61168 = pi16 ? n46546 : ~n61167;
  assign n61169 = pi15 ? n20660 : n61168;
  assign n61170 = pi14 ? n61165 : n61169;
  assign n61171 = pi16 ? n46555 : ~n3788;
  assign n61172 = pi15 ? n46441 : n61171;
  assign n61173 = pi14 ? n61172 : n46563;
  assign n61174 = pi13 ? n61170 : n61173;
  assign n61175 = pi15 ? n61094 : n46662;
  assign n61176 = pi14 ? n46573 : n61175;
  assign n61177 = pi17 ? n46401 : n3333;
  assign n61178 = pi16 ? n60924 : ~n61177;
  assign n61179 = pi15 ? n61178 : n61105;
  assign n61180 = pi15 ? n72 : n20538;
  assign n61181 = pi14 ? n61179 : n61180;
  assign n61182 = pi13 ? n61176 : n61181;
  assign n61183 = pi12 ? n61174 : n61182;
  assign n61184 = pi11 ? n61164 : n61183;
  assign n61185 = pi10 ? n61142 : n61184;
  assign n61186 = pi09 ? n61120 : n61185;
  assign n61187 = pi08 ? n61114 : n61186;
  assign n61188 = pi07 ? n61027 : n61187;
  assign n61189 = pi06 ? n60845 : n61188;
  assign n61190 = pi18 ? n880 : ~n6405;
  assign n61191 = pi17 ? n61190 : ~n2618;
  assign n61192 = pi16 ? n32 : n61191;
  assign n61193 = pi15 ? n24543 : n61192;
  assign n61194 = pi14 ? n32 : n61193;
  assign n61195 = pi13 ? n32 : n61194;
  assign n61196 = pi12 ? n32 : n61195;
  assign n61197 = pi11 ? n32 : n61196;
  assign n61198 = pi10 ? n32 : n61197;
  assign n61199 = pi18 ? n32 : n41276;
  assign n61200 = pi19 ? n19151 : ~n247;
  assign n61201 = pi19 ? n11899 : n32;
  assign n61202 = pi18 ? n61200 : ~n61201;
  assign n61203 = pi17 ? n61199 : ~n61202;
  assign n61204 = pi16 ? n32 : n61203;
  assign n61205 = pi18 ? n32584 : ~n595;
  assign n61206 = pi17 ? n32 : n61205;
  assign n61207 = pi16 ? n32 : n61206;
  assign n61208 = pi15 ? n61204 : n61207;
  assign n61209 = pi14 ? n61208 : n33236;
  assign n61210 = pi16 ? n28030 : ~n2629;
  assign n61211 = pi15 ? n61210 : n61123;
  assign n61212 = pi19 ? n18408 : ~n8064;
  assign n61213 = pi18 ? n18831 : ~n61212;
  assign n61214 = pi17 ? n32 : n61213;
  assign n61215 = pi16 ? n61214 : n32;
  assign n61216 = pi15 ? n61215 : n32;
  assign n61217 = pi14 ? n61211 : n61216;
  assign n61218 = pi13 ? n61209 : n61217;
  assign n61219 = pi15 ? n21853 : n648;
  assign n61220 = pi15 ? n648 : n33493;
  assign n61221 = pi14 ? n61219 : n61220;
  assign n61222 = pi13 ? n47691 : n61221;
  assign n61223 = pi12 ? n61218 : n61222;
  assign n61224 = pi15 ? n14394 : n21853;
  assign n61225 = pi14 ? n61224 : n22133;
  assign n61226 = pi14 ? n21687 : n21464;
  assign n61227 = pi13 ? n61225 : n61226;
  assign n61228 = pi12 ? n46731 : n61227;
  assign n61229 = pi11 ? n61223 : n61228;
  assign n61230 = pi18 ? n33278 : ~n532;
  assign n61231 = pi17 ? n32 : n61230;
  assign n61232 = pi16 ? n32 : n61231;
  assign n61233 = pi18 ? n33282 : ~n605;
  assign n61234 = pi17 ? n32 : n61233;
  assign n61235 = pi16 ? n32 : n61234;
  assign n61236 = pi15 ? n61232 : n61235;
  assign n61237 = pi14 ? n21217 : n61236;
  assign n61238 = pi16 ? n1233 : ~n2756;
  assign n61239 = pi15 ? n61238 : n60190;
  assign n61240 = pi14 ? n61238 : n61239;
  assign n61241 = pi13 ? n61237 : n61240;
  assign n61242 = pi17 ? n46740 : n45638;
  assign n61243 = pi16 ? n568 : n61242;
  assign n61244 = pi17 ? n46740 : n22165;
  assign n61245 = pi16 ? n568 : n61244;
  assign n61246 = pi15 ? n61243 : n61245;
  assign n61247 = pi14 ? n61246 : n22163;
  assign n61248 = pi15 ? n22174 : n21232;
  assign n61249 = pi14 ? n22171 : n61248;
  assign n61250 = pi13 ? n61247 : n61249;
  assign n61251 = pi12 ? n61241 : n61250;
  assign n61252 = pi19 ? n2358 : ~n6139;
  assign n61253 = pi18 ? n268 : ~n61252;
  assign n61254 = pi17 ? n32 : n61253;
  assign n61255 = pi19 ? n57838 : n246;
  assign n61256 = pi20 ? n266 : ~n287;
  assign n61257 = pi19 ? n61256 : n39181;
  assign n61258 = pi18 ? n61255 : n61257;
  assign n61259 = pi19 ? n43354 : ~n236;
  assign n61260 = pi18 ? n61259 : n13945;
  assign n61261 = pi17 ? n61258 : n61260;
  assign n61262 = pi16 ? n61254 : n61261;
  assign n61263 = pi20 ? n357 : n243;
  assign n61264 = pi19 ? n61263 : ~n32;
  assign n61265 = pi18 ? n32 : n61264;
  assign n61266 = pi17 ? n32 : n61265;
  assign n61267 = pi16 ? n46770 : ~n61266;
  assign n61268 = pi15 ? n61262 : n61267;
  assign n61269 = pi14 ? n31717 : n61268;
  assign n61270 = pi15 ? n46441 : n46774;
  assign n61271 = pi14 ? n61270 : n46782;
  assign n61272 = pi13 ? n61269 : n61271;
  assign n61273 = pi16 ? n33623 : ~n3788;
  assign n61274 = pi15 ? n61273 : n33459;
  assign n61275 = pi18 ? n209 : ~n28433;
  assign n61276 = pi17 ? n32 : n61275;
  assign n61277 = pi16 ? n61276 : ~n3625;
  assign n61278 = pi15 ? n33361 : n61277;
  assign n61279 = pi14 ? n61274 : n61278;
  assign n61280 = pi18 ? n366 : ~n32570;
  assign n61281 = pi17 ? n32 : n61280;
  assign n61282 = pi16 ? n61281 : ~n3625;
  assign n61283 = pi18 ? n6071 : n177;
  assign n61284 = pi17 ? n32 : n61283;
  assign n61285 = pi16 ? n32 : n61284;
  assign n61286 = pi15 ? n61282 : n61285;
  assign n61287 = pi16 ? n129 : n19867;
  assign n61288 = pi15 ? n180 : n61287;
  assign n61289 = pi14 ? n61286 : n61288;
  assign n61290 = pi13 ? n61279 : n61289;
  assign n61291 = pi12 ? n61272 : n61290;
  assign n61292 = pi11 ? n61251 : n61291;
  assign n61293 = pi10 ? n61229 : n61292;
  assign n61294 = pi09 ? n61198 : n61293;
  assign n61295 = pi15 ? n19172 : n33236;
  assign n61296 = pi14 ? n61208 : n61295;
  assign n61297 = pi16 ? n28030 : ~n3946;
  assign n61298 = pi16 ? n59546 : ~n3946;
  assign n61299 = pi15 ? n61297 : n61298;
  assign n61300 = pi19 ? n18173 : ~n5614;
  assign n61301 = pi18 ? n19082 : ~n61300;
  assign n61302 = pi17 ? n32 : n61301;
  assign n61303 = pi16 ? n61302 : n32;
  assign n61304 = pi15 ? n61303 : n32;
  assign n61305 = pi14 ? n61299 : n61304;
  assign n61306 = pi13 ? n61296 : n61305;
  assign n61307 = pi14 ? n32 : n15267;
  assign n61308 = pi15 ? n14790 : n15263;
  assign n61309 = pi20 ? n206 : n7880;
  assign n61310 = pi19 ? n61309 : n32;
  assign n61311 = pi18 ? n32 : n61310;
  assign n61312 = pi17 ? n32 : n61311;
  assign n61313 = pi16 ? n32 : n61312;
  assign n61314 = pi15 ? n15263 : n61313;
  assign n61315 = pi14 ? n61308 : n61314;
  assign n61316 = pi13 ? n61307 : n61315;
  assign n61317 = pi12 ? n61306 : n61316;
  assign n61318 = pi19 ? n40989 : ~n32;
  assign n61319 = pi18 ? n940 : ~n61318;
  assign n61320 = pi17 ? n32 : n61319;
  assign n61321 = pi16 ? n32 : n61320;
  assign n61322 = pi15 ? n33246 : n61321;
  assign n61323 = pi14 ? n61322 : n46716;
  assign n61324 = pi13 ? n61323 : n46837;
  assign n61325 = pi14 ? n21790 : n32;
  assign n61326 = pi13 ? n61225 : n61325;
  assign n61327 = pi12 ? n61324 : n61326;
  assign n61328 = pi11 ? n61317 : n61327;
  assign n61329 = pi16 ? n1135 : ~n2518;
  assign n61330 = pi15 ? n61329 : n60189;
  assign n61331 = pi14 ? n61329 : n61330;
  assign n61332 = pi13 ? n61237 : n61331;
  assign n61333 = pi17 ? n46740 : n11421;
  assign n61334 = pi16 ? n919 : n61333;
  assign n61335 = pi16 ? n919 : n61242;
  assign n61336 = pi15 ? n61334 : n61335;
  assign n61337 = pi14 ? n61336 : n22163;
  assign n61338 = pi15 ? n22174 : n13943;
  assign n61339 = pi14 ? n22171 : n61338;
  assign n61340 = pi13 ? n61337 : n61339;
  assign n61341 = pi12 ? n61332 : n61340;
  assign n61342 = pi20 ? n357 : n207;
  assign n61343 = pi19 ? n61342 : ~n32;
  assign n61344 = pi18 ? n32 : n61343;
  assign n61345 = pi17 ? n32 : n61344;
  assign n61346 = pi16 ? n46770 : ~n61345;
  assign n61347 = pi15 ? n61262 : n61346;
  assign n61348 = pi14 ? n45139 : n61347;
  assign n61349 = pi14 ? n46992 : n46879;
  assign n61350 = pi13 ? n61348 : n61349;
  assign n61351 = pi16 ? n61276 : ~n3788;
  assign n61352 = pi15 ? n33361 : n61351;
  assign n61353 = pi14 ? n46883 : n61352;
  assign n61354 = pi16 ? n61281 : ~n3788;
  assign n61355 = pi15 ? n61354 : n13392;
  assign n61356 = pi14 ? n61355 : n19982;
  assign n61357 = pi13 ? n61353 : n61356;
  assign n61358 = pi12 ? n61350 : n61357;
  assign n61359 = pi11 ? n61341 : n61358;
  assign n61360 = pi10 ? n61328 : n61359;
  assign n61361 = pi09 ? n61198 : n61360;
  assign n61362 = pi08 ? n61294 : n61361;
  assign n61363 = pi19 ? n7642 : n246;
  assign n61364 = pi18 ? n268 : n61363;
  assign n61365 = pi18 ? n31385 : ~n4098;
  assign n61366 = pi17 ? n61364 : n61365;
  assign n61367 = pi16 ? n32 : n61366;
  assign n61368 = pi17 ? n61190 : ~n4099;
  assign n61369 = pi16 ? n32 : n61368;
  assign n61370 = pi15 ? n61367 : n61369;
  assign n61371 = pi14 ? n32 : n61370;
  assign n61372 = pi13 ? n32 : n61371;
  assign n61373 = pi12 ? n32 : n61372;
  assign n61374 = pi11 ? n32 : n61373;
  assign n61375 = pi10 ? n32 : n61374;
  assign n61376 = pi19 ? n4342 : n342;
  assign n61377 = pi18 ? n4380 : n61376;
  assign n61378 = pi18 ? n61200 : n508;
  assign n61379 = pi17 ? n61377 : ~n61378;
  assign n61380 = pi16 ? n32 : n61379;
  assign n61381 = pi19 ? n20555 : ~n176;
  assign n61382 = pi18 ? n61381 : n47144;
  assign n61383 = pi17 ? n32 : ~n61382;
  assign n61384 = pi16 ? n32 : n61383;
  assign n61385 = pi15 ? n61380 : n61384;
  assign n61386 = pi20 ? n207 : ~n175;
  assign n61387 = pi19 ? n61386 : ~n32;
  assign n61388 = pi18 ? n32 : ~n61387;
  assign n61389 = pi17 ? n32 : n61388;
  assign n61390 = pi16 ? n32 : n61389;
  assign n61391 = pi14 ? n61385 : n61390;
  assign n61392 = pi16 ? n1471 : ~n3946;
  assign n61393 = pi18 ? n2197 : n237;
  assign n61394 = pi17 ? n32 : n61393;
  assign n61395 = pi16 ? n61394 : ~n3946;
  assign n61396 = pi15 ? n61392 : n61395;
  assign n61397 = pi14 ? n61396 : n32;
  assign n61398 = pi13 ? n61391 : n61397;
  assign n61399 = pi15 ? n15123 : n46926;
  assign n61400 = pi14 ? n22252 : n61399;
  assign n61401 = pi13 ? n33386 : n61400;
  assign n61402 = pi12 ? n61398 : n61401;
  assign n61403 = pi20 ? n321 : ~n14968;
  assign n61404 = pi19 ? n61403 : ~n32;
  assign n61405 = pi18 ? n32 : ~n61404;
  assign n61406 = pi17 ? n32 : n61405;
  assign n61407 = pi16 ? n32 : n61406;
  assign n61408 = pi18 ? n863 : n13623;
  assign n61409 = pi17 ? n32 : n61408;
  assign n61410 = pi16 ? n32 : n61409;
  assign n61411 = pi15 ? n61407 : n61410;
  assign n61412 = pi14 ? n46938 : n61411;
  assign n61413 = pi13 ? n61412 : n46967;
  assign n61414 = pi15 ? n14147 : n648;
  assign n61415 = pi14 ? n61414 : n649;
  assign n61416 = pi14 ? n21854 : n21543;
  assign n61417 = pi13 ? n61415 : n61416;
  assign n61418 = pi12 ? n61413 : n61417;
  assign n61419 = pi11 ? n61402 : n61418;
  assign n61420 = pi20 ? n9641 : n749;
  assign n61421 = pi19 ? n61420 : ~n32;
  assign n61422 = pi18 ? n697 : ~n61421;
  assign n61423 = pi17 ? n32 : n61422;
  assign n61424 = pi16 ? n32 : n61423;
  assign n61425 = pi15 ? n33557 : n61424;
  assign n61426 = pi14 ? n21217 : n61425;
  assign n61427 = pi13 ? n61426 : n61331;
  assign n61428 = pi18 ? n702 : ~n22299;
  assign n61429 = pi17 ? n46740 : n61428;
  assign n61430 = pi16 ? n919 : n61429;
  assign n61431 = pi15 ? n61334 : n61430;
  assign n61432 = pi14 ? n61431 : n22303;
  assign n61433 = pi15 ? n32 : n21226;
  assign n61434 = pi14 ? n22314 : n61433;
  assign n61435 = pi13 ? n61432 : n61434;
  assign n61436 = pi12 ? n61427 : n61435;
  assign n61437 = pi21 ? n14520 : n32;
  assign n61438 = pi20 ? n32 : n61437;
  assign n61439 = pi19 ? n61438 : n32;
  assign n61440 = pi18 ? n32 : n61439;
  assign n61441 = pi17 ? n32 : n61440;
  assign n61442 = pi16 ? n32 : n61441;
  assign n61443 = pi15 ? n61442 : n20831;
  assign n61444 = pi18 ? n18183 : ~n663;
  assign n61445 = pi17 ? n46997 : ~n61444;
  assign n61446 = pi16 ? n46995 : n61445;
  assign n61447 = pi16 ? n47001 : ~n2120;
  assign n61448 = pi15 ? n61446 : n61447;
  assign n61449 = pi14 ? n61443 : n61448;
  assign n61450 = pi14 ? n46992 : n47017;
  assign n61451 = pi13 ? n61449 : n61450;
  assign n61452 = pi16 ? n33623 : ~n2654;
  assign n61453 = pi17 ? n18395 : n21601;
  assign n61454 = pi16 ? n32 : n61453;
  assign n61455 = pi15 ? n61452 : n61454;
  assign n61456 = pi15 ? n33630 : n58837;
  assign n61457 = pi14 ? n61455 : n61456;
  assign n61458 = pi19 ? n266 : n1248;
  assign n61459 = pi18 ? n43189 : n61458;
  assign n61460 = pi17 ? n32 : n61459;
  assign n61461 = pi19 ? n18489 : n342;
  assign n61462 = pi19 ? n47025 : n247;
  assign n61463 = pi18 ? n61461 : n61462;
  assign n61464 = pi18 ? n47029 : ~n3786;
  assign n61465 = pi17 ? n61463 : ~n61464;
  assign n61466 = pi16 ? n61460 : ~n61465;
  assign n61467 = pi15 ? n61466 : n13392;
  assign n61468 = pi14 ? n61467 : n61288;
  assign n61469 = pi13 ? n61457 : n61468;
  assign n61470 = pi12 ? n61451 : n61469;
  assign n61471 = pi11 ? n61436 : n61470;
  assign n61472 = pi10 ? n61419 : n61471;
  assign n61473 = pi09 ? n61375 : n61472;
  assign n61474 = pi16 ? n1471 : ~n4100;
  assign n61475 = pi15 ? n61474 : n61395;
  assign n61476 = pi14 ? n61475 : n32;
  assign n61477 = pi13 ? n61391 : n61476;
  assign n61478 = pi14 ? n22424 : n22350;
  assign n61479 = pi15 ? n22347 : n47062;
  assign n61480 = pi14 ? n22348 : n61479;
  assign n61481 = pi13 ? n61478 : n61480;
  assign n61482 = pi12 ? n61477 : n61481;
  assign n61483 = pi20 ? n246 : n9641;
  assign n61484 = pi19 ? n61483 : ~n32;
  assign n61485 = pi18 ? n940 : ~n61484;
  assign n61486 = pi17 ? n32 : n61485;
  assign n61487 = pi16 ? n32 : n61486;
  assign n61488 = pi15 ? n20608 : n61487;
  assign n61489 = pi14 ? n61488 : n61411;
  assign n61490 = pi13 ? n61489 : n47084;
  assign n61491 = pi15 ? n40394 : n32;
  assign n61492 = pi14 ? n61414 : n61491;
  assign n61493 = pi14 ? n34408 : n21543;
  assign n61494 = pi13 ? n61492 : n61493;
  assign n61495 = pi12 ? n61490 : n61494;
  assign n61496 = pi11 ? n61482 : n61495;
  assign n61497 = pi15 ? n22087 : n32;
  assign n61498 = pi20 ? n1817 : n59970;
  assign n61499 = pi19 ? n61498 : ~n32;
  assign n61500 = pi18 ? n697 : ~n61499;
  assign n61501 = pi17 ? n32 : n61500;
  assign n61502 = pi16 ? n32 : n61501;
  assign n61503 = pi15 ? n33557 : n61502;
  assign n61504 = pi14 ? n61497 : n61503;
  assign n61505 = pi16 ? n1233 : ~n2749;
  assign n61506 = pi16 ? n1233 : ~n2518;
  assign n61507 = pi15 ? n61505 : n61506;
  assign n61508 = pi14 ? n61507 : n61506;
  assign n61509 = pi13 ? n61504 : n61508;
  assign n61510 = pi17 ? n46740 : n11416;
  assign n61511 = pi16 ? n568 : n61510;
  assign n61512 = pi18 ? n702 : ~n1333;
  assign n61513 = pi17 ? n46740 : n61512;
  assign n61514 = pi16 ? n568 : n61513;
  assign n61515 = pi15 ? n61511 : n61514;
  assign n61516 = pi14 ? n61515 : n22393;
  assign n61517 = pi20 ? n32 : n30091;
  assign n61518 = pi19 ? n61517 : n32;
  assign n61519 = pi18 ? n32 : n61518;
  assign n61520 = pi17 ? n32 : n61519;
  assign n61521 = pi16 ? n32 : n61520;
  assign n61522 = pi15 ? n20836 : n61521;
  assign n61523 = pi14 ? n22314 : n61522;
  assign n61524 = pi13 ? n61516 : n61523;
  assign n61525 = pi12 ? n61509 : n61524;
  assign n61526 = pi15 ? n61521 : n20836;
  assign n61527 = pi18 ? n18183 : ~n20828;
  assign n61528 = pi17 ? n46997 : ~n61527;
  assign n61529 = pi16 ? n47103 : n61528;
  assign n61530 = pi16 ? n47106 : ~n2120;
  assign n61531 = pi15 ? n61529 : n61530;
  assign n61532 = pi14 ? n61526 : n61531;
  assign n61533 = pi15 ? n36601 : n46991;
  assign n61534 = pi14 ? n61533 : n47017;
  assign n61535 = pi13 ? n61532 : n61534;
  assign n61536 = pi16 ? n33354 : ~n2654;
  assign n61537 = pi15 ? n61536 : n61454;
  assign n61538 = pi18 ? n323 : ~n35365;
  assign n61539 = pi17 ? n18395 : n61538;
  assign n61540 = pi16 ? n32 : n61539;
  assign n61541 = pi15 ? n61540 : n46655;
  assign n61542 = pi14 ? n61537 : n61541;
  assign n61543 = pi15 ? n61466 : n19972;
  assign n61544 = pi15 ? n13392 : n20531;
  assign n61545 = pi14 ? n61543 : n61544;
  assign n61546 = pi13 ? n61542 : n61545;
  assign n61547 = pi12 ? n61535 : n61546;
  assign n61548 = pi11 ? n61525 : n61547;
  assign n61549 = pi10 ? n61496 : n61548;
  assign n61550 = pi09 ? n61375 : n61549;
  assign n61551 = pi08 ? n61473 : n61550;
  assign n61552 = pi07 ? n61362 : n61551;
  assign n61553 = pi18 ? n24306 : n9012;
  assign n61554 = pi17 ? n32 : n61553;
  assign n61555 = pi16 ? n32 : n61554;
  assign n61556 = pi15 ? n32 : n61555;
  assign n61557 = pi16 ? n2958 : ~n2860;
  assign n61558 = pi16 ? n2860 : ~n2860;
  assign n61559 = pi15 ? n61557 : n61558;
  assign n61560 = pi14 ? n61556 : n61559;
  assign n61561 = pi13 ? n32 : n61560;
  assign n61562 = pi12 ? n32 : n61561;
  assign n61563 = pi11 ? n32 : n61562;
  assign n61564 = pi10 ? n32 : n61563;
  assign n61565 = pi18 ? n1758 : ~n41667;
  assign n61566 = pi18 ? n36162 : n323;
  assign n61567 = pi17 ? n61565 : ~n61566;
  assign n61568 = pi16 ? n32 : n61567;
  assign n61569 = pi17 ? n32 : n8820;
  assign n61570 = pi18 ? n16847 : n702;
  assign n61571 = pi17 ? n32 : n61570;
  assign n61572 = pi16 ? n61569 : ~n61571;
  assign n61573 = pi15 ? n61568 : n61572;
  assign n61574 = pi19 ? n18502 : ~n11107;
  assign n61575 = pi19 ? n266 : n60089;
  assign n61576 = pi18 ? n61574 : ~n61575;
  assign n61577 = pi20 ? n501 : n266;
  assign n61578 = pi19 ? n14463 : n61577;
  assign n61579 = pi18 ? n61578 : n595;
  assign n61580 = pi17 ? n61576 : n61579;
  assign n61581 = pi16 ? n16391 : ~n61580;
  assign n61582 = pi19 ? n5855 : n246;
  assign n61583 = pi18 ? n20172 : n61582;
  assign n61584 = pi20 ? n206 : n2358;
  assign n61585 = pi19 ? n61584 : ~n22652;
  assign n61586 = pi20 ? n206 : n101;
  assign n61587 = pi19 ? n61586 : ~n32;
  assign n61588 = pi18 ? n61585 : n61587;
  assign n61589 = pi17 ? n61583 : ~n61588;
  assign n61590 = pi16 ? n32 : n61589;
  assign n61591 = pi15 ? n61581 : n61590;
  assign n61592 = pi14 ? n61573 : n61591;
  assign n61593 = pi18 ? n18402 : n618;
  assign n61594 = pi17 ? n32 : n61593;
  assign n61595 = pi16 ? n61594 : ~n3946;
  assign n61596 = pi20 ? n206 : ~n11107;
  assign n61597 = pi19 ? n61596 : n32;
  assign n61598 = pi18 ? n32 : ~n61597;
  assign n61599 = pi17 ? n35241 : n61598;
  assign n61600 = pi16 ? n59546 : ~n61599;
  assign n61601 = pi15 ? n61595 : n61600;
  assign n61602 = pi14 ? n61601 : n15389;
  assign n61603 = pi13 ? n61592 : n61602;
  assign n61604 = pi14 ? n22424 : n15390;
  assign n61605 = pi15 ? n15123 : n15389;
  assign n61606 = pi18 ? n863 : ~n47144;
  assign n61607 = pi17 ? n32 : n61606;
  assign n61608 = pi16 ? n32 : n61607;
  assign n61609 = pi15 ? n61608 : n47175;
  assign n61610 = pi14 ? n61605 : n61609;
  assign n61611 = pi13 ? n61604 : n61610;
  assign n61612 = pi12 ? n61603 : n61611;
  assign n61613 = pi14 ? n22252 : n15127;
  assign n61614 = pi15 ? n33498 : n21928;
  assign n61615 = pi15 ? n32 : n22381;
  assign n61616 = pi14 ? n61614 : n61615;
  assign n61617 = pi13 ? n61613 : n61616;
  assign n61618 = pi12 ? n47218 : n61617;
  assign n61619 = pi11 ? n61612 : n61618;
  assign n61620 = pi18 ? n33787 : n7221;
  assign n61621 = pi17 ? n33785 : n61620;
  assign n61622 = pi16 ? n32 : n61621;
  assign n61623 = pi15 ? n21686 : n61622;
  assign n61624 = pi18 ? n33792 : n6059;
  assign n61625 = pi17 ? n32 : n61624;
  assign n61626 = pi16 ? n32 : n61625;
  assign n61627 = pi15 ? n61626 : n11848;
  assign n61628 = pi14 ? n61623 : n61627;
  assign n61629 = pi16 ? n1135 : ~n2749;
  assign n61630 = pi15 ? n61629 : n61329;
  assign n61631 = pi14 ? n61630 : n61329;
  assign n61632 = pi13 ? n61628 : n61631;
  assign n61633 = pi17 ? n46740 : n11849;
  assign n61634 = pi16 ? n919 : n61633;
  assign n61635 = pi15 ? n61634 : n22484;
  assign n61636 = pi14 ? n61635 : n22495;
  assign n61637 = pi18 ? n1379 : n34189;
  assign n61638 = pi17 ? n32 : n61637;
  assign n61639 = pi16 ? n32 : n61638;
  assign n61640 = pi15 ? n22505 : n61639;
  assign n61641 = pi15 ? n20836 : n21703;
  assign n61642 = pi14 ? n61640 : n61641;
  assign n61643 = pi13 ? n61636 : n61642;
  assign n61644 = pi12 ? n61632 : n61643;
  assign n61645 = pi18 ? n880 : n33824;
  assign n61646 = pi17 ? n32 : n61645;
  assign n61647 = pi16 ? n47258 : ~n61646;
  assign n61648 = pi15 ? n61521 : n61647;
  assign n61649 = pi18 ? n32 : n32381;
  assign n61650 = pi17 ? n32 : n61649;
  assign n61651 = pi16 ? n1214 : ~n61650;
  assign n61652 = pi15 ? n61651 : n47256;
  assign n61653 = pi14 ? n61648 : n61652;
  assign n61654 = pi15 ? n47256 : n46441;
  assign n61655 = pi15 ? n47264 : n46991;
  assign n61656 = pi14 ? n61654 : n61655;
  assign n61657 = pi13 ? n61653 : n61656;
  assign n61658 = pi18 ? n32 : n21749;
  assign n61659 = pi17 ? n32 : n61658;
  assign n61660 = pi16 ? n1214 : ~n61659;
  assign n61661 = pi15 ? n61660 : n33870;
  assign n61662 = pi19 ? n4982 : n1757;
  assign n61663 = pi18 ? n728 : ~n61662;
  assign n61664 = pi17 ? n32 : n61663;
  assign n61665 = pi18 ? n4380 : n1349;
  assign n61666 = pi17 ? n32 : n61665;
  assign n61667 = pi16 ? n61664 : ~n61666;
  assign n61668 = pi15 ? n11429 : n61667;
  assign n61669 = pi14 ? n61661 : n61668;
  assign n61670 = pi17 ? n16450 : n13682;
  assign n61671 = pi16 ? n129 : n61670;
  assign n61672 = pi15 ? n61671 : n20048;
  assign n61673 = pi15 ? n19969 : n47814;
  assign n61674 = pi14 ? n61672 : n61673;
  assign n61675 = pi13 ? n61669 : n61674;
  assign n61676 = pi12 ? n61657 : n61675;
  assign n61677 = pi11 ? n61644 : n61676;
  assign n61678 = pi10 ? n61619 : n61677;
  assign n61679 = pi09 ? n61564 : n61678;
  assign n61680 = pi16 ? n61594 : ~n2860;
  assign n61681 = pi15 ? n61680 : n61600;
  assign n61682 = pi14 ? n61681 : n32;
  assign n61683 = pi13 ? n61592 : n61682;
  assign n61684 = pi14 ? n22541 : n22543;
  assign n61685 = pi15 ? n15123 : n22540;
  assign n61686 = pi18 ? n863 : ~n2684;
  assign n61687 = pi17 ? n32 : n61686;
  assign n61688 = pi16 ? n32 : n61687;
  assign n61689 = pi15 ? n61688 : n47306;
  assign n61690 = pi14 ? n61685 : n61689;
  assign n61691 = pi13 ? n61684 : n61690;
  assign n61692 = pi12 ? n61683 : n61691;
  assign n61693 = pi15 ? n47184 : n13035;
  assign n61694 = pi14 ? n61693 : n47192;
  assign n61695 = pi13 ? n61694 : n47317;
  assign n61696 = pi14 ? n649 : n61615;
  assign n61697 = pi13 ? n61613 : n61696;
  assign n61698 = pi12 ? n61695 : n61697;
  assign n61699 = pi11 ? n61692 : n61698;
  assign n61700 = pi19 ? n17918 : ~n23806;
  assign n61701 = pi18 ? n33924 : n61700;
  assign n61702 = pi17 ? n61701 : n61620;
  assign n61703 = pi16 ? n32 : n61702;
  assign n61704 = pi15 ? n21543 : n61703;
  assign n61705 = pi18 ? n496 : ~n508;
  assign n61706 = pi17 ? n32 : n61705;
  assign n61707 = pi16 ? n32 : n61706;
  assign n61708 = pi15 ? n61626 : n61707;
  assign n61709 = pi14 ? n61704 : n61708;
  assign n61710 = pi16 ? n1233 : ~n2513;
  assign n61711 = pi15 ? n61710 : n61505;
  assign n61712 = pi14 ? n61711 : n61505;
  assign n61713 = pi13 ? n61709 : n61712;
  assign n61714 = pi19 ? n32 : n6158;
  assign n61715 = pi18 ? n61714 : ~n520;
  assign n61716 = pi17 ? n46740 : n61715;
  assign n61717 = pi16 ? n568 : n61716;
  assign n61718 = pi15 ? n61717 : n22588;
  assign n61719 = pi14 ? n61718 : n22495;
  assign n61720 = pi19 ? n41918 : n32;
  assign n61721 = pi18 ? n863 : n61720;
  assign n61722 = pi17 ? n32 : n61721;
  assign n61723 = pi16 ? n32 : n61722;
  assign n61724 = pi15 ? n22505 : n61723;
  assign n61725 = pi15 ? n14397 : n32361;
  assign n61726 = pi14 ? n61724 : n61725;
  assign n61727 = pi13 ? n61719 : n61726;
  assign n61728 = pi12 ? n61713 : n61727;
  assign n61729 = pi20 ? n246 : ~n7487;
  assign n61730 = pi19 ? n61729 : ~n32;
  assign n61731 = pi18 ? n880 : n61730;
  assign n61732 = pi17 ? n32 : n61731;
  assign n61733 = pi16 ? n47258 : ~n61732;
  assign n61734 = pi15 ? n20660 : n61733;
  assign n61735 = pi16 ? n1214 : ~n59711;
  assign n61736 = pi15 ? n61735 : n59560;
  assign n61737 = pi14 ? n61734 : n61736;
  assign n61738 = pi15 ? n60402 : n46991;
  assign n61739 = pi14 ? n61738 : n47342;
  assign n61740 = pi13 ? n61737 : n61739;
  assign n61741 = pi18 ? n33867 : ~n21749;
  assign n61742 = pi17 ? n33866 : n61741;
  assign n61743 = pi16 ? n32 : n61742;
  assign n61744 = pi15 ? n47261 : n61743;
  assign n61745 = pi15 ? n44870 : n61667;
  assign n61746 = pi14 ? n61744 : n61745;
  assign n61747 = pi17 ? n16450 : n20299;
  assign n61748 = pi16 ? n129 : n61747;
  assign n61749 = pi15 ? n61748 : n13684;
  assign n61750 = pi16 ? n129 : n13391;
  assign n61751 = pi15 ? n20048 : n61750;
  assign n61752 = pi14 ? n61749 : n61751;
  assign n61753 = pi13 ? n61746 : n61752;
  assign n61754 = pi12 ? n61740 : n61753;
  assign n61755 = pi11 ? n61728 : n61754;
  assign n61756 = pi10 ? n61699 : n61755;
  assign n61757 = pi09 ? n61564 : n61756;
  assign n61758 = pi08 ? n61679 : n61757;
  assign n61759 = pi20 ? n175 : ~n274;
  assign n61760 = pi19 ? n61759 : ~n531;
  assign n61761 = pi18 ? n61760 : n6163;
  assign n61762 = pi17 ? n32 : n61761;
  assign n61763 = pi16 ? n32 : n61762;
  assign n61764 = pi15 ? n32 : n61763;
  assign n61765 = pi16 ? n2958 : ~n2624;
  assign n61766 = pi19 ? n18741 : ~n32;
  assign n61767 = pi18 ? n32 : n61766;
  assign n61768 = pi17 ? n32 : n61767;
  assign n61769 = pi16 ? n61768 : ~n2624;
  assign n61770 = pi15 ? n61765 : n61769;
  assign n61771 = pi14 ? n61764 : n61770;
  assign n61772 = pi13 ? n32 : n61771;
  assign n61773 = pi12 ? n32 : n61772;
  assign n61774 = pi11 ? n32 : n61773;
  assign n61775 = pi10 ? n32 : n61774;
  assign n61776 = pi19 ? n32 : n58598;
  assign n61777 = pi18 ? n32 : n61776;
  assign n61778 = pi17 ? n32 : n61777;
  assign n61779 = pi19 ? n18782 : n56577;
  assign n61780 = pi20 ? n274 : n6822;
  assign n61781 = pi19 ? n61780 : n18282;
  assign n61782 = pi18 ? n61779 : ~n61781;
  assign n61783 = pi19 ? n9169 : ~n501;
  assign n61784 = pi18 ? n61783 : n323;
  assign n61785 = pi17 ? n61782 : ~n61784;
  assign n61786 = pi16 ? n61778 : n61785;
  assign n61787 = pi18 ? n36415 : n7519;
  assign n61788 = pi17 ? n32 : n61787;
  assign n61789 = pi16 ? n2745 : ~n61788;
  assign n61790 = pi15 ? n61786 : n61789;
  assign n61791 = pi20 ? n1076 : n9488;
  assign n61792 = pi19 ? n32 : n61791;
  assign n61793 = pi18 ? n32 : n61792;
  assign n61794 = pi17 ? n32 : n61793;
  assign n61795 = pi19 ? n36181 : ~n207;
  assign n61796 = pi18 ? n61795 : ~n18891;
  assign n61797 = pi19 ? n1490 : n247;
  assign n61798 = pi18 ? n61797 : n702;
  assign n61799 = pi17 ? n61796 : n61798;
  assign n61800 = pi16 ? n61794 : ~n61799;
  assign n61801 = pi19 ? n32 : ~n220;
  assign n61802 = pi19 ? n531 : n28686;
  assign n61803 = pi18 ? n61801 : ~n61802;
  assign n61804 = pi20 ? n1331 : n321;
  assign n61805 = pi19 ? n61804 : n19598;
  assign n61806 = pi18 ? n61805 : n28421;
  assign n61807 = pi17 ? n61803 : ~n61806;
  assign n61808 = pi16 ? n32 : n61807;
  assign n61809 = pi15 ? n61800 : n61808;
  assign n61810 = pi14 ? n61790 : n61809;
  assign n61811 = pi16 ? n2326 : ~n2860;
  assign n61812 = pi15 ? n61811 : n22540;
  assign n61813 = pi14 ? n61812 : n32;
  assign n61814 = pi13 ? n61810 : n61813;
  assign n61815 = pi20 ? n5854 : ~n260;
  assign n61816 = pi19 ? n61815 : n32;
  assign n61817 = pi18 ? n32 : n61816;
  assign n61818 = pi17 ? n32 : n61817;
  assign n61819 = pi16 ? n32 : n61818;
  assign n61820 = pi15 ? n32 : n61819;
  assign n61821 = pi17 ? n32 : n47296;
  assign n61822 = pi16 ? n32 : n61821;
  assign n61823 = pi15 ? n61822 : n47407;
  assign n61824 = pi14 ? n61820 : n61823;
  assign n61825 = pi13 ? n61684 : n61824;
  assign n61826 = pi12 ? n61814 : n61825;
  assign n61827 = pi19 ? n56386 : ~n32;
  assign n61828 = pi18 ? n47419 : ~n61827;
  assign n61829 = pi17 ? n16450 : n61828;
  assign n61830 = pi16 ? n32 : n61829;
  assign n61831 = pi15 ? n12756 : n61830;
  assign n61832 = pi14 ? n47415 : n61831;
  assign n61833 = pi18 ? n47429 : ~n47144;
  assign n61834 = pi17 ? n47428 : n61833;
  assign n61835 = pi16 ? n16391 : n61834;
  assign n61836 = pi15 ? n61835 : n47434;
  assign n61837 = pi15 ? n35650 : n47407;
  assign n61838 = pi14 ? n61836 : n61837;
  assign n61839 = pi13 ? n61832 : n61838;
  assign n61840 = pi15 ? n14967 : n648;
  assign n61841 = pi14 ? n61840 : n659;
  assign n61842 = pi13 ? n15391 : n61841;
  assign n61843 = pi12 ? n61839 : n61842;
  assign n61844 = pi11 ? n61826 : n61843;
  assign n61845 = pi19 ? n349 : ~n4670;
  assign n61846 = pi18 ? n32 : n61845;
  assign n61847 = pi17 ? n32 : n61846;
  assign n61848 = pi18 ? n47750 : ~n32;
  assign n61849 = pi17 ? n17346 : n61848;
  assign n61850 = pi16 ? n61847 : ~n61849;
  assign n61851 = pi15 ? n14397 : n61850;
  assign n61852 = pi19 ? n48234 : n342;
  assign n61853 = pi19 ? n20923 : n19280;
  assign n61854 = pi18 ? n61852 : n61853;
  assign n61855 = pi19 ? n18478 : n1757;
  assign n61856 = pi18 ? n61855 : n508;
  assign n61857 = pi17 ? n61854 : ~n61856;
  assign n61858 = pi16 ? n23573 : n61857;
  assign n61859 = pi19 ? n34319 : ~n236;
  assign n61860 = pi18 ? n863 : n61859;
  assign n61861 = pi17 ? n32 : n61860;
  assign n61862 = pi18 ? n44068 : n61853;
  assign n61863 = pi18 ? n19192 : n508;
  assign n61864 = pi17 ? n61862 : ~n61863;
  assign n61865 = pi16 ? n61861 : n61864;
  assign n61866 = pi15 ? n61858 : n61865;
  assign n61867 = pi14 ? n61851 : n61866;
  assign n61868 = pi16 ? n1135 : ~n2513;
  assign n61869 = pi15 ? n61868 : n61329;
  assign n61870 = pi14 ? n61869 : n61329;
  assign n61871 = pi13 ? n61867 : n61870;
  assign n61872 = pi18 ? n496 : ~n520;
  assign n61873 = pi17 ? n46740 : n61872;
  assign n61874 = pi16 ? n919 : n61873;
  assign n61875 = pi15 ? n61874 : n22669;
  assign n61876 = pi14 ? n61875 : n22681;
  assign n61877 = pi15 ? n22687 : n32;
  assign n61878 = pi14 ? n61877 : n21322;
  assign n61879 = pi13 ? n61876 : n61878;
  assign n61880 = pi12 ? n61871 : n61879;
  assign n61881 = pi20 ? n339 : n7487;
  assign n61882 = pi19 ? n61881 : n32;
  assign n61883 = pi18 ? n4380 : ~n61882;
  assign n61884 = pi17 ? n32 : n61883;
  assign n61885 = pi16 ? n47468 : ~n61884;
  assign n61886 = pi15 ? n32 : n61885;
  assign n61887 = pi16 ? n1214 : ~n2415;
  assign n61888 = pi15 ? n34146 : n61887;
  assign n61889 = pi14 ? n61886 : n61888;
  assign n61890 = pi20 ? n32 : n10446;
  assign n61891 = pi19 ? n61890 : ~n32;
  assign n61892 = pi18 ? n32 : n61891;
  assign n61893 = pi17 ? n32 : n61892;
  assign n61894 = pi16 ? n1214 : ~n61893;
  assign n61895 = pi15 ? n61894 : n47264;
  assign n61896 = pi17 ? n14395 : n2119;
  assign n61897 = pi16 ? n1214 : ~n61896;
  assign n61898 = pi17 ? n17119 : n2119;
  assign n61899 = pi16 ? n1214 : ~n61898;
  assign n61900 = pi15 ? n61897 : n61899;
  assign n61901 = pi14 ? n61895 : n61900;
  assign n61902 = pi13 ? n61889 : n61901;
  assign n61903 = pi18 ? n34087 : n2424;
  assign n61904 = pi17 ? n34086 : ~n61903;
  assign n61905 = pi16 ? n47483 : n61904;
  assign n61906 = pi15 ? n46441 : n61905;
  assign n61907 = pi18 ? n702 : ~n21749;
  assign n61908 = pi17 ? n32 : n61907;
  assign n61909 = pi16 ? n32 : n61908;
  assign n61910 = pi19 ? n34092 : n7399;
  assign n61911 = pi18 ? n917 : ~n61910;
  assign n61912 = pi17 ? n32 : n61911;
  assign n61913 = pi20 ? n339 : n12882;
  assign n61914 = pi19 ? n61913 : ~n22698;
  assign n61915 = pi18 ? n22696 : ~n61914;
  assign n61916 = pi18 ? n22703 : n6059;
  assign n61917 = pi17 ? n61915 : ~n61916;
  assign n61918 = pi16 ? n61912 : ~n61917;
  assign n61919 = pi15 ? n61909 : n61918;
  assign n61920 = pi14 ? n61906 : n61919;
  assign n61921 = pi17 ? n15845 : n13950;
  assign n61922 = pi16 ? n1014 : n61921;
  assign n61923 = pi15 ? n61922 : n20779;
  assign n61924 = pi16 ? n1014 : n19968;
  assign n61925 = pi15 ? n19972 : n61924;
  assign n61926 = pi14 ? n61923 : n61925;
  assign n61927 = pi13 ? n61920 : n61926;
  assign n61928 = pi12 ? n61902 : n61927;
  assign n61929 = pi11 ? n61880 : n61928;
  assign n61930 = pi10 ? n61844 : n61929;
  assign n61931 = pi09 ? n61775 : n61930;
  assign n61932 = pi19 ? n7363 : ~n1053;
  assign n61933 = pi19 ? n502 : ~n1105;
  assign n61934 = pi18 ? n61932 : n61933;
  assign n61935 = pi17 ? n32 : n61934;
  assign n61936 = pi16 ? n32 : n61935;
  assign n61937 = pi15 ? n32 : n61936;
  assign n61938 = pi16 ? n3946 : ~n2624;
  assign n61939 = pi15 ? n61765 : n61938;
  assign n61940 = pi14 ? n61937 : n61939;
  assign n61941 = pi13 ? n32 : n61940;
  assign n61942 = pi12 ? n32 : n61941;
  assign n61943 = pi11 ? n32 : n61942;
  assign n61944 = pi10 ? n32 : n61943;
  assign n61945 = pi19 ? n29527 : n18281;
  assign n61946 = pi18 ? n49467 : ~n61945;
  assign n61947 = pi17 ? n61946 : ~n61784;
  assign n61948 = pi16 ? n61778 : n61947;
  assign n61949 = pi15 ? n61948 : n61789;
  assign n61950 = pi14 ? n61949 : n61809;
  assign n61951 = pi16 ? n2326 : ~n3946;
  assign n61952 = pi15 ? n61951 : n22540;
  assign n61953 = pi14 ? n61952 : n32;
  assign n61954 = pi13 ? n61950 : n61953;
  assign n61955 = pi14 ? n1110 : n22812;
  assign n61956 = pi20 ? n5854 : ~n354;
  assign n61957 = pi19 ? n61956 : ~n1105;
  assign n61958 = pi18 ? n32 : n61957;
  assign n61959 = pi17 ? n32 : n61958;
  assign n61960 = pi16 ? n32 : n61959;
  assign n61961 = pi15 ? n1109 : n61960;
  assign n61962 = pi15 ? n13028 : n13904;
  assign n61963 = pi14 ? n61961 : n61962;
  assign n61964 = pi13 ? n61955 : n61963;
  assign n61965 = pi12 ? n61954 : n61964;
  assign n61966 = pi18 ? n32 : ~n2684;
  assign n61967 = pi17 ? n32 : n61966;
  assign n61968 = pi16 ? n32 : n61967;
  assign n61969 = pi15 ? n35668 : n61968;
  assign n61970 = pi14 ? n61969 : n61831;
  assign n61971 = pi13 ? n61970 : n61838;
  assign n61972 = pi15 ? n14967 : n32;
  assign n61973 = pi14 ? n61972 : n21320;
  assign n61974 = pi13 ? n15391 : n61973;
  assign n61975 = pi12 ? n61971 : n61974;
  assign n61976 = pi11 ? n61965 : n61975;
  assign n61977 = pi18 ? n61855 : n2627;
  assign n61978 = pi17 ? n61854 : ~n61977;
  assign n61979 = pi16 ? n23573 : n61978;
  assign n61980 = pi18 ? n19192 : n2627;
  assign n61981 = pi17 ? n61862 : ~n61980;
  assign n61982 = pi16 ? n61861 : n61981;
  assign n61983 = pi15 ? n61979 : n61982;
  assign n61984 = pi14 ? n61851 : n61983;
  assign n61985 = pi14 ? n61710 : n61711;
  assign n61986 = pi13 ? n61984 : n61985;
  assign n61987 = pi17 ? n46740 : n11846;
  assign n61988 = pi16 ? n568 : n61987;
  assign n61989 = pi15 ? n61988 : n22669;
  assign n61990 = pi18 ? n209 : ~n28193;
  assign n61991 = pi17 ? n32 : n61990;
  assign n61992 = pi16 ? n32 : n61991;
  assign n61993 = pi15 ? n22675 : n61992;
  assign n61994 = pi14 ? n61989 : n61993;
  assign n61995 = pi18 ? n17848 : n13945;
  assign n61996 = pi17 ? n32 : n61995;
  assign n61997 = pi16 ? n32 : n61996;
  assign n61998 = pi15 ? n61997 : n21464;
  assign n61999 = pi15 ? n21389 : n14397;
  assign n62000 = pi14 ? n61998 : n61999;
  assign n62001 = pi13 ? n61994 : n62000;
  assign n62002 = pi12 ? n61986 : n62001;
  assign n62003 = pi20 ? n339 : n266;
  assign n62004 = pi19 ? n62003 : n32;
  assign n62005 = pi18 ? n4380 : ~n62004;
  assign n62006 = pi17 ? n32 : n62005;
  assign n62007 = pi16 ? n47468 : ~n62006;
  assign n62008 = pi15 ? n32 : n62007;
  assign n62009 = pi16 ? n19652 : ~n2409;
  assign n62010 = pi15 ? n60814 : n62009;
  assign n62011 = pi14 ? n62008 : n62010;
  assign n62012 = pi13 ? n62011 : n61901;
  assign n62013 = pi18 ? n34087 : n605;
  assign n62014 = pi17 ? n34086 : ~n62013;
  assign n62015 = pi16 ? n47560 : n62014;
  assign n62016 = pi15 ? n46441 : n62015;
  assign n62017 = pi18 ? n702 : ~n805;
  assign n62018 = pi17 ? n32 : n62017;
  assign n62019 = pi16 ? n32 : n62018;
  assign n62020 = pi18 ? n566 : ~n61910;
  assign n62021 = pi17 ? n32 : n62020;
  assign n62022 = pi19 ? n22701 : ~n47564;
  assign n62023 = pi18 ? n62022 : n6059;
  assign n62024 = pi17 ? n61915 : ~n62023;
  assign n62025 = pi16 ? n62021 : ~n62024;
  assign n62026 = pi15 ? n62019 : n62025;
  assign n62027 = pi14 ? n62016 : n62026;
  assign n62028 = pi17 ? n15845 : n20475;
  assign n62029 = pi16 ? n465 : n62028;
  assign n62030 = pi15 ? n62029 : n13671;
  assign n62031 = pi16 ? n465 : n19968;
  assign n62032 = pi15 ? n19972 : n62031;
  assign n62033 = pi14 ? n62030 : n62032;
  assign n62034 = pi13 ? n62027 : n62033;
  assign n62035 = pi12 ? n62012 : n62034;
  assign n62036 = pi11 ? n62002 : n62035;
  assign n62037 = pi10 ? n61976 : n62036;
  assign n62038 = pi09 ? n61944 : n62037;
  assign n62039 = pi08 ? n61931 : n62038;
  assign n62040 = pi07 ? n61758 : n62039;
  assign n62041 = pi06 ? n61552 : n62040;
  assign n62042 = pi05 ? n61189 : n62041;
  assign n62043 = pi18 ? n32 : n49060;
  assign n62044 = pi17 ? n32 : n62043;
  assign n62045 = pi18 ? n28164 : n9012;
  assign n62046 = pi17 ? n62045 : n2855;
  assign n62047 = pi16 ? n62044 : ~n62046;
  assign n62048 = pi15 ? n32 : n62047;
  assign n62049 = pi17 ? n32 : n3621;
  assign n62050 = pi16 ? n62049 : ~n2856;
  assign n62051 = pi16 ? n3769 : ~n2860;
  assign n62052 = pi15 ? n62050 : n62051;
  assign n62053 = pi14 ? n62048 : n62052;
  assign n62054 = pi13 ? n32 : n62053;
  assign n62055 = pi12 ? n32 : n62054;
  assign n62056 = pi11 ? n32 : n62055;
  assign n62057 = pi10 ? n32 : n62056;
  assign n62058 = pi16 ? n2513 : ~n2860;
  assign n62059 = pi16 ? n2745 : ~n2856;
  assign n62060 = pi15 ? n62058 : n62059;
  assign n62061 = pi16 ? n2530 : ~n2860;
  assign n62062 = pi20 ? n428 : n9194;
  assign n62063 = pi20 ? n5854 : n342;
  assign n62064 = pi19 ? n62062 : ~n62063;
  assign n62065 = pi18 ? n32 : n62064;
  assign n62066 = pi17 ? n32 : n62065;
  assign n62067 = pi19 ? n9007 : ~n18677;
  assign n62068 = pi18 ? n62067 : n9012;
  assign n62069 = pi17 ? n62068 : n2623;
  assign n62070 = pi16 ? n62066 : ~n62069;
  assign n62071 = pi15 ? n62061 : n62070;
  assign n62072 = pi14 ? n62060 : n62071;
  assign n62073 = pi17 ? n32 : n2880;
  assign n62074 = pi16 ? n62073 : ~n2860;
  assign n62075 = pi15 ? n62074 : n1109;
  assign n62076 = pi14 ? n62075 : n32;
  assign n62077 = pi13 ? n62072 : n62076;
  assign n62078 = pi19 ? n358 : n1105;
  assign n62079 = pi18 ? n863 : ~n62078;
  assign n62080 = pi17 ? n32 : n62079;
  assign n62081 = pi16 ? n32 : n62080;
  assign n62082 = pi15 ? n32 : n62081;
  assign n62083 = pi15 ? n35947 : n25846;
  assign n62084 = pi14 ? n62082 : n62083;
  assign n62085 = pi13 ? n61955 : n62084;
  assign n62086 = pi12 ? n62077 : n62085;
  assign n62087 = pi15 ? n14156 : n22817;
  assign n62088 = pi14 ? n47687 : n62087;
  assign n62089 = pi13 ? n47678 : n62088;
  assign n62090 = pi14 ? n48187 : n32;
  assign n62091 = pi14 ? n24193 : n34217;
  assign n62092 = pi13 ? n62090 : n62091;
  assign n62093 = pi12 ? n62089 : n62092;
  assign n62094 = pi11 ? n62086 : n62093;
  assign n62095 = pi20 ? n10644 : ~n4279;
  assign n62096 = pi19 ? n62095 : n32;
  assign n62097 = pi18 ? n936 : ~n62096;
  assign n62098 = pi17 ? n32 : n62097;
  assign n62099 = pi16 ? n28804 : ~n62098;
  assign n62100 = pi15 ? n34224 : n62099;
  assign n62101 = pi16 ? n1471 : ~n2629;
  assign n62102 = pi16 ? n1214 : ~n2629;
  assign n62103 = pi15 ? n62101 : n62102;
  assign n62104 = pi14 ? n62100 : n62103;
  assign n62105 = pi17 ? n16848 : n12281;
  assign n62106 = pi16 ? n890 : n62105;
  assign n62107 = pi17 ? n16848 : n32883;
  assign n62108 = pi16 ? n890 : n62107;
  assign n62109 = pi15 ? n62106 : n62108;
  assign n62110 = pi14 ? n61868 : n62109;
  assign n62111 = pi13 ? n62104 : n62110;
  assign n62112 = pi15 ? n32 : n21695;
  assign n62113 = pi14 ? n62112 : n60801;
  assign n62114 = pi13 ? n22877 : n62113;
  assign n62115 = pi12 ? n62111 : n62114;
  assign n62116 = pi19 ? n342 : n274;
  assign n62117 = pi20 ? n274 : n4279;
  assign n62118 = pi20 ? n7939 : n2358;
  assign n62119 = pi19 ? n62117 : ~n62118;
  assign n62120 = pi18 ? n62116 : n62119;
  assign n62121 = pi20 ? n2358 : ~n6621;
  assign n62122 = pi20 ? n310 : ~n342;
  assign n62123 = pi19 ? n62121 : n62122;
  assign n62124 = pi18 ? n62123 : ~n43881;
  assign n62125 = pi17 ? n62120 : ~n62124;
  assign n62126 = pi16 ? n32 : n62125;
  assign n62127 = pi16 ? n47741 : ~n3769;
  assign n62128 = pi15 ? n62126 : n62127;
  assign n62129 = pi17 ? n47747 : n2292;
  assign n62130 = pi16 ? n47746 : ~n62129;
  assign n62131 = pi18 ? n47756 : n797;
  assign n62132 = pi17 ? n47755 : n62131;
  assign n62133 = pi16 ? n47752 : ~n62132;
  assign n62134 = pi15 ? n62130 : n62133;
  assign n62135 = pi14 ? n62128 : n62134;
  assign n62136 = pi18 ? n47782 : n2413;
  assign n62137 = pi17 ? n47781 : n62136;
  assign n62138 = pi16 ? n34526 : ~n62137;
  assign n62139 = pi18 ? n248 : n532;
  assign n62140 = pi17 ? n47792 : ~n62139;
  assign n62141 = pi16 ? n47788 : n62140;
  assign n62142 = pi15 ? n62138 : n62141;
  assign n62143 = pi14 ? n47899 : n62142;
  assign n62144 = pi13 ? n62135 : n62143;
  assign n62145 = pi18 ? n34305 : n605;
  assign n62146 = pi17 ? n34303 : ~n62145;
  assign n62147 = pi16 ? n32 : n62146;
  assign n62148 = pi15 ? n47810 : n62147;
  assign n62149 = pi18 ? n10078 : ~n34229;
  assign n62150 = pi17 ? n32 : n62149;
  assign n62151 = pi16 ? n32 : n62150;
  assign n62152 = pi18 ? n56127 : n34315;
  assign n62153 = pi17 ? n32 : n62152;
  assign n62154 = pi19 ? n19728 : ~n1817;
  assign n62155 = pi20 ? n1817 : ~n220;
  assign n62156 = pi20 ? n206 : ~n274;
  assign n62157 = pi19 ? n62155 : ~n62156;
  assign n62158 = pi18 ? n62154 : ~n62157;
  assign n62159 = pi20 ? n7939 : ~n6621;
  assign n62160 = pi19 ? n62159 : ~n3507;
  assign n62161 = pi18 ? n62160 : n32;
  assign n62162 = pi17 ? n62158 : n62161;
  assign n62163 = pi16 ? n62153 : n62162;
  assign n62164 = pi15 ? n62151 : n62163;
  assign n62165 = pi14 ? n62148 : n62164;
  assign n62166 = pi16 ? n568 : n20476;
  assign n62167 = pi15 ? n62166 : n20301;
  assign n62168 = pi15 ? n20048 : n47814;
  assign n62169 = pi14 ? n62167 : n62168;
  assign n62170 = pi13 ? n62165 : n62169;
  assign n62171 = pi12 ? n62144 : n62170;
  assign n62172 = pi11 ? n62115 : n62171;
  assign n62173 = pi10 ? n62094 : n62172;
  assign n62174 = pi09 ? n62057 : n62173;
  assign n62175 = pi16 ? n3625 : ~n2860;
  assign n62176 = pi17 ? n62068 : n2750;
  assign n62177 = pi16 ? n62066 : ~n62176;
  assign n62178 = pi15 ? n62175 : n62177;
  assign n62179 = pi14 ? n62060 : n62178;
  assign n62180 = pi17 ? n32 : n3509;
  assign n62181 = pi16 ? n62180 : ~n2624;
  assign n62182 = pi16 ? n17884 : n1108;
  assign n62183 = pi15 ? n62181 : n62182;
  assign n62184 = pi14 ? n62183 : n32;
  assign n62185 = pi13 ? n62179 : n62184;
  assign n62186 = pi15 ? n22923 : n62081;
  assign n62187 = pi14 ? n62186 : n47856;
  assign n62188 = pi13 ? n34349 : n62187;
  assign n62189 = pi12 ? n62185 : n62188;
  assign n62190 = pi19 ? n20006 : n1105;
  assign n62191 = pi18 ? n47659 : n62190;
  assign n62192 = pi17 ? n47658 : ~n62191;
  assign n62193 = pi16 ? n32 : n62192;
  assign n62194 = pi15 ? n22817 : n62193;
  assign n62195 = pi14 ? n62194 : n47677;
  assign n62196 = pi14 ? n47866 : n62087;
  assign n62197 = pi13 ? n62195 : n62196;
  assign n62198 = pi15 ? n22817 : n15389;
  assign n62199 = pi14 ? n62198 : n32;
  assign n62200 = pi14 ? n23771 : n34363;
  assign n62201 = pi13 ? n62199 : n62200;
  assign n62202 = pi12 ? n62197 : n62201;
  assign n62203 = pi11 ? n62189 : n62202;
  assign n62204 = pi20 ? n10644 : ~n428;
  assign n62205 = pi19 ? n62204 : n32;
  assign n62206 = pi18 ? n32 : ~n62205;
  assign n62207 = pi17 ? n32 : n62206;
  assign n62208 = pi16 ? n28677 : ~n62207;
  assign n62209 = pi15 ? n34224 : n62208;
  assign n62210 = pi16 ? n1214 : ~n3946;
  assign n62211 = pi15 ? n61392 : n62210;
  assign n62212 = pi14 ? n62209 : n62211;
  assign n62213 = pi16 ? n1135 : ~n2629;
  assign n62214 = pi16 ? n1233 : ~n2629;
  assign n62215 = pi15 ? n62213 : n62214;
  assign n62216 = pi17 ? n16848 : n46621;
  assign n62217 = pi16 ? n960 : n62216;
  assign n62218 = pi16 ? n960 : n62105;
  assign n62219 = pi15 ? n62217 : n62218;
  assign n62220 = pi14 ? n62215 : n62219;
  assign n62221 = pi13 ? n62212 : n62220;
  assign n62222 = pi15 ? n32 : n14394;
  assign n62223 = pi15 ? n14394 : n32;
  assign n62224 = pi14 ? n62222 : n62223;
  assign n62225 = pi13 ? n22969 : n62224;
  assign n62226 = pi12 ? n62221 : n62225;
  assign n62227 = pi16 ? n47741 : ~n2756;
  assign n62228 = pi15 ? n62126 : n62227;
  assign n62229 = pi17 ? n47747 : n2519;
  assign n62230 = pi16 ? n47746 : ~n62229;
  assign n62231 = pi18 ? n47756 : n2291;
  assign n62232 = pi17 ? n47755 : n62231;
  assign n62233 = pi16 ? n47752 : ~n62232;
  assign n62234 = pi15 ? n62230 : n62233;
  assign n62235 = pi14 ? n62228 : n62234;
  assign n62236 = pi17 ? n47765 : ~n2408;
  assign n62237 = pi16 ? n47764 : n62236;
  assign n62238 = pi15 ? n62237 : n47898;
  assign n62239 = pi16 ? n47901 : n62140;
  assign n62240 = pi15 ? n47785 : n62239;
  assign n62241 = pi14 ? n62238 : n62240;
  assign n62242 = pi13 ? n62235 : n62241;
  assign n62243 = pi18 ? n4492 : n32381;
  assign n62244 = pi17 ? n47807 : n62243;
  assign n62245 = pi16 ? n47803 : ~n62244;
  assign n62246 = pi18 ? n34305 : n2413;
  assign n62247 = pi17 ? n34303 : ~n62246;
  assign n62248 = pi16 ? n32 : n62247;
  assign n62249 = pi15 ? n62245 : n62248;
  assign n62250 = pi14 ? n62249 : n62164;
  assign n62251 = pi16 ? n568 : n13947;
  assign n62252 = pi15 ? n62251 : n21968;
  assign n62253 = pi16 ? n129 : n60268;
  assign n62254 = pi15 ? n13684 : n62253;
  assign n62255 = pi14 ? n62252 : n62254;
  assign n62256 = pi13 ? n62250 : n62255;
  assign n62257 = pi12 ? n62242 : n62256;
  assign n62258 = pi11 ? n62226 : n62257;
  assign n62259 = pi10 ? n62203 : n62258;
  assign n62260 = pi09 ? n62057 : n62259;
  assign n62261 = pi08 ? n62174 : n62260;
  assign n62262 = pi19 ? n18678 : n267;
  assign n62263 = pi19 ? n5707 : n349;
  assign n62264 = pi18 ? n62262 : n62263;
  assign n62265 = pi17 ? n62264 : ~n2616;
  assign n62266 = pi16 ? n17347 : n62265;
  assign n62267 = pi15 ? n32 : n62266;
  assign n62268 = pi16 ? n2958 : ~n2617;
  assign n62269 = pi16 ? n3061 : ~n2856;
  assign n62270 = pi15 ? n62268 : n62269;
  assign n62271 = pi14 ? n62267 : n62270;
  assign n62272 = pi13 ? n32 : n62271;
  assign n62273 = pi12 ? n32 : n62272;
  assign n62274 = pi11 ? n32 : n62273;
  assign n62275 = pi10 ? n32 : n62274;
  assign n62276 = pi19 ? n4670 : ~n18478;
  assign n62277 = pi19 ? n2025 : ~n220;
  assign n62278 = pi18 ? n62276 : ~n62277;
  assign n62279 = pi18 ? n1151 : n702;
  assign n62280 = pi17 ? n62278 : ~n62279;
  assign n62281 = pi16 ? n26461 : n62280;
  assign n62282 = pi17 ? n32 : n8653;
  assign n62283 = pi16 ? n62282 : ~n2617;
  assign n62284 = pi15 ? n62281 : n62283;
  assign n62285 = pi16 ? n2860 : ~n2624;
  assign n62286 = pi19 ? n1757 : n246;
  assign n62287 = pi18 ? n32 : n62286;
  assign n62288 = pi20 ? n220 : ~n220;
  assign n62289 = pi19 ? n62288 : n32;
  assign n62290 = pi18 ? n236 : ~n62289;
  assign n62291 = pi17 ? n62287 : ~n62290;
  assign n62292 = pi16 ? n32 : n62291;
  assign n62293 = pi15 ? n62285 : n62292;
  assign n62294 = pi14 ? n62284 : n62293;
  assign n62295 = pi19 ? n315 : ~n1331;
  assign n62296 = pi18 ? n16981 : ~n62295;
  assign n62297 = pi20 ? n17652 : ~n17665;
  assign n62298 = pi20 ? n18073 : n17669;
  assign n62299 = pi19 ? n62297 : ~n62298;
  assign n62300 = pi20 ? n310 : ~n260;
  assign n62301 = pi19 ? n62300 : n5635;
  assign n62302 = pi18 ? n62299 : ~n62301;
  assign n62303 = pi17 ? n62296 : ~n62302;
  assign n62304 = pi16 ? n32 : n62303;
  assign n62305 = pi15 ? n62304 : n24274;
  assign n62306 = pi14 ? n62305 : n32;
  assign n62307 = pi13 ? n62294 : n62306;
  assign n62308 = pi19 ? n10568 : ~n617;
  assign n62309 = pi18 ? n32 : n62308;
  assign n62310 = pi17 ? n32 : n62309;
  assign n62311 = pi16 ? n32 : n62310;
  assign n62312 = pi19 ? n6158 : ~n1105;
  assign n62313 = pi18 ? n32 : n62312;
  assign n62314 = pi17 ? n32 : n62313;
  assign n62315 = pi16 ? n32 : n62314;
  assign n62316 = pi15 ? n62311 : n62315;
  assign n62317 = pi15 ? n13913 : n15119;
  assign n62318 = pi14 ? n62316 : n62317;
  assign n62319 = pi13 ? n23089 : n62318;
  assign n62320 = pi12 ? n62307 : n62319;
  assign n62321 = pi14 ? n47968 : n1110;
  assign n62322 = pi13 ? n47967 : n62321;
  assign n62323 = pi14 ? n48187 : n34363;
  assign n62324 = pi13 ? n32 : n62323;
  assign n62325 = pi12 ? n62322 : n62324;
  assign n62326 = pi11 ? n62320 : n62325;
  assign n62327 = pi19 ? n207 : n236;
  assign n62328 = pi18 ? n41321 : n62327;
  assign n62329 = pi17 ? n32 : n62328;
  assign n62330 = pi18 ? n56104 : n18941;
  assign n62331 = pi18 ? n16449 : ~n32;
  assign n62332 = pi17 ? n62330 : n62331;
  assign n62333 = pi16 ? n62329 : ~n62332;
  assign n62334 = pi17 ? n32 : ~n10237;
  assign n62335 = pi16 ? n31252 : ~n62334;
  assign n62336 = pi15 ? n62333 : n62335;
  assign n62337 = pi16 ? n20208 : ~n3946;
  assign n62338 = pi16 ? n36009 : ~n2629;
  assign n62339 = pi15 ? n62337 : n62338;
  assign n62340 = pi14 ? n62336 : n62339;
  assign n62341 = pi17 ? n32 : n9428;
  assign n62342 = pi16 ? n1135 : ~n62341;
  assign n62343 = pi15 ? n62102 : n62342;
  assign n62344 = pi16 ? n890 : n62216;
  assign n62345 = pi15 ? n62344 : n62106;
  assign n62346 = pi14 ? n62343 : n62345;
  assign n62347 = pi13 ? n62340 : n62346;
  assign n62348 = pi15 ? n23056 : n32;
  assign n62349 = pi14 ? n23054 : n62348;
  assign n62350 = pi14 ? n21681 : n14398;
  assign n62351 = pi13 ? n62349 : n62350;
  assign n62352 = pi12 ? n62347 : n62351;
  assign n62353 = pi18 ? n48026 : ~n5436;
  assign n62354 = pi17 ? n48025 : n62353;
  assign n62355 = pi16 ? n32 : n62354;
  assign n62356 = pi17 ? n1028 : ~n2755;
  assign n62357 = pi16 ? n48033 : n62356;
  assign n62358 = pi15 ? n62355 : n62357;
  assign n62359 = pi20 ? n32 : n7479;
  assign n62360 = pi19 ? n62359 : ~n32;
  assign n62361 = pi18 ? n32 : n62360;
  assign n62362 = pi17 ? n47747 : n62361;
  assign n62363 = pi16 ? n48038 : ~n62362;
  assign n62364 = pi15 ? n62363 : n48050;
  assign n62365 = pi14 ? n62358 : n62364;
  assign n62366 = pi18 ? n28162 : n797;
  assign n62367 = pi17 ? n48065 : n62366;
  assign n62368 = pi16 ? n47770 : ~n62367;
  assign n62369 = pi15 ? n48062 : n62368;
  assign n62370 = pi14 ? n62369 : n48087;
  assign n62371 = pi13 ? n62365 : n62370;
  assign n62372 = pi15 ? n34576 : n11860;
  assign n62373 = pi17 ? n15832 : n1697;
  assign n62374 = pi16 ? n1233 : ~n62373;
  assign n62375 = pi15 ? n32 : n62374;
  assign n62376 = pi14 ? n62372 : n62375;
  assign n62377 = pi16 ? n30460 : n13947;
  assign n62378 = pi15 ? n62377 : n20477;
  assign n62379 = pi18 ? n32 : n18770;
  assign n62380 = pi17 ? n32 : n62379;
  assign n62381 = pi16 ? n129 : n62380;
  assign n62382 = pi15 ? n146 : n62381;
  assign n62383 = pi14 ? n62378 : n62382;
  assign n62384 = pi13 ? n62376 : n62383;
  assign n62385 = pi12 ? n62371 : n62384;
  assign n62386 = pi11 ? n62352 : n62385;
  assign n62387 = pi10 ? n62326 : n62386;
  assign n62388 = pi09 ? n62275 : n62387;
  assign n62389 = pi18 ? n1151 : n8884;
  assign n62390 = pi17 ? n62278 : ~n62389;
  assign n62391 = pi16 ? n26461 : n62390;
  assign n62392 = pi15 ? n62391 : n62283;
  assign n62393 = pi15 ? n61558 : n62292;
  assign n62394 = pi14 ? n62392 : n62393;
  assign n62395 = pi19 ? n358 : n50722;
  assign n62396 = pi20 ? n1331 : n428;
  assign n62397 = pi19 ? n62396 : ~n617;
  assign n62398 = pi18 ? n62395 : n62397;
  assign n62399 = pi17 ? n48400 : n62398;
  assign n62400 = pi16 ? n32 : n62399;
  assign n62401 = pi15 ? n62400 : n22923;
  assign n62402 = pi14 ? n62401 : n32;
  assign n62403 = pi13 ? n62394 : n62402;
  assign n62404 = pi14 ? n23828 : n23582;
  assign n62405 = pi19 ? n10568 : ~n2614;
  assign n62406 = pi18 ? n32 : n62405;
  assign n62407 = pi17 ? n32 : n62406;
  assign n62408 = pi16 ? n32 : n62407;
  assign n62409 = pi19 ? n6158 : ~n617;
  assign n62410 = pi18 ? n32 : n62409;
  assign n62411 = pi17 ? n32 : n62410;
  assign n62412 = pi16 ? n32 : n62411;
  assign n62413 = pi15 ? n62408 : n62412;
  assign n62414 = pi14 ? n62413 : n62317;
  assign n62415 = pi13 ? n62404 : n62414;
  assign n62416 = pi12 ? n62403 : n62415;
  assign n62417 = pi19 ? n5741 : n617;
  assign n62418 = pi18 ? n32 : ~n62417;
  assign n62419 = pi17 ? n32 : n62418;
  assign n62420 = pi16 ? n32 : n62419;
  assign n62421 = pi15 ? n22817 : n62420;
  assign n62422 = pi18 ? n1613 : ~n47667;
  assign n62423 = pi17 ? n32 : n62422;
  assign n62424 = pi16 ? n32 : n62423;
  assign n62425 = pi15 ? n62424 : n47965;
  assign n62426 = pi14 ? n62421 : n62425;
  assign n62427 = pi13 ? n62426 : n62321;
  assign n62428 = pi12 ? n62427 : n62324;
  assign n62429 = pi11 ? n62416 : n62428;
  assign n62430 = pi18 ? n237 : ~n4098;
  assign n62431 = pi17 ? n32 : ~n62430;
  assign n62432 = pi16 ? n31252 : ~n62431;
  assign n62433 = pi15 ? n62333 : n62432;
  assign n62434 = pi16 ? n20208 : ~n4100;
  assign n62435 = pi16 ? n36009 : ~n3946;
  assign n62436 = pi15 ? n62434 : n62435;
  assign n62437 = pi14 ? n62433 : n62436;
  assign n62438 = pi21 ? n100 : n405;
  assign n62439 = pi20 ? n32 : n62438;
  assign n62440 = pi19 ? n62439 : ~n32;
  assign n62441 = pi18 ? n32 : n62440;
  assign n62442 = pi17 ? n32 : n62441;
  assign n62443 = pi16 ? n1135 : ~n62442;
  assign n62444 = pi15 ? n62210 : n62443;
  assign n62445 = pi17 ? n16848 : n47164;
  assign n62446 = pi16 ? n890 : n62445;
  assign n62447 = pi15 ? n62446 : n62344;
  assign n62448 = pi14 ? n62444 : n62447;
  assign n62449 = pi13 ? n62437 : n62448;
  assign n62450 = pi15 ? n23127 : n23054;
  assign n62451 = pi14 ? n62450 : n62348;
  assign n62452 = pi15 ? n32 : n21686;
  assign n62453 = pi14 ? n62452 : n14398;
  assign n62454 = pi13 ? n62451 : n62453;
  assign n62455 = pi12 ? n62449 : n62454;
  assign n62456 = pi18 ? n48026 : ~n23291;
  assign n62457 = pi17 ? n48025 : n62456;
  assign n62458 = pi16 ? n32 : n62457;
  assign n62459 = pi16 ? n48033 : n34657;
  assign n62460 = pi15 ? n62458 : n62459;
  assign n62461 = pi17 ? n47747 : n61066;
  assign n62462 = pi16 ? n48038 : ~n62461;
  assign n62463 = pi18 ? n48047 : n32919;
  assign n62464 = pi17 ? n48046 : n62463;
  assign n62465 = pi16 ? n48042 : ~n62464;
  assign n62466 = pi15 ? n62462 : n62465;
  assign n62467 = pi14 ? n62460 : n62466;
  assign n62468 = pi18 ? n48083 : n797;
  assign n62469 = pi17 ? n48081 : ~n62468;
  assign n62470 = pi16 ? n48078 : n62469;
  assign n62471 = pi15 ? n48168 : n62470;
  assign n62472 = pi14 ? n48165 : n62471;
  assign n62473 = pi13 ? n62467 : n62472;
  assign n62474 = pi14 ? n34580 : n62375;
  assign n62475 = pi16 ? n30460 : n21231;
  assign n62476 = pi15 ? n62475 : n20477;
  assign n62477 = pi16 ? n32 : n62380;
  assign n62478 = pi15 ? n146 : n62477;
  assign n62479 = pi14 ? n62476 : n62478;
  assign n62480 = pi13 ? n62474 : n62479;
  assign n62481 = pi12 ? n62473 : n62480;
  assign n62482 = pi11 ? n62455 : n62481;
  assign n62483 = pi10 ? n62429 : n62482;
  assign n62484 = pi09 ? n62275 : n62483;
  assign n62485 = pi08 ? n62388 : n62484;
  assign n62486 = pi07 ? n62261 : n62485;
  assign n62487 = pi17 ? n36579 : ~n2736;
  assign n62488 = pi16 ? n32 : n62487;
  assign n62489 = pi15 ? n32 : n62488;
  assign n62490 = pi17 ? n2531 : ~n2736;
  assign n62491 = pi16 ? n32 : n62490;
  assign n62492 = pi17 ? n36006 : ~n2855;
  assign n62493 = pi16 ? n32 : n62492;
  assign n62494 = pi15 ? n62491 : n62493;
  assign n62495 = pi14 ? n62489 : n62494;
  assign n62496 = pi13 ? n32 : n62495;
  assign n62497 = pi12 ? n32 : n62496;
  assign n62498 = pi11 ? n32 : n62497;
  assign n62499 = pi10 ? n32 : n62498;
  assign n62500 = pi19 ? n18211 : n32336;
  assign n62501 = pi18 ? n268 : n62500;
  assign n62502 = pi17 ? n62501 : ~n2736;
  assign n62503 = pi16 ? n32 : n62502;
  assign n62504 = pi15 ? n10455 : n62503;
  assign n62505 = pi20 ? n175 : ~n246;
  assign n62506 = pi19 ? n32 : n62505;
  assign n62507 = pi18 ? n32 : n62506;
  assign n62508 = pi17 ? n32 : n62507;
  assign n62509 = pi18 ? n31850 : n18668;
  assign n62510 = pi18 ? n618 : ~n702;
  assign n62511 = pi17 ? n62509 : ~n62510;
  assign n62512 = pi16 ? n62508 : ~n62511;
  assign n62513 = pi19 ? n32848 : n18489;
  assign n62514 = pi20 ? n206 : ~n1817;
  assign n62515 = pi19 ? n62514 : ~n617;
  assign n62516 = pi18 ? n62513 : n62515;
  assign n62517 = pi17 ? n32 : n62516;
  assign n62518 = pi16 ? n32 : n62517;
  assign n62519 = pi15 ? n62512 : n62518;
  assign n62520 = pi14 ? n62504 : n62519;
  assign n62521 = pi13 ? n62520 : n23256;
  assign n62522 = pi15 ? n32 : n24185;
  assign n62523 = pi14 ? n23160 : n62522;
  assign n62524 = pi15 ? n48548 : n34616;
  assign n62525 = pi14 ? n62524 : n48198;
  assign n62526 = pi13 ? n62523 : n62525;
  assign n62527 = pi12 ? n62521 : n62526;
  assign n62528 = pi14 ? n48219 : n34348;
  assign n62529 = pi13 ? n48214 : n62528;
  assign n62530 = pi14 ? n48187 : n1110;
  assign n62531 = pi19 ? n1574 : ~n1105;
  assign n62532 = pi18 ? n32 : n62531;
  assign n62533 = pi17 ? n32 : n62532;
  assign n62534 = pi16 ? n32 : n62533;
  assign n62535 = pi15 ? n62534 : n32;
  assign n62536 = pi14 ? n62535 : n34625;
  assign n62537 = pi13 ? n62530 : n62536;
  assign n62538 = pi12 ? n62529 : n62537;
  assign n62539 = pi11 ? n62527 : n62538;
  assign n62540 = pi18 ? n6145 : n4098;
  assign n62541 = pi17 ? n1219 : ~n62540;
  assign n62542 = pi16 ? n32 : n62541;
  assign n62543 = pi18 ? n19232 : n4098;
  assign n62544 = pi17 ? n1219 : ~n62543;
  assign n62545 = pi16 ? n17434 : n62544;
  assign n62546 = pi15 ? n62542 : n62545;
  assign n62547 = pi18 ? n32 : n47144;
  assign n62548 = pi17 ? n32 : n62547;
  assign n62549 = pi16 ? n1808 : ~n62548;
  assign n62550 = pi16 ? n1808 : ~n3946;
  assign n62551 = pi15 ? n62549 : n62550;
  assign n62552 = pi14 ? n62546 : n62551;
  assign n62553 = pi15 ? n62210 : n61392;
  assign n62554 = pi18 ? n1395 : ~n496;
  assign n62555 = pi17 ? n32 : n62554;
  assign n62556 = pi17 ? n32 : n47164;
  assign n62557 = pi16 ? n62555 : n62556;
  assign n62558 = pi19 ? n8644 : n349;
  assign n62559 = pi18 ? n276 : ~n62558;
  assign n62560 = pi17 ? n32 : n62559;
  assign n62561 = pi16 ? n62560 : n23188;
  assign n62562 = pi15 ? n62557 : n62561;
  assign n62563 = pi14 ? n62553 : n62562;
  assign n62564 = pi13 ? n62552 : n62563;
  assign n62565 = pi15 ? n23203 : n32;
  assign n62566 = pi14 ? n23198 : n62565;
  assign n62567 = pi18 ? n12811 : n9578;
  assign n62568 = pi17 ? n1978 : n62567;
  assign n62569 = pi16 ? n32 : n62568;
  assign n62570 = pi19 ? n5707 : n4126;
  assign n62571 = pi20 ? n321 : ~n501;
  assign n62572 = pi19 ? n62571 : n32;
  assign n62573 = pi18 ? n62570 : ~n62572;
  assign n62574 = pi17 ? n1978 : ~n62573;
  assign n62575 = pi16 ? n32 : n62574;
  assign n62576 = pi15 ? n62569 : n62575;
  assign n62577 = pi14 ? n60592 : n62576;
  assign n62578 = pi13 ? n62566 : n62577;
  assign n62579 = pi12 ? n62564 : n62578;
  assign n62580 = pi19 ? n53174 : ~n32;
  assign n62581 = pi18 ? n496 : ~n62580;
  assign n62582 = pi17 ? n16450 : n62581;
  assign n62583 = pi16 ? n32 : n62582;
  assign n62584 = pi17 ? n48271 : ~n2517;
  assign n62585 = pi16 ? n32 : n62584;
  assign n62586 = pi15 ? n62583 : n62585;
  assign n62587 = pi20 ? n32 : n16168;
  assign n62588 = pi19 ? n62587 : ~n32;
  assign n62589 = pi18 ? n880 : ~n62588;
  assign n62590 = pi17 ? n1219 : ~n62589;
  assign n62591 = pi16 ? n48276 : ~n62590;
  assign n62592 = pi15 ? n62591 : n48358;
  assign n62593 = pi14 ? n62586 : n62592;
  assign n62594 = pi15 ? n48362 : n48286;
  assign n62595 = pi18 ? n6063 : ~n797;
  assign n62596 = pi17 ? n48292 : n62595;
  assign n62597 = pi16 ? n32 : n62596;
  assign n62598 = pi15 ? n48290 : n62597;
  assign n62599 = pi14 ? n62594 : n62598;
  assign n62600 = pi13 ? n62593 : n62599;
  assign n62601 = pi17 ? n34706 : ~n2408;
  assign n62602 = pi16 ? n32 : n62601;
  assign n62603 = pi15 ? n62602 : n20831;
  assign n62604 = pi19 ? n5004 : ~n32;
  assign n62605 = pi18 ? n62604 : ~n32;
  assign n62606 = pi17 ? n34711 : n62605;
  assign n62607 = pi16 ? n1233 : ~n62606;
  assign n62608 = pi15 ? n32 : n62607;
  assign n62609 = pi14 ? n62603 : n62608;
  assign n62610 = pi19 ? n25120 : n507;
  assign n62611 = pi18 ? n56696 : ~n62610;
  assign n62612 = pi17 ? n32 : n62611;
  assign n62613 = pi18 ? n34720 : ~n22604;
  assign n62614 = pi17 ? n34719 : n62613;
  assign n62615 = pi16 ? n62612 : ~n62614;
  assign n62616 = pi15 ? n62615 : n20477;
  assign n62617 = pi16 ? n465 : n145;
  assign n62618 = pi16 ? n1014 : n19971;
  assign n62619 = pi15 ? n62617 : n62618;
  assign n62620 = pi14 ? n62616 : n62619;
  assign n62621 = pi13 ? n62609 : n62620;
  assign n62622 = pi12 ? n62600 : n62621;
  assign n62623 = pi11 ? n62579 : n62622;
  assign n62624 = pi10 ? n62539 : n62623;
  assign n62625 = pi09 ? n62499 : n62624;
  assign n62626 = pi18 ? n237 : ~n702;
  assign n62627 = pi17 ? n62509 : ~n62626;
  assign n62628 = pi16 ? n49781 : ~n62627;
  assign n62629 = pi15 ? n62628 : n62518;
  assign n62630 = pi14 ? n62504 : n62629;
  assign n62631 = pi13 ? n62630 : n23163;
  assign n62632 = pi19 ? n4126 : ~n236;
  assign n62633 = pi18 ? n32 : n62632;
  assign n62634 = pi17 ? n32 : n62633;
  assign n62635 = pi16 ? n32 : n62634;
  assign n62636 = pi15 ? n32 : n62635;
  assign n62637 = pi14 ? n23250 : n62636;
  assign n62638 = pi15 ? n48389 : n23836;
  assign n62639 = pi14 ? n62638 : n34537;
  assign n62640 = pi13 ? n62637 : n62639;
  assign n62641 = pi12 ? n62631 : n62640;
  assign n62642 = pi19 ? n48202 : ~n2614;
  assign n62643 = pi18 ? n6118 : n62642;
  assign n62644 = pi17 ? n2954 : n62643;
  assign n62645 = pi16 ? n32 : n62644;
  assign n62646 = pi15 ? n22923 : n62645;
  assign n62647 = pi14 ? n62646 : n48213;
  assign n62648 = pi14 ? n48325 : n22923;
  assign n62649 = pi13 ? n62647 : n62648;
  assign n62650 = pi19 ? n857 : ~n1105;
  assign n62651 = pi18 ? n32 : n62650;
  assign n62652 = pi17 ? n32 : n62651;
  assign n62653 = pi16 ? n32 : n62652;
  assign n62654 = pi15 ? n23011 : n62653;
  assign n62655 = pi14 ? n62654 : n32;
  assign n62656 = pi14 ? n22812 : n34625;
  assign n62657 = pi13 ? n62655 : n62656;
  assign n62658 = pi12 ? n62649 : n62657;
  assign n62659 = pi11 ? n62641 : n62658;
  assign n62660 = pi18 ? n6145 : n702;
  assign n62661 = pi17 ? n1219 : ~n62660;
  assign n62662 = pi16 ? n32 : n62661;
  assign n62663 = pi17 ? n1219 : ~n49416;
  assign n62664 = pi16 ? n17434 : n62663;
  assign n62665 = pi15 ? n62662 : n62664;
  assign n62666 = pi17 ? n32 : n2861;
  assign n62667 = pi16 ? n1808 : ~n62666;
  assign n62668 = pi16 ? n1808 : ~n4100;
  assign n62669 = pi15 ? n62667 : n62668;
  assign n62670 = pi14 ? n62665 : n62669;
  assign n62671 = pi16 ? n1214 : ~n4100;
  assign n62672 = pi15 ? n62671 : n61474;
  assign n62673 = pi16 ? n586 : n12270;
  assign n62674 = pi19 ? n785 : n502;
  assign n62675 = pi18 ? n32 : ~n62674;
  assign n62676 = pi17 ? n32 : n62675;
  assign n62677 = pi16 ? n62676 : n23036;
  assign n62678 = pi15 ? n62673 : n62677;
  assign n62679 = pi14 ? n62672 : n62678;
  assign n62680 = pi13 ? n62670 : n62679;
  assign n62681 = pi15 ? n19172 : n476;
  assign n62682 = pi14 ? n23275 : n62681;
  assign n62683 = pi15 ? n476 : n21786;
  assign n62684 = pi18 ? n12811 : n21683;
  assign n62685 = pi17 ? n1978 : n62684;
  assign n62686 = pi16 ? n32 : n62685;
  assign n62687 = pi20 ? n321 : ~n10889;
  assign n62688 = pi19 ? n62687 : n32;
  assign n62689 = pi18 ? n62570 : ~n62688;
  assign n62690 = pi17 ? n1978 : ~n62689;
  assign n62691 = pi16 ? n32 : n62690;
  assign n62692 = pi15 ? n62686 : n62691;
  assign n62693 = pi14 ? n62683 : n62692;
  assign n62694 = pi13 ? n62682 : n62693;
  assign n62695 = pi12 ? n62680 : n62694;
  assign n62696 = pi19 ? n56061 : ~n32;
  assign n62697 = pi18 ? n496 : ~n62696;
  assign n62698 = pi17 ? n16450 : n62697;
  assign n62699 = pi16 ? n32 : n62698;
  assign n62700 = pi17 ? n48271 : ~n2748;
  assign n62701 = pi16 ? n32 : n62700;
  assign n62702 = pi15 ? n62699 : n62701;
  assign n62703 = pi17 ? n1219 : ~n12081;
  assign n62704 = pi16 ? n48276 : ~n62703;
  assign n62705 = pi15 ? n62704 : n48588;
  assign n62706 = pi14 ? n62702 : n62705;
  assign n62707 = pi18 ? n6063 : ~n2291;
  assign n62708 = pi17 ? n48292 : n62707;
  assign n62709 = pi16 ? n32 : n62708;
  assign n62710 = pi15 ? n48290 : n62709;
  assign n62711 = pi14 ? n48365 : n62710;
  assign n62712 = pi13 ? n62706 : n62711;
  assign n62713 = pi17 ? n34706 : ~n2292;
  assign n62714 = pi16 ? n32 : n62713;
  assign n62715 = pi15 ? n62714 : n32;
  assign n62716 = pi18 ? n62604 : ~n5158;
  assign n62717 = pi17 ? n34711 : n62716;
  assign n62718 = pi16 ? n1233 : ~n62717;
  assign n62719 = pi15 ? n32 : n62718;
  assign n62720 = pi14 ? n62715 : n62719;
  assign n62721 = pi18 ? n34720 : ~n13940;
  assign n62722 = pi17 ? n34719 : n62721;
  assign n62723 = pi16 ? n62612 : ~n62722;
  assign n62724 = pi15 ? n62723 : n13948;
  assign n62725 = pi16 ? n1014 : n670;
  assign n62726 = pi15 ? n62725 : n62618;
  assign n62727 = pi14 ? n62724 : n62726;
  assign n62728 = pi13 ? n62720 : n62727;
  assign n62729 = pi12 ? n62712 : n62728;
  assign n62730 = pi11 ? n62695 : n62729;
  assign n62731 = pi10 ? n62659 : n62730;
  assign n62732 = pi09 ? n62499 : n62731;
  assign n62733 = pi08 ? n62625 : n62732;
  assign n62734 = pi18 ? n32 : n33878;
  assign n62735 = pi17 ? n62734 : ~n2731;
  assign n62736 = pi16 ? n32 : n62735;
  assign n62737 = pi15 ? n32 : n62736;
  assign n62738 = pi19 ? n531 : ~n1757;
  assign n62739 = pi18 ? n32 : n62738;
  assign n62740 = pi17 ? n62739 : ~n2736;
  assign n62741 = pi16 ? n32 : n62740;
  assign n62742 = pi15 ? n62491 : n62741;
  assign n62743 = pi14 ? n62737 : n62742;
  assign n62744 = pi13 ? n32 : n62743;
  assign n62745 = pi12 ? n32 : n62744;
  assign n62746 = pi11 ? n32 : n62745;
  assign n62747 = pi10 ? n32 : n62746;
  assign n62748 = pi19 ? n221 : n4406;
  assign n62749 = pi18 ? n32 : n62748;
  assign n62750 = pi19 ? n32 : n10447;
  assign n62751 = pi18 ? n32 : n62750;
  assign n62752 = pi17 ? n62749 : ~n62751;
  assign n62753 = pi16 ? n32 : n62752;
  assign n62754 = pi19 ? n4982 : n236;
  assign n62755 = pi18 ? n32 : n62754;
  assign n62756 = pi17 ? n62755 : ~n2731;
  assign n62757 = pi16 ? n32 : n62756;
  assign n62758 = pi15 ? n62753 : n62757;
  assign n62759 = pi19 ? n5748 : ~n6050;
  assign n62760 = pi18 ? n32 : n62759;
  assign n62761 = pi18 ? n56198 : n1750;
  assign n62762 = pi17 ? n62760 : ~n62761;
  assign n62763 = pi16 ? n32 : n62762;
  assign n62764 = pi19 ? n18741 : n1757;
  assign n62765 = pi20 ? n3523 : ~n5854;
  assign n62766 = pi19 ? n62765 : n32;
  assign n62767 = pi18 ? n62764 : n62766;
  assign n62768 = pi17 ? n32 : n62767;
  assign n62769 = pi16 ? n32 : n62768;
  assign n62770 = pi15 ? n62763 : n62769;
  assign n62771 = pi14 ? n62758 : n62770;
  assign n62772 = pi13 ? n62771 : n23253;
  assign n62773 = pi19 ? n1740 : ~n236;
  assign n62774 = pi18 ? n32 : n62773;
  assign n62775 = pi17 ? n32 : n62774;
  assign n62776 = pi16 ? n32 : n62775;
  assign n62777 = pi15 ? n32 : n62776;
  assign n62778 = pi14 ? n23326 : n62777;
  assign n62779 = pi19 ? n349 : ~n56769;
  assign n62780 = pi18 ? n32 : n62779;
  assign n62781 = pi17 ? n32 : n62780;
  assign n62782 = pi16 ? n32 : n62781;
  assign n62783 = pi19 ? n343 : n5626;
  assign n62784 = pi18 ? n32 : n62783;
  assign n62785 = pi17 ? n32 : n62784;
  assign n62786 = pi16 ? n32 : n62785;
  assign n62787 = pi15 ? n62782 : n62786;
  assign n62788 = pi14 ? n62787 : n48385;
  assign n62789 = pi13 ? n62778 : n62788;
  assign n62790 = pi12 ? n62772 : n62789;
  assign n62791 = pi14 ? n48325 : n23160;
  assign n62792 = pi13 ? n48424 : n62791;
  assign n62793 = pi14 ? n15127 : n24327;
  assign n62794 = pi19 ? n857 : n422;
  assign n62795 = pi18 ? n858 : n62794;
  assign n62796 = pi19 ? n59860 : n47141;
  assign n62797 = pi18 ? n62796 : ~n702;
  assign n62798 = pi17 ? n62795 : n62797;
  assign n62799 = pi16 ? n32 : n62798;
  assign n62800 = pi15 ? n22437 : n62799;
  assign n62801 = pi14 ? n22925 : n62800;
  assign n62802 = pi13 ? n62793 : n62801;
  assign n62803 = pi12 ? n62792 : n62802;
  assign n62804 = pi11 ? n62790 : n62803;
  assign n62805 = pi17 ? n1219 : ~n2750;
  assign n62806 = pi16 ? n32 : n62805;
  assign n62807 = pi17 ? n1219 : ~n31241;
  assign n62808 = pi16 ? n32 : n62807;
  assign n62809 = pi15 ? n62806 : n62808;
  assign n62810 = pi16 ? n1808 : ~n2860;
  assign n62811 = pi15 ? n62810 : n62668;
  assign n62812 = pi14 ? n62809 : n62811;
  assign n62813 = pi16 ? n1135 : ~n3946;
  assign n62814 = pi15 ? n62813 : n61868;
  assign n62815 = pi16 ? n890 : n12270;
  assign n62816 = pi15 ? n62815 : n23359;
  assign n62817 = pi14 ? n62814 : n62816;
  assign n62818 = pi13 ? n62812 : n62817;
  assign n62819 = pi14 ? n23370 : n21929;
  assign n62820 = pi15 ? n62686 : n48459;
  assign n62821 = pi14 ? n22213 : n62820;
  assign n62822 = pi13 ? n62819 : n62821;
  assign n62823 = pi12 ? n62818 : n62822;
  assign n62824 = pi21 ? n100 : n242;
  assign n62825 = pi20 ? n32 : n62824;
  assign n62826 = pi19 ? n62825 : ~n32;
  assign n62827 = pi18 ? n32 : n62826;
  assign n62828 = pi17 ? n48271 : ~n62827;
  assign n62829 = pi16 ? n32 : n62828;
  assign n62830 = pi15 ? n48465 : n62829;
  assign n62831 = pi17 ? n1219 : ~n12287;
  assign n62832 = pi16 ? n16396 : ~n62831;
  assign n62833 = pi15 ? n62832 : n48588;
  assign n62834 = pi14 ? n62830 : n62833;
  assign n62835 = pi13 ? n62834 : n48487;
  assign n62836 = pi18 ? n366 : ~n6071;
  assign n62837 = pi17 ? n32 : n62836;
  assign n62838 = pi19 ? n34907 : ~n32;
  assign n62839 = pi18 ? n62838 : ~n21030;
  assign n62840 = pi17 ? n34906 : n62839;
  assign n62841 = pi16 ? n62837 : ~n62840;
  assign n62842 = pi15 ? n20836 : n62841;
  assign n62843 = pi14 ? n34903 : n62842;
  assign n62844 = pi20 ? n314 : ~n3843;
  assign n62845 = pi19 ? n32 : ~n62844;
  assign n62846 = pi18 ? n127 : n62845;
  assign n62847 = pi17 ? n32 : n62846;
  assign n62848 = pi20 ? n3843 : ~n18415;
  assign n62849 = pi20 ? n9488 : n18073;
  assign n62850 = pi19 ? n62848 : n62849;
  assign n62851 = pi19 ? n9641 : n47025;
  assign n62852 = pi18 ? n62850 : n62851;
  assign n62853 = pi20 ? n3843 : n175;
  assign n62854 = pi19 ? n62853 : ~n617;
  assign n62855 = pi18 ? n62854 : n21548;
  assign n62856 = pi17 ? n62852 : n62855;
  assign n62857 = pi16 ? n62847 : n62856;
  assign n62858 = pi15 ? n62857 : n13948;
  assign n62859 = pi15 ? n20486 : n130;
  assign n62860 = pi14 ? n62858 : n62859;
  assign n62861 = pi13 ? n62843 : n62860;
  assign n62862 = pi12 ? n62835 : n62861;
  assign n62863 = pi11 ? n62823 : n62862;
  assign n62864 = pi10 ? n62804 : n62863;
  assign n62865 = pi09 ? n62747 : n62864;
  assign n62866 = pi19 ? n32 : n49001;
  assign n62867 = pi18 ? n32 : n62866;
  assign n62868 = pi17 ? n62749 : ~n62867;
  assign n62869 = pi16 ? n32 : n62868;
  assign n62870 = pi15 ? n62869 : n62757;
  assign n62871 = pi19 ? n5748 : ~n29457;
  assign n62872 = pi18 ? n32 : n62871;
  assign n62873 = pi17 ? n62872 : ~n62761;
  assign n62874 = pi16 ? n32 : n62873;
  assign n62875 = pi18 ? n5657 : n62766;
  assign n62876 = pi17 ? n32 : n62875;
  assign n62877 = pi16 ? n32 : n62876;
  assign n62878 = pi15 ? n62874 : n62877;
  assign n62879 = pi14 ? n62870 : n62878;
  assign n62880 = pi13 ? n62879 : n23327;
  assign n62881 = pi19 ? n1740 : ~n1941;
  assign n62882 = pi18 ? n32 : n62881;
  assign n62883 = pi17 ? n32 : n62882;
  assign n62884 = pi16 ? n32 : n62883;
  assign n62885 = pi15 ? n32 : n62884;
  assign n62886 = pi14 ? n16110 : n62885;
  assign n62887 = pi15 ? n37592 : n48535;
  assign n62888 = pi14 ? n62887 : n15655;
  assign n62889 = pi13 ? n62886 : n62888;
  assign n62890 = pi12 ? n62880 : n62889;
  assign n62891 = pi19 ? n6018 : ~n236;
  assign n62892 = pi18 ? n32 : n62891;
  assign n62893 = pi17 ? n32 : n62892;
  assign n62894 = pi16 ? n32 : n62893;
  assign n62895 = pi15 ? n34950 : n62894;
  assign n62896 = pi15 ? n34616 : n48548;
  assign n62897 = pi14 ? n62895 : n62896;
  assign n62898 = pi13 ? n62897 : n62791;
  assign n62899 = pi15 ? n24274 : n32;
  assign n62900 = pi20 ? n357 : n9194;
  assign n62901 = pi19 ? n32 : n62900;
  assign n62902 = pi20 ? n9194 : ~n32;
  assign n62903 = pi19 ? n41328 : n62902;
  assign n62904 = pi18 ? n62901 : n62903;
  assign n62905 = pi20 ? n18261 : n428;
  assign n62906 = pi19 ? n59860 : ~n62905;
  assign n62907 = pi18 ? n62906 : ~n2622;
  assign n62908 = pi17 ? n62904 : n62907;
  assign n62909 = pi16 ? n32 : n62908;
  assign n62910 = pi15 ? n22437 : n62909;
  assign n62911 = pi14 ? n62899 : n62910;
  assign n62912 = pi13 ? n15128 : n62911;
  assign n62913 = pi12 ? n62898 : n62912;
  assign n62914 = pi11 ? n62890 : n62913;
  assign n62915 = pi17 ? n1219 : ~n2623;
  assign n62916 = pi16 ? n32 : n62915;
  assign n62917 = pi18 ? n20615 : n2622;
  assign n62918 = pi17 ? n1219 : ~n62917;
  assign n62919 = pi16 ? n32 : n62918;
  assign n62920 = pi15 ? n62916 : n62919;
  assign n62921 = pi14 ? n62920 : n62810;
  assign n62922 = pi16 ? n1135 : ~n2860;
  assign n62923 = pi18 ? n880 : ~n702;
  assign n62924 = pi17 ? n32 : n62923;
  assign n62925 = pi16 ? n890 : n62924;
  assign n62926 = pi15 ? n62925 : n23356;
  assign n62927 = pi14 ? n62922 : n62926;
  assign n62928 = pi13 ? n62921 : n62927;
  assign n62929 = pi15 ? n23457 : n23369;
  assign n62930 = pi14 ? n62929 : n32;
  assign n62931 = pi18 ? n12811 : n384;
  assign n62932 = pi17 ? n1978 : n62931;
  assign n62933 = pi16 ? n32 : n62932;
  assign n62934 = pi15 ? n62933 : n48577;
  assign n62935 = pi14 ? n33672 : n62934;
  assign n62936 = pi13 ? n62930 : n62935;
  assign n62937 = pi12 ? n62928 : n62936;
  assign n62938 = pi18 ? n496 : ~n1166;
  assign n62939 = pi17 ? n16802 : n62938;
  assign n62940 = pi16 ? n32 : n62939;
  assign n62941 = pi17 ? n48271 : ~n2512;
  assign n62942 = pi16 ? n32 : n62941;
  assign n62943 = pi15 ? n62940 : n62942;
  assign n62944 = pi14 ? n62943 : n62833;
  assign n62945 = pi17 ? n48479 : n2519;
  assign n62946 = pi16 ? n16605 : ~n62945;
  assign n62947 = pi18 ? n22705 : ~n323;
  assign n62948 = pi17 ? n48596 : n62947;
  assign n62949 = pi16 ? n32 : n62948;
  assign n62950 = pi15 ? n62946 : n62949;
  assign n62951 = pi14 ? n48594 : n62950;
  assign n62952 = pi13 ? n62944 : n62951;
  assign n62953 = pi16 ? n129 : n21550;
  assign n62954 = pi15 ? n62953 : n13948;
  assign n62955 = pi14 ? n62954 : n32;
  assign n62956 = pi13 ? n62843 : n62955;
  assign n62957 = pi12 ? n62952 : n62956;
  assign n62958 = pi11 ? n62937 : n62957;
  assign n62959 = pi10 ? n62914 : n62958;
  assign n62960 = pi09 ? n62747 : n62959;
  assign n62961 = pi08 ? n62865 : n62960;
  assign n62962 = pi07 ? n62733 : n62961;
  assign n62963 = pi06 ? n62486 : n62962;
  assign n62964 = pi20 ? n17652 : n339;
  assign n62965 = pi19 ? n62964 : ~n32;
  assign n62966 = pi18 ? n32 : n62965;
  assign n62967 = pi17 ? n62966 : ~n2724;
  assign n62968 = pi16 ? n32 : n62967;
  assign n62969 = pi15 ? n32 : n62968;
  assign n62970 = pi17 ? n1470 : ~n2736;
  assign n62971 = pi16 ? n32 : n62970;
  assign n62972 = pi14 ? n62969 : n62971;
  assign n62973 = pi13 ? n32 : n62972;
  assign n62974 = pi12 ? n32 : n62973;
  assign n62975 = pi11 ? n32 : n62974;
  assign n62976 = pi10 ? n32 : n62975;
  assign n62977 = pi19 ? n3692 : n813;
  assign n62978 = pi18 ? n32 : n62977;
  assign n62979 = pi17 ? n2519 : ~n62978;
  assign n62980 = pi16 ? n32 : n62979;
  assign n62981 = pi17 ? n3100 : ~n2736;
  assign n62982 = pi16 ? n32 : n62981;
  assign n62983 = pi15 ? n62980 : n62982;
  assign n62984 = pi17 ? n1219 : ~n2736;
  assign n62985 = pi16 ? n32 : n62984;
  assign n62986 = pi15 ? n62985 : n32;
  assign n62987 = pi14 ? n62983 : n62986;
  assign n62988 = pi14 ? n16110 : n23421;
  assign n62989 = pi13 ? n62987 : n62988;
  assign n62990 = pi15 ? n23443 : n24179;
  assign n62991 = pi14 ? n16110 : n62990;
  assign n62992 = pi19 ? n343 : n53;
  assign n62993 = pi18 ? n32 : n62992;
  assign n62994 = pi17 ? n32 : n62993;
  assign n62995 = pi16 ? n32 : n62994;
  assign n62996 = pi19 ? n5694 : ~n236;
  assign n62997 = pi18 ? n32 : n62996;
  assign n62998 = pi17 ? n32 : n62997;
  assign n62999 = pi16 ? n32 : n62998;
  assign n63000 = pi15 ? n62995 : n62999;
  assign n63001 = pi15 ? n22923 : n35023;
  assign n63002 = pi14 ? n63000 : n63001;
  assign n63003 = pi13 ? n62991 : n63002;
  assign n63004 = pi12 ? n62989 : n63003;
  assign n63005 = pi14 ? n21558 : n23484;
  assign n63006 = pi13 ? n48675 : n63005;
  assign n63007 = pi14 ? n22925 : n23582;
  assign n63008 = pi15 ? n15518 : n1109;
  assign n63009 = pi17 ? n1500 : ~n2750;
  assign n63010 = pi16 ? n32 : n63009;
  assign n63011 = pi15 ? n35049 : n63010;
  assign n63012 = pi14 ? n63008 : n63011;
  assign n63013 = pi13 ? n63007 : n63012;
  assign n63014 = pi12 ? n63006 : n63013;
  assign n63015 = pi11 ? n63004 : n63014;
  assign n63016 = pi18 ? n20193 : ~n14153;
  assign n63017 = pi17 ? n63016 : ~n2623;
  assign n63018 = pi16 ? n32 : n63017;
  assign n63019 = pi18 ? n20193 : n33312;
  assign n63020 = pi18 ? n5158 : n2622;
  assign n63021 = pi17 ? n63019 : ~n63020;
  assign n63022 = pi16 ? n32 : n63021;
  assign n63023 = pi15 ? n63018 : n63022;
  assign n63024 = pi16 ? n1471 : ~n2860;
  assign n63025 = pi16 ? n59546 : ~n2860;
  assign n63026 = pi15 ? n63024 : n63025;
  assign n63027 = pi14 ? n63023 : n63026;
  assign n63028 = pi16 ? n19652 : ~n62666;
  assign n63029 = pi19 ? n18865 : ~n32;
  assign n63030 = pi18 ? n32 : n63029;
  assign n63031 = pi17 ? n32 : n63030;
  assign n63032 = pi16 ? n1808 : ~n63031;
  assign n63033 = pi15 ? n63028 : n63032;
  assign n63034 = pi19 ? n18502 : ~n247;
  assign n63035 = pi18 ? n209 : n63034;
  assign n63036 = pi17 ? n32 : n63035;
  assign n63037 = pi17 ? n18482 : n47296;
  assign n63038 = pi16 ? n63036 : n63037;
  assign n63039 = pi18 ? n940 : n23514;
  assign n63040 = pi17 ? n32 : n63039;
  assign n63041 = pi16 ? n32 : n63040;
  assign n63042 = pi15 ? n63038 : n63041;
  assign n63043 = pi14 ? n63033 : n63042;
  assign n63044 = pi13 ? n63027 : n63043;
  assign n63045 = pi15 ? n21928 : n14973;
  assign n63046 = pi20 ? n246 : ~n287;
  assign n63047 = pi19 ? n63046 : n32;
  assign n63048 = pi18 ? n4983 : ~n63047;
  assign n63049 = pi17 ? n8859 : ~n63048;
  assign n63050 = pi16 ? n32 : n63049;
  assign n63051 = pi15 ? n63050 : n48719;
  assign n63052 = pi14 ? n63045 : n63051;
  assign n63053 = pi13 ? n23530 : n63052;
  assign n63054 = pi12 ? n63044 : n63053;
  assign n63055 = pi19 ? n55229 : ~n32;
  assign n63056 = pi18 ? n880 : ~n63055;
  assign n63057 = pi17 ? n17346 : n63056;
  assign n63058 = pi16 ? n32 : n63057;
  assign n63059 = pi18 ? n20164 : n2627;
  assign n63060 = pi17 ? n48726 : ~n63059;
  assign n63061 = pi16 ? n32 : n63060;
  assign n63062 = pi15 ? n63058 : n63061;
  assign n63063 = pi20 ? n339 : ~n1319;
  assign n63064 = pi19 ? n63063 : n32;
  assign n63065 = pi18 ? n48732 : n63064;
  assign n63066 = pi17 ? n48731 : ~n63065;
  assign n63067 = pi16 ? n3165 : ~n63066;
  assign n63068 = pi15 ? n63067 : n48814;
  assign n63069 = pi14 ? n63062 : n63068;
  assign n63070 = pi13 ? n63069 : n48755;
  assign n63071 = pi18 ? n366 : ~n19082;
  assign n63072 = pi17 ? n32 : n63071;
  assign n63073 = pi17 ? n35156 : ~n14395;
  assign n63074 = pi16 ? n63072 : ~n63073;
  assign n63075 = pi15 ? n14156 : n63074;
  assign n63076 = pi14 ? n32 : n63075;
  assign n63077 = pi15 ? n21551 : n13948;
  assign n63078 = pi19 ? n22652 : n28191;
  assign n63079 = pi18 ? n30779 : n63078;
  assign n63080 = pi19 ? n28134 : ~n349;
  assign n63081 = pi18 ? n63080 : n32;
  assign n63082 = pi17 ? n63079 : ~n63081;
  assign n63083 = pi16 ? n19652 : ~n63082;
  assign n63084 = pi15 ? n130 : n63083;
  assign n63085 = pi14 ? n63077 : n63084;
  assign n63086 = pi13 ? n63076 : n63085;
  assign n63087 = pi12 ? n63070 : n63086;
  assign n63088 = pi11 ? n63054 : n63087;
  assign n63089 = pi10 ? n63015 : n63088;
  assign n63090 = pi09 ? n62976 : n63089;
  assign n63091 = pi14 ? n16110 : n23570;
  assign n63092 = pi13 ? n62987 : n63091;
  assign n63093 = pi15 ? n23443 : n35701;
  assign n63094 = pi14 ? n35174 : n63093;
  assign n63095 = pi19 ? n343 : n5614;
  assign n63096 = pi18 ? n32 : n63095;
  assign n63097 = pi17 ? n32 : n63096;
  assign n63098 = pi16 ? n32 : n63097;
  assign n63099 = pi15 ? n63098 : n23999;
  assign n63100 = pi15 ? n32 : n35023;
  assign n63101 = pi14 ? n63099 : n63100;
  assign n63102 = pi13 ? n63094 : n63101;
  assign n63103 = pi12 ? n63092 : n63102;
  assign n63104 = pi18 ? n48660 : n48864;
  assign n63105 = pi17 ? n32 : n63104;
  assign n63106 = pi16 ? n32 : n63105;
  assign n63107 = pi15 ? n35393 : n63106;
  assign n63108 = pi14 ? n63107 : n48792;
  assign n63109 = pi13 ? n63108 : n63005;
  assign n63110 = pi17 ? n1500 : ~n2855;
  assign n63111 = pi16 ? n32 : n63110;
  assign n63112 = pi15 ? n35049 : n63111;
  assign n63113 = pi14 ? n23085 : n63112;
  assign n63114 = pi13 ? n23086 : n63113;
  assign n63115 = pi12 ? n63109 : n63114;
  assign n63116 = pi11 ? n63103 : n63115;
  assign n63117 = pi17 ? n63016 : ~n2855;
  assign n63118 = pi16 ? n32 : n63117;
  assign n63119 = pi18 ? n5158 : n1750;
  assign n63120 = pi17 ? n63019 : ~n63119;
  assign n63121 = pi16 ? n32 : n63120;
  assign n63122 = pi15 ? n63118 : n63121;
  assign n63123 = pi16 ? n1471 : ~n2856;
  assign n63124 = pi16 ? n59546 : ~n2624;
  assign n63125 = pi15 ? n63123 : n63124;
  assign n63126 = pi14 ? n63122 : n63125;
  assign n63127 = pi16 ? n1214 : ~n2624;
  assign n63128 = pi16 ? n1808 : ~n35573;
  assign n63129 = pi15 ? n63127 : n63128;
  assign n63130 = pi17 ? n18482 : n13026;
  assign n63131 = pi16 ? n63036 : n63130;
  assign n63132 = pi15 ? n63131 : n63041;
  assign n63133 = pi14 ? n63129 : n63132;
  assign n63134 = pi13 ? n63126 : n63133;
  assign n63135 = pi14 ? n23529 : n22205;
  assign n63136 = pi14 ? n14974 : n63051;
  assign n63137 = pi13 ? n63135 : n63136;
  assign n63138 = pi12 ? n63134 : n63137;
  assign n63139 = pi17 ? n48751 : ~n2755;
  assign n63140 = pi16 ? n17434 : n63139;
  assign n63141 = pi18 ? n14153 : n2754;
  assign n63142 = pi17 ? n2519 : ~n63141;
  assign n63143 = pi16 ? n32 : n63142;
  assign n63144 = pi15 ? n63140 : n63143;
  assign n63145 = pi14 ? n48748 : n63144;
  assign n63146 = pi13 ? n63069 : n63145;
  assign n63147 = pi12 ? n63146 : n63086;
  assign n63148 = pi11 ? n63138 : n63147;
  assign n63149 = pi10 ? n63116 : n63148;
  assign n63150 = pi09 ? n62976 : n63149;
  assign n63151 = pi08 ? n63090 : n63150;
  assign n63152 = pi17 ? n1470 : ~n4245;
  assign n63153 = pi16 ? n32 : n63152;
  assign n63154 = pi15 ? n32 : n63153;
  assign n63155 = pi17 ? n1470 : ~n2724;
  assign n63156 = pi16 ? n32 : n63155;
  assign n63157 = pi14 ? n63154 : n63156;
  assign n63158 = pi13 ? n32 : n63157;
  assign n63159 = pi12 ? n32 : n63158;
  assign n63160 = pi11 ? n32 : n63159;
  assign n63161 = pi10 ? n32 : n63160;
  assign n63162 = pi20 ? n60202 : ~n32;
  assign n63163 = pi19 ? n3692 : n63162;
  assign n63164 = pi18 ? n32 : n63163;
  assign n63165 = pi17 ? n2519 : ~n63164;
  assign n63166 = pi16 ? n32 : n63165;
  assign n63167 = pi18 ? n6145 : n237;
  assign n63168 = pi17 ? n63167 : ~n2724;
  assign n63169 = pi16 ? n32 : n63168;
  assign n63170 = pi15 ? n63166 : n63169;
  assign n63171 = pi17 ? n2355 : ~n2731;
  assign n63172 = pi16 ? n32 : n63171;
  assign n63173 = pi15 ? n63172 : n32;
  assign n63174 = pi14 ? n63170 : n63173;
  assign n63175 = pi14 ? n35174 : n23623;
  assign n63176 = pi13 ? n63174 : n63175;
  assign n63177 = pi14 ? n23576 : n63093;
  assign n63178 = pi15 ? n63098 : n54357;
  assign n63179 = pi15 ? n23484 : n14570;
  assign n63180 = pi14 ? n63178 : n63179;
  assign n63181 = pi13 ? n63177 : n63180;
  assign n63182 = pi12 ? n63176 : n63181;
  assign n63183 = pi14 ? n23421 : n16110;
  assign n63184 = pi13 ? n48873 : n63183;
  assign n63185 = pi15 ? n32 : n25888;
  assign n63186 = pi14 ? n32 : n63185;
  assign n63187 = pi19 ? n18571 : ~n35248;
  assign n63188 = pi20 ? n19731 : ~n2180;
  assign n63189 = pi19 ? n63188 : ~n18173;
  assign n63190 = pi18 ? n63187 : n63189;
  assign n63191 = pi20 ? n1331 : n1076;
  assign n63192 = pi20 ? n428 : n357;
  assign n63193 = pi19 ? n63191 : n63192;
  assign n63194 = pi18 ? n63193 : n1750;
  assign n63195 = pi17 ? n63190 : n63194;
  assign n63196 = pi16 ? n59450 : ~n63195;
  assign n63197 = pi15 ? n63196 : n63111;
  assign n63198 = pi14 ? n38992 : n63197;
  assign n63199 = pi13 ? n63186 : n63198;
  assign n63200 = pi12 ? n63184 : n63199;
  assign n63201 = pi11 ? n63182 : n63200;
  assign n63202 = pi19 ? n4721 : n4670;
  assign n63203 = pi18 ? n20193 : ~n63202;
  assign n63204 = pi17 ? n63203 : ~n2750;
  assign n63205 = pi16 ? n32 : n63204;
  assign n63206 = pi18 ? n20020 : n1750;
  assign n63207 = pi17 ? n5766 : ~n63206;
  assign n63208 = pi16 ? n32 : n63207;
  assign n63209 = pi15 ? n63205 : n63208;
  assign n63210 = pi16 ? n2326 : ~n2856;
  assign n63211 = pi16 ? n1808 : ~n2856;
  assign n63212 = pi15 ? n63210 : n63211;
  assign n63213 = pi14 ? n63209 : n63212;
  assign n63214 = pi17 ? n32 : n3812;
  assign n63215 = pi16 ? n1581 : ~n63214;
  assign n63216 = pi15 ? n63215 : n63211;
  assign n63217 = pi19 ? n321 : ~n5688;
  assign n63218 = pi18 ? n63217 : n2622;
  assign n63219 = pi17 ? n32 : ~n63218;
  assign n63220 = pi16 ? n32 : n63219;
  assign n63221 = pi15 ? n13025 : n63220;
  assign n63222 = pi14 ? n63216 : n63221;
  assign n63223 = pi13 ? n63213 : n63222;
  assign n63224 = pi14 ? n23674 : n22252;
  assign n63225 = pi15 ? n15123 : n21928;
  assign n63226 = pi18 ? n48912 : n976;
  assign n63227 = pi17 ? n8859 : ~n63226;
  assign n63228 = pi16 ? n32 : n63227;
  assign n63229 = pi15 ? n48911 : n63228;
  assign n63230 = pi14 ? n63225 : n63229;
  assign n63231 = pi13 ? n63224 : n63230;
  assign n63232 = pi12 ? n63223 : n63231;
  assign n63233 = pi18 ? n880 : ~n1326;
  assign n63234 = pi17 ? n23052 : n63233;
  assign n63235 = pi16 ? n32 : n63234;
  assign n63236 = pi15 ? n63235 : n63061;
  assign n63237 = pi18 ? n48732 : ~n2747;
  assign n63238 = pi17 ? n48731 : ~n63237;
  assign n63239 = pi16 ? n3165 : ~n63238;
  assign n63240 = pi15 ? n63239 : n48931;
  assign n63241 = pi14 ? n63236 : n63240;
  assign n63242 = pi16 ? n32 : n48951;
  assign n63243 = pi15 ? n48949 : n63242;
  assign n63244 = pi14 ? n48940 : n63243;
  assign n63245 = pi13 ? n63241 : n63244;
  assign n63246 = pi15 ? n466 : n21464;
  assign n63247 = pi18 ? n35348 : ~n21798;
  assign n63248 = pi17 ? n35347 : n63247;
  assign n63249 = pi16 ? n1135 : ~n63248;
  assign n63250 = pi17 ? n35354 : ~n14395;
  assign n63251 = pi16 ? n1233 : ~n63250;
  assign n63252 = pi15 ? n63249 : n63251;
  assign n63253 = pi14 ? n63246 : n63252;
  assign n63254 = pi15 ? n21551 : n20660;
  assign n63255 = pi18 ? n17391 : n32;
  assign n63256 = pi17 ? n32 : n63255;
  assign n63257 = pi16 ? n63256 : n13951;
  assign n63258 = pi17 ? n23711 : n1682;
  assign n63259 = pi16 ? n1233 : ~n63258;
  assign n63260 = pi15 ? n63257 : n63259;
  assign n63261 = pi14 ? n63254 : n63260;
  assign n63262 = pi13 ? n63253 : n63261;
  assign n63263 = pi12 ? n63245 : n63262;
  assign n63264 = pi11 ? n63232 : n63263;
  assign n63265 = pi10 ? n63201 : n63264;
  assign n63266 = pi09 ? n63161 : n63265;
  assign n63267 = pi19 ? n3692 : n1812;
  assign n63268 = pi18 ? n32 : n63267;
  assign n63269 = pi17 ? n2519 : ~n63268;
  assign n63270 = pi16 ? n32 : n63269;
  assign n63271 = pi15 ? n63270 : n63169;
  assign n63272 = pi17 ? n2355 : ~n2736;
  assign n63273 = pi16 ? n32 : n63272;
  assign n63274 = pi15 ? n63273 : n32;
  assign n63275 = pi14 ? n63271 : n63274;
  assign n63276 = pi14 ? n23576 : n23726;
  assign n63277 = pi13 ? n63275 : n63276;
  assign n63278 = pi15 ? n23443 : n14339;
  assign n63279 = pi14 ? n23794 : n63278;
  assign n63280 = pi19 ? n343 : n7488;
  assign n63281 = pi18 ? n32 : n63280;
  assign n63282 = pi17 ? n32 : n63281;
  assign n63283 = pi16 ? n32 : n63282;
  assign n63284 = pi15 ? n63283 : n23802;
  assign n63285 = pi14 ? n63284 : n63179;
  assign n63286 = pi13 ? n63279 : n63285;
  assign n63287 = pi12 ? n63277 : n63286;
  assign n63288 = pi19 ? n6173 : ~n813;
  assign n63289 = pi18 ? n48863 : n63288;
  assign n63290 = pi17 ? n32 : n63289;
  assign n63291 = pi16 ? n32 : n63290;
  assign n63292 = pi15 ? n48997 : n63291;
  assign n63293 = pi14 ? n63292 : n49006;
  assign n63294 = pi15 ? n15836 : n16108;
  assign n63295 = pi14 ? n63294 : n16110;
  assign n63296 = pi13 ? n63293 : n63295;
  assign n63297 = pi15 ? n32 : n25932;
  assign n63298 = pi14 ? n23252 : n63297;
  assign n63299 = pi15 ? n23749 : n32;
  assign n63300 = pi19 ? n18778 : ~n19426;
  assign n63301 = pi20 ? n18129 : n448;
  assign n63302 = pi19 ? n63301 : ~n339;
  assign n63303 = pi18 ? n63300 : n63302;
  assign n63304 = pi19 ? n18741 : n4491;
  assign n63305 = pi18 ? n63304 : n2615;
  assign n63306 = pi17 ? n63303 : n63305;
  assign n63307 = pi16 ? n59332 : ~n63306;
  assign n63308 = pi17 ? n1500 : ~n2616;
  assign n63309 = pi16 ? n32 : n63308;
  assign n63310 = pi15 ? n63307 : n63309;
  assign n63311 = pi14 ? n63299 : n63310;
  assign n63312 = pi13 ? n63298 : n63311;
  assign n63313 = pi12 ? n63296 : n63312;
  assign n63314 = pi11 ? n63287 : n63313;
  assign n63315 = pi17 ? n63203 : ~n8885;
  assign n63316 = pi16 ? n32 : n63315;
  assign n63317 = pi18 ? n20020 : n2615;
  assign n63318 = pi17 ? n5766 : ~n63317;
  assign n63319 = pi16 ? n32 : n63318;
  assign n63320 = pi15 ? n63316 : n63319;
  assign n63321 = pi14 ? n63320 : n63212;
  assign n63322 = pi16 ? n465 : n63219;
  assign n63323 = pi15 ? n13025 : n63322;
  assign n63324 = pi14 ? n63216 : n63323;
  assign n63325 = pi13 ? n63321 : n63324;
  assign n63326 = pi21 ? n206 : n9326;
  assign n63327 = pi20 ? n8943 : ~n63326;
  assign n63328 = pi19 ? n63327 : n32;
  assign n63329 = pi18 ? n32 : n63328;
  assign n63330 = pi17 ? n32 : n63329;
  assign n63331 = pi16 ? n32 : n63330;
  assign n63332 = pi15 ? n63331 : n32;
  assign n63333 = pi14 ? n63332 : n22348;
  assign n63334 = pi15 ? n22347 : n21928;
  assign n63335 = pi14 ? n63334 : n63229;
  assign n63336 = pi13 ? n63333 : n63335;
  assign n63337 = pi12 ? n63325 : n63336;
  assign n63338 = pi18 ? n880 : ~n976;
  assign n63339 = pi17 ? n23052 : n63338;
  assign n63340 = pi16 ? n32 : n63339;
  assign n63341 = pi15 ? n63340 : n63061;
  assign n63342 = pi14 ? n63341 : n63240;
  assign n63343 = pi18 ? n20020 : n520;
  assign n63344 = pi17 ? n19886 : n63343;
  assign n63345 = pi16 ? n1214 : ~n63344;
  assign n63346 = pi15 ? n48936 : n63345;
  assign n63347 = pi18 ? n5502 : n520;
  assign n63348 = pi17 ? n49033 : ~n63347;
  assign n63349 = pi16 ? n32 : n63348;
  assign n63350 = pi15 ? n63349 : n63242;
  assign n63351 = pi14 ? n63346 : n63350;
  assign n63352 = pi13 ? n63342 : n63351;
  assign n63353 = pi16 ? n1233 : ~n63248;
  assign n63354 = pi17 ? n35354 : ~n22085;
  assign n63355 = pi16 ? n1233 : ~n63354;
  assign n63356 = pi15 ? n63353 : n63355;
  assign n63357 = pi14 ? n63246 : n63356;
  assign n63358 = pi18 ? n56696 : n32;
  assign n63359 = pi17 ? n32 : n63358;
  assign n63360 = pi16 ? n63359 : n13951;
  assign n63361 = pi18 ? n32 : ~n7221;
  assign n63362 = pi17 ? n23711 : n63361;
  assign n63363 = pi16 ? n1233 : ~n63362;
  assign n63364 = pi15 ? n63360 : n63363;
  assign n63365 = pi14 ? n63254 : n63364;
  assign n63366 = pi13 ? n63357 : n63365;
  assign n63367 = pi12 ? n63352 : n63366;
  assign n63368 = pi11 ? n63337 : n63367;
  assign n63369 = pi10 ? n63314 : n63368;
  assign n63370 = pi09 ? n63161 : n63369;
  assign n63371 = pi08 ? n63266 : n63370;
  assign n63372 = pi07 ? n63151 : n63371;
  assign n63373 = pi15 ? n32 : n6591;
  assign n63374 = pi17 ? n1704 : ~n2724;
  assign n63375 = pi16 ? n32 : n63374;
  assign n63376 = pi15 ? n63375 : n62971;
  assign n63377 = pi14 ? n63373 : n63376;
  assign n63378 = pi13 ? n32 : n63377;
  assign n63379 = pi12 ? n32 : n63378;
  assign n63380 = pi11 ? n32 : n63379;
  assign n63381 = pi10 ? n32 : n63380;
  assign n63382 = pi17 ? n4685 : ~n2724;
  assign n63383 = pi16 ? n32 : n63382;
  assign n63384 = pi15 ? n6591 : n63383;
  assign n63385 = pi14 ? n63384 : n32;
  assign n63386 = pi14 ? n23794 : n23726;
  assign n63387 = pi13 ? n63385 : n63386;
  assign n63388 = pi19 ? n531 : n7488;
  assign n63389 = pi18 ? n32 : n63388;
  assign n63390 = pi17 ? n32 : n63389;
  assign n63391 = pi16 ? n32 : n63390;
  assign n63392 = pi15 ? n49078 : n63391;
  assign n63393 = pi14 ? n23794 : n63392;
  assign n63394 = pi19 ? n531 : ~n20022;
  assign n63395 = pi18 ? n32 : n63394;
  assign n63396 = pi17 ? n32 : n63395;
  assign n63397 = pi16 ? n32 : n63396;
  assign n63398 = pi15 ? n63397 : n24256;
  assign n63399 = pi14 ? n63398 : n49086;
  assign n63400 = pi13 ? n63393 : n63399;
  assign n63401 = pi12 ? n63387 : n63400;
  assign n63402 = pi13 ? n49105 : n48618;
  assign n63403 = pi15 ? n23741 : n23340;
  assign n63404 = pi16 ? n3068 : ~n2617;
  assign n63405 = pi19 ? n32 : ~n176;
  assign n63406 = pi18 ? n32 : n63405;
  assign n63407 = pi17 ? n32 : n63406;
  assign n63408 = pi17 ? n32 : n8885;
  assign n63409 = pi16 ? n63407 : ~n63408;
  assign n63410 = pi15 ? n63404 : n63409;
  assign n63411 = pi14 ? n63403 : n63410;
  assign n63412 = pi13 ? n23627 : n63411;
  assign n63413 = pi12 ? n63402 : n63412;
  assign n63414 = pi11 ? n63401 : n63413;
  assign n63415 = pi16 ? n44190 : ~n63408;
  assign n63416 = pi19 ? n507 : n7089;
  assign n63417 = pi18 ? n63416 : ~n13945;
  assign n63418 = pi18 ? n1541 : n2615;
  assign n63419 = pi17 ? n63417 : ~n63418;
  assign n63420 = pi16 ? n32 : n63419;
  assign n63421 = pi15 ? n63415 : n63420;
  assign n63422 = pi16 ? n2860 : ~n2617;
  assign n63423 = pi14 ? n63421 : n63422;
  assign n63424 = pi18 ? n863 : n423;
  assign n63425 = pi17 ? n32 : n63424;
  assign n63426 = pi16 ? n63425 : ~n2617;
  assign n63427 = pi17 ? n10723 : n48108;
  assign n63428 = pi16 ? n32 : n63427;
  assign n63429 = pi15 ? n63426 : n63428;
  assign n63430 = pi16 ? n18325 : n23850;
  assign n63431 = pi15 ? n23847 : n63430;
  assign n63432 = pi14 ? n63429 : n63431;
  assign n63433 = pi13 ? n63423 : n63432;
  assign n63434 = pi14 ? n32 : n23179;
  assign n63435 = pi17 ? n48315 : n35666;
  assign n63436 = pi16 ? n32 : n63435;
  assign n63437 = pi15 ? n15123 : n63436;
  assign n63438 = pi18 ? n6384 : n47144;
  assign n63439 = pi17 ? n2959 : ~n63438;
  assign n63440 = pi16 ? n32 : n63439;
  assign n63441 = pi21 ? n32 : ~n7478;
  assign n63442 = pi20 ? n32 : ~n63441;
  assign n63443 = pi19 ? n63442 : ~n32;
  assign n63444 = pi18 ? n49140 : n63443;
  assign n63445 = pi17 ? n32 : ~n63444;
  assign n63446 = pi16 ? n32 : n63445;
  assign n63447 = pi15 ? n63440 : n63446;
  assign n63448 = pi14 ? n63437 : n63447;
  assign n63449 = pi13 ? n63434 : n63448;
  assign n63450 = pi12 ? n63433 : n63449;
  assign n63451 = pi18 ? n237 : n1326;
  assign n63452 = pi17 ? n32 : ~n63451;
  assign n63453 = pi16 ? n32 : n63452;
  assign n63454 = pi18 ? n6163 : n2627;
  assign n63455 = pi17 ? n3164 : ~n63454;
  assign n63456 = pi16 ? n32 : n63455;
  assign n63457 = pi15 ? n63453 : n63456;
  assign n63458 = pi15 ? n49349 : n49157;
  assign n63459 = pi14 ? n63457 : n63458;
  assign n63460 = pi15 ? n49171 : n32;
  assign n63461 = pi14 ? n49167 : n63460;
  assign n63462 = pi13 ? n63459 : n63461;
  assign n63463 = pi16 ? n49181 : n21542;
  assign n63464 = pi15 ? n63463 : n21543;
  assign n63465 = pi18 ? n35581 : n21692;
  assign n63466 = pi17 ? n35580 : ~n63465;
  assign n63467 = pi16 ? n1233 : ~n63466;
  assign n63468 = pi18 ? n5694 : n14153;
  assign n63469 = pi17 ? n35586 : ~n63468;
  assign n63470 = pi16 ? n1233 : ~n63469;
  assign n63471 = pi15 ? n63467 : n63470;
  assign n63472 = pi14 ? n63464 : n63471;
  assign n63473 = pi15 ? n21033 : n32;
  assign n63474 = pi21 ? n1009 : ~n174;
  assign n63475 = pi20 ? n32 : n63474;
  assign n63476 = pi19 ? n32 : n63475;
  assign n63477 = pi19 ? n236 : ~n23644;
  assign n63478 = pi18 ? n63476 : ~n63477;
  assign n63479 = pi17 ? n32 : n63478;
  assign n63480 = pi19 ? n4670 : n45905;
  assign n63481 = pi18 ? n63480 : n1757;
  assign n63482 = pi18 ? n38787 : n32;
  assign n63483 = pi17 ? n63481 : n63482;
  assign n63484 = pi16 ? n63479 : n63483;
  assign n63485 = pi18 ? n63476 : ~n32;
  assign n63486 = pi17 ? n32 : n63485;
  assign n63487 = pi16 ? n63486 : ~n35611;
  assign n63488 = pi15 ? n63484 : n63487;
  assign n63489 = pi14 ? n63473 : n63488;
  assign n63490 = pi13 ? n63472 : n63489;
  assign n63491 = pi12 ? n63462 : n63490;
  assign n63492 = pi11 ? n63450 : n63491;
  assign n63493 = pi10 ? n63414 : n63492;
  assign n63494 = pi09 ? n63381 : n63493;
  assign n63495 = pi14 ? n63384 : n23726;
  assign n63496 = pi14 ? n23794 : n23924;
  assign n63497 = pi13 ? n63495 : n63496;
  assign n63498 = pi19 ? n531 : n1757;
  assign n63499 = pi18 ? n32 : n63498;
  assign n63500 = pi17 ? n32 : n63499;
  assign n63501 = pi16 ? n32 : n63500;
  assign n63502 = pi15 ? n49078 : n63501;
  assign n63503 = pi14 ? n16321 : n63502;
  assign n63504 = pi19 ? n531 : ~n502;
  assign n63505 = pi18 ? n32 : n63504;
  assign n63506 = pi17 ? n32 : n63505;
  assign n63507 = pi16 ? n32 : n63506;
  assign n63508 = pi15 ? n63507 : n25331;
  assign n63509 = pi14 ? n63508 : n49217;
  assign n63510 = pi13 ? n63503 : n63509;
  assign n63511 = pi12 ? n63497 : n63510;
  assign n63512 = pi17 ? n34522 : ~n4245;
  assign n63513 = pi16 ? n32 : n63512;
  assign n63514 = pi15 ? n49095 : n63513;
  assign n63515 = pi14 ? n63514 : n49226;
  assign n63516 = pi13 ? n63515 : n48618;
  assign n63517 = pi15 ? n23574 : n25888;
  assign n63518 = pi16 ? n3068 : ~n2745;
  assign n63519 = pi17 ? n32 : n3070;
  assign n63520 = pi16 ? n63407 : ~n63519;
  assign n63521 = pi15 ? n63518 : n63520;
  assign n63522 = pi14 ? n63517 : n63521;
  assign n63523 = pi13 ? n50045 : n63522;
  assign n63524 = pi12 ? n63516 : n63523;
  assign n63525 = pi11 ? n63511 : n63524;
  assign n63526 = pi19 ? n32 : n274;
  assign n63527 = pi18 ? n32 : n63526;
  assign n63528 = pi17 ? n63527 : n3070;
  assign n63529 = pi16 ? n44190 : ~n63528;
  assign n63530 = pi18 ? n1541 : n697;
  assign n63531 = pi17 ? n63417 : ~n63530;
  assign n63532 = pi16 ? n32 : n63531;
  assign n63533 = pi15 ? n63529 : n63532;
  assign n63534 = pi16 ? n2860 : ~n2856;
  assign n63535 = pi14 ? n63533 : n63534;
  assign n63536 = pi18 ? n863 : n532;
  assign n63537 = pi17 ? n32 : n63536;
  assign n63538 = pi16 ? n63537 : ~n2617;
  assign n63539 = pi15 ? n63538 : n63428;
  assign n63540 = pi14 ? n63539 : n63431;
  assign n63541 = pi13 ? n63535 : n63540;
  assign n63542 = pi14 ? n32 : n23264;
  assign n63543 = pi13 ? n63542 : n63448;
  assign n63544 = pi12 ? n63541 : n63543;
  assign n63545 = pi14 ? n63457 : n49158;
  assign n63546 = pi16 ? n49162 : ~n2749;
  assign n63547 = pi16 ? n49165 : ~n2749;
  assign n63548 = pi15 ? n63546 : n63547;
  assign n63549 = pi14 ? n63548 : n63460;
  assign n63550 = pi13 ? n63545 : n63549;
  assign n63551 = pi18 ? n56696 : ~n63477;
  assign n63552 = pi17 ? n32 : n63551;
  assign n63553 = pi18 ? n38787 : n20828;
  assign n63554 = pi17 ? n63481 : n63553;
  assign n63555 = pi16 ? n63552 : n63554;
  assign n63556 = pi20 ? n749 : ~n52;
  assign n63557 = pi19 ? n63556 : ~n32;
  assign n63558 = pi18 ? n16432 : ~n63557;
  assign n63559 = pi17 ? n23912 : ~n63558;
  assign n63560 = pi16 ? n63486 : ~n63559;
  assign n63561 = pi15 ? n63555 : n63560;
  assign n63562 = pi14 ? n63473 : n63561;
  assign n63563 = pi13 ? n63472 : n63562;
  assign n63564 = pi12 ? n63550 : n63563;
  assign n63565 = pi11 ? n63544 : n63564;
  assign n63566 = pi10 ? n63525 : n63565;
  assign n63567 = pi09 ? n63381 : n63566;
  assign n63568 = pi08 ? n63494 : n63567;
  assign n63569 = pi17 ? n1470 : ~n2850;
  assign n63570 = pi16 ? n32 : n63569;
  assign n63571 = pi15 ? n32 : n63570;
  assign n63572 = pi17 ? n2670 : ~n2724;
  assign n63573 = pi16 ? n32 : n63572;
  assign n63574 = pi15 ? n7034 : n63573;
  assign n63575 = pi14 ? n63571 : n63574;
  assign n63576 = pi13 ? n32 : n63575;
  assign n63577 = pi12 ? n32 : n63576;
  assign n63578 = pi11 ? n32 : n63577;
  assign n63579 = pi10 ? n32 : n63578;
  assign n63580 = pi17 ? n1213 : ~n2852;
  assign n63581 = pi16 ? n32 : n63580;
  assign n63582 = pi15 ? n63570 : n63581;
  assign n63583 = pi14 ? n63582 : n23924;
  assign n63584 = pi14 ? n35691 : n23982;
  assign n63585 = pi13 ? n63583 : n63584;
  assign n63586 = pi15 ? n49292 : n63501;
  assign n63587 = pi14 ? n35691 : n63586;
  assign n63588 = pi18 ? n49295 : n35698;
  assign n63589 = pi17 ? n32 : n63588;
  assign n63590 = pi16 ? n32 : n63589;
  assign n63591 = pi15 ? n63590 : n14917;
  assign n63592 = pi14 ? n63591 : n49303;
  assign n63593 = pi13 ? n63587 : n63592;
  assign n63594 = pi12 ? n63585 : n63593;
  assign n63595 = pi17 ? n48166 : ~n3067;
  assign n63596 = pi16 ? n32 : n63595;
  assign n63597 = pi15 ? n49311 : n63596;
  assign n63598 = pi15 ? n23725 : n23574;
  assign n63599 = pi14 ? n63597 : n63598;
  assign n63600 = pi14 ? n23576 : n63598;
  assign n63601 = pi13 ? n63599 : n63600;
  assign n63602 = pi15 ? n16108 : n23484;
  assign n63603 = pi16 ? n2745 : ~n2745;
  assign n63604 = pi15 ? n63518 : n63603;
  assign n63605 = pi14 ? n63602 : n63604;
  assign n63606 = pi13 ? n50045 : n63605;
  assign n63607 = pi12 ? n63601 : n63606;
  assign n63608 = pi11 ? n63594 : n63607;
  assign n63609 = pi16 ? n3068 : ~n63519;
  assign n63610 = pi15 ? n63609 : n63603;
  assign n63611 = pi16 ? n2860 : ~n2745;
  assign n63612 = pi14 ? n63610 : n63611;
  assign n63613 = pi16 ? n3769 : ~n2745;
  assign n63614 = pi18 ? n20172 : n13945;
  assign n63615 = pi17 ? n63614 : n23840;
  assign n63616 = pi16 ? n32 : n63615;
  assign n63617 = pi15 ? n63613 : n63616;
  assign n63618 = pi14 ? n63617 : n24022;
  assign n63619 = pi13 ? n63612 : n63618;
  assign n63620 = pi14 ? n32 : n22817;
  assign n63621 = pi15 ? n32 : n49135;
  assign n63622 = pi18 ? n6669 : n702;
  assign n63623 = pi17 ? n2959 : ~n63622;
  assign n63624 = pi16 ? n32 : n63623;
  assign n63625 = pi19 ? n6355 : ~n32;
  assign n63626 = pi18 ? n49337 : n63625;
  assign n63627 = pi17 ? n32 : ~n63626;
  assign n63628 = pi16 ? n32 : n63627;
  assign n63629 = pi15 ? n63624 : n63628;
  assign n63630 = pi14 ? n63621 : n63629;
  assign n63631 = pi13 ? n63620 : n63630;
  assign n63632 = pi12 ? n63619 : n63631;
  assign n63633 = pi19 ? n56516 : ~n32;
  assign n63634 = pi18 ? n32 : ~n63633;
  assign n63635 = pi17 ? n32 : n63634;
  assign n63636 = pi16 ? n32 : n63635;
  assign n63637 = pi18 ? n6163 : n595;
  assign n63638 = pi17 ? n3164 : ~n63637;
  assign n63639 = pi16 ? n32 : n63638;
  assign n63640 = pi15 ? n63636 : n63639;
  assign n63641 = pi14 ? n63640 : n49349;
  assign n63642 = pi15 ? n49359 : n32;
  assign n63643 = pi14 ? n49355 : n63642;
  assign n63644 = pi13 ? n63641 : n63643;
  assign n63645 = pi16 ? n17850 : n2095;
  assign n63646 = pi15 ? n63645 : n21686;
  assign n63647 = pi18 ? n46739 : n5351;
  assign n63648 = pi17 ? n35797 : ~n63647;
  assign n63649 = pi16 ? n1233 : ~n63648;
  assign n63650 = pi18 ? n35804 : n21798;
  assign n63651 = pi17 ? n35803 : ~n63650;
  assign n63652 = pi16 ? n1233 : ~n63651;
  assign n63653 = pi15 ? n63649 : n63652;
  assign n63654 = pi14 ? n63646 : n63653;
  assign n63655 = pi19 ? n29613 : n18678;
  assign n63656 = pi18 ? n29316 : ~n63655;
  assign n63657 = pi17 ? n32 : n63656;
  assign n63658 = pi19 ? n9007 : n18678;
  assign n63659 = pi18 ? n63658 : ~n24064;
  assign n63660 = pi17 ? n63659 : ~n35821;
  assign n63661 = pi16 ? n63657 : ~n63660;
  assign n63662 = pi16 ? n29318 : ~n35827;
  assign n63663 = pi15 ? n63661 : n63662;
  assign n63664 = pi14 ? n21217 : n63663;
  assign n63665 = pi13 ? n63654 : n63664;
  assign n63666 = pi12 ? n63644 : n63665;
  assign n63667 = pi11 ? n63632 : n63666;
  assign n63668 = pi10 ? n63608 : n63667;
  assign n63669 = pi09 ? n63579 : n63668;
  assign n63670 = pi17 ? n2670 : ~n4245;
  assign n63671 = pi16 ? n32 : n63670;
  assign n63672 = pi15 ? n7034 : n63671;
  assign n63673 = pi14 ? n63571 : n63672;
  assign n63674 = pi13 ? n32 : n63673;
  assign n63675 = pi12 ? n32 : n63674;
  assign n63676 = pi11 ? n32 : n63675;
  assign n63677 = pi10 ? n32 : n63676;
  assign n63678 = pi17 ? n1213 : ~n2736;
  assign n63679 = pi16 ? n32 : n63678;
  assign n63680 = pi15 ? n63570 : n63679;
  assign n63681 = pi14 ? n63680 : n23982;
  assign n63682 = pi13 ? n63681 : n32;
  assign n63683 = pi14 ? n16377 : n63586;
  assign n63684 = pi19 ? n531 : ~n9668;
  assign n63685 = pi18 ? n49295 : n63684;
  assign n63686 = pi17 ? n32 : n63685;
  assign n63687 = pi16 ? n32 : n63686;
  assign n63688 = pi15 ? n63687 : n14917;
  assign n63689 = pi14 ? n63688 : n49303;
  assign n63690 = pi13 ? n63683 : n63689;
  assign n63691 = pi12 ? n63682 : n63690;
  assign n63692 = pi14 ? n23576 : n23623;
  assign n63693 = pi13 ? n63599 : n63692;
  assign n63694 = pi14 ? n32 : n63598;
  assign n63695 = pi15 ? n23569 : n23749;
  assign n63696 = pi16 ? n3068 : ~n2732;
  assign n63697 = pi16 ? n2745 : ~n2732;
  assign n63698 = pi15 ? n63696 : n63697;
  assign n63699 = pi14 ? n63695 : n63698;
  assign n63700 = pi13 ? n63694 : n63699;
  assign n63701 = pi12 ? n63693 : n63700;
  assign n63702 = pi11 ? n63691 : n63701;
  assign n63703 = pi19 ? n32 : ~n7502;
  assign n63704 = pi18 ? n32 : n63703;
  assign n63705 = pi17 ? n32 : n63704;
  assign n63706 = pi16 ? n3068 : ~n63705;
  assign n63707 = pi15 ? n63706 : n63603;
  assign n63708 = pi14 ? n63707 : n63611;
  assign n63709 = pi15 ? n23847 : n1109;
  assign n63710 = pi14 ? n63617 : n63709;
  assign n63711 = pi13 ? n63708 : n63710;
  assign n63712 = pi14 ? n32 : n24189;
  assign n63713 = pi20 ? n32 : ~n34841;
  assign n63714 = pi19 ? n63713 : ~n32;
  assign n63715 = pi18 ? n49337 : n63714;
  assign n63716 = pi17 ? n32 : ~n63715;
  assign n63717 = pi16 ? n32 : n63716;
  assign n63718 = pi15 ? n63624 : n63717;
  assign n63719 = pi14 ? n63621 : n63718;
  assign n63720 = pi13 ? n63712 : n63719;
  assign n63721 = pi12 ? n63711 : n63720;
  assign n63722 = pi18 ? n32 : ~n1326;
  assign n63723 = pi17 ? n32 : n63722;
  assign n63724 = pi16 ? n32 : n63723;
  assign n63725 = pi15 ? n63724 : n63456;
  assign n63726 = pi14 ? n63725 : n49155;
  assign n63727 = pi16 ? n2860 : ~n2513;
  assign n63728 = pi15 ? n63727 : n49428;
  assign n63729 = pi14 ? n63728 : n63642;
  assign n63730 = pi13 ? n63726 : n63729;
  assign n63731 = pi16 ? n49432 : n2095;
  assign n63732 = pi15 ? n63731 : n21543;
  assign n63733 = pi18 ? n46739 : n21692;
  assign n63734 = pi17 ? n35797 : ~n63733;
  assign n63735 = pi16 ? n1233 : ~n63734;
  assign n63736 = pi18 ? n35804 : n14153;
  assign n63737 = pi17 ? n35803 : ~n63736;
  assign n63738 = pi16 ? n1233 : ~n63737;
  assign n63739 = pi15 ? n63735 : n63738;
  assign n63740 = pi14 ? n63732 : n63739;
  assign n63741 = pi20 ? n287 : n266;
  assign n63742 = pi19 ? n63741 : n18678;
  assign n63743 = pi18 ? n29316 : ~n63742;
  assign n63744 = pi17 ? n32 : n63743;
  assign n63745 = pi17 ? n63659 : ~n35864;
  assign n63746 = pi16 ? n63744 : ~n63745;
  assign n63747 = pi16 ? n29318 : ~n35870;
  assign n63748 = pi15 ? n63746 : n63747;
  assign n63749 = pi14 ? n21035 : n63748;
  assign n63750 = pi13 ? n63740 : n63749;
  assign n63751 = pi12 ? n63730 : n63750;
  assign n63752 = pi11 ? n63721 : n63751;
  assign n63753 = pi10 ? n63702 : n63752;
  assign n63754 = pi09 ? n63677 : n63753;
  assign n63755 = pi08 ? n63669 : n63754;
  assign n63756 = pi07 ? n63568 : n63755;
  assign n63757 = pi06 ? n63372 : n63756;
  assign n63758 = pi05 ? n62963 : n63757;
  assign n63759 = pi04 ? n62042 : n63758;
  assign n63760 = pi19 ? n176 : n589;
  assign n63761 = pi18 ? n1353 : ~n63760;
  assign n63762 = pi17 ? n30283 : n63761;
  assign n63763 = pi16 ? n32 : n63762;
  assign n63764 = pi15 ? n32 : n63763;
  assign n63765 = pi18 ? n268 : n940;
  assign n63766 = pi17 ? n63765 : ~n2839;
  assign n63767 = pi16 ? n32 : n63766;
  assign n63768 = pi20 ? n10889 : n207;
  assign n63769 = pi19 ? n63768 : ~n32;
  assign n63770 = pi18 ? n32 : n63769;
  assign n63771 = pi17 ? n63770 : ~n3067;
  assign n63772 = pi16 ? n32 : n63771;
  assign n63773 = pi15 ? n63767 : n63772;
  assign n63774 = pi14 ? n63764 : n63773;
  assign n63775 = pi13 ? n32 : n63774;
  assign n63776 = pi12 ? n32 : n63775;
  assign n63777 = pi11 ? n32 : n63776;
  assign n63778 = pi10 ? n32 : n63777;
  assign n63779 = pi20 ? n1324 : n9491;
  assign n63780 = pi20 ? n9488 : ~n5854;
  assign n63781 = pi19 ? n63779 : n63780;
  assign n63782 = pi18 ? n32 : n63781;
  assign n63783 = pi19 ? n42535 : n358;
  assign n63784 = pi19 ? n247 : ~n10662;
  assign n63785 = pi18 ? n63783 : n63784;
  assign n63786 = pi17 ? n63782 : ~n63785;
  assign n63787 = pi16 ? n32 : n63786;
  assign n63788 = pi15 ? n63787 : n32;
  assign n63789 = pi16 ? n32 : n44666;
  assign n63790 = pi15 ? n63789 : n32;
  assign n63791 = pi14 ? n63788 : n63790;
  assign n63792 = pi13 ? n63791 : n32;
  assign n63793 = pi15 ? n24382 : n49496;
  assign n63794 = pi15 ? n49501 : n24382;
  assign n63795 = pi14 ? n63793 : n63794;
  assign n63796 = pi15 ? n16377 : n35889;
  assign n63797 = pi14 ? n63796 : n49505;
  assign n63798 = pi13 ? n63795 : n63797;
  assign n63799 = pi12 ? n63792 : n63798;
  assign n63800 = pi19 ? n17194 : n7693;
  assign n63801 = pi18 ? n23571 : n63800;
  assign n63802 = pi17 ? n32 : n63801;
  assign n63803 = pi16 ? n32 : n63802;
  assign n63804 = pi15 ? n49512 : n63803;
  assign n63805 = pi14 ? n63804 : n32;
  assign n63806 = pi15 ? n24247 : n23725;
  assign n63807 = pi14 ? n36285 : n63806;
  assign n63808 = pi13 ? n63805 : n63807;
  assign n63809 = pi14 ? n23726 : n23794;
  assign n63810 = pi16 ? n3165 : ~n2732;
  assign n63811 = pi15 ? n23933 : n63810;
  assign n63812 = pi17 ? n18718 : n2731;
  assign n63813 = pi16 ? n44945 : ~n63812;
  assign n63814 = pi18 ? n32 : n36042;
  assign n63815 = pi17 ? n32 : n63814;
  assign n63816 = pi16 ? n4578 : ~n63815;
  assign n63817 = pi15 ? n63813 : n63816;
  assign n63818 = pi14 ? n63811 : n63817;
  assign n63819 = pi13 ? n63809 : n63818;
  assign n63820 = pi12 ? n63808 : n63819;
  assign n63821 = pi11 ? n63799 : n63820;
  assign n63822 = pi16 ? n49529 : ~n2732;
  assign n63823 = pi16 ? n2958 : ~n2732;
  assign n63824 = pi15 ? n63822 : n63823;
  assign n63825 = pi18 ? n32 : n37593;
  assign n63826 = pi17 ? n32 : n63825;
  assign n63827 = pi16 ? n3068 : ~n63826;
  assign n63828 = pi18 ? n940 : n62604;
  assign n63829 = pi17 ? n63828 : ~n2731;
  assign n63830 = pi16 ? n32 : n63829;
  assign n63831 = pi15 ? n63827 : n63830;
  assign n63832 = pi14 ? n63824 : n63831;
  assign n63833 = pi16 ? n49581 : ~n2732;
  assign n63834 = pi16 ? n3165 : n24017;
  assign n63835 = pi15 ? n63833 : n63834;
  assign n63836 = pi14 ? n63835 : n24186;
  assign n63837 = pi13 ? n63832 : n63836;
  assign n63838 = pi14 ? n32 : n23503;
  assign n63839 = pi18 ? n23539 : n702;
  assign n63840 = pi17 ? n48248 : ~n63839;
  assign n63841 = pi16 ? n32 : n63840;
  assign n63842 = pi15 ? n63841 : n49563;
  assign n63843 = pi19 ? n857 : n1105;
  assign n63844 = pi18 ? n35966 : n63843;
  assign n63845 = pi17 ? n32 : ~n63844;
  assign n63846 = pi16 ? n32 : n63845;
  assign n63847 = pi18 ? n35970 : ~n702;
  assign n63848 = pi17 ? n32 : n63847;
  assign n63849 = pi16 ? n32 : n63848;
  assign n63850 = pi15 ? n63846 : n63849;
  assign n63851 = pi14 ? n63842 : n63850;
  assign n63852 = pi13 ? n63838 : n63851;
  assign n63853 = pi12 ? n63837 : n63852;
  assign n63854 = pi19 ? n4670 : n1740;
  assign n63855 = pi18 ? n32 : n63854;
  assign n63856 = pi17 ? n32 : n63855;
  assign n63857 = pi17 ? n49570 : n2618;
  assign n63858 = pi16 ? n63856 : ~n63857;
  assign n63859 = pi15 ? n13035 : n63858;
  assign n63860 = pi14 ? n63859 : n49579;
  assign n63861 = pi17 ? n32 : n9347;
  assign n63862 = pi16 ? n63861 : n21852;
  assign n63863 = pi15 ? n32 : n63862;
  assign n63864 = pi14 ? n49583 : n63863;
  assign n63865 = pi13 ? n63860 : n63864;
  assign n63866 = pi19 ? n44258 : n32;
  assign n63867 = pi18 ? n32 : ~n63866;
  assign n63868 = pi17 ? n32 : n63867;
  assign n63869 = pi16 ? n1233 : ~n63868;
  assign n63870 = pi20 ? n342 : ~n2102;
  assign n63871 = pi19 ? n63870 : ~n32;
  assign n63872 = pi18 ? n32 : n63871;
  assign n63873 = pi17 ? n32 : n63872;
  assign n63874 = pi16 ? n1233 : ~n63873;
  assign n63875 = pi15 ? n63869 : n63874;
  assign n63876 = pi14 ? n22136 : n63875;
  assign n63877 = pi16 ? n12787 : n21318;
  assign n63878 = pi16 ? n12787 : n32;
  assign n63879 = pi15 ? n63877 : n63878;
  assign n63880 = pi18 ? n366 : ~n5715;
  assign n63881 = pi17 ? n32 : n63880;
  assign n63882 = pi16 ? n63881 : ~n36016;
  assign n63883 = pi19 ? n4391 : n1844;
  assign n63884 = pi18 ? n29316 : ~n63883;
  assign n63885 = pi17 ? n32 : n63884;
  assign n63886 = pi16 ? n63885 : ~n2120;
  assign n63887 = pi15 ? n63882 : n63886;
  assign n63888 = pi14 ? n63879 : n63887;
  assign n63889 = pi13 ? n63876 : n63888;
  assign n63890 = pi12 ? n63865 : n63889;
  assign n63891 = pi11 ? n63853 : n63890;
  assign n63892 = pi10 ? n63821 : n63891;
  assign n63893 = pi09 ? n63778 : n63892;
  assign n63894 = pi20 ? n518 : n207;
  assign n63895 = pi19 ? n63894 : ~n32;
  assign n63896 = pi18 ? n32 : n63895;
  assign n63897 = pi17 ? n63896 : ~n3067;
  assign n63898 = pi16 ? n32 : n63897;
  assign n63899 = pi15 ? n63767 : n63898;
  assign n63900 = pi14 ? n63764 : n63899;
  assign n63901 = pi13 ? n32 : n63900;
  assign n63902 = pi12 ? n32 : n63901;
  assign n63903 = pi11 ? n32 : n63902;
  assign n63904 = pi10 ? n32 : n63903;
  assign n63905 = pi19 ? n247 : ~n19136;
  assign n63906 = pi18 ? n63783 : n63905;
  assign n63907 = pi17 ? n63782 : ~n63906;
  assign n63908 = pi16 ? n32 : n63907;
  assign n63909 = pi15 ? n63908 : n32;
  assign n63910 = pi14 ? n63909 : n63790;
  assign n63911 = pi13 ? n63910 : n32;
  assign n63912 = pi15 ? n24511 : n36100;
  assign n63913 = pi15 ? n49501 : n24511;
  assign n63914 = pi14 ? n63912 : n63913;
  assign n63915 = pi15 ? n24237 : n35889;
  assign n63916 = pi14 ? n63915 : n49505;
  assign n63917 = pi13 ? n63914 : n63916;
  assign n63918 = pi12 ? n63911 : n63917;
  assign n63919 = pi19 ? n9007 : n7693;
  assign n63920 = pi18 ? n32 : n63919;
  assign n63921 = pi17 ? n32 : n63920;
  assign n63922 = pi16 ? n32 : n63921;
  assign n63923 = pi15 ? n49512 : n63922;
  assign n63924 = pi14 ? n63923 : n32;
  assign n63925 = pi14 ? n36285 : n38876;
  assign n63926 = pi13 ? n63924 : n63925;
  assign n63927 = pi14 ? n23924 : n16321;
  assign n63928 = pi16 ? n3165 : ~n2725;
  assign n63929 = pi15 ? n23933 : n63928;
  assign n63930 = pi17 ? n18718 : n2724;
  assign n63931 = pi16 ? n3438 : ~n63930;
  assign n63932 = pi17 ? n32 : n8260;
  assign n63933 = pi16 ? n4578 : ~n63932;
  assign n63934 = pi15 ? n63931 : n63933;
  assign n63935 = pi14 ? n63929 : n63934;
  assign n63936 = pi13 ? n63927 : n63935;
  assign n63937 = pi12 ? n63926 : n63936;
  assign n63938 = pi11 ? n63918 : n63937;
  assign n63939 = pi16 ? n4578 : ~n2725;
  assign n63940 = pi15 ? n63939 : n63823;
  assign n63941 = pi17 ? n32 : n6685;
  assign n63942 = pi16 ? n63941 : ~n63826;
  assign n63943 = pi15 ? n63942 : n63830;
  assign n63944 = pi14 ? n63940 : n63943;
  assign n63945 = pi19 ? n857 : n6298;
  assign n63946 = pi18 ? n32 : n63945;
  assign n63947 = pi17 ? n32 : n63946;
  assign n63948 = pi16 ? n63947 : ~n2732;
  assign n63949 = pi19 ? n32 : ~n6800;
  assign n63950 = pi18 ? n32 : n63949;
  assign n63951 = pi17 ? n32 : n63950;
  assign n63952 = pi16 ? n63951 : n24017;
  assign n63953 = pi15 ? n63948 : n63952;
  assign n63954 = pi16 ? n22539 : n24266;
  assign n63955 = pi15 ? n63954 : n22923;
  assign n63956 = pi14 ? n63953 : n63955;
  assign n63957 = pi13 ? n63944 : n63956;
  assign n63958 = pi14 ? n55548 : n26341;
  assign n63959 = pi18 ? n49653 : ~n7519;
  assign n63960 = pi17 ? n36054 : n63959;
  assign n63961 = pi16 ? n32 : n63960;
  assign n63962 = pi15 ? n63841 : n63961;
  assign n63963 = pi14 ? n63962 : n63850;
  assign n63964 = pi13 ? n63958 : n63963;
  assign n63965 = pi12 ? n63957 : n63964;
  assign n63966 = pi17 ? n49575 : n2628;
  assign n63967 = pi16 ? n49568 : ~n63966;
  assign n63968 = pi16 ? n2958 : ~n2629;
  assign n63969 = pi15 ? n63967 : n63968;
  assign n63970 = pi14 ? n63859 : n63969;
  assign n63971 = pi13 ? n63970 : n63864;
  assign n63972 = pi16 ? n20835 : n21852;
  assign n63973 = pi15 ? n63972 : n21686;
  assign n63974 = pi18 ? n32 : ~n5351;
  assign n63975 = pi17 ? n32 : n63974;
  assign n63976 = pi16 ? n1233 : ~n63975;
  assign n63977 = pi20 ? n342 : ~n16309;
  assign n63978 = pi19 ? n63977 : ~n32;
  assign n63979 = pi18 ? n32 : n63978;
  assign n63980 = pi17 ? n32 : n63979;
  assign n63981 = pi16 ? n1233 : ~n63980;
  assign n63982 = pi15 ? n63976 : n63981;
  assign n63983 = pi14 ? n63973 : n63982;
  assign n63984 = pi18 ? n366 : ~n6147;
  assign n63985 = pi17 ? n32 : n63984;
  assign n63986 = pi16 ? n63985 : ~n36016;
  assign n63987 = pi19 ? n4391 : ~n6683;
  assign n63988 = pi18 ? n29316 : ~n63987;
  assign n63989 = pi17 ? n32 : n63988;
  assign n63990 = pi16 ? n63989 : ~n2120;
  assign n63991 = pi15 ? n63986 : n63990;
  assign n63992 = pi14 ? n63879 : n63991;
  assign n63993 = pi13 ? n63983 : n63992;
  assign n63994 = pi12 ? n63971 : n63993;
  assign n63995 = pi11 ? n63965 : n63994;
  assign n63996 = pi10 ? n63938 : n63995;
  assign n63997 = pi09 ? n63904 : n63996;
  assign n63998 = pi08 ? n63893 : n63997;
  assign n63999 = pi19 ? n4670 : n2317;
  assign n64000 = pi18 ? n5856 : n63999;
  assign n64001 = pi17 ? n3296 : ~n64000;
  assign n64002 = pi16 ? n32 : n64001;
  assign n64003 = pi15 ? n32 : n64002;
  assign n64004 = pi17 ? n45014 : ~n2836;
  assign n64005 = pi16 ? n32 : n64004;
  assign n64006 = pi17 ? n35983 : ~n3067;
  assign n64007 = pi16 ? n32 : n64006;
  assign n64008 = pi15 ? n64005 : n64007;
  assign n64009 = pi14 ? n64003 : n64008;
  assign n64010 = pi13 ? n32 : n64009;
  assign n64011 = pi12 ? n32 : n64010;
  assign n64012 = pi11 ? n32 : n64011;
  assign n64013 = pi10 ? n32 : n64012;
  assign n64014 = pi19 ? n32 : n28041;
  assign n64015 = pi19 ? n23895 : n19317;
  assign n64016 = pi18 ? n64014 : n64015;
  assign n64017 = pi17 ? n32 : n64016;
  assign n64018 = pi16 ? n32 : n64017;
  assign n64019 = pi15 ? n64018 : n24237;
  assign n64020 = pi14 ? n64019 : n24370;
  assign n64021 = pi13 ? n64020 : n32;
  assign n64022 = pi14 ? n63912 : n37789;
  assign n64023 = pi15 ? n24237 : n36095;
  assign n64024 = pi14 ? n64023 : n49716;
  assign n64025 = pi13 ? n64022 : n64024;
  assign n64026 = pi12 ? n64021 : n64025;
  assign n64027 = pi15 ? n49722 : n24237;
  assign n64028 = pi14 ? n64027 : n36285;
  assign n64029 = pi21 ? n7107 : n140;
  assign n64030 = pi20 ? n64029 : ~n32;
  assign n64031 = pi19 ? n32 : ~n64030;
  assign n64032 = pi18 ? n32 : n64031;
  assign n64033 = pi17 ? n32 : n64032;
  assign n64034 = pi16 ? n32 : n64033;
  assign n64035 = pi15 ? n64034 : n32;
  assign n64036 = pi14 ? n35688 : n64035;
  assign n64037 = pi13 ? n64028 : n64036;
  assign n64038 = pi14 ? n23924 : n36111;
  assign n64039 = pi17 ? n18482 : n2724;
  assign n64040 = pi16 ? n32 : ~n64039;
  assign n64041 = pi15 ? n23933 : n64040;
  assign n64042 = pi17 ? n1219 : ~n2724;
  assign n64043 = pi16 ? n32 : n64042;
  assign n64044 = pi19 ? n4670 : ~n3692;
  assign n64045 = pi18 ? n64044 : ~n32;
  assign n64046 = pi17 ? n64045 : ~n8260;
  assign n64047 = pi16 ? n32 : n64046;
  assign n64048 = pi15 ? n64043 : n64047;
  assign n64049 = pi14 ? n64041 : n64048;
  assign n64050 = pi13 ? n64038 : n64049;
  assign n64051 = pi12 ? n64037 : n64050;
  assign n64052 = pi11 ? n64026 : n64051;
  assign n64053 = pi19 ? n349 : ~n1248;
  assign n64054 = pi19 ? n4670 : n19598;
  assign n64055 = pi18 ? n64053 : ~n64054;
  assign n64056 = pi19 ? n15923 : n267;
  assign n64057 = pi18 ? n64056 : n8259;
  assign n64058 = pi17 ? n64055 : ~n64057;
  assign n64059 = pi16 ? n32 : n64058;
  assign n64060 = pi18 ? n32 : n1509;
  assign n64061 = pi17 ? n32 : n64060;
  assign n64062 = pi17 ? n37886 : n2724;
  assign n64063 = pi16 ? n64061 : ~n64062;
  assign n64064 = pi15 ? n64059 : n64063;
  assign n64065 = pi19 ? n23644 : n1740;
  assign n64066 = pi18 ? n64065 : ~n32;
  assign n64067 = pi19 ? n13069 : n813;
  assign n64068 = pi18 ? n20172 : n64067;
  assign n64069 = pi17 ? n64066 : ~n64068;
  assign n64070 = pi16 ? n32 : n64069;
  assign n64071 = pi17 ? n2750 : ~n2724;
  assign n64072 = pi16 ? n32 : n64071;
  assign n64073 = pi15 ? n64070 : n64072;
  assign n64074 = pi14 ? n64064 : n64073;
  assign n64075 = pi19 ? n44373 : ~n1817;
  assign n64076 = pi18 ? n41285 : ~n64075;
  assign n64077 = pi20 ? n17671 : n274;
  assign n64078 = pi19 ? n275 : n64077;
  assign n64079 = pi19 ? n1757 : n813;
  assign n64080 = pi18 ? n64078 : n64079;
  assign n64081 = pi17 ? n64076 : n64080;
  assign n64082 = pi16 ? n3165 : ~n64081;
  assign n64083 = pi16 ? n34460 : n24322;
  assign n64084 = pi15 ? n64082 : n64083;
  assign n64085 = pi16 ? n24236 : n23249;
  assign n64086 = pi15 ? n64085 : n32;
  assign n64087 = pi14 ? n64084 : n64086;
  assign n64088 = pi13 ? n64074 : n64087;
  assign n64089 = pi15 ? n22923 : n22817;
  assign n64090 = pi14 ? n32 : n64089;
  assign n64091 = pi18 ? n222 : ~n7921;
  assign n64092 = pi17 ? n32 : n64091;
  assign n64093 = pi16 ? n32 : n64092;
  assign n64094 = pi15 ? n49762 : n64093;
  assign n64095 = pi18 ? n14873 : n1750;
  assign n64096 = pi17 ? n32 : ~n64095;
  assign n64097 = pi16 ? n32 : n64096;
  assign n64098 = pi15 ? n64097 : n12509;
  assign n64099 = pi14 ? n64094 : n64098;
  assign n64100 = pi13 ? n64090 : n64099;
  assign n64101 = pi12 ? n64088 : n64100;
  assign n64102 = pi19 ? n38795 : ~n32;
  assign n64103 = pi18 ? n262 : ~n64102;
  assign n64104 = pi17 ? n32 : n64103;
  assign n64105 = pi17 ? n49771 : ~n4099;
  assign n64106 = pi16 ? n64104 : n64105;
  assign n64107 = pi15 ? n61968 : n64106;
  assign n64108 = pi14 ? n64107 : n49779;
  assign n64109 = pi21 ? n206 : ~n173;
  assign n64110 = pi20 ? n64109 : ~n32;
  assign n64111 = pi19 ? n32 : n64110;
  assign n64112 = pi18 ? n32 : n64111;
  assign n64113 = pi17 ? n32 : n64112;
  assign n64114 = pi16 ? n64113 : n14789;
  assign n64115 = pi15 ? n648 : n64114;
  assign n64116 = pi14 ? n49783 : n64115;
  assign n64117 = pi13 ? n64108 : n64116;
  assign n64118 = pi18 ? n32 : ~n22003;
  assign n64119 = pi17 ? n32 : n64118;
  assign n64120 = pi16 ? n1233 : ~n64119;
  assign n64121 = pi20 ? n342 : ~n1685;
  assign n64122 = pi19 ? n64121 : ~n32;
  assign n64123 = pi18 ? n32 : n64122;
  assign n64124 = pi17 ? n32 : n64123;
  assign n64125 = pi16 ? n1233 : ~n64124;
  assign n64126 = pi15 ? n64120 : n64125;
  assign n64127 = pi14 ? n21853 : n64126;
  assign n64128 = pi16 ? n12787 : n21388;
  assign n64129 = pi15 ? n64128 : n63878;
  assign n64130 = pi19 ? n1464 : n36510;
  assign n64131 = pi18 ? n366 : ~n64130;
  assign n64132 = pi17 ? n32 : n64131;
  assign n64133 = pi16 ? n64132 : ~n36220;
  assign n64134 = pi19 ? n349 : ~n6327;
  assign n64135 = pi18 ? n29325 : ~n64134;
  assign n64136 = pi17 ? n32 : n64135;
  assign n64137 = pi16 ? n64136 : ~n2409;
  assign n64138 = pi15 ? n64133 : n64137;
  assign n64139 = pi14 ? n64129 : n64138;
  assign n64140 = pi13 ? n64127 : n64139;
  assign n64141 = pi12 ? n64117 : n64140;
  assign n64142 = pi11 ? n64101 : n64141;
  assign n64143 = pi10 ? n64052 : n64142;
  assign n64144 = pi09 ? n64013 : n64143;
  assign n64145 = pi19 ? n32 : ~n14552;
  assign n64146 = pi18 ? n32 : n64145;
  assign n64147 = pi17 ? n32 : n64146;
  assign n64148 = pi16 ? n32 : n64147;
  assign n64149 = pi15 ? n64148 : n36100;
  assign n64150 = pi15 ? n24511 : n24640;
  assign n64151 = pi14 ? n64149 : n64150;
  assign n64152 = pi15 ? n24367 : n36095;
  assign n64153 = pi14 ? n64152 : n49716;
  assign n64154 = pi13 ? n64151 : n64153;
  assign n64155 = pi12 ? n64021 : n64154;
  assign n64156 = pi14 ? n49723 : n24292;
  assign n64157 = pi15 ? n38371 : n32;
  assign n64158 = pi14 ? n32 : n64157;
  assign n64159 = pi13 ? n64156 : n64158;
  assign n64160 = pi15 ? n24289 : n38371;
  assign n64161 = pi14 ? n35688 : n64160;
  assign n64162 = pi17 ? n18482 : n4245;
  assign n64163 = pi16 ? n32 : ~n64162;
  assign n64164 = pi15 ? n24097 : n64163;
  assign n64165 = pi17 ? n1219 : ~n4245;
  assign n64166 = pi16 ? n32 : n64165;
  assign n64167 = pi19 ? n32 : ~n6230;
  assign n64168 = pi18 ? n32 : n64167;
  assign n64169 = pi17 ? n64045 : ~n64168;
  assign n64170 = pi16 ? n32 : n64169;
  assign n64171 = pi15 ? n64166 : n64170;
  assign n64172 = pi14 ? n64164 : n64171;
  assign n64173 = pi13 ? n64161 : n64172;
  assign n64174 = pi12 ? n64159 : n64173;
  assign n64175 = pi11 ? n64155 : n64174;
  assign n64176 = pi20 ? n428 : n18762;
  assign n64177 = pi19 ? n4670 : n64176;
  assign n64178 = pi18 ? n64053 : ~n64177;
  assign n64179 = pi19 ? n58603 : n267;
  assign n64180 = pi18 ? n64179 : n7703;
  assign n64181 = pi17 ? n64178 : ~n64180;
  assign n64182 = pi16 ? n32 : n64181;
  assign n64183 = pi20 ? n32 : ~n333;
  assign n64184 = pi19 ? n32 : n64183;
  assign n64185 = pi18 ? n32 : n64184;
  assign n64186 = pi17 ? n32 : n64185;
  assign n64187 = pi16 ? n64186 : ~n64039;
  assign n64188 = pi15 ? n64182 : n64187;
  assign n64189 = pi14 ? n64188 : n64073;
  assign n64190 = pi20 ? n310 : n287;
  assign n64191 = pi19 ? n64190 : ~n1817;
  assign n64192 = pi18 ? n37954 : ~n64191;
  assign n64193 = pi20 ? n12884 : ~n6621;
  assign n64194 = pi19 ? n275 : ~n64193;
  assign n64195 = pi18 ? n64194 : n64079;
  assign n64196 = pi17 ? n64192 : n64195;
  assign n64197 = pi16 ? n45017 : ~n64196;
  assign n64198 = pi20 ? n342 : ~n1331;
  assign n64199 = pi19 ? n32 : n64198;
  assign n64200 = pi18 ? n32 : n64199;
  assign n64201 = pi17 ? n32 : n64200;
  assign n64202 = pi16 ? n64201 : n24322;
  assign n64203 = pi15 ? n64197 : n64202;
  assign n64204 = pi14 ? n64203 : n64086;
  assign n64205 = pi13 ? n64189 : n64204;
  assign n64206 = pi14 ? n23160 : n64089;
  assign n64207 = pi13 ? n64206 : n64099;
  assign n64208 = pi12 ? n64205 : n64207;
  assign n64209 = pi14 ? n64107 : n49847;
  assign n64210 = pi13 ? n64209 : n64116;
  assign n64211 = pi18 ? n366 : ~n41052;
  assign n64212 = pi17 ? n32 : n64211;
  assign n64213 = pi16 ? n64212 : ~n36220;
  assign n64214 = pi19 ? n349 : ~n208;
  assign n64215 = pi18 ? n940 : ~n64214;
  assign n64216 = pi17 ? n32 : n64215;
  assign n64217 = pi16 ? n64216 : ~n2293;
  assign n64218 = pi15 ? n64213 : n64217;
  assign n64219 = pi14 ? n64129 : n64218;
  assign n64220 = pi13 ? n64127 : n64219;
  assign n64221 = pi12 ? n64210 : n64220;
  assign n64222 = pi11 ? n64208 : n64221;
  assign n64223 = pi10 ? n64175 : n64222;
  assign n64224 = pi09 ? n64013 : n64223;
  assign n64225 = pi08 ? n64144 : n64224;
  assign n64226 = pi07 ? n63998 : n64225;
  assign n64227 = pi18 ? n28164 : n684;
  assign n64228 = pi17 ? n23052 : ~n64227;
  assign n64229 = pi16 ? n32 : n64228;
  assign n64230 = pi15 ? n32 : n64229;
  assign n64231 = pi17 ? n7039 : ~n2836;
  assign n64232 = pi16 ? n32 : n64231;
  assign n64233 = pi15 ? n64232 : n7568;
  assign n64234 = pi14 ? n64230 : n64233;
  assign n64235 = pi13 ? n32 : n64234;
  assign n64236 = pi12 ? n32 : n64235;
  assign n64237 = pi11 ? n32 : n64236;
  assign n64238 = pi10 ? n32 : n64237;
  assign n64239 = pi18 ? n463 : n16449;
  assign n64240 = pi17 ? n32 : n64239;
  assign n64241 = pi16 ? n32 : n64240;
  assign n64242 = pi15 ? n64241 : n32;
  assign n64243 = pi14 ? n64242 : n24498;
  assign n64244 = pi14 ? n24368 : n32;
  assign n64245 = pi13 ? n64243 : n64244;
  assign n64246 = pi15 ? n24237 : n24712;
  assign n64247 = pi14 ? n49885 : n64246;
  assign n64248 = pi15 ? n25155 : n24640;
  assign n64249 = pi14 ? n64248 : n24640;
  assign n64250 = pi13 ? n64247 : n64249;
  assign n64251 = pi12 ? n64245 : n64250;
  assign n64252 = pi14 ? n26994 : n24239;
  assign n64253 = pi13 ? n49896 : n64252;
  assign n64254 = pi14 ? n35688 : n24383;
  assign n64255 = pi19 ? n20884 : ~n287;
  assign n64256 = pi18 ? n37815 : n64255;
  assign n64257 = pi22 ? n84 : n34;
  assign n64258 = pi21 ? n64257 : ~n32;
  assign n64259 = pi20 ? n64258 : ~n32;
  assign n64260 = pi19 ? n33674 : n64259;
  assign n64261 = pi18 ? n20611 : n64260;
  assign n64262 = pi17 ? n64256 : ~n64261;
  assign n64263 = pi16 ? n32 : n64262;
  assign n64264 = pi17 ? n1682 : ~n2724;
  assign n64265 = pi16 ? n32 : n64264;
  assign n64266 = pi15 ? n64263 : n64265;
  assign n64267 = pi19 ? n2386 : ~n4670;
  assign n64268 = pi18 ? n64267 : ~n32;
  assign n64269 = pi19 ? n32 : n20022;
  assign n64270 = pi18 ? n32 : n64269;
  assign n64271 = pi17 ? n64268 : ~n64270;
  assign n64272 = pi16 ? n32 : n64271;
  assign n64273 = pi15 ? n6614 : n64272;
  assign n64274 = pi14 ? n64266 : n64273;
  assign n64275 = pi13 ? n64254 : n64274;
  assign n64276 = pi12 ? n64253 : n64275;
  assign n64277 = pi11 ? n64251 : n64276;
  assign n64278 = pi19 ? n42107 : ~n32;
  assign n64279 = pi18 ? n64278 : ~n32;
  assign n64280 = pi17 ? n64279 : ~n4245;
  assign n64281 = pi16 ? n32 : n64280;
  assign n64282 = pi20 ? n207 : n439;
  assign n64283 = pi19 ? n64282 : n32;
  assign n64284 = pi18 ? n64283 : n32;
  assign n64285 = pi19 ? n5694 : n18728;
  assign n64286 = pi19 ? n4342 : n1812;
  assign n64287 = pi18 ? n64285 : n64286;
  assign n64288 = pi17 ? n64284 : n64287;
  assign n64289 = pi16 ? n32 : ~n64288;
  assign n64290 = pi15 ? n64281 : n64289;
  assign n64291 = pi19 ? n6342 : n1812;
  assign n64292 = pi18 ? n268 : n64291;
  assign n64293 = pi17 ? n5010 : ~n64292;
  assign n64294 = pi16 ? n32 : n64293;
  assign n64295 = pi15 ? n64294 : n50986;
  assign n64296 = pi14 ? n64290 : n64295;
  assign n64297 = pi17 ? n1028 : ~n24455;
  assign n64298 = pi16 ? n3165 : ~n64297;
  assign n64299 = pi17 ? n1124 : n1527;
  assign n64300 = pi16 ? n3165 : n64299;
  assign n64301 = pi15 ? n64298 : n64300;
  assign n64302 = pi14 ? n64301 : n23252;
  assign n64303 = pi13 ? n64296 : n64302;
  assign n64304 = pi19 ? n4126 : ~n617;
  assign n64305 = pi18 ? n32 : n64304;
  assign n64306 = pi17 ? n32 : n64305;
  assign n64307 = pi16 ? n32 : n64306;
  assign n64308 = pi18 ? n42558 : ~n702;
  assign n64309 = pi17 ? n32 : n64308;
  assign n64310 = pi16 ? n32 : n64309;
  assign n64311 = pi15 ? n64307 : n64310;
  assign n64312 = pi14 ? n23582 : n64311;
  assign n64313 = pi18 ? n49948 : n8884;
  assign n64314 = pi17 ? n49947 : ~n64313;
  assign n64315 = pi16 ? n32 : n64314;
  assign n64316 = pi19 ? n507 : n2614;
  assign n64317 = pi18 ? n32 : ~n64316;
  assign n64318 = pi17 ? n32 : n64317;
  assign n64319 = pi16 ? n32 : n64318;
  assign n64320 = pi15 ? n64315 : n64319;
  assign n64321 = pi18 ? n36360 : ~n7921;
  assign n64322 = pi17 ? n32 : n64321;
  assign n64323 = pi16 ? n32 : n64322;
  assign n64324 = pi18 ? n36364 : ~n63843;
  assign n64325 = pi17 ? n32 : n64324;
  assign n64326 = pi16 ? n32 : n64325;
  assign n64327 = pi15 ? n64323 : n64326;
  assign n64328 = pi14 ? n64320 : n64327;
  assign n64329 = pi13 ? n64312 : n64328;
  assign n64330 = pi12 ? n64303 : n64329;
  assign n64331 = pi20 ? n18762 : n342;
  assign n64332 = pi19 ? n64331 : ~n12854;
  assign n64333 = pi18 ? n209 : ~n64332;
  assign n64334 = pi17 ? n32 : n64333;
  assign n64335 = pi18 ? n49956 : ~n2684;
  assign n64336 = pi17 ? n32 : n64335;
  assign n64337 = pi16 ? n64334 : n64336;
  assign n64338 = pi18 ? n49963 : ~n4098;
  assign n64339 = pi17 ? n49961 : n64338;
  assign n64340 = pi16 ? n882 : n64339;
  assign n64341 = pi15 ? n64337 : n64340;
  assign n64342 = pi18 ? n49975 : ~n508;
  assign n64343 = pi17 ? n49973 : n64342;
  assign n64344 = pi16 ? n32 : n64343;
  assign n64345 = pi15 ? n64344 : n49983;
  assign n64346 = pi14 ? n64341 : n64345;
  assign n64347 = pi16 ? n48707 : n647;
  assign n64348 = pi15 ? n32 : n64347;
  assign n64349 = pi14 ? n49991 : n64348;
  assign n64350 = pi13 ? n64346 : n64349;
  assign n64351 = pi18 ? n24025 : ~n21683;
  assign n64352 = pi17 ? n32 : n64351;
  assign n64353 = pi16 ? n1233 : ~n64352;
  assign n64354 = pi19 ? n208 : n16002;
  assign n64355 = pi18 ? n323 : ~n64354;
  assign n64356 = pi19 ? n4721 : ~n13069;
  assign n64357 = pi18 ? n64356 : ~n9578;
  assign n64358 = pi17 ? n64355 : n64357;
  assign n64359 = pi16 ? n1233 : ~n64358;
  assign n64360 = pi15 ? n64353 : n64359;
  assign n64361 = pi14 ? n22261 : n64360;
  assign n64362 = pi18 ? n14429 : n32;
  assign n64363 = pi17 ? n64362 : n14395;
  assign n64364 = pi16 ? n10984 : n64363;
  assign n64365 = pi16 ? n1046 : n50004;
  assign n64366 = pi15 ? n64364 : n64365;
  assign n64367 = pi17 ? n1028 : ~n2653;
  assign n64368 = pi16 ? n1243 : n64367;
  assign n64369 = pi17 ? n1500 : ~n2408;
  assign n64370 = pi16 ? n11695 : n64369;
  assign n64371 = pi15 ? n64368 : n64370;
  assign n64372 = pi14 ? n64366 : n64371;
  assign n64373 = pi13 ? n64361 : n64372;
  assign n64374 = pi12 ? n64350 : n64373;
  assign n64375 = pi11 ? n64330 : n64374;
  assign n64376 = pi10 ? n64277 : n64375;
  assign n64377 = pi09 ? n64238 : n64376;
  assign n64378 = pi17 ? n7039 : ~n2839;
  assign n64379 = pi16 ? n32 : n64378;
  assign n64380 = pi15 ? n64379 : n7568;
  assign n64381 = pi14 ? n64230 : n64380;
  assign n64382 = pi13 ? n32 : n64381;
  assign n64383 = pi12 ? n32 : n64382;
  assign n64384 = pi11 ? n32 : n64383;
  assign n64385 = pi10 ? n32 : n64384;
  assign n64386 = pi14 ? n32 : n24496;
  assign n64387 = pi13 ? n64243 : n64386;
  assign n64388 = pi15 ? n24237 : n16101;
  assign n64389 = pi14 ? n50036 : n64388;
  assign n64390 = pi15 ? n25301 : n24640;
  assign n64391 = pi14 ? n64390 : n64150;
  assign n64392 = pi13 ? n64389 : n64391;
  assign n64393 = pi12 ? n64387 : n64392;
  assign n64394 = pi13 ? n50043 : n64252;
  assign n64395 = pi14 ? n26994 : n25924;
  assign n64396 = pi20 ? n2019 : ~n274;
  assign n64397 = pi19 ? n64396 : n19731;
  assign n64398 = pi18 ? n37872 : ~n64397;
  assign n64399 = pi20 ? n19731 : n32;
  assign n64400 = pi19 ? n64399 : n32;
  assign n64401 = pi19 ? n23193 : n349;
  assign n64402 = pi18 ? n64400 : n64401;
  assign n64403 = pi17 ? n64398 : ~n64402;
  assign n64404 = pi16 ? n32 : n64403;
  assign n64405 = pi15 ? n64404 : n6985;
  assign n64406 = pi19 ? n507 : ~n4670;
  assign n64407 = pi18 ? n64406 : ~n32;
  assign n64408 = pi17 ? n64407 : ~n2852;
  assign n64409 = pi16 ? n32 : n64408;
  assign n64410 = pi15 ? n7051 : n64409;
  assign n64411 = pi14 ? n64405 : n64410;
  assign n64412 = pi13 ? n64395 : n64411;
  assign n64413 = pi12 ? n64394 : n64412;
  assign n64414 = pi11 ? n64393 : n64413;
  assign n64415 = pi18 ? n10710 : ~n32;
  assign n64416 = pi19 ? n32 : n63162;
  assign n64417 = pi18 ? n32 : n64416;
  assign n64418 = pi17 ? n64415 : ~n64417;
  assign n64419 = pi16 ? n32 : n64418;
  assign n64420 = pi18 ? n13058 : n32;
  assign n64421 = pi17 ? n64420 : n64287;
  assign n64422 = pi16 ? n32 : ~n64421;
  assign n64423 = pi15 ? n64419 : n64422;
  assign n64424 = pi19 ? n6342 : n813;
  assign n64425 = pi18 ? n268 : n64424;
  assign n64426 = pi17 ? n5010 : ~n64425;
  assign n64427 = pi16 ? n32 : n64426;
  assign n64428 = pi15 ? n64427 : n50986;
  assign n64429 = pi14 ? n64423 : n64428;
  assign n64430 = pi17 ? n1354 : ~n24455;
  assign n64431 = pi16 ? n3165 : ~n64430;
  assign n64432 = pi17 ? n1124 : n23572;
  assign n64433 = pi16 ? n3165 : n64432;
  assign n64434 = pi15 ? n64431 : n64433;
  assign n64435 = pi14 ? n64434 : n24522;
  assign n64436 = pi13 ? n64429 : n64435;
  assign n64437 = pi15 ? n64307 : n50267;
  assign n64438 = pi14 ? n23582 : n64437;
  assign n64439 = pi18 ? n32 : ~n7510;
  assign n64440 = pi17 ? n32 : n64439;
  assign n64441 = pi16 ? n32 : n64440;
  assign n64442 = pi15 ? n64315 : n64441;
  assign n64443 = pi19 ? n18982 : n617;
  assign n64444 = pi18 ? n36364 : ~n64443;
  assign n64445 = pi17 ? n32 : n64444;
  assign n64446 = pi16 ? n32 : n64445;
  assign n64447 = pi15 ? n64323 : n64446;
  assign n64448 = pi14 ? n64442 : n64447;
  assign n64449 = pi13 ? n64438 : n64448;
  assign n64450 = pi12 ? n64436 : n64449;
  assign n64451 = pi19 ? n428 : ~n12854;
  assign n64452 = pi18 ? n1395 : ~n64451;
  assign n64453 = pi17 ? n32 : n64452;
  assign n64454 = pi18 ? n49956 : ~n2622;
  assign n64455 = pi17 ? n32 : n64454;
  assign n64456 = pi16 ? n64453 : n64455;
  assign n64457 = pi18 ? n49963 : ~n702;
  assign n64458 = pi17 ? n49961 : n64457;
  assign n64459 = pi16 ? n1059 : n64458;
  assign n64460 = pi15 ? n64456 : n64459;
  assign n64461 = pi16 ? n32 : n50076;
  assign n64462 = pi15 ? n64461 : n50080;
  assign n64463 = pi14 ? n64460 : n64462;
  assign n64464 = pi20 ? n342 : n310;
  assign n64465 = pi19 ? n32 : n64464;
  assign n64466 = pi18 ? n32 : n64465;
  assign n64467 = pi17 ? n32 : n64466;
  assign n64468 = pi16 ? n64467 : n15122;
  assign n64469 = pi15 ? n15123 : n64468;
  assign n64470 = pi14 ? n50084 : n64469;
  assign n64471 = pi13 ? n64463 : n64470;
  assign n64472 = pi18 ? n24025 : ~n39579;
  assign n64473 = pi17 ? n32 : n64472;
  assign n64474 = pi16 ? n1233 : ~n64473;
  assign n64475 = pi18 ? n64356 : ~n384;
  assign n64476 = pi17 ? n64355 : n64475;
  assign n64477 = pi16 ? n1233 : ~n64476;
  assign n64478 = pi15 ? n64474 : n64477;
  assign n64479 = pi14 ? n14790 : n64478;
  assign n64480 = pi17 ? n64362 : n21693;
  assign n64481 = pi16 ? n10984 : n64480;
  assign n64482 = pi16 ? n1243 : n50089;
  assign n64483 = pi15 ? n64481 : n64482;
  assign n64484 = pi18 ? n32 : n60983;
  assign n64485 = pi17 ? n1354 : ~n64484;
  assign n64486 = pi16 ? n1243 : n64485;
  assign n64487 = pi16 ? n11695 : n38281;
  assign n64488 = pi15 ? n64486 : n64487;
  assign n64489 = pi14 ? n64483 : n64488;
  assign n64490 = pi13 ? n64479 : n64489;
  assign n64491 = pi12 ? n64471 : n64490;
  assign n64492 = pi11 ? n64450 : n64491;
  assign n64493 = pi10 ? n64414 : n64492;
  assign n64494 = pi09 ? n64385 : n64493;
  assign n64495 = pi08 ? n64377 : n64494;
  assign n64496 = pi19 ? n3495 : n2303;
  assign n64497 = pi18 ? n222 : ~n64496;
  assign n64498 = pi17 ? n32 : n64497;
  assign n64499 = pi16 ? n32 : n64498;
  assign n64500 = pi15 ? n32 : n64499;
  assign n64501 = pi18 ? n880 : ~n684;
  assign n64502 = pi17 ? n32 : n64501;
  assign n64503 = pi16 ? n32 : n64502;
  assign n64504 = pi15 ? n64503 : n9335;
  assign n64505 = pi14 ? n64500 : n64504;
  assign n64506 = pi13 ? n32 : n64505;
  assign n64507 = pi12 ? n32 : n64506;
  assign n64508 = pi11 ? n32 : n64507;
  assign n64509 = pi10 ? n32 : n64508;
  assign n64510 = pi14 ? n25965 : n16840;
  assign n64511 = pi14 ? n16606 : n24563;
  assign n64512 = pi13 ? n64510 : n64511;
  assign n64513 = pi14 ? n50121 : n64388;
  assign n64514 = pi13 ? n64513 : n24700;
  assign n64515 = pi12 ? n64512 : n64514;
  assign n64516 = pi14 ? n24633 : n24237;
  assign n64517 = pi14 ? n36807 : n24370;
  assign n64518 = pi13 ? n64516 : n64517;
  assign n64519 = pi14 ? n26994 : n24512;
  assign n64520 = pi19 ? n18396 : ~n32;
  assign n64521 = pi18 ? n4380 : n64520;
  assign n64522 = pi17 ? n64521 : ~n2724;
  assign n64523 = pi16 ? n32 : n64522;
  assign n64524 = pi15 ? n64523 : n6985;
  assign n64525 = pi14 ? n64524 : n7051;
  assign n64526 = pi13 ? n64519 : n64525;
  assign n64527 = pi12 ? n64518 : n64526;
  assign n64528 = pi11 ? n64515 : n64527;
  assign n64529 = pi18 ? n10923 : ~n32;
  assign n64530 = pi17 ? n64529 : ~n3067;
  assign n64531 = pi16 ? n32 : n64530;
  assign n64532 = pi19 ? n11374 : n617;
  assign n64533 = pi18 ? n64532 : ~n32;
  assign n64534 = pi19 ? n4721 : n18728;
  assign n64535 = pi19 ? n36510 : n349;
  assign n64536 = pi18 ? n64534 : n64535;
  assign n64537 = pi17 ? n64533 : ~n64536;
  assign n64538 = pi16 ? n32 : n64537;
  assign n64539 = pi15 ? n64531 : n64538;
  assign n64540 = pi19 ? n247 : n349;
  assign n64541 = pi18 ? n24775 : n64540;
  assign n64542 = pi17 ? n5010 : ~n64541;
  assign n64543 = pi16 ? n32 : n64542;
  assign n64544 = pi15 ? n64543 : n8587;
  assign n64545 = pi14 ? n64539 : n64544;
  assign n64546 = pi19 ? n9208 : ~n32;
  assign n64547 = pi18 ? n64546 : ~n32;
  assign n64548 = pi17 ? n64547 : ~n24602;
  assign n64549 = pi16 ? n3165 : ~n64548;
  assign n64550 = pi17 ? n18718 : n23572;
  assign n64551 = pi16 ? n3165 : n64550;
  assign n64552 = pi15 ? n64549 : n64551;
  assign n64553 = pi14 ? n64552 : n23632;
  assign n64554 = pi13 ? n64545 : n64553;
  assign n64555 = pi15 ? n36533 : n50267;
  assign n64556 = pi14 ? n23582 : n64555;
  assign n64557 = pi15 ? n50167 : n64441;
  assign n64558 = pi18 ? n6581 : ~n64316;
  assign n64559 = pi17 ? n32 : n64558;
  assign n64560 = pi16 ? n32 : n64559;
  assign n64561 = pi18 ? n6145 : ~n776;
  assign n64562 = pi17 ? n32 : n64561;
  assign n64563 = pi16 ? n32 : n64562;
  assign n64564 = pi15 ? n64560 : n64563;
  assign n64565 = pi14 ? n64557 : n64564;
  assign n64566 = pi13 ? n64556 : n64565;
  assign n64567 = pi12 ? n64554 : n64566;
  assign n64568 = pi19 ? n32 : n33796;
  assign n64569 = pi18 ? n366 : ~n64568;
  assign n64570 = pi17 ? n32 : n64569;
  assign n64571 = pi18 ? n6145 : ~n2622;
  assign n64572 = pi17 ? n32 : n64571;
  assign n64573 = pi16 ? n64570 : n64572;
  assign n64574 = pi18 ? n21274 : ~n702;
  assign n64575 = pi17 ? n8617 : n64574;
  assign n64576 = pi16 ? n11462 : n64575;
  assign n64577 = pi15 ? n64573 : n64576;
  assign n64578 = pi14 ? n64577 : n50184;
  assign n64579 = pi14 ? n50188 : n15123;
  assign n64580 = pi13 ? n64578 : n64579;
  assign n64581 = pi18 ? n36574 : ~n20020;
  assign n64582 = pi17 ? n36573 : n64581;
  assign n64583 = pi16 ? n1233 : ~n64582;
  assign n64584 = pi18 ? n366 : ~n50192;
  assign n64585 = pi17 ? n32 : n64584;
  assign n64586 = pi17 ? n1124 : n21541;
  assign n64587 = pi16 ? n64585 : n64586;
  assign n64588 = pi15 ? n64583 : n64587;
  assign n64589 = pi14 ? n22260 : n64588;
  assign n64590 = pi16 ? n1046 : n64480;
  assign n64591 = pi16 ? n1243 : n50206;
  assign n64592 = pi15 ? n64590 : n64591;
  assign n64593 = pi17 ? n36590 : ~n2519;
  assign n64594 = pi16 ? n1243 : n64593;
  assign n64595 = pi20 ? n321 : ~n448;
  assign n64596 = pi19 ? n64595 : ~n32;
  assign n64597 = pi18 ? n64596 : ~n32;
  assign n64598 = pi20 ? n32 : n15930;
  assign n64599 = pi19 ? n64598 : ~n32;
  assign n64600 = pi18 ? n32 : n64599;
  assign n64601 = pi17 ? n64597 : ~n64600;
  assign n64602 = pi16 ? n11695 : n64601;
  assign n64603 = pi15 ? n64594 : n64602;
  assign n64604 = pi14 ? n64592 : n64603;
  assign n64605 = pi13 ? n64589 : n64604;
  assign n64606 = pi12 ? n64580 : n64605;
  assign n64607 = pi11 ? n64567 : n64606;
  assign n64608 = pi10 ? n64528 : n64607;
  assign n64609 = pi09 ? n64509 : n64608;
  assign n64610 = pi14 ? n16607 : n16840;
  assign n64611 = pi14 ? n32 : n24627;
  assign n64612 = pi13 ? n64610 : n64611;
  assign n64613 = pi15 ? n24237 : n25044;
  assign n64614 = pi14 ? n50239 : n64613;
  assign n64615 = pi15 ? n50341 : n24700;
  assign n64616 = pi14 ? n64615 : n24700;
  assign n64617 = pi13 ? n64614 : n64616;
  assign n64618 = pi12 ? n64612 : n64617;
  assign n64619 = pi14 ? n24567 : n24573;
  assign n64620 = pi14 ? n26994 : n32;
  assign n64621 = pi13 ? n64619 : n64620;
  assign n64622 = pi14 ? n36807 : n51985;
  assign n64623 = pi17 ? n64521 : ~n2850;
  assign n64624 = pi16 ? n32 : n64623;
  assign n64625 = pi17 ? n1682 : ~n2850;
  assign n64626 = pi16 ? n32 : n64625;
  assign n64627 = pi15 ? n64624 : n64626;
  assign n64628 = pi14 ? n64627 : n7051;
  assign n64629 = pi13 ? n64622 : n64628;
  assign n64630 = pi12 ? n64621 : n64629;
  assign n64631 = pi11 ? n64618 : n64630;
  assign n64632 = pi19 ? n9864 : n617;
  assign n64633 = pi18 ? n64632 : ~n32;
  assign n64634 = pi17 ? n64633 : ~n64536;
  assign n64635 = pi16 ? n32 : n64634;
  assign n64636 = pi15 ? n64531 : n64635;
  assign n64637 = pi14 ? n64636 : n64544;
  assign n64638 = pi19 ? n25120 : ~n32;
  assign n64639 = pi18 ? n64638 : ~n32;
  assign n64640 = pi19 ? n24600 : n6230;
  assign n64641 = pi18 ? n24647 : n64640;
  assign n64642 = pi17 ? n64639 : ~n64641;
  assign n64643 = pi16 ? n3165 : ~n64642;
  assign n64644 = pi19 ? n18111 : n32;
  assign n64645 = pi18 ? n64644 : n32;
  assign n64646 = pi17 ? n64645 : n23723;
  assign n64647 = pi16 ? n3165 : n64646;
  assign n64648 = pi15 ? n64643 : n64647;
  assign n64649 = pi14 ? n64648 : n24654;
  assign n64650 = pi13 ? n64637 : n64649;
  assign n64651 = pi15 ? n36631 : n50267;
  assign n64652 = pi14 ? n23250 : n64651;
  assign n64653 = pi18 ? n50164 : n772;
  assign n64654 = pi17 ? n15845 : ~n64653;
  assign n64655 = pi16 ? n32 : n64654;
  assign n64656 = pi18 ? n32 : ~n5983;
  assign n64657 = pi17 ? n32 : n64656;
  assign n64658 = pi16 ? n32 : n64657;
  assign n64659 = pi15 ? n64655 : n64658;
  assign n64660 = pi18 ? n6145 : ~n9960;
  assign n64661 = pi17 ? n32 : n64660;
  assign n64662 = pi16 ? n32 : n64661;
  assign n64663 = pi15 ? n64560 : n64662;
  assign n64664 = pi14 ? n64659 : n64663;
  assign n64665 = pi13 ? n64652 : n64664;
  assign n64666 = pi12 ? n64650 : n64665;
  assign n64667 = pi18 ? n341 : ~n64568;
  assign n64668 = pi17 ? n32 : n64667;
  assign n64669 = pi18 ? n6145 : ~n1750;
  assign n64670 = pi17 ? n32 : n64669;
  assign n64671 = pi16 ? n64668 : n64670;
  assign n64672 = pi15 ? n64671 : n64576;
  assign n64673 = pi14 ? n64672 : n50277;
  assign n64674 = pi17 ? n50279 : n2080;
  assign n64675 = pi16 ? n32 : n64674;
  assign n64676 = pi15 ? n50187 : n64675;
  assign n64677 = pi14 ? n64676 : n24193;
  assign n64678 = pi13 ? n64673 : n64677;
  assign n64679 = pi17 ? n50279 : n15121;
  assign n64680 = pi16 ? n32 : n64679;
  assign n64681 = pi15 ? n64680 : n14790;
  assign n64682 = pi15 ? n64583 : n21686;
  assign n64683 = pi14 ? n64681 : n64682;
  assign n64684 = pi17 ? n64362 : n14392;
  assign n64685 = pi16 ? n1046 : n64684;
  assign n64686 = pi17 ? n50295 : n2279;
  assign n64687 = pi16 ? n1243 : n64686;
  assign n64688 = pi15 ? n64685 : n64687;
  assign n64689 = pi17 ? n36647 : ~n2755;
  assign n64690 = pi16 ? n1243 : n64689;
  assign n64691 = pi18 ? n22486 : ~n32;
  assign n64692 = pi17 ? n64691 : ~n61066;
  assign n64693 = pi16 ? n11695 : n64692;
  assign n64694 = pi15 ? n64690 : n64693;
  assign n64695 = pi14 ? n64688 : n64694;
  assign n64696 = pi13 ? n64683 : n64695;
  assign n64697 = pi12 ? n64678 : n64696;
  assign n64698 = pi11 ? n64666 : n64697;
  assign n64699 = pi10 ? n64631 : n64698;
  assign n64700 = pi09 ? n64509 : n64699;
  assign n64701 = pi08 ? n64609 : n64700;
  assign n64702 = pi07 ? n64495 : n64701;
  assign n64703 = pi06 ? n64226 : n64702;
  assign n64704 = pi18 ? n940 : ~n48595;
  assign n64705 = pi17 ? n32 : n64704;
  assign n64706 = pi16 ? n32 : n64705;
  assign n64707 = pi15 ? n32 : n64706;
  assign n64708 = pi19 ? n6057 : n343;
  assign n64709 = pi18 ? n880 : ~n64708;
  assign n64710 = pi17 ? n32 : n64709;
  assign n64711 = pi16 ? n32 : n64710;
  assign n64712 = pi20 ? n32 : ~n18255;
  assign n64713 = pi20 ? n266 : n29457;
  assign n64714 = pi19 ? n64712 : n64713;
  assign n64715 = pi20 ? n6822 : n21111;
  assign n64716 = pi19 ? n64715 : n12885;
  assign n64717 = pi18 ? n64714 : n64716;
  assign n64718 = pi17 ? n32 : n64717;
  assign n64719 = pi16 ? n32 : n64718;
  assign n64720 = pi15 ? n64711 : n64719;
  assign n64721 = pi14 ? n64707 : n64720;
  assign n64722 = pi13 ? n32 : n64721;
  assign n64723 = pi12 ? n32 : n64722;
  assign n64724 = pi11 ? n32 : n64723;
  assign n64725 = pi10 ? n32 : n64724;
  assign n64726 = pi18 ? n32 : n48732;
  assign n64727 = pi17 ? n32 : n64726;
  assign n64728 = pi16 ? n32 : n64727;
  assign n64729 = pi15 ? n64728 : n50335;
  assign n64730 = pi14 ? n16840 : n64729;
  assign n64731 = pi13 ? n24799 : n64730;
  assign n64732 = pi18 ? n49295 : n50233;
  assign n64733 = pi17 ? n32 : n64732;
  assign n64734 = pi16 ? n32 : n64733;
  assign n64735 = pi15 ? n50345 : n64734;
  assign n64736 = pi14 ? n50342 : n64735;
  assign n64737 = pi15 ? n50341 : n25044;
  assign n64738 = pi14 ? n64737 : n50357;
  assign n64739 = pi13 ? n64736 : n64738;
  assign n64740 = pi12 ? n64731 : n64739;
  assign n64741 = pi14 ? n16606 : n32;
  assign n64742 = pi13 ? n16841 : n64741;
  assign n64743 = pi15 ? n32 : n24712;
  assign n64744 = pi19 ? n322 : ~n9724;
  assign n64745 = pi18 ? n863 : ~n64744;
  assign n64746 = pi17 ? n32 : n64745;
  assign n64747 = pi16 ? n32 : n64746;
  assign n64748 = pi15 ? n24712 : n64747;
  assign n64749 = pi14 ? n64743 : n64748;
  assign n64750 = pi17 ? n1807 : ~n9670;
  assign n64751 = pi16 ? n32 : n64750;
  assign n64752 = pi15 ? n7904 : n64751;
  assign n64753 = pi17 ? n24786 : ~n3067;
  assign n64754 = pi16 ? n32 : n64753;
  assign n64755 = pi15 ? n6559 : n64754;
  assign n64756 = pi14 ? n64752 : n64755;
  assign n64757 = pi13 ? n64749 : n64756;
  assign n64758 = pi12 ? n64742 : n64757;
  assign n64759 = pi11 ? n64740 : n64758;
  assign n64760 = pi19 ? n343 : n349;
  assign n64761 = pi18 ? n32 : n64760;
  assign n64762 = pi17 ? n1933 : ~n64761;
  assign n64763 = pi16 ? n32 : n64762;
  assign n64764 = pi20 ? n18762 : n2358;
  assign n64765 = pi19 ? n32 : n64764;
  assign n64766 = pi18 ? n64765 : ~n32;
  assign n64767 = pi17 ? n64766 : ~n3067;
  assign n64768 = pi16 ? n32 : n64767;
  assign n64769 = pi15 ? n64763 : n64768;
  assign n64770 = pi17 ? n2531 : n50873;
  assign n64771 = pi16 ? n32 : n64770;
  assign n64772 = pi15 ? n64771 : n24734;
  assign n64773 = pi14 ? n64769 : n64772;
  assign n64774 = pi17 ? n20200 : n16103;
  assign n64775 = pi16 ? n32 : n64774;
  assign n64776 = pi15 ? n64775 : n23725;
  assign n64777 = pi14 ? n64776 : n24654;
  assign n64778 = pi13 ? n64773 : n64777;
  assign n64779 = pi15 ? n50558 : n50385;
  assign n64780 = pi14 ? n23484 : n64779;
  assign n64781 = pi18 ? n36720 : n48314;
  assign n64782 = pi17 ? n32 : n64781;
  assign n64783 = pi16 ? n32 : n64782;
  assign n64784 = pi18 ? n36726 : n5725;
  assign n64785 = pi17 ? n32 : n64784;
  assign n64786 = pi16 ? n32 : n64785;
  assign n64787 = pi15 ? n64783 : n64786;
  assign n64788 = pi19 ? n813 : n5626;
  assign n64789 = pi18 ? n36731 : n64788;
  assign n64790 = pi17 ? n32 : n64789;
  assign n64791 = pi16 ? n32 : n64790;
  assign n64792 = pi19 ? n813 : ~n2614;
  assign n64793 = pi18 ? n16041 : n64792;
  assign n64794 = pi17 ? n32 : n64793;
  assign n64795 = pi16 ? n32 : n64794;
  assign n64796 = pi15 ? n64791 : n64795;
  assign n64797 = pi14 ? n64787 : n64796;
  assign n64798 = pi13 ? n64780 : n64797;
  assign n64799 = pi12 ? n64778 : n64798;
  assign n64800 = pi18 ? n15844 : n48117;
  assign n64801 = pi17 ? n32 : n64800;
  assign n64802 = pi16 ? n31463 : n64801;
  assign n64803 = pi16 ? n31463 : n7354;
  assign n64804 = pi15 ? n64802 : n64803;
  assign n64805 = pi14 ? n64804 : n50407;
  assign n64806 = pi14 ? n22424 : n23771;
  assign n64807 = pi13 ? n64805 : n64806;
  assign n64808 = pi19 ? n28481 : n1844;
  assign n64809 = pi18 ? n19245 : n64808;
  assign n64810 = pi19 ? n17737 : n32;
  assign n64811 = pi20 ? n339 : ~n7880;
  assign n64812 = pi19 ? n64811 : ~n32;
  assign n64813 = pi18 ? n64810 : ~n64812;
  assign n64814 = pi17 ? n64809 : n64813;
  assign n64815 = pi16 ? n32 : n64814;
  assign n64816 = pi15 ? n15123 : n64815;
  assign n64817 = pi18 ? n13080 : n32584;
  assign n64818 = pi17 ? n32 : ~n64817;
  assign n64819 = pi16 ? n1233 : ~n64818;
  assign n64820 = pi15 ? n64819 : n21786;
  assign n64821 = pi14 ? n64816 : n64820;
  assign n64822 = pi18 ? n14429 : ~n32;
  assign n64823 = pi19 ? n33526 : ~n32;
  assign n64824 = pi18 ? n16847 : ~n64823;
  assign n64825 = pi17 ? n64822 : ~n64824;
  assign n64826 = pi16 ? n1135 : ~n64825;
  assign n64827 = pi17 ? n36789 : n2755;
  assign n64828 = pi16 ? n19652 : ~n64827;
  assign n64829 = pi15 ? n64826 : n64828;
  assign n64830 = pi18 ? n127 : ~n532;
  assign n64831 = pi17 ? n32 : n64830;
  assign n64832 = pi18 ? n8988 : ~n32;
  assign n64833 = pi17 ? n64832 : ~n2755;
  assign n64834 = pi16 ? n64831 : n64833;
  assign n64835 = pi18 ? n917 : ~n532;
  assign n64836 = pi17 ? n32 : n64835;
  assign n64837 = pi18 ? n31033 : ~n32;
  assign n64838 = pi17 ? n64837 : ~n2755;
  assign n64839 = pi16 ? n64836 : n64838;
  assign n64840 = pi15 ? n64834 : n64839;
  assign n64841 = pi14 ? n64829 : n64840;
  assign n64842 = pi13 ? n64821 : n64841;
  assign n64843 = pi12 ? n64807 : n64842;
  assign n64844 = pi11 ? n64799 : n64843;
  assign n64845 = pi10 ? n64759 : n64844;
  assign n64846 = pi09 ? n64725 : n64845;
  assign n64847 = pi19 ? n6727 : n28889;
  assign n64848 = pi20 ? n3523 : n5854;
  assign n64849 = pi19 ? n64848 : n9169;
  assign n64850 = pi18 ? n64847 : n64849;
  assign n64851 = pi17 ? n32 : n64850;
  assign n64852 = pi16 ? n32 : n64851;
  assign n64853 = pi15 ? n64711 : n64852;
  assign n64854 = pi14 ? n64707 : n64853;
  assign n64855 = pi13 ? n32 : n64854;
  assign n64856 = pi12 ? n32 : n64855;
  assign n64857 = pi11 ? n32 : n64856;
  assign n64858 = pi10 ? n32 : n64857;
  assign n64859 = pi19 ? n321 : ~n6042;
  assign n64860 = pi18 ? n32 : n64859;
  assign n64861 = pi17 ? n32 : n64860;
  assign n64862 = pi16 ? n32 : n64861;
  assign n64863 = pi15 ? n64862 : n50447;
  assign n64864 = pi14 ? n32 : n64863;
  assign n64865 = pi13 ? n24799 : n64864;
  assign n64866 = pi18 ? n49295 : n14892;
  assign n64867 = pi17 ? n32 : n64866;
  assign n64868 = pi16 ? n32 : n64867;
  assign n64869 = pi15 ? n50345 : n64868;
  assign n64870 = pi14 ? n27529 : n64869;
  assign n64871 = pi15 ? n27528 : n25044;
  assign n64872 = pi14 ? n64871 : n50357;
  assign n64873 = pi13 ? n64870 : n64872;
  assign n64874 = pi12 ? n64865 : n64873;
  assign n64875 = pi14 ? n16840 : n24370;
  assign n64876 = pi13 ? n64875 : n32;
  assign n64877 = pi15 ? n16606 : n16101;
  assign n64878 = pi19 ? n322 : ~n7468;
  assign n64879 = pi18 ? n863 : ~n64878;
  assign n64880 = pi17 ? n32 : n64879;
  assign n64881 = pi16 ? n32 : n64880;
  assign n64882 = pi15 ? n24712 : n64881;
  assign n64883 = pi14 ? n64877 : n64882;
  assign n64884 = pi17 ? n1807 : ~n2839;
  assign n64885 = pi16 ? n32 : n64884;
  assign n64886 = pi17 ? n1807 : ~n3763;
  assign n64887 = pi16 ? n32 : n64886;
  assign n64888 = pi15 ? n64885 : n64887;
  assign n64889 = pi17 ? n24786 : ~n2850;
  assign n64890 = pi16 ? n32 : n64889;
  assign n64891 = pi15 ? n7904 : n64890;
  assign n64892 = pi14 ? n64888 : n64891;
  assign n64893 = pi13 ? n64883 : n64892;
  assign n64894 = pi12 ? n64876 : n64893;
  assign n64895 = pi11 ? n64874 : n64894;
  assign n64896 = pi19 ? n343 : n2848;
  assign n64897 = pi18 ? n32 : n64896;
  assign n64898 = pi17 ? n1933 : ~n64897;
  assign n64899 = pi16 ? n32 : n64898;
  assign n64900 = pi20 ? n18762 : n321;
  assign n64901 = pi19 ? n32 : n64900;
  assign n64902 = pi18 ? n64901 : ~n32;
  assign n64903 = pi17 ? n64902 : ~n2850;
  assign n64904 = pi16 ? n32 : n64903;
  assign n64905 = pi15 ? n64899 : n64904;
  assign n64906 = pi17 ? n2531 : n51119;
  assign n64907 = pi16 ? n32 : n64906;
  assign n64908 = pi15 ? n64907 : n24829;
  assign n64909 = pi14 ? n64905 : n64908;
  assign n64910 = pi18 ? n21425 : n32;
  assign n64911 = pi17 ? n64910 : n16103;
  assign n64912 = pi16 ? n32 : n64911;
  assign n64913 = pi15 ? n64912 : n16319;
  assign n64914 = pi15 ? n23730 : n16108;
  assign n64915 = pi14 ? n64913 : n64914;
  assign n64916 = pi13 ? n64909 : n64915;
  assign n64917 = pi19 ? n349 : n53;
  assign n64918 = pi18 ? n50382 : n64917;
  assign n64919 = pi17 ? n32 : n64918;
  assign n64920 = pi16 ? n32 : n64919;
  assign n64921 = pi15 ? n50558 : n64920;
  assign n64922 = pi14 ? n24909 : n64921;
  assign n64923 = pi18 ? n36720 : n48634;
  assign n64924 = pi17 ? n32 : n64923;
  assign n64925 = pi16 ? n32 : n64924;
  assign n64926 = pi15 ? n64925 : n64786;
  assign n64927 = pi19 ? n813 : n358;
  assign n64928 = pi18 ? n36731 : n64927;
  assign n64929 = pi17 ? n32 : n64928;
  assign n64930 = pi16 ? n32 : n64929;
  assign n64931 = pi15 ? n64930 : n64795;
  assign n64932 = pi14 ? n64926 : n64931;
  assign n64933 = pi13 ? n64922 : n64932;
  assign n64934 = pi12 ? n64916 : n64933;
  assign n64935 = pi16 ? n31463 : n7724;
  assign n64936 = pi15 ? n64802 : n64935;
  assign n64937 = pi15 ? n50469 : n22540;
  assign n64938 = pi14 ? n64936 : n64937;
  assign n64939 = pi15 ? n22540 : n50281;
  assign n64940 = pi14 ? n64939 : n23179;
  assign n64941 = pi13 ? n64938 : n64940;
  assign n64942 = pi18 ? n19245 : n36827;
  assign n64943 = pi19 ? n36768 : n32;
  assign n64944 = pi20 ? n287 : ~n7880;
  assign n64945 = pi19 ? n64944 : ~n32;
  assign n64946 = pi18 ? n64943 : ~n64945;
  assign n64947 = pi17 ? n64942 : n64946;
  assign n64948 = pi16 ? n32 : n64947;
  assign n64949 = pi15 ? n64680 : n64948;
  assign n64950 = pi15 ? n64819 : n21928;
  assign n64951 = pi14 ? n64949 : n64950;
  assign n64952 = pi18 ? n16847 : ~n46501;
  assign n64953 = pi17 ? n64822 : ~n64952;
  assign n64954 = pi16 ? n1135 : ~n64953;
  assign n64955 = pi17 ? n31079 : n2517;
  assign n64956 = pi16 ? n19652 : ~n64955;
  assign n64957 = pi15 ? n64954 : n64956;
  assign n64958 = pi19 ? n322 : ~n1844;
  assign n64959 = pi18 ? n64958 : ~n32;
  assign n64960 = pi17 ? n64959 : ~n61145;
  assign n64961 = pi16 ? n64836 : n64960;
  assign n64962 = pi15 ? n64834 : n64961;
  assign n64963 = pi14 ? n64957 : n64962;
  assign n64964 = pi13 ? n64951 : n64963;
  assign n64965 = pi12 ? n64941 : n64964;
  assign n64966 = pi11 ? n64934 : n64965;
  assign n64967 = pi10 ? n64895 : n64966;
  assign n64968 = pi09 ? n64858 : n64967;
  assign n64969 = pi08 ? n64846 : n64968;
  assign n64970 = pi19 ? n1464 : n2297;
  assign n64971 = pi18 ? n940 : ~n64970;
  assign n64972 = pi17 ? n32 : n64971;
  assign n64973 = pi16 ? n32 : n64972;
  assign n64974 = pi15 ? n32 : n64973;
  assign n64975 = pi18 ? n880 : ~n1965;
  assign n64976 = pi17 ? n32 : n64975;
  assign n64977 = pi16 ? n32 : n64976;
  assign n64978 = pi15 ? n64977 : n32;
  assign n64979 = pi14 ? n64974 : n64978;
  assign n64980 = pi13 ? n32 : n64979;
  assign n64981 = pi12 ? n32 : n64980;
  assign n64982 = pi11 ? n32 : n64981;
  assign n64983 = pi10 ? n32 : n64982;
  assign n64984 = pi15 ? n16973 : n36851;
  assign n64985 = pi14 ? n25138 : n64984;
  assign n64986 = pi15 ? n64728 : n50505;
  assign n64987 = pi14 ? n40800 : n64986;
  assign n64988 = pi13 ? n64985 : n64987;
  assign n64989 = pi12 ? n64988 : n50522;
  assign n64990 = pi15 ? n16837 : n16606;
  assign n64991 = pi14 ? n64990 : n24627;
  assign n64992 = pi13 ? n64991 : n32;
  assign n64993 = pi15 ? n32 : n16101;
  assign n64994 = pi18 ? n344 : ~n2835;
  assign n64995 = pi17 ? n32 : n64994;
  assign n64996 = pi16 ? n32 : n64995;
  assign n64997 = pi15 ? n16298 : n64996;
  assign n64998 = pi14 ? n64993 : n64997;
  assign n64999 = pi17 ? n1933 : ~n2839;
  assign n65000 = pi16 ? n32 : n64999;
  assign n65001 = pi15 ? n65000 : n64885;
  assign n65002 = pi18 ? n32 : n23543;
  assign n65003 = pi17 ? n65002 : ~n2850;
  assign n65004 = pi16 ? n32 : n65003;
  assign n65005 = pi15 ? n7904 : n65004;
  assign n65006 = pi14 ? n65001 : n65005;
  assign n65007 = pi13 ? n64998 : n65006;
  assign n65008 = pi12 ? n64992 : n65007;
  assign n65009 = pi11 ? n64989 : n65008;
  assign n65010 = pi19 ? n4406 : n349;
  assign n65011 = pi18 ? n36879 : n65010;
  assign n65012 = pi17 ? n1933 : ~n65011;
  assign n65013 = pi16 ? n32 : n65012;
  assign n65014 = pi18 ? n6071 : n350;
  assign n65015 = pi17 ? n65014 : ~n3067;
  assign n65016 = pi16 ? n32 : n65015;
  assign n65017 = pi15 ? n65013 : n65016;
  assign n65018 = pi15 ? n64907 : n24289;
  assign n65019 = pi14 ? n65017 : n65018;
  assign n65020 = pi19 ? n32 : n8044;
  assign n65021 = pi18 ? n65020 : n32;
  assign n65022 = pi17 ? n65021 : n16103;
  assign n65023 = pi16 ? n32 : n65022;
  assign n65024 = pi18 ? n28579 : n32;
  assign n65025 = pi17 ? n65024 : n16103;
  assign n65026 = pi16 ? n32 : n65025;
  assign n65027 = pi15 ? n65023 : n65026;
  assign n65028 = pi15 ? n24905 : n16108;
  assign n65029 = pi14 ? n65027 : n65028;
  assign n65030 = pi13 ? n65019 : n65029;
  assign n65031 = pi19 ? n32 : ~n56769;
  assign n65032 = pi18 ? n32 : n65031;
  assign n65033 = pi17 ? n32 : n65032;
  assign n65034 = pi16 ? n32 : n65033;
  assign n65035 = pi15 ? n16108 : n65034;
  assign n65036 = pi19 ? n1757 : ~n53;
  assign n65037 = pi18 ? n50559 : ~n65036;
  assign n65038 = pi17 ? n32 : n65037;
  assign n65039 = pi16 ? n32 : n65038;
  assign n65040 = pi15 ? n50558 : n65039;
  assign n65041 = pi14 ? n65035 : n65040;
  assign n65042 = pi19 ? n358 : n1941;
  assign n65043 = pi18 ? n36911 : ~n65042;
  assign n65044 = pi17 ? n32 : n65043;
  assign n65045 = pi16 ? n32 : n65044;
  assign n65046 = pi18 ? n36917 : ~n37418;
  assign n65047 = pi17 ? n32 : n65046;
  assign n65048 = pi16 ? n32 : n65047;
  assign n65049 = pi15 ? n65045 : n65048;
  assign n65050 = pi19 ? n343 : ~n40268;
  assign n65051 = pi18 ? n15844 : n65050;
  assign n65052 = pi17 ? n32 : n65051;
  assign n65053 = pi16 ? n32 : n65052;
  assign n65054 = pi18 ? n15844 : n24015;
  assign n65055 = pi17 ? n32 : n65054;
  assign n65056 = pi16 ? n32 : n65055;
  assign n65057 = pi15 ? n65053 : n65056;
  assign n65058 = pi14 ? n65049 : n65057;
  assign n65059 = pi13 ? n65041 : n65058;
  assign n65060 = pi12 ? n65030 : n65059;
  assign n65061 = pi19 ? n343 : n5635;
  assign n65062 = pi18 ? n15844 : n65061;
  assign n65063 = pi17 ? n32 : n65062;
  assign n65064 = pi16 ? n31463 : n65063;
  assign n65065 = pi15 ? n65064 : n7725;
  assign n65066 = pi14 ? n65065 : n50586;
  assign n65067 = pi17 ? n28638 : n22538;
  assign n65068 = pi16 ? n32 : n65067;
  assign n65069 = pi14 ? n65068 : n22347;
  assign n65070 = pi13 ? n65066 : n65069;
  assign n65071 = pi17 ? n28638 : n22345;
  assign n65072 = pi16 ? n32 : n65071;
  assign n65073 = pi20 ? n246 : n10878;
  assign n65074 = pi19 ? n65073 : n32;
  assign n65075 = pi18 ? n32 : n65074;
  assign n65076 = pi17 ? n36944 : ~n65075;
  assign n65077 = pi16 ? n1233 : ~n65076;
  assign n65078 = pi15 ? n65072 : n65077;
  assign n65079 = pi18 ? n13080 : n20020;
  assign n65080 = pi17 ? n32 : ~n65079;
  assign n65081 = pi16 ? n1233 : ~n65080;
  assign n65082 = pi15 ? n65081 : n21853;
  assign n65083 = pi14 ? n65078 : n65082;
  assign n65084 = pi20 ? n246 : n20265;
  assign n65085 = pi19 ? n65084 : ~n32;
  assign n65086 = pi18 ? n36955 : n65085;
  assign n65087 = pi17 ? n64822 : n65086;
  assign n65088 = pi16 ? n1233 : ~n65087;
  assign n65089 = pi17 ? n36960 : n2517;
  assign n65090 = pi16 ? n1233 : ~n65089;
  assign n65091 = pi15 ? n65088 : n65090;
  assign n65092 = pi17 ? n64832 : ~n2517;
  assign n65093 = pi16 ? n64831 : n65092;
  assign n65094 = pi18 ? n268 : ~n532;
  assign n65095 = pi17 ? n32 : n65094;
  assign n65096 = pi19 ? n322 : ~n266;
  assign n65097 = pi18 ? n65096 : ~n32;
  assign n65098 = pi17 ? n65097 : ~n61145;
  assign n65099 = pi16 ? n65095 : n65098;
  assign n65100 = pi15 ? n65093 : n65099;
  assign n65101 = pi14 ? n65091 : n65100;
  assign n65102 = pi13 ? n65083 : n65101;
  assign n65103 = pi12 ? n65070 : n65102;
  assign n65104 = pi11 ? n65060 : n65103;
  assign n65105 = pi10 ? n65009 : n65104;
  assign n65106 = pi09 ? n64983 : n65105;
  assign n65107 = pi18 ? n880 : ~n2962;
  assign n65108 = pi17 ? n32 : n65107;
  assign n65109 = pi16 ? n32 : n65108;
  assign n65110 = pi15 ? n65109 : n32;
  assign n65111 = pi14 ? n64974 : n65110;
  assign n65112 = pi13 ? n32 : n65111;
  assign n65113 = pi12 ? n32 : n65112;
  assign n65114 = pi11 ? n32 : n65113;
  assign n65115 = pi10 ? n32 : n65114;
  assign n65116 = pi19 ? n321 : ~n22911;
  assign n65117 = pi18 ? n32 : n65116;
  assign n65118 = pi17 ? n32 : n65117;
  assign n65119 = pi16 ? n32 : n65118;
  assign n65120 = pi15 ? n65119 : n50631;
  assign n65121 = pi14 ? n32 : n65120;
  assign n65122 = pi13 ? n16974 : n65121;
  assign n65123 = pi15 ? n50513 : n14909;
  assign n65124 = pi14 ? n50639 : n65123;
  assign n65125 = pi13 ? n65124 : n50521;
  assign n65126 = pi12 ? n65122 : n65125;
  assign n65127 = pi14 ? n24799 : n24627;
  assign n65128 = pi13 ? n65127 : n32;
  assign n65129 = pi15 ? n16298 : n10084;
  assign n65130 = pi14 ? n64993 : n65129;
  assign n65131 = pi17 ? n1933 : ~n2836;
  assign n65132 = pi16 ? n32 : n65131;
  assign n65133 = pi15 ? n65132 : n64885;
  assign n65134 = pi17 ? n65002 : ~n2839;
  assign n65135 = pi16 ? n32 : n65134;
  assign n65136 = pi15 ? n64885 : n65135;
  assign n65137 = pi14 ? n65133 : n65136;
  assign n65138 = pi13 ? n65130 : n65137;
  assign n65139 = pi12 ? n65128 : n65138;
  assign n65140 = pi11 ? n65126 : n65139;
  assign n65141 = pi19 ? n4406 : n589;
  assign n65142 = pi18 ? n36879 : n65141;
  assign n65143 = pi17 ? n1933 : ~n65142;
  assign n65144 = pi16 ? n32 : n65143;
  assign n65145 = pi17 ? n65014 : ~n2839;
  assign n65146 = pi16 ? n32 : n65145;
  assign n65147 = pi15 ? n65144 : n65146;
  assign n65148 = pi18 ? n350 : ~n590;
  assign n65149 = pi17 ? n2531 : n65148;
  assign n65150 = pi16 ? n32 : n65149;
  assign n65151 = pi15 ? n65150 : n16105;
  assign n65152 = pi14 ? n65147 : n65151;
  assign n65153 = pi17 ? n65021 : n24287;
  assign n65154 = pi16 ? n32 : n65153;
  assign n65155 = pi17 ? n28638 : n16103;
  assign n65156 = pi16 ? n32 : n65155;
  assign n65157 = pi15 ? n65154 : n65156;
  assign n65158 = pi14 ? n65157 : n48969;
  assign n65159 = pi13 ? n65152 : n65158;
  assign n65160 = pi19 ? n349 : n5614;
  assign n65161 = pi18 ? n20020 : n65160;
  assign n65162 = pi17 ? n32 : n65161;
  assign n65163 = pi16 ? n32 : n65162;
  assign n65164 = pi15 ? n65163 : n50562;
  assign n65165 = pi14 ? n48385 : n65164;
  assign n65166 = pi19 ? n358 : n236;
  assign n65167 = pi18 ? n36911 : ~n65166;
  assign n65168 = pi17 ? n32 : n65167;
  assign n65169 = pi16 ? n32 : n65168;
  assign n65170 = pi19 ? n4342 : n1941;
  assign n65171 = pi18 ? n36917 : ~n65170;
  assign n65172 = pi17 ? n32 : n65171;
  assign n65173 = pi16 ? n32 : n65172;
  assign n65174 = pi15 ? n65169 : n65173;
  assign n65175 = pi18 ? n15844 : n23833;
  assign n65176 = pi17 ? n32 : n65175;
  assign n65177 = pi16 ? n32 : n65176;
  assign n65178 = pi15 ? n65056 : n65177;
  assign n65179 = pi14 ? n65174 : n65178;
  assign n65180 = pi13 ? n65165 : n65179;
  assign n65181 = pi12 ? n65159 : n65180;
  assign n65182 = pi16 ? n31463 : n50579;
  assign n65183 = pi17 ? n1807 : ~n2855;
  assign n65184 = pi16 ? n32 : n65183;
  assign n65185 = pi15 ? n65182 : n65184;
  assign n65186 = pi17 ? n36981 : n1107;
  assign n65187 = pi16 ? n32 : n65186;
  assign n65188 = pi15 ? n50583 : n65187;
  assign n65189 = pi14 ? n65185 : n65188;
  assign n65190 = pi14 ? n65068 : n22829;
  assign n65191 = pi13 ? n65189 : n65190;
  assign n65192 = pi17 ? n28638 : n15121;
  assign n65193 = pi16 ? n32 : n65192;
  assign n65194 = pi20 ? n246 : n7839;
  assign n65195 = pi19 ? n65194 : n32;
  assign n65196 = pi18 ? n32 : n65195;
  assign n65197 = pi17 ? n37006 : ~n65196;
  assign n65198 = pi16 ? n1233 : ~n65197;
  assign n65199 = pi15 ? n65193 : n65198;
  assign n65200 = pi18 ? n13080 : n14787;
  assign n65201 = pi17 ? n32 : ~n65200;
  assign n65202 = pi16 ? n1233 : ~n65201;
  assign n65203 = pi15 ? n65202 : n21853;
  assign n65204 = pi14 ? n65199 : n65203;
  assign n65205 = pi17 ? n37014 : n2517;
  assign n65206 = pi16 ? n1233 : ~n65205;
  assign n65207 = pi15 ? n65088 : n65206;
  assign n65208 = pi16 ? n12787 : n65092;
  assign n65209 = pi19 ? n322 : ~n17769;
  assign n65210 = pi18 ? n65209 : ~n32;
  assign n65211 = pi19 ? n1378 : ~n32;
  assign n65212 = pi18 ? n32 : n65211;
  assign n65213 = pi17 ? n65210 : ~n65212;
  assign n65214 = pi16 ? n65095 : n65213;
  assign n65215 = pi15 ? n65208 : n65214;
  assign n65216 = pi14 ? n65207 : n65215;
  assign n65217 = pi13 ? n65204 : n65216;
  assign n65218 = pi12 ? n65191 : n65217;
  assign n65219 = pi11 ? n65181 : n65218;
  assign n65220 = pi10 ? n65140 : n65219;
  assign n65221 = pi09 ? n65115 : n65220;
  assign n65222 = pi08 ? n65106 : n65221;
  assign n65223 = pi07 ? n64969 : n65222;
  assign n65224 = pi15 ? n32 : n11463;
  assign n65225 = pi20 ? n357 : n206;
  assign n65226 = pi19 ? n65225 : ~n429;
  assign n65227 = pi18 ? n863 : n65226;
  assign n65228 = pi17 ? n32 : n65227;
  assign n65229 = pi16 ? n32 : n65228;
  assign n65230 = pi15 ? n65229 : n32;
  assign n65231 = pi14 ? n65224 : n65230;
  assign n65232 = pi13 ? n32 : n65231;
  assign n65233 = pi12 ? n32 : n65232;
  assign n65234 = pi11 ? n32 : n65233;
  assign n65235 = pi10 ? n32 : n65234;
  assign n65236 = pi14 ? n25133 : n26164;
  assign n65237 = pi14 ? n24962 : n27071;
  assign n65238 = pi13 ? n65236 : n65237;
  assign n65239 = pi14 ? n52240 : n50737;
  assign n65240 = pi13 ? n50729 : n65239;
  assign n65241 = pi12 ? n65238 : n65240;
  assign n65242 = pi13 ? n50313 : n32;
  assign n65243 = pi15 ? n16101 : n9121;
  assign n65244 = pi14 ? n25452 : n65243;
  assign n65245 = pi17 ? n2750 : ~n2836;
  assign n65246 = pi16 ? n32 : n65245;
  assign n65247 = pi17 ? n3067 : ~n2839;
  assign n65248 = pi16 ? n32 : n65247;
  assign n65249 = pi15 ? n65246 : n65248;
  assign n65250 = pi17 ? n2519 : ~n2839;
  assign n65251 = pi16 ? n32 : n65250;
  assign n65252 = pi19 ? n4126 : n589;
  assign n65253 = pi18 ? n32 : n65252;
  assign n65254 = pi17 ? n3067 : ~n65253;
  assign n65255 = pi16 ? n32 : n65254;
  assign n65256 = pi15 ? n65251 : n65255;
  assign n65257 = pi14 ? n65249 : n65256;
  assign n65258 = pi13 ? n65244 : n65257;
  assign n65259 = pi12 ? n65242 : n65258;
  assign n65260 = pi11 ? n65241 : n65259;
  assign n65261 = pi19 ? n32 : n31647;
  assign n65262 = pi19 ? n5004 : ~n9724;
  assign n65263 = pi18 ? n65261 : n65262;
  assign n65264 = pi17 ? n32 : ~n65263;
  assign n65265 = pi16 ? n32 : n65264;
  assign n65266 = pi18 ? n32 : n31033;
  assign n65267 = pi19 ? n9007 : ~n9724;
  assign n65268 = pi18 ? n20164 : n65267;
  assign n65269 = pi17 ? n65266 : ~n65268;
  assign n65270 = pi16 ? n32 : n65269;
  assign n65271 = pi15 ? n65265 : n65270;
  assign n65272 = pi15 ? n25066 : n32;
  assign n65273 = pi14 ? n65271 : n65272;
  assign n65274 = pi17 ? n17901 : n3243;
  assign n65275 = pi16 ? n32 : n65274;
  assign n65276 = pi15 ? n65275 : n25070;
  assign n65277 = pi14 ? n65276 : n63598;
  assign n65278 = pi13 ? n65273 : n65277;
  assign n65279 = pi18 ? n34208 : ~n8259;
  assign n65280 = pi17 ? n32 : n65279;
  assign n65281 = pi16 ? n32 : n65280;
  assign n65282 = pi15 ? n12056 : n65281;
  assign n65283 = pi14 ? n26656 : n65282;
  assign n65284 = pi18 ? n702 : ~n2730;
  assign n65285 = pi17 ? n32 : n65284;
  assign n65286 = pi16 ? n32 : n65285;
  assign n65287 = pi15 ? n50789 : n65286;
  assign n65288 = pi18 ? n9346 : ~n2730;
  assign n65289 = pi17 ? n32 : n65288;
  assign n65290 = pi16 ? n32 : n65289;
  assign n65291 = pi18 ? n7038 : n6132;
  assign n65292 = pi17 ? n32 : n65291;
  assign n65293 = pi16 ? n1059 : n65292;
  assign n65294 = pi15 ? n65290 : n65293;
  assign n65295 = pi14 ? n65287 : n65294;
  assign n65296 = pi13 ? n65283 : n65295;
  assign n65297 = pi12 ? n65278 : n65296;
  assign n65298 = pi17 ? n32 : n50808;
  assign n65299 = pi16 ? n1014 : n65298;
  assign n65300 = pi17 ? n35572 : ~n2855;
  assign n65301 = pi16 ? n32 : n65300;
  assign n65302 = pi15 ? n65299 : n65301;
  assign n65303 = pi14 ? n65302 : n48800;
  assign n65304 = pi17 ? n50815 : n1107;
  assign n65305 = pi16 ? n32 : n65304;
  assign n65306 = pi19 ? n19306 : n32;
  assign n65307 = pi18 ? n16981 : n65306;
  assign n65308 = pi17 ? n65307 : n32;
  assign n65309 = pi16 ? n32 : n65308;
  assign n65310 = pi15 ? n65305 : n65309;
  assign n65311 = pi14 ? n65310 : n33897;
  assign n65312 = pi13 ? n65303 : n65311;
  assign n65313 = pi17 ? n50815 : n22345;
  assign n65314 = pi16 ? n32 : n65313;
  assign n65315 = pi17 ? n36742 : ~n1787;
  assign n65316 = pi16 ? n1233 : ~n65315;
  assign n65317 = pi15 ? n65314 : n65316;
  assign n65318 = pi18 ? n605 : ~n645;
  assign n65319 = pi17 ? n32 : n65318;
  assign n65320 = pi16 ? n1233 : ~n65319;
  assign n65321 = pi16 ? n12897 : n33568;
  assign n65322 = pi15 ? n65320 : n65321;
  assign n65323 = pi14 ? n65317 : n65322;
  assign n65324 = pi18 ? n50825 : ~n508;
  assign n65325 = pi17 ? n35126 : ~n65324;
  assign n65326 = pi16 ? n18981 : ~n65325;
  assign n65327 = pi17 ? n19071 : n2748;
  assign n65328 = pi16 ? n2958 : ~n65327;
  assign n65329 = pi15 ? n65326 : n65328;
  assign n65330 = pi20 ? n32 : n54153;
  assign n65331 = pi19 ? n65330 : ~n32;
  assign n65332 = pi18 ? n32 : n65331;
  assign n65333 = pi17 ? n1470 : ~n65332;
  assign n65334 = pi16 ? n882 : n65333;
  assign n65335 = pi18 ? n940 : ~n4689;
  assign n65336 = pi17 ? n65335 : ~n2517;
  assign n65337 = pi16 ? n32 : n65336;
  assign n65338 = pi15 ? n65334 : n65337;
  assign n65339 = pi14 ? n65329 : n65338;
  assign n65340 = pi13 ? n65323 : n65339;
  assign n65341 = pi12 ? n65312 : n65340;
  assign n65342 = pi11 ? n65297 : n65341;
  assign n65343 = pi10 ? n65260 : n65342;
  assign n65344 = pi09 ? n65235 : n65343;
  assign n65345 = pi15 ? n50943 : n15847;
  assign n65346 = pi14 ? n26163 : n65345;
  assign n65347 = pi13 ? n25133 : n65346;
  assign n65348 = pi15 ? n16837 : n15847;
  assign n65349 = pi19 ? n5694 : n2297;
  assign n65350 = pi18 ? n50723 : ~n65349;
  assign n65351 = pi17 ? n32 : n65350;
  assign n65352 = pi16 ? n32 : n65351;
  assign n65353 = pi15 ? n15403 : n65352;
  assign n65354 = pi14 ? n65348 : n65353;
  assign n65355 = pi14 ? n52240 : n32;
  assign n65356 = pi13 ? n65354 : n65355;
  assign n65357 = pi12 ? n65347 : n65356;
  assign n65358 = pi14 ? n16974 : n16837;
  assign n65359 = pi14 ? n24627 : n16840;
  assign n65360 = pi13 ? n65358 : n65359;
  assign n65361 = pi17 ? n3067 : ~n2831;
  assign n65362 = pi16 ? n32 : n65361;
  assign n65363 = pi15 ? n25044 : n65362;
  assign n65364 = pi14 ? n25452 : n65363;
  assign n65365 = pi17 ? n3067 : ~n2836;
  assign n65366 = pi16 ? n32 : n65365;
  assign n65367 = pi15 ? n7570 : n65366;
  assign n65368 = pi17 ? n2519 : ~n2836;
  assign n65369 = pi16 ? n32 : n65368;
  assign n65370 = pi19 ? n4126 : n2317;
  assign n65371 = pi18 ? n32 : n65370;
  assign n65372 = pi17 ? n3067 : ~n65371;
  assign n65373 = pi16 ? n32 : n65372;
  assign n65374 = pi15 ? n65369 : n65373;
  assign n65375 = pi14 ? n65367 : n65374;
  assign n65376 = pi13 ? n65364 : n65375;
  assign n65377 = pi12 ? n65360 : n65376;
  assign n65378 = pi11 ? n65357 : n65377;
  assign n65379 = pi19 ? n5004 : ~n7468;
  assign n65380 = pi18 ? n65261 : n65379;
  assign n65381 = pi17 ? n32 : ~n65380;
  assign n65382 = pi16 ? n32 : n65381;
  assign n65383 = pi19 ? n9007 : ~n7468;
  assign n65384 = pi18 ? n20164 : n65383;
  assign n65385 = pi17 ? n65266 : ~n65384;
  assign n65386 = pi16 ? n32 : n65385;
  assign n65387 = pi15 ? n65382 : n65386;
  assign n65388 = pi14 ? n65387 : n25165;
  assign n65389 = pi17 ? n17901 : n3497;
  assign n65390 = pi16 ? n32 : n65389;
  assign n65391 = pi15 ? n65390 : n16377;
  assign n65392 = pi14 ? n65391 : n26367;
  assign n65393 = pi13 ? n65388 : n65392;
  assign n65394 = pi15 ? n23933 : n24388;
  assign n65395 = pi18 ? n496 : ~n64269;
  assign n65396 = pi17 ? n32 : n65395;
  assign n65397 = pi16 ? n32 : n65396;
  assign n65398 = pi15 ? n65397 : n65281;
  assign n65399 = pi14 ? n65394 : n65398;
  assign n65400 = pi18 ? n702 : ~n962;
  assign n65401 = pi17 ? n32 : n65400;
  assign n65402 = pi16 ? n32 : n65401;
  assign n65403 = pi15 ? n50789 : n65402;
  assign n65404 = pi16 ? n11695 : n65292;
  assign n65405 = pi15 ? n65290 : n65404;
  assign n65406 = pi14 ? n65403 : n65405;
  assign n65407 = pi13 ? n65399 : n65406;
  assign n65408 = pi12 ? n65393 : n65407;
  assign n65409 = pi16 ? n32 : n65298;
  assign n65410 = pi17 ? n35572 : ~n2616;
  assign n65411 = pi16 ? n32 : n65410;
  assign n65412 = pi15 ? n65409 : n65411;
  assign n65413 = pi15 ? n22923 : n21853;
  assign n65414 = pi14 ? n65412 : n65413;
  assign n65415 = pi18 ? n16981 : n13945;
  assign n65416 = pi17 ? n65415 : n32;
  assign n65417 = pi16 ? n32 : n65416;
  assign n65418 = pi15 ? n50589 : n65417;
  assign n65419 = pi15 ? n22728 : n22733;
  assign n65420 = pi14 ? n65418 : n65419;
  assign n65421 = pi13 ? n65414 : n65420;
  assign n65422 = pi17 ? n37203 : ~n32;
  assign n65423 = pi16 ? n1705 : ~n65422;
  assign n65424 = pi15 ? n65072 : n65423;
  assign n65425 = pi18 ? n605 : ~n8106;
  assign n65426 = pi17 ? n32 : n65425;
  assign n65427 = pi16 ? n1972 : ~n65426;
  assign n65428 = pi20 ? n32 : ~n16008;
  assign n65429 = pi19 ? n65428 : n32;
  assign n65430 = pi18 ? n268 : n65429;
  assign n65431 = pi17 ? n32 : n65430;
  assign n65432 = pi16 ? n12897 : n65431;
  assign n65433 = pi15 ? n65427 : n65432;
  assign n65434 = pi14 ? n65424 : n65433;
  assign n65435 = pi18 ? n1477 : ~n16389;
  assign n65436 = pi17 ? n32 : n65435;
  assign n65437 = pi16 ? n65436 : ~n65325;
  assign n65438 = pi15 ? n65437 : n65328;
  assign n65439 = pi17 ? n1470 : ~n2748;
  assign n65440 = pi16 ? n11454 : n65439;
  assign n65441 = pi18 ? n940 : ~n248;
  assign n65442 = pi17 ? n65441 : ~n2748;
  assign n65443 = pi16 ? n32 : n65442;
  assign n65444 = pi15 ? n65440 : n65443;
  assign n65445 = pi14 ? n65438 : n65444;
  assign n65446 = pi13 ? n65434 : n65445;
  assign n65447 = pi12 ? n65421 : n65446;
  assign n65448 = pi11 ? n65408 : n65447;
  assign n65449 = pi10 ? n65378 : n65448;
  assign n65450 = pi09 ? n65235 : n65449;
  assign n65451 = pi08 ? n65344 : n65450;
  assign n65452 = pi18 ? n12368 : ~n880;
  assign n65453 = pi17 ? n32 : n65452;
  assign n65454 = pi16 ? n32 : n65453;
  assign n65455 = pi15 ? n32 : n65454;
  assign n65456 = pi14 ? n65455 : n17273;
  assign n65457 = pi13 ? n32 : n65456;
  assign n65458 = pi12 ? n32 : n65457;
  assign n65459 = pi11 ? n32 : n65458;
  assign n65460 = pi10 ? n32 : n65459;
  assign n65461 = pi14 ? n25133 : n17070;
  assign n65462 = pi14 ? n26163 : n50944;
  assign n65463 = pi13 ? n65461 : n65462;
  assign n65464 = pi19 ? n507 : n4342;
  assign n65465 = pi18 ? n32 : n65464;
  assign n65466 = pi17 ? n32 : n65465;
  assign n65467 = pi16 ? n32 : n65466;
  assign n65468 = pi15 ? n22817 : n65467;
  assign n65469 = pi19 ? n50956 : ~n11561;
  assign n65470 = pi18 ? n32 : n65469;
  assign n65471 = pi17 ? n32 : n65470;
  assign n65472 = pi16 ? n32 : n65471;
  assign n65473 = pi15 ? n51091 : n65472;
  assign n65474 = pi14 ? n65468 : n65473;
  assign n65475 = pi19 ? n6398 : ~n11561;
  assign n65476 = pi18 ? n32 : n65475;
  assign n65477 = pi17 ? n32 : n65476;
  assign n65478 = pi16 ? n32 : n65477;
  assign n65479 = pi15 ? n65478 : n15403;
  assign n65480 = pi14 ? n65479 : n16974;
  assign n65481 = pi13 ? n65474 : n65480;
  assign n65482 = pi12 ? n65463 : n65481;
  assign n65483 = pi13 ? n25036 : n32;
  assign n65484 = pi18 ? n63034 : ~n2830;
  assign n65485 = pi17 ? n2959 : n65484;
  assign n65486 = pi16 ? n32 : n65485;
  assign n65487 = pi15 ? n65486 : n65362;
  assign n65488 = pi14 ? n24874 : n65487;
  assign n65489 = pi15 ? n8598 : n65248;
  assign n65490 = pi19 ? n32 : n14552;
  assign n65491 = pi18 ? n32 : n65490;
  assign n65492 = pi17 ? n2750 : ~n65491;
  assign n65493 = pi16 ? n32 : n65492;
  assign n65494 = pi19 ? n22525 : n14552;
  assign n65495 = pi18 ? n32 : n65494;
  assign n65496 = pi17 ? n3067 : ~n65495;
  assign n65497 = pi16 ? n32 : n65496;
  assign n65498 = pi15 ? n65493 : n65497;
  assign n65499 = pi14 ? n65489 : n65498;
  assign n65500 = pi13 ? n65488 : n65499;
  assign n65501 = pi12 ? n65483 : n65500;
  assign n65502 = pi11 ? n65482 : n65501;
  assign n65503 = pi19 ? n507 : n22864;
  assign n65504 = pi18 ? n32 : n65503;
  assign n65505 = pi19 ? n4670 : n589;
  assign n65506 = pi18 ? n32 : n65505;
  assign n65507 = pi17 ? n65504 : ~n65506;
  assign n65508 = pi16 ? n32 : n65507;
  assign n65509 = pi18 ? n32 : n64958;
  assign n65510 = pi18 ? n20164 : n2835;
  assign n65511 = pi17 ? n65509 : ~n65510;
  assign n65512 = pi16 ? n32 : n65511;
  assign n65513 = pi15 ? n65508 : n65512;
  assign n65514 = pi14 ? n65513 : n24430;
  assign n65515 = pi17 ? n18395 : n3497;
  assign n65516 = pi16 ? n32 : n65515;
  assign n65517 = pi15 ? n65516 : n24237;
  assign n65518 = pi14 ? n65517 : n25726;
  assign n65519 = pi13 ? n65514 : n65518;
  assign n65520 = pi18 ? n34208 : ~n64269;
  assign n65521 = pi17 ? n32 : n65520;
  assign n65522 = pi16 ? n32 : n65521;
  assign n65523 = pi15 ? n51136 : n65522;
  assign n65524 = pi14 ? n37282 : n65523;
  assign n65525 = pi18 ? n684 : ~n962;
  assign n65526 = pi17 ? n32 : n65525;
  assign n65527 = pi16 ? n32 : n65526;
  assign n65528 = pi20 ? n9641 : n266;
  assign n65529 = pi19 ? n65528 : n32;
  assign n65530 = pi18 ? n32 : n65529;
  assign n65531 = pi18 ? n37293 : ~n967;
  assign n65532 = pi17 ? n65530 : n65531;
  assign n65533 = pi16 ? n32 : n65532;
  assign n65534 = pi15 ? n65527 : n65533;
  assign n65535 = pi18 ? n880 : ~n2730;
  assign n65536 = pi17 ? n32 : n65535;
  assign n65537 = pi16 ? n32 : n65536;
  assign n65538 = pi18 ? n7038 : n37589;
  assign n65539 = pi17 ? n32 : n65538;
  assign n65540 = pi16 ? n11692 : n65539;
  assign n65541 = pi15 ? n65537 : n65540;
  assign n65542 = pi14 ? n65534 : n65541;
  assign n65543 = pi13 ? n65524 : n65542;
  assign n65544 = pi12 ? n65519 : n65543;
  assign n65545 = pi17 ? n32 : n51015;
  assign n65546 = pi16 ? n32 : n65545;
  assign n65547 = pi18 ? n32 : n64316;
  assign n65548 = pi17 ? n2750 : ~n65547;
  assign n65549 = pi16 ? n32 : n65548;
  assign n65550 = pi15 ? n65546 : n65549;
  assign n65551 = pi21 ? n32 : ~n8275;
  assign n65552 = pi20 ? n32 : n65551;
  assign n65553 = pi19 ? n65552 : ~n617;
  assign n65554 = pi18 ? n32 : n65553;
  assign n65555 = pi17 ? n32 : n65554;
  assign n65556 = pi16 ? n32 : n65555;
  assign n65557 = pi15 ? n15123 : n65556;
  assign n65558 = pi14 ? n65550 : n65557;
  assign n65559 = pi17 ? n28818 : n1542;
  assign n65560 = pi16 ? n32 : n65559;
  assign n65561 = pi18 ? n32 : n65306;
  assign n65562 = pi17 ? n65561 : n62532;
  assign n65563 = pi16 ? n32 : n65562;
  assign n65564 = pi15 ? n65560 : n65563;
  assign n65565 = pi14 ? n65564 : n24533;
  assign n65566 = pi13 ? n65558 : n65565;
  assign n65567 = pi17 ? n28818 : n2080;
  assign n65568 = pi16 ? n32 : n65567;
  assign n65569 = pi17 ? n37337 : ~n22345;
  assign n65570 = pi16 ? n1323 : ~n65569;
  assign n65571 = pi15 ? n65568 : n65570;
  assign n65572 = pi19 ? n12821 : ~n32;
  assign n65573 = pi18 ? n323 : n65572;
  assign n65574 = pi17 ? n32 : n65573;
  assign n65575 = pi16 ? n1594 : ~n65574;
  assign n65576 = pi18 ? n22885 : n4983;
  assign n65577 = pi17 ? n32 : n65576;
  assign n65578 = pi16 ? n11886 : n65577;
  assign n65579 = pi15 ? n65575 : n65578;
  assign n65580 = pi14 ? n65571 : n65579;
  assign n65581 = pi18 ? n20193 : n22752;
  assign n65582 = pi17 ? n35126 : ~n65581;
  assign n65583 = pi16 ? n1577 : ~n65582;
  assign n65584 = pi17 ? n19071 : n2512;
  assign n65585 = pi16 ? n2958 : ~n65584;
  assign n65586 = pi15 ? n65583 : n65585;
  assign n65587 = pi18 ? n940 : ~n6145;
  assign n65588 = pi18 ? n32 : n62696;
  assign n65589 = pi17 ? n65587 : ~n65588;
  assign n65590 = pi16 ? n11684 : n65589;
  assign n65591 = pi18 ? n940 : ~n34142;
  assign n65592 = pi17 ? n65591 : ~n2748;
  assign n65593 = pi16 ? n32 : n65592;
  assign n65594 = pi15 ? n65590 : n65593;
  assign n65595 = pi14 ? n65586 : n65594;
  assign n65596 = pi13 ? n65580 : n65595;
  assign n65597 = pi12 ? n65566 : n65596;
  assign n65598 = pi11 ? n65544 : n65597;
  assign n65599 = pi10 ? n65502 : n65598;
  assign n65600 = pi09 ? n65460 : n65599;
  assign n65601 = pi14 ? n17273 : n51076;
  assign n65602 = pi13 ? n65461 : n65601;
  assign n65603 = pi19 ? n507 : n13376;
  assign n65604 = pi18 ? n32 : n65603;
  assign n65605 = pi17 ? n32 : n65604;
  assign n65606 = pi16 ? n32 : n65605;
  assign n65607 = pi15 ? n51082 : n65606;
  assign n65608 = pi20 ? n266 : n141;
  assign n65609 = pi19 ? n50951 : ~n65608;
  assign n65610 = pi18 ? n1819 : n65609;
  assign n65611 = pi17 ? n32 : n65610;
  assign n65612 = pi16 ? n32 : n65611;
  assign n65613 = pi15 ? n65612 : n51095;
  assign n65614 = pi14 ? n65607 : n65613;
  assign n65615 = pi13 ? n65614 : n51103;
  assign n65616 = pi12 ? n65602 : n65615;
  assign n65617 = pi14 ? n25133 : n16973;
  assign n65618 = pi13 ? n65617 : n32;
  assign n65619 = pi18 ? n63034 : ~n1965;
  assign n65620 = pi17 ? n2959 : n65619;
  assign n65621 = pi16 ? n32 : n65620;
  assign n65622 = pi17 ? n3067 : ~n3182;
  assign n65623 = pi16 ? n32 : n65622;
  assign n65624 = pi15 ? n65621 : n65623;
  assign n65625 = pi14 ? n24874 : n65624;
  assign n65626 = pi15 ? n8598 : n9121;
  assign n65627 = pi17 ? n2750 : ~n8639;
  assign n65628 = pi16 ? n32 : n65627;
  assign n65629 = pi19 ? n22525 : n1077;
  assign n65630 = pi18 ? n32 : n65629;
  assign n65631 = pi17 ? n3067 : ~n65630;
  assign n65632 = pi16 ? n32 : n65631;
  assign n65633 = pi15 ? n65628 : n65632;
  assign n65634 = pi14 ? n65626 : n65633;
  assign n65635 = pi13 ? n65625 : n65634;
  assign n65636 = pi12 ? n65618 : n65635;
  assign n65637 = pi11 ? n65616 : n65636;
  assign n65638 = pi19 ? n4670 : n343;
  assign n65639 = pi18 ? n32 : n65638;
  assign n65640 = pi17 ? n65504 : ~n65639;
  assign n65641 = pi16 ? n32 : n65640;
  assign n65642 = pi18 ? n20164 : n684;
  assign n65643 = pi17 ? n65266 : ~n65642;
  assign n65644 = pi16 ? n32 : n65643;
  assign n65645 = pi15 ? n65641 : n65644;
  assign n65646 = pi15 ? n24237 : n24367;
  assign n65647 = pi14 ? n65645 : n65646;
  assign n65648 = pi17 ? n18395 : n25317;
  assign n65649 = pi16 ? n32 : n65648;
  assign n65650 = pi15 ? n65649 : n16374;
  assign n65651 = pi14 ? n65650 : n49389;
  assign n65652 = pi13 ? n65647 : n65651;
  assign n65653 = pi19 ? n1818 : ~n349;
  assign n65654 = pi18 ? n32 : n65653;
  assign n65655 = pi17 ? n32 : n65654;
  assign n65656 = pi16 ? n32 : n65655;
  assign n65657 = pi15 ? n65656 : n15834;
  assign n65658 = pi14 ? n65657 : n51140;
  assign n65659 = pi18 ? n684 : ~n4244;
  assign n65660 = pi17 ? n32 : n65659;
  assign n65661 = pi16 ? n32 : n65660;
  assign n65662 = pi19 ? n32 : n13587;
  assign n65663 = pi18 ? n37293 : ~n65662;
  assign n65664 = pi17 ? n52185 : n65663;
  assign n65665 = pi16 ? n32 : n65664;
  assign n65666 = pi15 ? n65661 : n65665;
  assign n65667 = pi18 ? n880 : ~n962;
  assign n65668 = pi17 ? n32 : n65667;
  assign n65669 = pi16 ? n51150 : n65668;
  assign n65670 = pi16 ? n11886 : n65539;
  assign n65671 = pi15 ? n65669 : n65670;
  assign n65672 = pi14 ? n65666 : n65671;
  assign n65673 = pi13 ? n65658 : n65672;
  assign n65674 = pi12 ? n65652 : n65673;
  assign n65675 = pi18 ? n22885 : ~n37418;
  assign n65676 = pi17 ? n32 : n65675;
  assign n65677 = pi16 ? n32 : n65676;
  assign n65678 = pi19 ? n2141 : n236;
  assign n65679 = pi18 ? n32 : n65678;
  assign n65680 = pi17 ? n2750 : ~n65679;
  assign n65681 = pi16 ? n32 : n65680;
  assign n65682 = pi15 ? n65677 : n65681;
  assign n65683 = pi19 ? n1369 : ~n617;
  assign n65684 = pi18 ? n32 : n65683;
  assign n65685 = pi17 ? n32 : n65684;
  assign n65686 = pi16 ? n32 : n65685;
  assign n65687 = pi15 ? n15263 : n65686;
  assign n65688 = pi14 ? n65682 : n65687;
  assign n65689 = pi17 ? n20658 : n1542;
  assign n65690 = pi16 ? n32 : n65689;
  assign n65691 = pi17 ? n13946 : n1542;
  assign n65692 = pi16 ? n32 : n65691;
  assign n65693 = pi15 ? n65690 : n65692;
  assign n65694 = pi14 ? n65693 : n26288;
  assign n65695 = pi13 ? n65688 : n65694;
  assign n65696 = pi17 ? n20658 : n22538;
  assign n65697 = pi16 ? n32 : n65696;
  assign n65698 = pi16 ? n3352 : ~n65569;
  assign n65699 = pi15 ? n65697 : n65698;
  assign n65700 = pi18 ? n323 : n47421;
  assign n65701 = pi17 ? n32 : n65700;
  assign n65702 = pi16 ? n3356 : ~n65701;
  assign n65703 = pi20 ? n32 : ~n13674;
  assign n65704 = pi19 ? n65703 : n32;
  assign n65705 = pi18 ? n22885 : n65704;
  assign n65706 = pi17 ? n32 : n65705;
  assign n65707 = pi16 ? n11886 : n65706;
  assign n65708 = pi15 ? n65702 : n65707;
  assign n65709 = pi14 ? n65699 : n65708;
  assign n65710 = pi16 ? n2326 : ~n65582;
  assign n65711 = pi16 ? n51177 : ~n65584;
  assign n65712 = pi15 ? n65710 : n65711;
  assign n65713 = pi19 ? n813 : ~n531;
  assign n65714 = pi18 ? n32 : n65713;
  assign n65715 = pi17 ? n32 : n65714;
  assign n65716 = pi17 ? n65587 : ~n52550;
  assign n65717 = pi16 ? n65715 : n65716;
  assign n65718 = pi18 ? n940 : ~n34040;
  assign n65719 = pi17 ? n65718 : ~n2748;
  assign n65720 = pi16 ? n32 : n65719;
  assign n65721 = pi15 ? n65717 : n65720;
  assign n65722 = pi14 ? n65712 : n65721;
  assign n65723 = pi13 ? n65709 : n65722;
  assign n65724 = pi12 ? n65695 : n65723;
  assign n65725 = pi11 ? n65674 : n65724;
  assign n65726 = pi10 ? n65637 : n65725;
  assign n65727 = pi09 ? n65460 : n65726;
  assign n65728 = pi08 ? n65600 : n65727;
  assign n65729 = pi07 ? n65451 : n65728;
  assign n65730 = pi06 ? n65223 : n65729;
  assign n65731 = pi05 ? n64703 : n65730;
  assign n65732 = pi19 ? n519 : n13376;
  assign n65733 = pi18 ? n32 : n65732;
  assign n65734 = pi17 ? n32 : n65733;
  assign n65735 = pi16 ? n32 : n65734;
  assign n65736 = pi15 ? n32 : n65735;
  assign n65737 = pi14 ? n65736 : n17111;
  assign n65738 = pi13 ? n32 : n65737;
  assign n65739 = pi12 ? n32 : n65738;
  assign n65740 = pi11 ? n32 : n65739;
  assign n65741 = pi10 ? n32 : n65740;
  assign n65742 = pi14 ? n17189 : n17188;
  assign n65743 = pi14 ? n15848 : n51219;
  assign n65744 = pi13 ? n65742 : n65743;
  assign n65745 = pi20 ? n1385 : ~n141;
  assign n65746 = pi19 ? n32 : n65745;
  assign n65747 = pi18 ? n32 : n65746;
  assign n65748 = pi17 ? n32 : n65747;
  assign n65749 = pi16 ? n32 : n65748;
  assign n65750 = pi15 ? n16392 : n65749;
  assign n65751 = pi20 ? n10644 : ~n141;
  assign n65752 = pi19 ? n594 : n65751;
  assign n65753 = pi18 ? n32 : n65752;
  assign n65754 = pi17 ? n32 : n65753;
  assign n65755 = pi16 ? n32 : n65754;
  assign n65756 = pi15 ? n65755 : n51230;
  assign n65757 = pi14 ? n65750 : n65756;
  assign n65758 = pi13 ? n65757 : n51234;
  assign n65759 = pi12 ? n65744 : n65758;
  assign n65760 = pi14 ? n32 : n17039;
  assign n65761 = pi19 ? n23193 : ~n11561;
  assign n65762 = pi18 ? n32 : n65761;
  assign n65763 = pi17 ? n32 : n65762;
  assign n65764 = pi16 ? n32 : n65763;
  assign n65765 = pi15 ? n16452 : n65764;
  assign n65766 = pi14 ? n32 : n65765;
  assign n65767 = pi13 ? n65760 : n65766;
  assign n65768 = pi18 ? n19613 : ~n1965;
  assign n65769 = pi17 ? n32 : n65768;
  assign n65770 = pi16 ? n32 : n65769;
  assign n65771 = pi18 ? n45480 : ~n1965;
  assign n65772 = pi17 ? n3282 : n65771;
  assign n65773 = pi16 ? n32 : n65772;
  assign n65774 = pi15 ? n65770 : n65773;
  assign n65775 = pi14 ? n25384 : n65774;
  assign n65776 = pi17 ? n32 : ~n2733;
  assign n65777 = pi16 ? n32 : n65776;
  assign n65778 = pi18 ? n4671 : n684;
  assign n65779 = pi17 ? n3164 : ~n65778;
  assign n65780 = pi16 ? n32 : n65779;
  assign n65781 = pi15 ? n65777 : n65780;
  assign n65782 = pi19 ? n32 : ~n6338;
  assign n65783 = pi18 ? n32 : n65782;
  assign n65784 = pi20 ? n18834 : n32;
  assign n65785 = pi20 ? n6050 : ~n32;
  assign n65786 = pi19 ? n65784 : ~n65785;
  assign n65787 = pi19 ? n1464 : ~n3692;
  assign n65788 = pi18 ? n65786 : n65787;
  assign n65789 = pi17 ? n65783 : ~n65788;
  assign n65790 = pi16 ? n32 : n65789;
  assign n65791 = pi20 ? n974 : n17652;
  assign n65792 = pi19 ? n65791 : n6683;
  assign n65793 = pi19 ? n1464 : ~n247;
  assign n65794 = pi18 ? n65792 : ~n65793;
  assign n65795 = pi17 ? n26094 : n65794;
  assign n65796 = pi16 ? n32 : n65795;
  assign n65797 = pi15 ? n65790 : n65796;
  assign n65798 = pi14 ? n65781 : n65797;
  assign n65799 = pi13 ? n65775 : n65798;
  assign n65800 = pi12 ? n65767 : n65799;
  assign n65801 = pi11 ? n65759 : n65800;
  assign n65802 = pi19 ? n507 : n975;
  assign n65803 = pi18 ? n32 : n65802;
  assign n65804 = pi19 ? n32 : ~n16294;
  assign n65805 = pi18 ? n359 : n65804;
  assign n65806 = pi17 ? n65803 : ~n65805;
  assign n65807 = pi16 ? n32 : n65806;
  assign n65808 = pi19 ? n32 : ~n8907;
  assign n65809 = pi18 ? n32 : n65808;
  assign n65810 = pi20 ? n5854 : n18415;
  assign n65811 = pi19 ? n32 : n65810;
  assign n65812 = pi20 ? n2358 : n439;
  assign n65813 = pi19 ? n65812 : n247;
  assign n65814 = pi18 ? n65811 : ~n65813;
  assign n65815 = pi17 ? n65809 : ~n65814;
  assign n65816 = pi16 ? n32 : n65815;
  assign n65817 = pi15 ? n65807 : n65816;
  assign n65818 = pi17 ? n23572 : n16604;
  assign n65819 = pi16 ? n32 : n65818;
  assign n65820 = pi15 ? n65819 : n24367;
  assign n65821 = pi14 ? n65817 : n65820;
  assign n65822 = pi15 ? n16377 : n24582;
  assign n65823 = pi14 ? n24573 : n65822;
  assign n65824 = pi13 ? n65821 : n65823;
  assign n65825 = pi17 ? n32 : ~n51277;
  assign n65826 = pi16 ? n32 : n65825;
  assign n65827 = pi15 ? n62999 : n65826;
  assign n65828 = pi19 ? n24218 : ~n502;
  assign n65829 = pi18 ? n51281 : n65828;
  assign n65830 = pi17 ? n32 : n65829;
  assign n65831 = pi16 ? n32 : n65830;
  assign n65832 = pi18 ? n4380 : n6669;
  assign n65833 = pi17 ? n32 : n65832;
  assign n65834 = pi16 ? n32 : n65833;
  assign n65835 = pi15 ? n65831 : n65834;
  assign n65836 = pi14 ? n65827 : n65835;
  assign n65837 = pi18 ? n1819 : n48972;
  assign n65838 = pi17 ? n32 : n65837;
  assign n65839 = pi16 ? n32 : n65838;
  assign n65840 = pi19 ? n1757 : n1812;
  assign n65841 = pi18 ? n12368 : ~n65840;
  assign n65842 = pi17 ? n2637 : ~n65841;
  assign n65843 = pi16 ? n1808 : ~n65842;
  assign n65844 = pi15 ? n65839 : n65843;
  assign n65845 = pi19 ? n28926 : ~n507;
  assign n65846 = pi18 ? n32 : n65845;
  assign n65847 = pi17 ? n32 : n65846;
  assign n65848 = pi19 ? n343 : ~n1941;
  assign n65849 = pi18 ? n32 : n65848;
  assign n65850 = pi17 ? n32 : n65849;
  assign n65851 = pi16 ? n65847 : n65850;
  assign n65852 = pi20 ? n1385 : ~n342;
  assign n65853 = pi19 ? n65852 : n5694;
  assign n65854 = pi18 ? n32 : n65853;
  assign n65855 = pi17 ? n32 : n65854;
  assign n65856 = pi18 ? n4127 : n14572;
  assign n65857 = pi17 ? n32 : n65856;
  assign n65858 = pi16 ? n65855 : n65857;
  assign n65859 = pi15 ? n65851 : n65858;
  assign n65860 = pi14 ? n65844 : n65859;
  assign n65861 = pi13 ? n65836 : n65860;
  assign n65862 = pi12 ? n65824 : n65861;
  assign n65863 = pi15 ? n51310 : n23484;
  assign n65864 = pi19 ? n1818 : n5626;
  assign n65865 = pi18 ? n32 : n65864;
  assign n65866 = pi17 ? n32 : n65865;
  assign n65867 = pi16 ? n32 : n65866;
  assign n65868 = pi15 ? n15123 : n65867;
  assign n65869 = pi14 ? n65863 : n65868;
  assign n65870 = pi17 ? n20658 : n23158;
  assign n65871 = pi16 ? n32 : n65870;
  assign n65872 = pi15 ? n65871 : n65690;
  assign n65873 = pi14 ? n65872 : n64089;
  assign n65874 = pi13 ? n65869 : n65873;
  assign n65875 = pi19 ? n19116 : ~n32;
  assign n65876 = pi18 ? n32 : n65875;
  assign n65877 = pi17 ? n65876 : ~n19886;
  assign n65878 = pi16 ? n2860 : ~n65877;
  assign n65879 = pi18 ? n684 : ~n2079;
  assign n65880 = pi17 ? n32 : n65879;
  assign n65881 = pi16 ? n1808 : ~n65880;
  assign n65882 = pi15 ? n65878 : n65881;
  assign n65883 = pi20 ? n266 : ~n34841;
  assign n65884 = pi19 ? n65883 : ~n32;
  assign n65885 = pi18 ? n12368 : n65884;
  assign n65886 = pi17 ? n32 : n65885;
  assign n65887 = pi16 ? n1815 : ~n65886;
  assign n65888 = pi18 ? n12368 : n13324;
  assign n65889 = pi17 ? n32 : n65888;
  assign n65890 = pi16 ? n2320 : n65889;
  assign n65891 = pi15 ? n65887 : n65890;
  assign n65892 = pi14 ? n65882 : n65891;
  assign n65893 = pi18 ? n237 : ~n29978;
  assign n65894 = pi18 ? n17118 : n595;
  assign n65895 = pi17 ? n65893 : ~n65894;
  assign n65896 = pi16 ? n2320 : n65895;
  assign n65897 = pi16 ? n1934 : ~n2513;
  assign n65898 = pi15 ? n65896 : n65897;
  assign n65899 = pi20 ? n1319 : n220;
  assign n65900 = pi19 ? n65899 : n32;
  assign n65901 = pi18 ? n32 : n65900;
  assign n65902 = pi17 ? n32 : n65901;
  assign n65903 = pi18 ? n32 : n41364;
  assign n65904 = pi17 ? n65903 : ~n52550;
  assign n65905 = pi16 ? n65902 : n65904;
  assign n65906 = pi18 ? n32 : n41425;
  assign n65907 = pi17 ? n65906 : ~n2748;
  assign n65908 = pi16 ? n32 : n65907;
  assign n65909 = pi15 ? n65905 : n65908;
  assign n65910 = pi14 ? n65898 : n65909;
  assign n65911 = pi13 ? n65892 : n65910;
  assign n65912 = pi12 ? n65874 : n65911;
  assign n65913 = pi11 ? n65862 : n65912;
  assign n65914 = pi10 ? n65801 : n65913;
  assign n65915 = pi09 ? n65741 : n65914;
  assign n65916 = pi19 ? n519 : n4342;
  assign n65917 = pi18 ? n32 : n65916;
  assign n65918 = pi17 ? n32 : n65917;
  assign n65919 = pi16 ? n32 : n65918;
  assign n65920 = pi15 ? n32 : n65919;
  assign n65921 = pi14 ? n65920 : n16984;
  assign n65922 = pi13 ? n32 : n65921;
  assign n65923 = pi12 ? n32 : n65922;
  assign n65924 = pi11 ? n32 : n65923;
  assign n65925 = pi10 ? n32 : n65924;
  assign n65926 = pi14 ? n38060 : n51345;
  assign n65927 = pi13 ? n40855 : n65926;
  assign n65928 = pi20 ? n1385 : n125;
  assign n65929 = pi19 ? n32 : n65928;
  assign n65930 = pi18 ? n32 : n65929;
  assign n65931 = pi17 ? n32 : n65930;
  assign n65932 = pi16 ? n32 : n65931;
  assign n65933 = pi15 ? n16832 : n65932;
  assign n65934 = pi20 ? n10644 : ~n339;
  assign n65935 = pi19 ? n594 : n65934;
  assign n65936 = pi18 ? n32 : n65935;
  assign n65937 = pi17 ? n32 : n65936;
  assign n65938 = pi16 ? n32 : n65937;
  assign n65939 = pi19 ? n594 : n13074;
  assign n65940 = pi18 ? n32 : n65939;
  assign n65941 = pi17 ? n32 : n65940;
  assign n65942 = pi16 ? n32 : n65941;
  assign n65943 = pi15 ? n65938 : n65942;
  assign n65944 = pi14 ? n65933 : n65943;
  assign n65945 = pi14 ? n25438 : n17189;
  assign n65946 = pi13 ? n65944 : n65945;
  assign n65947 = pi12 ? n65927 : n65946;
  assign n65948 = pi14 ? n17189 : n17039;
  assign n65949 = pi13 ? n65948 : n65766;
  assign n65950 = pi18 ? n1078 : ~n2962;
  assign n65951 = pi17 ? n32 : n65950;
  assign n65952 = pi16 ? n32 : n65951;
  assign n65953 = pi19 ? n8946 : ~n32;
  assign n65954 = pi18 ? n65953 : ~n2962;
  assign n65955 = pi17 ? n3282 : n65954;
  assign n65956 = pi16 ? n32 : n65955;
  assign n65957 = pi15 ? n65952 : n65956;
  assign n65958 = pi14 ? n25384 : n65957;
  assign n65959 = pi17 ? n32 : ~n3182;
  assign n65960 = pi16 ? n32 : n65959;
  assign n65961 = pi18 ? n4671 : n2830;
  assign n65962 = pi17 ? n3164 : ~n65961;
  assign n65963 = pi16 ? n32 : n65962;
  assign n65964 = pi15 ? n65960 : n65963;
  assign n65965 = pi19 ? n55424 : n65785;
  assign n65966 = pi19 ? n1464 : ~n7443;
  assign n65967 = pi18 ? n65965 : ~n65966;
  assign n65968 = pi17 ? n65783 : n65967;
  assign n65969 = pi16 ? n32 : n65968;
  assign n65970 = pi19 ? n1464 : ~n7881;
  assign n65971 = pi18 ? n65792 : ~n65970;
  assign n65972 = pi17 ? n32 : n65971;
  assign n65973 = pi16 ? n32 : n65972;
  assign n65974 = pi15 ? n65969 : n65973;
  assign n65975 = pi14 ? n65964 : n65974;
  assign n65976 = pi13 ? n65958 : n65975;
  assign n65977 = pi12 ? n65949 : n65976;
  assign n65978 = pi11 ? n65947 : n65977;
  assign n65979 = pi19 ? n32 : ~n25448;
  assign n65980 = pi18 ? n359 : n65979;
  assign n65981 = pi17 ? n19886 : ~n65980;
  assign n65982 = pi16 ? n32 : n65981;
  assign n65983 = pi20 ? n1324 : n274;
  assign n65984 = pi19 ? n65983 : n32;
  assign n65985 = pi18 ? n9346 : ~n65984;
  assign n65986 = pi17 ? n65809 : ~n65985;
  assign n65987 = pi16 ? n32 : n65986;
  assign n65988 = pi15 ? n65982 : n65987;
  assign n65989 = pi17 ? n23572 : n32;
  assign n65990 = pi16 ? n32 : n65989;
  assign n65991 = pi17 ? n16317 : n16604;
  assign n65992 = pi16 ? n32 : n65991;
  assign n65993 = pi15 ? n65990 : n65992;
  assign n65994 = pi14 ? n65988 : n65993;
  assign n65995 = pi15 ? n26885 : n37654;
  assign n65996 = pi14 ? n24633 : n65995;
  assign n65997 = pi13 ? n65994 : n65996;
  assign n65998 = pi19 ? n5694 : ~n7014;
  assign n65999 = pi18 ? n32 : n65998;
  assign n66000 = pi17 ? n32 : n65999;
  assign n66001 = pi16 ? n32 : n66000;
  assign n66002 = pi17 ? n32 : n51374;
  assign n66003 = pi16 ? n32 : n66002;
  assign n66004 = pi15 ? n66001 : n66003;
  assign n66005 = pi19 ? n24218 : ~n349;
  assign n66006 = pi18 ? n51281 : n66005;
  assign n66007 = pi17 ? n32 : n66006;
  assign n66008 = pi16 ? n32 : n66007;
  assign n66009 = pi15 ? n66008 : n65834;
  assign n66010 = pi14 ? n66004 : n66009;
  assign n66011 = pi19 ? n349 : ~n12245;
  assign n66012 = pi18 ? n1819 : n66011;
  assign n66013 = pi17 ? n32 : n66012;
  assign n66014 = pi16 ? n32 : n66013;
  assign n66015 = pi19 ? n1757 : n12245;
  assign n66016 = pi18 ? n12368 : ~n66015;
  assign n66017 = pi17 ? n2519 : ~n66016;
  assign n66018 = pi16 ? n2306 : ~n66017;
  assign n66019 = pi15 ? n66014 : n66018;
  assign n66020 = pi19 ? n51391 : ~n507;
  assign n66021 = pi18 ? n32 : n66020;
  assign n66022 = pi17 ? n32 : n66021;
  assign n66023 = pi19 ? n343 : ~n31155;
  assign n66024 = pi18 ? n32 : n66023;
  assign n66025 = pi17 ? n32 : n66024;
  assign n66026 = pi16 ? n66022 : n66025;
  assign n66027 = pi19 ? n4982 : n5694;
  assign n66028 = pi18 ? n32 : n66027;
  assign n66029 = pi17 ? n32 : n66028;
  assign n66030 = pi19 ? n208 : ~n31155;
  assign n66031 = pi18 ? n4127 : n66030;
  assign n66032 = pi17 ? n32 : n66031;
  assign n66033 = pi16 ? n66029 : n66032;
  assign n66034 = pi15 ? n66026 : n66033;
  assign n66035 = pi14 ? n66019 : n66034;
  assign n66036 = pi13 ? n66010 : n66035;
  assign n66037 = pi12 ? n65997 : n66036;
  assign n66038 = pi18 ? n863 : n54354;
  assign n66039 = pi17 ? n32 : n66038;
  assign n66040 = pi16 ? n32 : n66039;
  assign n66041 = pi15 ? n66040 : n23749;
  assign n66042 = pi14 ? n66041 : n21681;
  assign n66043 = pi17 ? n20658 : n15516;
  assign n66044 = pi16 ? n32 : n66043;
  assign n66045 = pi15 ? n65871 : n66044;
  assign n66046 = pi15 ? n24274 : n23011;
  assign n66047 = pi14 ? n66045 : n66046;
  assign n66048 = pi13 ? n66042 : n66047;
  assign n66049 = pi17 ? n65876 : ~n23009;
  assign n66050 = pi16 ? n2860 : ~n66049;
  assign n66051 = pi18 ? n684 : ~n6118;
  assign n66052 = pi17 ? n32 : n66051;
  assign n66053 = pi16 ? n2300 : ~n66052;
  assign n66054 = pi15 ? n66050 : n66053;
  assign n66055 = pi16 ? n2530 : ~n65886;
  assign n66056 = pi16 ? n3625 : n65889;
  assign n66057 = pi15 ? n66055 : n66056;
  assign n66058 = pi14 ? n66054 : n66057;
  assign n66059 = pi16 ? n3625 : n65895;
  assign n66060 = pi16 ? n2426 : ~n2629;
  assign n66061 = pi15 ? n66059 : n66060;
  assign n66062 = pi19 ? n32 : ~n15983;
  assign n66063 = pi18 ? n32 : n66062;
  assign n66064 = pi17 ? n66063 : ~n52550;
  assign n66065 = pi16 ? n14388 : n66064;
  assign n66066 = pi20 ? n974 : ~n207;
  assign n66067 = pi19 ? n322 : ~n66066;
  assign n66068 = pi18 ? n32 : n66067;
  assign n66069 = pi17 ? n66068 : ~n2748;
  assign n66070 = pi16 ? n32 : n66069;
  assign n66071 = pi15 ? n66065 : n66070;
  assign n66072 = pi14 ? n66061 : n66071;
  assign n66073 = pi13 ? n66058 : n66072;
  assign n66074 = pi12 ? n66048 : n66073;
  assign n66075 = pi11 ? n66037 : n66074;
  assign n66076 = pi10 ? n65978 : n66075;
  assign n66077 = pi09 ? n65925 : n66076;
  assign n66078 = pi08 ? n65915 : n66077;
  assign n66079 = pi14 ? n16985 : n25556;
  assign n66080 = pi13 ? n32 : n66079;
  assign n66081 = pi12 ? n32 : n66080;
  assign n66082 = pi11 ? n32 : n66081;
  assign n66083 = pi10 ? n32 : n66082;
  assign n66084 = pi14 ? n17412 : n37458;
  assign n66085 = pi15 ? n17188 : n25704;
  assign n66086 = pi14 ? n66085 : n26330;
  assign n66087 = pi13 ? n66084 : n66086;
  assign n66088 = pi14 ? n52908 : n26548;
  assign n66089 = pi14 ? n16838 : n51429;
  assign n66090 = pi13 ? n66088 : n66089;
  assign n66091 = pi12 ? n66087 : n66090;
  assign n66092 = pi14 ? n27934 : n51428;
  assign n66093 = pi18 ? n32 : n42092;
  assign n66094 = pi17 ? n32 : n66093;
  assign n66095 = pi16 ? n32 : n66094;
  assign n66096 = pi15 ? n15847 : n66095;
  assign n66097 = pi14 ? n32 : n66096;
  assign n66098 = pi13 ? n66092 : n66097;
  assign n66099 = pi18 ? n4428 : ~n2962;
  assign n66100 = pi17 ? n32 : n66099;
  assign n66101 = pi16 ? n32 : n66100;
  assign n66102 = pi15 ? n11725 : n66101;
  assign n66103 = pi14 ? n15847 : n66102;
  assign n66104 = pi18 ? n13070 : n1965;
  assign n66105 = pi17 ? n32 : ~n66104;
  assign n66106 = pi16 ? n32 : n66105;
  assign n66107 = pi18 ? n13080 : n684;
  assign n66108 = pi17 ? n3164 : ~n66107;
  assign n66109 = pi16 ? n32 : n66108;
  assign n66110 = pi15 ? n66106 : n66109;
  assign n66111 = pi19 ? n507 : n4721;
  assign n66112 = pi18 ? n66111 : ~n65966;
  assign n66113 = pi17 ? n32 : n66112;
  assign n66114 = pi16 ? n32 : n66113;
  assign n66115 = pi18 ? n22885 : ~n65966;
  assign n66116 = pi17 ? n32 : n66115;
  assign n66117 = pi16 ? n32 : n66116;
  assign n66118 = pi15 ? n66114 : n66117;
  assign n66119 = pi14 ? n66110 : n66118;
  assign n66120 = pi13 ? n66103 : n66119;
  assign n66121 = pi12 ? n66098 : n66120;
  assign n66122 = pi11 ? n66091 : n66121;
  assign n66123 = pi19 ? n32 : ~n25514;
  assign n66124 = pi18 ? n24205 : ~n66123;
  assign n66125 = pi17 ? n32 : n66124;
  assign n66126 = pi16 ? n32 : n66125;
  assign n66127 = pi18 ? n51208 : n16783;
  assign n66128 = pi17 ? n4111 : n66127;
  assign n66129 = pi16 ? n32 : n66128;
  assign n66130 = pi15 ? n66126 : n66129;
  assign n66131 = pi17 ? n2959 : n16784;
  assign n66132 = pi16 ? n32 : n66131;
  assign n66133 = pi15 ? n66132 : n16606;
  assign n66134 = pi14 ? n66130 : n66133;
  assign n66135 = pi15 ? n24237 : n37654;
  assign n66136 = pi14 ? n24633 : n66135;
  assign n66137 = pi13 ? n66134 : n66136;
  assign n66138 = pi15 ? n62999 : n51464;
  assign n66139 = pi19 ? n5688 : ~n9668;
  assign n66140 = pi18 ? n940 : n66139;
  assign n66141 = pi17 ? n32 : n66140;
  assign n66142 = pi16 ? n32 : n66141;
  assign n66143 = pi18 ? n32 : n63684;
  assign n66144 = pi17 ? n32 : n66143;
  assign n66145 = pi16 ? n32 : n66144;
  assign n66146 = pi15 ? n66142 : n66145;
  assign n66147 = pi14 ? n66138 : n66146;
  assign n66148 = pi18 ? n32 : n6628;
  assign n66149 = pi17 ? n32 : n66148;
  assign n66150 = pi16 ? n32 : n66149;
  assign n66151 = pi18 ? n4380 : n5747;
  assign n66152 = pi17 ? n2750 : ~n66151;
  assign n66153 = pi16 ? n2120 : ~n66152;
  assign n66154 = pi15 ? n66150 : n66153;
  assign n66155 = pi16 ? n2518 : n35700;
  assign n66156 = pi19 ? n5350 : n5694;
  assign n66157 = pi18 ? n32 : n66156;
  assign n66158 = pi17 ? n32 : n66157;
  assign n66159 = pi18 ? n863 : n14567;
  assign n66160 = pi17 ? n32 : n66159;
  assign n66161 = pi16 ? n66158 : n66160;
  assign n66162 = pi15 ? n66155 : n66161;
  assign n66163 = pi14 ? n66154 : n66162;
  assign n66164 = pi13 ? n66147 : n66163;
  assign n66165 = pi12 ? n66137 : n66164;
  assign n66166 = pi15 ? n14397 : n23749;
  assign n66167 = pi14 ? n66166 : n23484;
  assign n66168 = pi15 ? n23160 : n15665;
  assign n66169 = pi19 ? n244 : ~n5748;
  assign n66170 = pi18 ? n32 : n66169;
  assign n66171 = pi17 ? n32 : n66170;
  assign n66172 = pi16 ? n66171 : n1108;
  assign n66173 = pi15 ? n22923 : n66172;
  assign n66174 = pi14 ? n66168 : n66173;
  assign n66175 = pi13 ? n66167 : n66174;
  assign n66176 = pi18 ? n32 : n48270;
  assign n66177 = pi17 ? n66176 : ~n23009;
  assign n66178 = pi16 ? n2860 : ~n66177;
  assign n66179 = pi18 ? n209 : ~n6145;
  assign n66180 = pi17 ? n32 : n66179;
  assign n66181 = pi16 ? n2120 : ~n66180;
  assign n66182 = pi15 ? n66178 : n66181;
  assign n66183 = pi16 ? n2426 : ~n2860;
  assign n66184 = pi20 ? n749 : ~n101;
  assign n66185 = pi19 ? n66184 : n32;
  assign n66186 = pi18 ? n940 : n66185;
  assign n66187 = pi17 ? n1028 : ~n66186;
  assign n66188 = pi16 ? n2293 : ~n66187;
  assign n66189 = pi15 ? n66183 : n66188;
  assign n66190 = pi14 ? n66182 : n66189;
  assign n66191 = pi16 ? n2293 : ~n3946;
  assign n66192 = pi16 ? n3769 : ~n2629;
  assign n66193 = pi15 ? n66191 : n66192;
  assign n66194 = pi20 ? n32 : n9897;
  assign n66195 = pi19 ? n66194 : n32;
  assign n66196 = pi18 ? n32 : n66195;
  assign n66197 = pi17 ? n32 : n66196;
  assign n66198 = pi18 ? n32 : n33637;
  assign n66199 = pi18 ? n1548 : ~n508;
  assign n66200 = pi17 ? n66198 : n66199;
  assign n66201 = pi16 ? n66197 : n66200;
  assign n66202 = pi18 ? n32 : n18193;
  assign n66203 = pi20 ? n32 : n20265;
  assign n66204 = pi19 ? n66203 : ~n32;
  assign n66205 = pi18 ? n237 : ~n66204;
  assign n66206 = pi17 ? n66202 : n66205;
  assign n66207 = pi16 ? n32 : n66206;
  assign n66208 = pi15 ? n66201 : n66207;
  assign n66209 = pi14 ? n66193 : n66208;
  assign n66210 = pi13 ? n66190 : n66209;
  assign n66211 = pi12 ? n66175 : n66210;
  assign n66212 = pi11 ? n66165 : n66211;
  assign n66213 = pi10 ? n66122 : n66212;
  assign n66214 = pi09 ? n66083 : n66213;
  assign n66215 = pi15 ? n16984 : n25556;
  assign n66216 = pi14 ? n66215 : n17111;
  assign n66217 = pi15 ? n32 : n51510;
  assign n66218 = pi14 ? n66217 : n25815;
  assign n66219 = pi13 ? n66216 : n66218;
  assign n66220 = pi20 ? n428 : n481;
  assign n66221 = pi19 ? n32 : n66220;
  assign n66222 = pi18 ? n32 : n66221;
  assign n66223 = pi17 ? n32 : n66222;
  assign n66224 = pi16 ? n32 : n66223;
  assign n66225 = pi15 ? n32 : n66224;
  assign n66226 = pi15 ? n38071 : n25708;
  assign n66227 = pi14 ? n66225 : n66226;
  assign n66228 = pi19 ? n32 : n6106;
  assign n66229 = pi18 ? n32 : n66228;
  assign n66230 = pi17 ? n32 : n66229;
  assign n66231 = pi16 ? n32 : n66230;
  assign n66232 = pi15 ? n16392 : n66231;
  assign n66233 = pi14 ? n66232 : n17412;
  assign n66234 = pi13 ? n66227 : n66233;
  assign n66235 = pi12 ? n66219 : n66234;
  assign n66236 = pi18 ? n4428 : ~n880;
  assign n66237 = pi17 ? n32 : n66236;
  assign n66238 = pi16 ? n32 : n66237;
  assign n66239 = pi15 ? n11000 : n66238;
  assign n66240 = pi14 ? n16485 : n66239;
  assign n66241 = pi18 ? n46371 : n1965;
  assign n66242 = pi17 ? n3164 : ~n66241;
  assign n66243 = pi16 ? n32 : n66242;
  assign n66244 = pi15 ? n66106 : n66243;
  assign n66245 = pi19 ? n1464 : ~n10645;
  assign n66246 = pi18 ? n66111 : ~n66245;
  assign n66247 = pi17 ? n32 : n66246;
  assign n66248 = pi16 ? n32 : n66247;
  assign n66249 = pi18 ? n22885 : ~n66245;
  assign n66250 = pi17 ? n32 : n66249;
  assign n66251 = pi16 ? n32 : n66250;
  assign n66252 = pi15 ? n66248 : n66251;
  assign n66253 = pi14 ? n66244 : n66252;
  assign n66254 = pi13 ? n66240 : n66253;
  assign n66255 = pi12 ? n66098 : n66254;
  assign n66256 = pi11 ? n66235 : n66255;
  assign n66257 = pi18 ? n520 : ~n66123;
  assign n66258 = pi17 ? n32 : n66257;
  assign n66259 = pi16 ? n32 : n66258;
  assign n66260 = pi18 ? n51208 : n32;
  assign n66261 = pi17 ? n4111 : n66260;
  assign n66262 = pi16 ? n32 : n66261;
  assign n66263 = pi15 ? n66259 : n66262;
  assign n66264 = pi17 ? n2959 : n1124;
  assign n66265 = pi16 ? n32 : n66264;
  assign n66266 = pi15 ? n66265 : n16601;
  assign n66267 = pi14 ? n66263 : n66266;
  assign n66268 = pi19 ? n507 : n9724;
  assign n66269 = pi18 ? n32 : n66268;
  assign n66270 = pi17 ? n32 : n66269;
  assign n66271 = pi16 ? n32 : n66270;
  assign n66272 = pi15 ? n24572 : n66271;
  assign n66273 = pi14 ? n37574 : n66272;
  assign n66274 = pi13 ? n66267 : n66273;
  assign n66275 = pi19 ? n5694 : ~n288;
  assign n66276 = pi18 ? n32 : n66275;
  assign n66277 = pi17 ? n32 : n66276;
  assign n66278 = pi16 ? n32 : n66277;
  assign n66279 = pi15 ? n66278 : n51464;
  assign n66280 = pi15 ? n51469 : n66145;
  assign n66281 = pi14 ? n66279 : n66280;
  assign n66282 = pi19 ? n349 : ~n9368;
  assign n66283 = pi18 ? n32 : n66282;
  assign n66284 = pi17 ? n32 : n66283;
  assign n66285 = pi16 ? n32 : n66284;
  assign n66286 = pi16 ? n2756 : ~n66152;
  assign n66287 = pi15 ? n66285 : n66286;
  assign n66288 = pi16 ? n2756 : n14338;
  assign n66289 = pi18 ? n863 : n24440;
  assign n66290 = pi17 ? n32 : n66289;
  assign n66291 = pi16 ? n16849 : n66290;
  assign n66292 = pi15 ? n66288 : n66291;
  assign n66293 = pi14 ? n66287 : n66292;
  assign n66294 = pi13 ? n66281 : n66293;
  assign n66295 = pi12 ? n66274 : n66294;
  assign n66296 = pi15 ? n23802 : n23749;
  assign n66297 = pi14 ? n66296 : n23484;
  assign n66298 = pi19 ? n322 : ~n5748;
  assign n66299 = pi18 ? n32 : n66298;
  assign n66300 = pi17 ? n32 : n66299;
  assign n66301 = pi16 ? n66300 : n1543;
  assign n66302 = pi15 ? n22923 : n66301;
  assign n66303 = pi14 ? n24397 : n66302;
  assign n66304 = pi13 ? n66297 : n66303;
  assign n66305 = pi16 ? n2749 : ~n66180;
  assign n66306 = pi15 ? n66178 : n66305;
  assign n66307 = pi16 ? n2518 : ~n2860;
  assign n66308 = pi16 ? n2513 : ~n66187;
  assign n66309 = pi15 ? n66307 : n66308;
  assign n66310 = pi14 ? n66306 : n66309;
  assign n66311 = pi16 ? n2513 : ~n4100;
  assign n66312 = pi16 ? n4100 : ~n3946;
  assign n66313 = pi15 ? n66311 : n66312;
  assign n66314 = pi19 ? n32 : ~n39738;
  assign n66315 = pi18 ? n32 : n66314;
  assign n66316 = pi17 ? n66315 : n10700;
  assign n66317 = pi16 ? n32 : n66316;
  assign n66318 = pi19 ? n322 : ~n38520;
  assign n66319 = pi18 ? n32 : n66318;
  assign n66320 = pi18 ? n618 : ~n5778;
  assign n66321 = pi17 ? n66319 : n66320;
  assign n66322 = pi16 ? n32 : n66321;
  assign n66323 = pi15 ? n66317 : n66322;
  assign n66324 = pi14 ? n66313 : n66323;
  assign n66325 = pi13 ? n66310 : n66324;
  assign n66326 = pi12 ? n66304 : n66325;
  assign n66327 = pi11 ? n66295 : n66326;
  assign n66328 = pi10 ? n66256 : n66327;
  assign n66329 = pi09 ? n66083 : n66328;
  assign n66330 = pi08 ? n66214 : n66329;
  assign n66331 = pi07 ? n66078 : n66330;
  assign n66332 = pi14 ? n32 : n17435;
  assign n66333 = pi13 ? n32 : n66332;
  assign n66334 = pi12 ? n32 : n66333;
  assign n66335 = pi11 ? n32 : n66334;
  assign n66336 = pi10 ? n32 : n66335;
  assign n66337 = pi14 ? n17578 : n25867;
  assign n66338 = pi14 ? n25557 : n51560;
  assign n66339 = pi13 ? n66337 : n66338;
  assign n66340 = pi15 ? n16392 : n51644;
  assign n66341 = pi19 ? n32 : n7405;
  assign n66342 = pi18 ? n32 : n66341;
  assign n66343 = pi17 ? n32 : n66342;
  assign n66344 = pi16 ? n32 : n66343;
  assign n66345 = pi15 ? n51510 : n66344;
  assign n66346 = pi14 ? n66340 : n66345;
  assign n66347 = pi14 ? n16985 : n32;
  assign n66348 = pi13 ? n66346 : n66347;
  assign n66349 = pi12 ? n66339 : n66348;
  assign n66350 = pi14 ? n25625 : n16984;
  assign n66351 = pi14 ? n55556 : n55525;
  assign n66352 = pi13 ? n66350 : n66351;
  assign n66353 = pi18 ? n209 : ~n366;
  assign n66354 = pi17 ? n32 : n66353;
  assign n66355 = pi16 ? n32 : n66354;
  assign n66356 = pi15 ? n16629 : n66355;
  assign n66357 = pi18 ? n863 : ~n34633;
  assign n66358 = pi17 ? n32 : n66357;
  assign n66359 = pi16 ? n32 : n66358;
  assign n66360 = pi15 ? n66359 : n11696;
  assign n66361 = pi14 ? n66356 : n66360;
  assign n66362 = pi19 ? n267 : n531;
  assign n66363 = pi18 ? n66362 : ~n1965;
  assign n66364 = pi17 ? n32 : n66363;
  assign n66365 = pi16 ? n32 : n66364;
  assign n66366 = pi18 ? n8535 : ~n1965;
  assign n66367 = pi17 ? n32 : n66366;
  assign n66368 = pi16 ? n32 : n66367;
  assign n66369 = pi15 ? n66365 : n66368;
  assign n66370 = pi19 ? n507 : ~n176;
  assign n66371 = pi18 ? n863 : ~n66370;
  assign n66372 = pi17 ? n32 : n66371;
  assign n66373 = pi16 ? n32 : n66372;
  assign n66374 = pi19 ? n531 : ~n11546;
  assign n66375 = pi18 ? n32 : n66374;
  assign n66376 = pi17 ? n32 : n66375;
  assign n66377 = pi16 ? n32 : n66376;
  assign n66378 = pi15 ? n66373 : n66377;
  assign n66379 = pi14 ? n66369 : n66378;
  assign n66380 = pi13 ? n66361 : n66379;
  assign n66381 = pi12 ? n66352 : n66380;
  assign n66382 = pi11 ? n66349 : n66381;
  assign n66383 = pi19 ? n5614 : n247;
  assign n66384 = pi18 ? n17848 : n66383;
  assign n66385 = pi17 ? n32 : n66384;
  assign n66386 = pi16 ? n32 : n66385;
  assign n66387 = pi18 ? n9012 : n16834;
  assign n66388 = pi17 ? n32 : n66387;
  assign n66389 = pi16 ? n32 : n66388;
  assign n66390 = pi15 ? n66386 : n66389;
  assign n66391 = pi18 ? n5009 : n16834;
  assign n66392 = pi17 ? n32 : n66391;
  assign n66393 = pi16 ? n32 : n66392;
  assign n66394 = pi15 ? n66393 : n16520;
  assign n66395 = pi14 ? n66390 : n66394;
  assign n66396 = pi15 ? n16520 : n24237;
  assign n66397 = pi15 ? n24712 : n16105;
  assign n66398 = pi14 ? n66396 : n66397;
  assign n66399 = pi13 ? n66395 : n66398;
  assign n66400 = pi15 ? n37190 : n37501;
  assign n66401 = pi19 ? n208 : ~n766;
  assign n66402 = pi18 ? n32 : n66401;
  assign n66403 = pi17 ? n32 : n66402;
  assign n66404 = pi16 ? n32 : n66403;
  assign n66405 = pi19 ? n322 : ~n7014;
  assign n66406 = pi18 ? n32 : n66405;
  assign n66407 = pi17 ? n32 : n66406;
  assign n66408 = pi16 ? n32 : n66407;
  assign n66409 = pi15 ? n66404 : n66408;
  assign n66410 = pi14 ? n66400 : n66409;
  assign n66411 = pi17 ? n2726 : ~n39518;
  assign n66412 = pi16 ? n2725 : ~n66411;
  assign n66413 = pi17 ? n2726 : ~n37188;
  assign n66414 = pi16 ? n2624 : ~n66413;
  assign n66415 = pi15 ? n66412 : n66414;
  assign n66416 = pi16 ? n38771 : n37196;
  assign n66417 = pi20 ? n141 : n274;
  assign n66418 = pi19 ? n32 : n66417;
  assign n66419 = pi18 ? n32 : n66418;
  assign n66420 = pi17 ? n32 : n66419;
  assign n66421 = pi19 ? n507 : ~n20022;
  assign n66422 = pi18 ? n32 : n66421;
  assign n66423 = pi17 ? n19655 : n66422;
  assign n66424 = pi16 ? n66420 : n66423;
  assign n66425 = pi15 ? n66416 : n66424;
  assign n66426 = pi14 ? n66415 : n66425;
  assign n66427 = pi13 ? n66410 : n66426;
  assign n66428 = pi12 ? n66399 : n66427;
  assign n66429 = pi19 ? n6398 : n5614;
  assign n66430 = pi18 ? n32 : n66429;
  assign n66431 = pi17 ? n32 : n66430;
  assign n66432 = pi16 ? n32 : n66431;
  assign n66433 = pi15 ? n32 : n66432;
  assign n66434 = pi18 ? n51606 : n6114;
  assign n66435 = pi17 ? n32 : n66434;
  assign n66436 = pi16 ? n32 : n66435;
  assign n66437 = pi15 ? n16108 : n66436;
  assign n66438 = pi14 ? n66433 : n66437;
  assign n66439 = pi14 ? n24397 : n22923;
  assign n66440 = pi13 ? n66438 : n66439;
  assign n66441 = pi18 ? n5747 : ~n54506;
  assign n66442 = pi17 ? n58032 : n66441;
  assign n66443 = pi16 ? n32 : ~n66442;
  assign n66444 = pi15 ? n66443 : n62285;
  assign n66445 = pi19 ? n357 : n1105;
  assign n66446 = pi18 ? n51614 : n66445;
  assign n66447 = pi17 ? n32 : n66446;
  assign n66448 = pi16 ? n4100 : ~n66447;
  assign n66449 = pi20 ? n266 : n13084;
  assign n66450 = pi19 ? n66449 : n32;
  assign n66451 = pi18 ? n32 : n66450;
  assign n66452 = pi17 ? n2355 : ~n66451;
  assign n66453 = pi16 ? n2745 : ~n66452;
  assign n66454 = pi15 ? n66448 : n66453;
  assign n66455 = pi14 ? n66444 : n66454;
  assign n66456 = pi16 ? n2745 : ~n4100;
  assign n66457 = pi15 ? n66456 : n46804;
  assign n66458 = pi19 ? n38221 : n1740;
  assign n66459 = pi18 ? n66458 : ~n2627;
  assign n66460 = pi17 ? n64639 : ~n66459;
  assign n66461 = pi16 ? n3165 : ~n66460;
  assign n66462 = pi18 ? n62604 : ~n52549;
  assign n66463 = pi17 ? n32 : n66462;
  assign n66464 = pi16 ? n32 : n66463;
  assign n66465 = pi15 ? n66461 : n66464;
  assign n66466 = pi14 ? n66457 : n66465;
  assign n66467 = pi13 ? n66455 : n66466;
  assign n66468 = pi12 ? n66440 : n66467;
  assign n66469 = pi11 ? n66428 : n66468;
  assign n66470 = pi10 ? n66382 : n66469;
  assign n66471 = pi09 ? n66336 : n66470;
  assign n66472 = pi14 ? n32 : n25753;
  assign n66473 = pi13 ? n32 : n66472;
  assign n66474 = pi12 ? n32 : n66473;
  assign n66475 = pi11 ? n32 : n66474;
  assign n66476 = pi10 ? n32 : n66475;
  assign n66477 = pi15 ? n25556 : n17435;
  assign n66478 = pi15 ? n25556 : n16984;
  assign n66479 = pi14 ? n66477 : n66478;
  assign n66480 = pi14 ? n17578 : n51648;
  assign n66481 = pi13 ? n66479 : n66480;
  assign n66482 = pi18 ? n32 : n41030;
  assign n66483 = pi17 ? n32 : n66482;
  assign n66484 = pi16 ? n32 : n66483;
  assign n66485 = pi15 ? n16392 : n66484;
  assign n66486 = pi19 ? n32 : n21042;
  assign n66487 = pi18 ? n32 : n66486;
  assign n66488 = pi17 ? n32 : n66487;
  assign n66489 = pi16 ? n32 : n66488;
  assign n66490 = pi15 ? n16595 : n66489;
  assign n66491 = pi14 ? n66485 : n66490;
  assign n66492 = pi13 ? n66491 : n66347;
  assign n66493 = pi12 ? n66481 : n66492;
  assign n66494 = pi14 ? n15848 : n55525;
  assign n66495 = pi13 ? n66350 : n66494;
  assign n66496 = pi18 ? n209 : ~n341;
  assign n66497 = pi17 ? n32 : n66496;
  assign n66498 = pi16 ? n32 : n66497;
  assign n66499 = pi15 ? n25704 : n66498;
  assign n66500 = pi19 ? n1757 : n365;
  assign n66501 = pi18 ? n863 : ~n66500;
  assign n66502 = pi17 ? n32 : n66501;
  assign n66503 = pi16 ? n32 : n66502;
  assign n66504 = pi18 ? n940 : ~n366;
  assign n66505 = pi17 ? n32 : n66504;
  assign n66506 = pi16 ? n32 : n66505;
  assign n66507 = pi15 ? n66503 : n66506;
  assign n66508 = pi14 ? n66499 : n66507;
  assign n66509 = pi19 ? n311 : n531;
  assign n66510 = pi18 ? n66509 : ~n2962;
  assign n66511 = pi17 ? n32 : n66510;
  assign n66512 = pi16 ? n32 : n66511;
  assign n66513 = pi19 ? n30659 : n531;
  assign n66514 = pi18 ? n66513 : ~n2962;
  assign n66515 = pi17 ? n32 : n66514;
  assign n66516 = pi16 ? n32 : n66515;
  assign n66517 = pi15 ? n66512 : n66516;
  assign n66518 = pi19 ? n507 : ~n13388;
  assign n66519 = pi18 ? n863 : ~n66518;
  assign n66520 = pi17 ? n32 : n66519;
  assign n66521 = pi16 ? n32 : n66520;
  assign n66522 = pi19 ? n531 : ~n20517;
  assign n66523 = pi18 ? n32 : n66522;
  assign n66524 = pi17 ? n32 : n66523;
  assign n66525 = pi16 ? n32 : n66524;
  assign n66526 = pi15 ? n66521 : n66525;
  assign n66527 = pi14 ? n66517 : n66526;
  assign n66528 = pi13 ? n66508 : n66527;
  assign n66529 = pi12 ? n66495 : n66528;
  assign n66530 = pi11 ? n66493 : n66529;
  assign n66531 = pi18 ? n17848 : n16449;
  assign n66532 = pi17 ? n32 : n66531;
  assign n66533 = pi16 ? n32 : n66532;
  assign n66534 = pi15 ? n66533 : n66389;
  assign n66535 = pi18 ? n23871 : n16834;
  assign n66536 = pi17 ? n32 : n66535;
  assign n66537 = pi16 ? n32 : n66536;
  assign n66538 = pi15 ? n66537 : n24874;
  assign n66539 = pi14 ? n66534 : n66538;
  assign n66540 = pi15 ? n16101 : n25155;
  assign n66541 = pi14 ? n66396 : n66540;
  assign n66542 = pi13 ? n66539 : n66541;
  assign n66543 = pi18 ? n32 : n48641;
  assign n66544 = pi17 ? n32 : n66543;
  assign n66545 = pi16 ? n32 : n66544;
  assign n66546 = pi15 ? n66404 : n66545;
  assign n66547 = pi14 ? n66400 : n66546;
  assign n66548 = pi16 ? n2725 : ~n66413;
  assign n66549 = pi15 ? n66412 : n66548;
  assign n66550 = pi15 ? n14917 : n15248;
  assign n66551 = pi14 ? n66549 : n66550;
  assign n66552 = pi13 ? n66547 : n66551;
  assign n66553 = pi12 ? n66542 : n66552;
  assign n66554 = pi19 ? n6398 : n1630;
  assign n66555 = pi18 ? n32 : n66554;
  assign n66556 = pi17 ? n32 : n66555;
  assign n66557 = pi16 ? n32 : n66556;
  assign n66558 = pi15 ? n32 : n66557;
  assign n66559 = pi18 ? n51606 : n23738;
  assign n66560 = pi17 ? n32 : n66559;
  assign n66561 = pi16 ? n32 : n66560;
  assign n66562 = pi15 ? n32 : n66561;
  assign n66563 = pi14 ? n66558 : n66562;
  assign n66564 = pi15 ? n23741 : n23160;
  assign n66565 = pi15 ? n15665 : n22923;
  assign n66566 = pi14 ? n66564 : n66565;
  assign n66567 = pi13 ? n66563 : n66566;
  assign n66568 = pi15 ? n66443 : n49412;
  assign n66569 = pi19 ? n207 : ~n1105;
  assign n66570 = pi18 ? n51661 : ~n66569;
  assign n66571 = pi17 ? n32 : n66570;
  assign n66572 = pi16 ? n4246 : ~n66571;
  assign n66573 = pi19 ? n18200 : n32;
  assign n66574 = pi18 ? n32 : n66573;
  assign n66575 = pi17 ? n2355 : ~n66574;
  assign n66576 = pi16 ? n2851 : ~n66575;
  assign n66577 = pi15 ? n66572 : n66576;
  assign n66578 = pi14 ? n66568 : n66577;
  assign n66579 = pi16 ? n3061 : ~n4100;
  assign n66580 = pi15 ? n66579 : n46804;
  assign n66581 = pi19 ? n9007 : n1740;
  assign n66582 = pi18 ? n66581 : ~n2627;
  assign n66583 = pi17 ? n64639 : ~n66582;
  assign n66584 = pi16 ? n3165 : ~n66583;
  assign n66585 = pi20 ? n321 : ~n765;
  assign n66586 = pi19 ? n66585 : ~n32;
  assign n66587 = pi18 ? n66586 : ~n9427;
  assign n66588 = pi17 ? n32 : n66587;
  assign n66589 = pi16 ? n32 : n66588;
  assign n66590 = pi15 ? n66584 : n66589;
  assign n66591 = pi14 ? n66580 : n66590;
  assign n66592 = pi13 ? n66578 : n66591;
  assign n66593 = pi12 ? n66567 : n66592;
  assign n66594 = pi11 ? n66553 : n66593;
  assign n66595 = pi10 ? n66530 : n66594;
  assign n66596 = pi09 ? n66476 : n66595;
  assign n66597 = pi08 ? n66471 : n66596;
  assign n66598 = pi14 ? n32 : n17336;
  assign n66599 = pi13 ? n32 : n66598;
  assign n66600 = pi12 ? n32 : n66599;
  assign n66601 = pi11 ? n32 : n66600;
  assign n66602 = pi10 ? n32 : n66601;
  assign n66603 = pi14 ? n25861 : n25693;
  assign n66604 = pi14 ? n17271 : n51689;
  assign n66605 = pi13 ? n66603 : n66604;
  assign n66606 = pi20 ? n342 : ~n56768;
  assign n66607 = pi19 ? n32 : n66606;
  assign n66608 = pi18 ? n32 : n66607;
  assign n66609 = pi17 ? n32 : n66608;
  assign n66610 = pi16 ? n32 : n66609;
  assign n66611 = pi15 ? n25708 : n66610;
  assign n66612 = pi15 ? n25763 : n25814;
  assign n66613 = pi14 ? n66611 : n66612;
  assign n66614 = pi13 ? n66613 : n17413;
  assign n66615 = pi12 ? n66605 : n66614;
  assign n66616 = pi14 ? n39461 : n25556;
  assign n66617 = pi15 ? n32 : n25763;
  assign n66618 = pi14 ? n66617 : n26330;
  assign n66619 = pi13 ? n66616 : n66618;
  assign n66620 = pi19 ? n236 : ~n13543;
  assign n66621 = pi18 ? n863 : n66620;
  assign n66622 = pi17 ? n32 : n66621;
  assign n66623 = pi16 ? n32 : n66622;
  assign n66624 = pi15 ? n25704 : n66623;
  assign n66625 = pi20 ? n3523 : n141;
  assign n66626 = pi19 ? n349 : ~n66625;
  assign n66627 = pi18 ? n32 : n66626;
  assign n66628 = pi17 ? n32 : n66627;
  assign n66629 = pi16 ? n32 : n66628;
  assign n66630 = pi18 ? n32 : ~n366;
  assign n66631 = pi17 ? n32 : n66630;
  assign n66632 = pi16 ? n32 : n66631;
  assign n66633 = pi15 ? n66629 : n66632;
  assign n66634 = pi14 ? n66624 : n66633;
  assign n66635 = pi19 ? n267 : n1464;
  assign n66636 = pi18 ? n66635 : ~n2962;
  assign n66637 = pi17 ? n32 : n66636;
  assign n66638 = pi16 ? n32 : n66637;
  assign n66639 = pi19 ? n5694 : n4721;
  assign n66640 = pi18 ? n66639 : ~n2962;
  assign n66641 = pi17 ? n32 : n66640;
  assign n66642 = pi16 ? n32 : n66641;
  assign n66643 = pi15 ? n66638 : n66642;
  assign n66644 = pi18 ? n32 : ~n11562;
  assign n66645 = pi17 ? n32 : n66644;
  assign n66646 = pi16 ? n32 : n66645;
  assign n66647 = pi19 ? n531 : ~n6042;
  assign n66648 = pi18 ? n32 : n66647;
  assign n66649 = pi17 ? n32 : n66648;
  assign n66650 = pi16 ? n32 : n66649;
  assign n66651 = pi15 ? n66646 : n66650;
  assign n66652 = pi14 ? n66643 : n66651;
  assign n66653 = pi13 ? n66634 : n66652;
  assign n66654 = pi12 ? n66619 : n66653;
  assign n66655 = pi11 ? n66615 : n66654;
  assign n66656 = pi21 ? n32 : n57667;
  assign n66657 = pi20 ? n66656 : n32;
  assign n66658 = pi19 ? n32 : n66657;
  assign n66659 = pi18 ? n32 : n66658;
  assign n66660 = pi17 ? n32 : n66659;
  assign n66661 = pi16 ? n32 : n66660;
  assign n66662 = pi15 ? n66661 : n16973;
  assign n66663 = pi18 ? n5009 : n36848;
  assign n66664 = pi17 ? n32 : n66663;
  assign n66665 = pi16 ? n32 : n66664;
  assign n66666 = pi15 ? n66665 : n16837;
  assign n66667 = pi14 ? n66662 : n66666;
  assign n66668 = pi19 ? n32 : n7412;
  assign n66669 = pi18 ? n32 : n66668;
  assign n66670 = pi17 ? n32 : n66669;
  assign n66671 = pi16 ? n32 : n66670;
  assign n66672 = pi15 ? n66671 : n37931;
  assign n66673 = pi14 ? n37574 : n66672;
  assign n66674 = pi13 ? n66667 : n66673;
  assign n66675 = pi15 ? n14556 : n14923;
  assign n66676 = pi19 ? n208 : ~n589;
  assign n66677 = pi18 ? n32 : n66676;
  assign n66678 = pi17 ? n32 : n66677;
  assign n66679 = pi16 ? n32 : n66678;
  assign n66680 = pi15 ? n66679 : n66545;
  assign n66681 = pi14 ? n66675 : n66680;
  assign n66682 = pi19 ? n322 : n161;
  assign n66683 = pi18 ? n32 : n66682;
  assign n66684 = pi17 ? n2726 : ~n66683;
  assign n66685 = pi16 ? n2832 : ~n66684;
  assign n66686 = pi17 ? n2726 : ~n24657;
  assign n66687 = pi16 ? n3165 : ~n66686;
  assign n66688 = pi15 ? n66685 : n66687;
  assign n66689 = pi19 ? n507 : n1844;
  assign n66690 = pi18 ? n32 : n66689;
  assign n66691 = pi17 ? n32 : n66690;
  assign n66692 = pi16 ? n32 : n66691;
  assign n66693 = pi15 ? n14917 : n66692;
  assign n66694 = pi14 ? n66688 : n66693;
  assign n66695 = pi13 ? n66681 : n66694;
  assign n66696 = pi12 ? n66674 : n66695;
  assign n66697 = pi19 ? n975 : n32;
  assign n66698 = pi18 ? n32 : n66697;
  assign n66699 = pi17 ? n32 : n66698;
  assign n66700 = pi16 ? n32 : n66699;
  assign n66701 = pi19 ? n1464 : n53;
  assign n66702 = pi18 ? n51606 : n66701;
  assign n66703 = pi17 ? n32 : n66702;
  assign n66704 = pi16 ? n32 : n66703;
  assign n66705 = pi15 ? n66700 : n66704;
  assign n66706 = pi14 ? n25170 : n66705;
  assign n66707 = pi15 ? n23631 : n23484;
  assign n66708 = pi14 ? n66707 : n23160;
  assign n66709 = pi13 ? n66706 : n66708;
  assign n66710 = pi18 ? n5747 : ~n25244;
  assign n66711 = pi17 ? n58032 : n66710;
  assign n66712 = pi16 ? n32 : ~n66711;
  assign n66713 = pi16 ? n2832 : ~n2856;
  assign n66714 = pi15 ? n66712 : n66713;
  assign n66715 = pi19 ? n1757 : n1105;
  assign n66716 = pi18 ? n37954 : ~n66715;
  assign n66717 = pi17 ? n37953 : ~n66716;
  assign n66718 = pi16 ? n2958 : ~n66717;
  assign n66719 = pi17 ? n1718 : ~n24668;
  assign n66720 = pi16 ? n2958 : ~n66719;
  assign n66721 = pi15 ? n66718 : n66720;
  assign n66722 = pi14 ? n66714 : n66721;
  assign n66723 = pi16 ? n4578 : ~n4100;
  assign n66724 = pi17 ? n37965 : ~n4099;
  assign n66725 = pi16 ? n32 : n66724;
  assign n66726 = pi15 ? n66723 : n66725;
  assign n66727 = pi18 ? n46704 : ~n32;
  assign n66728 = pi18 ? n4519 : ~n2627;
  assign n66729 = pi17 ? n66727 : ~n66728;
  assign n66730 = pi16 ? n2958 : ~n66729;
  assign n66731 = pi19 ? n5004 : ~n247;
  assign n66732 = pi20 ? n32 : n8285;
  assign n66733 = pi19 ? n66732 : ~n32;
  assign n66734 = pi18 ? n66731 : ~n66733;
  assign n66735 = pi17 ? n32 : n66734;
  assign n66736 = pi16 ? n32 : n66735;
  assign n66737 = pi15 ? n66730 : n66736;
  assign n66738 = pi14 ? n66726 : n66737;
  assign n66739 = pi13 ? n66722 : n66738;
  assign n66740 = pi12 ? n66709 : n66739;
  assign n66741 = pi11 ? n66696 : n66740;
  assign n66742 = pi10 ? n66655 : n66741;
  assign n66743 = pi09 ? n66602 : n66742;
  assign n66744 = pi14 ? n25861 : n37902;
  assign n66745 = pi13 ? n66744 : n51743;
  assign n66746 = pi20 ? n342 : ~n10446;
  assign n66747 = pi19 ? n32 : n66746;
  assign n66748 = pi18 ? n32 : n66747;
  assign n66749 = pi17 ? n32 : n66748;
  assign n66750 = pi16 ? n32 : n66749;
  assign n66751 = pi15 ? n66750 : n16804;
  assign n66752 = pi14 ? n51745 : n66751;
  assign n66753 = pi13 ? n66752 : n17413;
  assign n66754 = pi12 ? n66745 : n66753;
  assign n66755 = pi14 ? n17178 : n25625;
  assign n66756 = pi13 ? n66755 : n66618;
  assign n66757 = pi19 ? n236 : ~n340;
  assign n66758 = pi18 ? n863 : n66757;
  assign n66759 = pi17 ? n32 : n66758;
  assign n66760 = pi16 ? n32 : n66759;
  assign n66761 = pi15 ? n25814 : n66760;
  assign n66762 = pi19 ? n349 : ~n340;
  assign n66763 = pi18 ? n32 : n66762;
  assign n66764 = pi17 ? n32 : n66763;
  assign n66765 = pi16 ? n32 : n66764;
  assign n66766 = pi19 ? n32 : n66625;
  assign n66767 = pi18 ? n32 : ~n66766;
  assign n66768 = pi17 ? n32 : n66767;
  assign n66769 = pi16 ? n32 : n66768;
  assign n66770 = pi15 ? n66765 : n66769;
  assign n66771 = pi14 ? n66761 : n66770;
  assign n66772 = pi18 ? n66635 : ~n880;
  assign n66773 = pi17 ? n32 : n66772;
  assign n66774 = pi16 ? n32 : n66773;
  assign n66775 = pi18 ? n66639 : ~n880;
  assign n66776 = pi17 ? n32 : n66775;
  assign n66777 = pi16 ? n32 : n66776;
  assign n66778 = pi15 ? n66774 : n66777;
  assign n66779 = pi18 ? n32 : ~n8819;
  assign n66780 = pi17 ? n32 : n66779;
  assign n66781 = pi16 ? n32 : n66780;
  assign n66782 = pi19 ? n531 : ~n12008;
  assign n66783 = pi18 ? n32 : n66782;
  assign n66784 = pi17 ? n32 : n66783;
  assign n66785 = pi16 ? n32 : n66784;
  assign n66786 = pi15 ? n66781 : n66785;
  assign n66787 = pi14 ? n66778 : n66786;
  assign n66788 = pi13 ? n66771 : n66787;
  assign n66789 = pi12 ? n66756 : n66788;
  assign n66790 = pi11 ? n66754 : n66789;
  assign n66791 = pi16 ? n32 : n46792;
  assign n66792 = pi15 ? n16837 : n66791;
  assign n66793 = pi18 ? n5009 : n16970;
  assign n66794 = pi17 ? n32 : n66793;
  assign n66795 = pi16 ? n32 : n66794;
  assign n66796 = pi15 ? n66795 : n16837;
  assign n66797 = pi14 ? n66792 : n66796;
  assign n66798 = pi15 ? n16452 : n16786;
  assign n66799 = pi15 ? n16101 : n38004;
  assign n66800 = pi14 ? n66798 : n66799;
  assign n66801 = pi13 ? n66797 : n66800;
  assign n66802 = pi15 ? n14556 : n14917;
  assign n66803 = pi19 ? n322 : ~n20266;
  assign n66804 = pi18 ? n32 : n66803;
  assign n66805 = pi17 ? n32 : n66804;
  assign n66806 = pi16 ? n32 : n66805;
  assign n66807 = pi15 ? n66679 : n66806;
  assign n66808 = pi14 ? n66802 : n66807;
  assign n66809 = pi17 ? n2726 : ~n23441;
  assign n66810 = pi16 ? n3293 : ~n66809;
  assign n66811 = pi17 ? n2726 : ~n66406;
  assign n66812 = pi16 ? n3165 : ~n66811;
  assign n66813 = pi15 ? n66810 : n66812;
  assign n66814 = pi15 ? n14917 : n22817;
  assign n66815 = pi14 ? n66813 : n66814;
  assign n66816 = pi13 ? n66808 : n66815;
  assign n66817 = pi12 ? n66801 : n66816;
  assign n66818 = pi15 ? n32 : n23730;
  assign n66819 = pi18 ? n51770 : n66701;
  assign n66820 = pi17 ? n32 : n66819;
  assign n66821 = pi16 ? n32 : n66820;
  assign n66822 = pi15 ? n66700 : n66821;
  assign n66823 = pi14 ? n66818 : n66822;
  assign n66824 = pi18 ? n32 : n1190;
  assign n66825 = pi17 ? n32 : n66824;
  assign n66826 = pi20 ? n357 : ~n749;
  assign n66827 = pi19 ? n66826 : n32;
  assign n66828 = pi18 ? n66827 : n32;
  assign n66829 = pi17 ? n66828 : n23248;
  assign n66830 = pi16 ? n66825 : n66829;
  assign n66831 = pi15 ? n66830 : n23250;
  assign n66832 = pi14 ? n63602 : n66831;
  assign n66833 = pi13 ? n66823 : n66832;
  assign n66834 = pi19 ? n322 : n15661;
  assign n66835 = pi18 ? n5747 : ~n66834;
  assign n66836 = pi17 ? n58032 : n66835;
  assign n66837 = pi16 ? n32 : ~n66836;
  assign n66838 = pi16 ? n4578 : ~n2856;
  assign n66839 = pi15 ? n66837 : n66838;
  assign n66840 = pi18 ? n4127 : ~n66715;
  assign n66841 = pi17 ? n37953 : ~n66840;
  assign n66842 = pi16 ? n3588 : ~n66841;
  assign n66843 = pi17 ? n1718 : ~n22823;
  assign n66844 = pi16 ? n3588 : ~n66843;
  assign n66845 = pi15 ? n66842 : n66844;
  assign n66846 = pi14 ? n66839 : n66845;
  assign n66847 = pi17 ? n38032 : ~n2750;
  assign n66848 = pi16 ? n32 : n66847;
  assign n66849 = pi17 ? n38037 : ~n4099;
  assign n66850 = pi16 ? n32 : n66849;
  assign n66851 = pi15 ? n66848 : n66850;
  assign n66852 = pi17 ? n66727 : ~n22937;
  assign n66853 = pi16 ? n3047 : ~n66852;
  assign n66854 = pi19 ? n5004 : ~n3495;
  assign n66855 = pi18 ? n66854 : ~n66733;
  assign n66856 = pi17 ? n32 : n66855;
  assign n66857 = pi16 ? n32 : n66856;
  assign n66858 = pi15 ? n66853 : n66857;
  assign n66859 = pi14 ? n66851 : n66858;
  assign n66860 = pi13 ? n66846 : n66859;
  assign n66861 = pi12 ? n66833 : n66860;
  assign n66862 = pi11 ? n66817 : n66861;
  assign n66863 = pi10 ? n66790 : n66862;
  assign n66864 = pi09 ? n66602 : n66863;
  assign n66865 = pi08 ? n66743 : n66864;
  assign n66866 = pi07 ? n66597 : n66865;
  assign n66867 = pi06 ? n66331 : n66866;
  assign n66868 = pi15 ? n32 : n25902;
  assign n66869 = pi14 ? n32 : n66868;
  assign n66870 = pi13 ? n32 : n66869;
  assign n66871 = pi12 ? n32 : n66870;
  assign n66872 = pi11 ? n32 : n66871;
  assign n66873 = pi10 ? n32 : n66872;
  assign n66874 = pi15 ? n17336 : n25904;
  assign n66875 = pi15 ? n17336 : n17298;
  assign n66876 = pi14 ? n66874 : n66875;
  assign n66877 = pi14 ? n17261 : n51742;
  assign n66878 = pi13 ? n66876 : n66877;
  assign n66879 = pi17 ? n32 : n47188;
  assign n66880 = pi16 ? n32 : n66879;
  assign n66881 = pi15 ? n25997 : n66880;
  assign n66882 = pi14 ? n27734 : n66881;
  assign n66883 = pi13 ? n66882 : n32;
  assign n66884 = pi12 ? n66878 : n66883;
  assign n66885 = pi15 ? n17336 : n17435;
  assign n66886 = pi15 ? n17121 : n17111;
  assign n66887 = pi14 ? n66885 : n66886;
  assign n66888 = pi22 ? n33 : ~n32;
  assign n66889 = pi21 ? n66888 : ~n32;
  assign n66890 = pi20 ? n321 : ~n66889;
  assign n66891 = pi19 ? n32 : n66890;
  assign n66892 = pi18 ? n32 : n66891;
  assign n66893 = pi17 ? n32 : n66892;
  assign n66894 = pi16 ? n32 : n66893;
  assign n66895 = pi15 ? n51644 : n66894;
  assign n66896 = pi14 ? n66895 : n25763;
  assign n66897 = pi13 ? n66887 : n66896;
  assign n66898 = pi19 ? n322 : ~n340;
  assign n66899 = pi18 ? n32 : n66898;
  assign n66900 = pi17 ? n32 : n66899;
  assign n66901 = pi16 ? n32 : n66900;
  assign n66902 = pi15 ? n66489 : n66901;
  assign n66903 = pi19 ? n531 : ~n340;
  assign n66904 = pi18 ? n32 : n66903;
  assign n66905 = pi17 ? n32 : n66904;
  assign n66906 = pi16 ? n32 : n66905;
  assign n66907 = pi19 ? n322 : ~n365;
  assign n66908 = pi18 ? n32 : n66907;
  assign n66909 = pi17 ? n32 : n66908;
  assign n66910 = pi16 ? n32 : n66909;
  assign n66911 = pi15 ? n66906 : n66910;
  assign n66912 = pi14 ? n66902 : n66911;
  assign n66913 = pi19 ? n50776 : ~n531;
  assign n66914 = pi18 ? n4380 : n66913;
  assign n66915 = pi17 ? n32 : n66914;
  assign n66916 = pi16 ? n32 : n66915;
  assign n66917 = pi19 ? n4406 : ~n531;
  assign n66918 = pi18 ? n4722 : n66917;
  assign n66919 = pi17 ? n32 : n66918;
  assign n66920 = pi16 ? n32 : n66919;
  assign n66921 = pi15 ? n66916 : n66920;
  assign n66922 = pi19 ? n1490 : ~n1386;
  assign n66923 = pi18 ? n32 : n66922;
  assign n66924 = pi17 ? n32 : n66923;
  assign n66925 = pi16 ? n32 : n66924;
  assign n66926 = pi19 ? n507 : n176;
  assign n66927 = pi18 ? n32 : n66926;
  assign n66928 = pi17 ? n32 : n66927;
  assign n66929 = pi16 ? n32 : n66928;
  assign n66930 = pi15 ? n66925 : n66929;
  assign n66931 = pi14 ? n66921 : n66930;
  assign n66932 = pi13 ? n66912 : n66931;
  assign n66933 = pi12 ? n66897 : n66932;
  assign n66934 = pi11 ? n66884 : n66933;
  assign n66935 = pi19 ? n236 : ~n16969;
  assign n66936 = pi18 ? n16847 : ~n66935;
  assign n66937 = pi17 ? n32 : n66936;
  assign n66938 = pi16 ? n32 : n66937;
  assign n66939 = pi15 ? n66938 : n16837;
  assign n66940 = pi14 ? n40562 : n66939;
  assign n66941 = pi15 ? n16655 : n16298;
  assign n66942 = pi21 ? n405 : ~n48999;
  assign n66943 = pi20 ? n66942 : n32;
  assign n66944 = pi19 ? n322 : n66943;
  assign n66945 = pi18 ? n32 : n66944;
  assign n66946 = pi17 ? n32 : n66945;
  assign n66947 = pi16 ? n32 : n66946;
  assign n66948 = pi15 ? n66947 : n14917;
  assign n66949 = pi14 ? n66941 : n66948;
  assign n66950 = pi13 ? n66940 : n66949;
  assign n66951 = pi21 ? n32 : n66888;
  assign n66952 = pi20 ? n66951 : ~n32;
  assign n66953 = pi19 ? n507 : ~n66952;
  assign n66954 = pi18 ? n32 : n66953;
  assign n66955 = pi17 ? n51844 : n66954;
  assign n66956 = pi16 ? n32 : n66955;
  assign n66957 = pi15 ? n15244 : n66956;
  assign n66958 = pi14 ? n37927 : n66957;
  assign n66959 = pi17 ? n64832 : ~n37499;
  assign n66960 = pi16 ? n32 : ~n66959;
  assign n66961 = pi20 ? n765 : ~n7839;
  assign n66962 = pi19 ? n66961 : ~n32;
  assign n66963 = pi18 ? n66962 : ~n32;
  assign n66964 = pi17 ? n66963 : ~n25655;
  assign n66965 = pi16 ? n4740 : ~n66964;
  assign n66966 = pi15 ? n66960 : n66965;
  assign n66967 = pi19 ? n507 : n161;
  assign n66968 = pi18 ? n32 : n66967;
  assign n66969 = pi17 ? n32 : n66968;
  assign n66970 = pi16 ? n26424 : n66969;
  assign n66971 = pi15 ? n66970 : n16319;
  assign n66972 = pi14 ? n66966 : n66971;
  assign n66973 = pi13 ? n66958 : n66972;
  assign n66974 = pi12 ? n66950 : n66973;
  assign n66975 = pi20 ? n321 : n448;
  assign n66976 = pi19 ? n32 : ~n66975;
  assign n66977 = pi19 ? n23123 : n32;
  assign n66978 = pi18 ? n66976 : n66977;
  assign n66979 = pi17 ? n32 : n66978;
  assign n66980 = pi16 ? n32 : n66979;
  assign n66981 = pi15 ? n32 : n66980;
  assign n66982 = pi14 ? n26367 : n66981;
  assign n66983 = pi19 ? n594 : n53;
  assign n66984 = pi18 ? n32 : n66983;
  assign n66985 = pi17 ? n32 : n66984;
  assign n66986 = pi16 ? n32 : n66985;
  assign n66987 = pi15 ? n66986 : n32;
  assign n66988 = pi19 ? n247 : ~n32;
  assign n66989 = pi18 ? n66988 : ~n32;
  assign n66990 = pi19 ? n5694 : n358;
  assign n66991 = pi18 ? n32 : n66990;
  assign n66992 = pi17 ? n66989 : ~n66991;
  assign n66993 = pi16 ? n3165 : ~n66992;
  assign n66994 = pi17 ? n36746 : n23158;
  assign n66995 = pi16 ? n32 : n66994;
  assign n66996 = pi15 ? n66993 : n66995;
  assign n66997 = pi14 ? n66987 : n66996;
  assign n66998 = pi13 ? n66982 : n66997;
  assign n66999 = pi18 ? n268 : n8992;
  assign n67000 = pi17 ? n32 : n66999;
  assign n67001 = pi16 ? n32 : ~n67000;
  assign n67002 = pi17 ? n32 : n49934;
  assign n67003 = pi16 ? n3161 : ~n67002;
  assign n67004 = pi15 ? n67001 : n67003;
  assign n67005 = pi18 ? n36119 : ~n25248;
  assign n67006 = pi17 ? n32 : n67005;
  assign n67007 = pi16 ? n3438 : ~n67006;
  assign n67008 = pi17 ? n38122 : ~n22823;
  assign n67009 = pi16 ? n3438 : ~n67008;
  assign n67010 = pi15 ? n67007 : n67009;
  assign n67011 = pi14 ? n67004 : n67010;
  assign n67012 = pi19 ? n56278 : ~n32;
  assign n67013 = pi18 ? n32 : n67012;
  assign n67014 = pi17 ? n38128 : ~n67013;
  assign n67015 = pi16 ? n32 : n67014;
  assign n67016 = pi18 ? n32 : n28019;
  assign n67017 = pi17 ? n32 : n67016;
  assign n67018 = pi16 ? n67017 : ~n4100;
  assign n67019 = pi15 ? n67015 : n67018;
  assign n67020 = pi19 ? n6988 : ~n32;
  assign n67021 = pi18 ? n67020 : ~n32;
  assign n67022 = pi18 ? n4380 : n24540;
  assign n67023 = pi17 ? n67021 : ~n67022;
  assign n67024 = pi16 ? n3438 : ~n67023;
  assign n67025 = pi20 ? n339 : n7880;
  assign n67026 = pi19 ? n67025 : n32;
  assign n67027 = pi18 ? n880 : n67026;
  assign n67028 = pi17 ? n32 : n67027;
  assign n67029 = pi16 ? n32 : n67028;
  assign n67030 = pi15 ? n67024 : n67029;
  assign n67031 = pi14 ? n67019 : n67030;
  assign n67032 = pi13 ? n67011 : n67031;
  assign n67033 = pi12 ? n66998 : n67032;
  assign n67034 = pi11 ? n66974 : n67033;
  assign n67035 = pi10 ? n66934 : n67034;
  assign n67036 = pi09 ? n66873 : n67035;
  assign n67037 = pi15 ? n32 : n25904;
  assign n67038 = pi14 ? n32 : n67037;
  assign n67039 = pi13 ? n32 : n67038;
  assign n67040 = pi12 ? n32 : n67039;
  assign n67041 = pi11 ? n32 : n67040;
  assign n67042 = pi10 ? n32 : n67041;
  assign n67043 = pi14 ? n67037 : n32;
  assign n67044 = pi14 ? n25948 : n51884;
  assign n67045 = pi13 ? n67043 : n67044;
  assign n67046 = pi20 ? n342 : n1629;
  assign n67047 = pi19 ? n32 : n67046;
  assign n67048 = pi18 ? n32 : n67047;
  assign n67049 = pi17 ? n32 : n67048;
  assign n67050 = pi16 ? n32 : n67049;
  assign n67051 = pi15 ? n26201 : n67050;
  assign n67052 = pi20 ? n246 : ~n1940;
  assign n67053 = pi19 ? n32 : n67052;
  assign n67054 = pi18 ? n32 : n67053;
  assign n67055 = pi17 ? n32 : n67054;
  assign n67056 = pi16 ? n32 : n67055;
  assign n67057 = pi15 ? n26479 : n67056;
  assign n67058 = pi14 ? n67051 : n67057;
  assign n67059 = pi14 ? n32 : n25805;
  assign n67060 = pi13 ? n67058 : n67059;
  assign n67061 = pi12 ? n67045 : n67060;
  assign n67062 = pi14 ? n66885 : n17122;
  assign n67063 = pi20 ? n2140 : n481;
  assign n67064 = pi19 ? n32 : n67063;
  assign n67065 = pi18 ? n32 : n67064;
  assign n67066 = pi17 ? n32 : n67065;
  assign n67067 = pi16 ? n32 : n67066;
  assign n67068 = pi15 ? n67067 : n39775;
  assign n67069 = pi14 ? n67068 : n25763;
  assign n67070 = pi13 ? n67062 : n67069;
  assign n67071 = pi15 ? n53803 : n14900;
  assign n67072 = pi19 ? n531 : ~n244;
  assign n67073 = pi18 ? n32 : n67072;
  assign n67074 = pi17 ? n32 : n67073;
  assign n67075 = pi16 ? n32 : n67074;
  assign n67076 = pi15 ? n67075 : n66901;
  assign n67077 = pi14 ? n67071 : n67076;
  assign n67078 = pi19 ? n1248 : ~n365;
  assign n67079 = pi18 ? n4380 : n67078;
  assign n67080 = pi17 ? n32 : n67079;
  assign n67081 = pi16 ? n32 : n67080;
  assign n67082 = pi19 ? n12801 : ~n365;
  assign n67083 = pi18 ? n4722 : n67082;
  assign n67084 = pi17 ? n32 : n67083;
  assign n67085 = pi16 ? n32 : n67084;
  assign n67086 = pi15 ? n67081 : n67085;
  assign n67087 = pi19 ? n1490 : ~n349;
  assign n67088 = pi18 ? n32 : n67087;
  assign n67089 = pi17 ? n32 : n67088;
  assign n67090 = pi16 ? n32 : n67089;
  assign n67091 = pi19 ? n507 : n4670;
  assign n67092 = pi18 ? n32 : n67091;
  assign n67093 = pi17 ? n32 : n67092;
  assign n67094 = pi16 ? n32 : n67093;
  assign n67095 = pi15 ? n67090 : n67094;
  assign n67096 = pi14 ? n67086 : n67095;
  assign n67097 = pi13 ? n67077 : n67096;
  assign n67098 = pi12 ? n67070 : n67097;
  assign n67099 = pi11 ? n67061 : n67098;
  assign n67100 = pi16 ? n32 : n36787;
  assign n67101 = pi15 ? n67100 : n16392;
  assign n67102 = pi14 ? n40562 : n67101;
  assign n67103 = pi15 ? n32 : n26880;
  assign n67104 = pi19 ? n322 : n25448;
  assign n67105 = pi18 ? n32 : n67104;
  assign n67106 = pi17 ? n32 : n67105;
  assign n67107 = pi16 ? n32 : n67106;
  assign n67108 = pi15 ? n67107 : n14917;
  assign n67109 = pi14 ? n67103 : n67108;
  assign n67110 = pi13 ? n67102 : n67109;
  assign n67111 = pi17 ? n51917 : ~n24703;
  assign n67112 = pi16 ? n3283 : ~n67111;
  assign n67113 = pi15 ? n15244 : n67112;
  assign n67114 = pi14 ? n50123 : n67113;
  assign n67115 = pi19 ? n322 : ~n2317;
  assign n67116 = pi18 ? n32 : n67115;
  assign n67117 = pi17 ? n64832 : ~n67116;
  assign n67118 = pi16 ? n32 : ~n67117;
  assign n67119 = pi15 ? n67118 : n25657;
  assign n67120 = pi17 ? n51923 : ~n55401;
  assign n67121 = pi16 ? n3283 : ~n67120;
  assign n67122 = pi15 ? n67121 : n16314;
  assign n67123 = pi14 ? n67119 : n67122;
  assign n67124 = pi13 ? n67114 : n67123;
  assign n67125 = pi12 ? n67110 : n67124;
  assign n67126 = pi19 ? n32 : ~n62571;
  assign n67127 = pi18 ? n67126 : n53495;
  assign n67128 = pi17 ? n32 : n67127;
  assign n67129 = pi16 ? n32 : n67128;
  assign n67130 = pi15 ? n32 : n67129;
  assign n67131 = pi14 ? n26367 : n67130;
  assign n67132 = pi15 ? n66986 : n16108;
  assign n67133 = pi19 ? n5694 : n37;
  assign n67134 = pi18 ? n32 : n67133;
  assign n67135 = pi17 ? n66989 : ~n67134;
  assign n67136 = pi16 ? n3156 : ~n67135;
  assign n67137 = pi19 ? n1818 : n358;
  assign n67138 = pi18 ? n32 : n67137;
  assign n67139 = pi17 ? n36746 : n67138;
  assign n67140 = pi16 ? n3570 : n67139;
  assign n67141 = pi15 ? n67136 : n67140;
  assign n67142 = pi14 ? n67132 : n67141;
  assign n67143 = pi13 ? n67131 : n67142;
  assign n67144 = pi19 ? n5694 : n2614;
  assign n67145 = pi18 ? n268 : n67144;
  assign n67146 = pi17 ? n32 : n67145;
  assign n67147 = pi16 ? n32 : ~n67146;
  assign n67148 = pi18 ? n268 : n2615;
  assign n67149 = pi17 ? n32 : n67148;
  assign n67150 = pi16 ? n32 : ~n67149;
  assign n67151 = pi15 ? n67147 : n67150;
  assign n67152 = pi18 ? n36119 : ~n6147;
  assign n67153 = pi17 ? n3557 : ~n67152;
  assign n67154 = pi16 ? n32 : n67153;
  assign n67155 = pi17 ? n38183 : n14578;
  assign n67156 = pi16 ? n32 : n67155;
  assign n67157 = pi15 ? n67154 : n67156;
  assign n67158 = pi14 ? n67151 : n67157;
  assign n67159 = pi18 ? n32 : n54054;
  assign n67160 = pi17 ? n38128 : ~n67159;
  assign n67161 = pi16 ? n32 : n67160;
  assign n67162 = pi17 ? n1028 : ~n4099;
  assign n67163 = pi16 ? n32 : n67162;
  assign n67164 = pi15 ? n67161 : n67163;
  assign n67165 = pi18 ? n48299 : n32;
  assign n67166 = pi17 ? n67165 : n67022;
  assign n67167 = pi16 ? n32 : n67166;
  assign n67168 = pi18 ? n880 : ~n7278;
  assign n67169 = pi17 ? n32 : n67168;
  assign n67170 = pi16 ? n32 : n67169;
  assign n67171 = pi15 ? n67167 : n67170;
  assign n67172 = pi14 ? n67164 : n67171;
  assign n67173 = pi13 ? n67158 : n67172;
  assign n67174 = pi12 ? n67143 : n67173;
  assign n67175 = pi11 ? n67125 : n67174;
  assign n67176 = pi10 ? n67099 : n67175;
  assign n67177 = pi09 ? n67042 : n67176;
  assign n67178 = pi08 ? n67036 : n67177;
  assign n67179 = pi15 ? n32 : n38209;
  assign n67180 = pi14 ? n32 : n67179;
  assign n67181 = pi13 ? n32 : n67180;
  assign n67182 = pi12 ? n32 : n67181;
  assign n67183 = pi11 ? n32 : n67182;
  assign n67184 = pi10 ? n32 : n67183;
  assign n67185 = pi15 ? n25904 : n25988;
  assign n67186 = pi14 ? n67185 : n38053;
  assign n67187 = pi15 ? n25948 : n17121;
  assign n67188 = pi14 ? n67187 : n51884;
  assign n67189 = pi13 ? n67186 : n67188;
  assign n67190 = pi15 ? n17121 : n40426;
  assign n67191 = pi15 ? n26479 : n17261;
  assign n67192 = pi14 ? n67190 : n67191;
  assign n67193 = pi13 ? n67192 : n51747;
  assign n67194 = pi12 ? n67189 : n67193;
  assign n67195 = pi15 ? n25904 : n17298;
  assign n67196 = pi14 ? n67195 : n25805;
  assign n67197 = pi14 ? n27733 : n16804;
  assign n67198 = pi13 ? n67196 : n67197;
  assign n67199 = pi15 ? n16044 : n14900;
  assign n67200 = pi15 ? n14900 : n66901;
  assign n67201 = pi14 ? n67199 : n67200;
  assign n67202 = pi19 ? n8818 : ~n365;
  assign n67203 = pi18 ? n4722 : n67202;
  assign n67204 = pi17 ? n32 : n67203;
  assign n67205 = pi16 ? n32 : n67204;
  assign n67206 = pi15 ? n66910 : n67205;
  assign n67207 = pi15 ? n15244 : n17036;
  assign n67208 = pi14 ? n67206 : n67207;
  assign n67209 = pi13 ? n67201 : n67208;
  assign n67210 = pi12 ? n67198 : n67209;
  assign n67211 = pi11 ? n67194 : n67210;
  assign n67212 = pi19 ? n236 : ~n4491;
  assign n67213 = pi18 ? n16847 : ~n67212;
  assign n67214 = pi17 ? n32 : n67213;
  assign n67215 = pi16 ? n32 : n67214;
  assign n67216 = pi15 ? n67215 : n17039;
  assign n67217 = pi14 ? n51428 : n67216;
  assign n67218 = pi15 ? n16899 : n16298;
  assign n67219 = pi19 ? n322 : n10879;
  assign n67220 = pi18 ? n32 : n67219;
  assign n67221 = pi17 ? n32 : n67220;
  assign n67222 = pi16 ? n32 : n67221;
  assign n67223 = pi19 ? n322 : ~n58188;
  assign n67224 = pi18 ? n32 : n67223;
  assign n67225 = pi17 ? n32 : n67224;
  assign n67226 = pi16 ? n32 : n67225;
  assign n67227 = pi15 ? n67222 : n67226;
  assign n67228 = pi14 ? n67218 : n67227;
  assign n67229 = pi13 ? n67217 : n67228;
  assign n67230 = pi19 ? n236 : ~n47180;
  assign n67231 = pi20 ? n1611 : ~n1331;
  assign n67232 = pi20 ? n1611 : n371;
  assign n67233 = pi19 ? n67231 : n67232;
  assign n67234 = pi18 ? n67230 : ~n67233;
  assign n67235 = pi17 ? n67234 : n24703;
  assign n67236 = pi16 ? n32 : n67235;
  assign n67237 = pi15 ? n24705 : n67236;
  assign n67238 = pi14 ? n64615 : n67237;
  assign n67239 = pi19 ? n507 : ~n14552;
  assign n67240 = pi18 ? n32 : n67239;
  assign n67241 = pi17 ? n36789 : n67240;
  assign n67242 = pi16 ? n32 : n67241;
  assign n67243 = pi15 ? n67242 : n15357;
  assign n67244 = pi19 ? n594 : n3495;
  assign n67245 = pi18 ? n32 : n67244;
  assign n67246 = pi17 ? n32 : n67245;
  assign n67247 = pi16 ? n32 : n67246;
  assign n67248 = pi15 ? n67247 : n16314;
  assign n67249 = pi14 ? n67243 : n67248;
  assign n67250 = pi13 ? n67238 : n67249;
  assign n67251 = pi12 ? n67229 : n67250;
  assign n67252 = pi19 ? n2141 : n1844;
  assign n67253 = pi18 ? n32 : n67252;
  assign n67254 = pi17 ? n32 : n67253;
  assign n67255 = pi16 ? n32 : n67254;
  assign n67256 = pi15 ? n16105 : n67255;
  assign n67257 = pi19 ? n644 : ~n813;
  assign n67258 = pi18 ? n51851 : n67257;
  assign n67259 = pi17 ? n32 : n67258;
  assign n67260 = pi16 ? n32 : n67259;
  assign n67261 = pi15 ? n23574 : n67260;
  assign n67262 = pi14 ? n67256 : n67261;
  assign n67263 = pi15 ? n23340 : n66986;
  assign n67264 = pi19 ? n589 : n3692;
  assign n67265 = pi18 ? n67264 : n32;
  assign n67266 = pi20 ? n32 : ~n1324;
  assign n67267 = pi19 ? n67266 : n53;
  assign n67268 = pi18 ? n32 : n67267;
  assign n67269 = pi17 ? n67265 : n67268;
  assign n67270 = pi16 ? n32 : n67269;
  assign n67271 = pi19 ? n4518 : ~n236;
  assign n67272 = pi18 ? n32 : n67271;
  assign n67273 = pi17 ? n36746 : n67272;
  assign n67274 = pi16 ? n32 : n67273;
  assign n67275 = pi15 ? n67270 : n67274;
  assign n67276 = pi14 ? n67263 : n67275;
  assign n67277 = pi13 ? n67262 : n67276;
  assign n67278 = pi17 ? n3715 : ~n8989;
  assign n67279 = pi16 ? n32 : n67278;
  assign n67280 = pi19 ? n4491 : n2614;
  assign n67281 = pi18 ? n32 : n67280;
  assign n67282 = pi17 ? n3715 : ~n67281;
  assign n67283 = pi16 ? n32 : n67282;
  assign n67284 = pi15 ? n67279 : n67283;
  assign n67285 = pi17 ? n3704 : ~n67152;
  assign n67286 = pi16 ? n32 : n67285;
  assign n67287 = pi15 ? n67286 : n14580;
  assign n67288 = pi14 ? n67284 : n67287;
  assign n67289 = pi19 ? n1464 : n1105;
  assign n67290 = pi18 ? n32 : n67289;
  assign n67291 = pi17 ? n1697 : ~n67290;
  assign n67292 = pi16 ? n32 : n67291;
  assign n67293 = pi20 ? n1368 : n266;
  assign n67294 = pi19 ? n67293 : ~n32;
  assign n67295 = pi18 ? n32 : n67294;
  assign n67296 = pi17 ? n4041 : ~n67295;
  assign n67297 = pi16 ? n32 : n67296;
  assign n67298 = pi15 ? n67292 : n67297;
  assign n67299 = pi17 ? n28440 : n24668;
  assign n67300 = pi16 ? n32 : n67299;
  assign n67301 = pi20 ? n321 : n1385;
  assign n67302 = pi19 ? n67301 : n32;
  assign n67303 = pi18 ? n880 : n67302;
  assign n67304 = pi17 ? n32 : n67303;
  assign n67305 = pi16 ? n32 : n67304;
  assign n67306 = pi15 ? n67300 : n67305;
  assign n67307 = pi14 ? n67298 : n67306;
  assign n67308 = pi13 ? n67288 : n67307;
  assign n67309 = pi12 ? n67277 : n67308;
  assign n67310 = pi11 ? n67251 : n67309;
  assign n67311 = pi10 ? n67211 : n67310;
  assign n67312 = pi09 ? n67184 : n67311;
  assign n67313 = pi15 ? n32 : n25984;
  assign n67314 = pi14 ? n32 : n67313;
  assign n67315 = pi13 ? n32 : n67314;
  assign n67316 = pi12 ? n32 : n67315;
  assign n67317 = pi11 ? n32 : n67316;
  assign n67318 = pi10 ? n32 : n67317;
  assign n67319 = pi14 ? n26031 : n67037;
  assign n67320 = pi14 ? n17216 : n52055;
  assign n67321 = pi13 ? n67319 : n67320;
  assign n67322 = pi15 ? n17121 : n40558;
  assign n67323 = pi15 ? n16824 : n25948;
  assign n67324 = pi14 ? n67322 : n67323;
  assign n67325 = pi13 ? n67324 : n51747;
  assign n67326 = pi12 ? n67321 : n67325;
  assign n67327 = pi19 ? n32 : n13062;
  assign n67328 = pi18 ? n32 : n67327;
  assign n67329 = pi17 ? n32 : n67328;
  assign n67330 = pi16 ? n32 : n67329;
  assign n67331 = pi15 ? n67330 : n14876;
  assign n67332 = pi14 ? n67331 : n14876;
  assign n67333 = pi19 ? n11108 : ~n340;
  assign n67334 = pi18 ? n4722 : n67333;
  assign n67335 = pi17 ? n32 : n67334;
  assign n67336 = pi16 ? n32 : n67335;
  assign n67337 = pi15 ? n66901 : n67336;
  assign n67338 = pi19 ? n507 : ~n7993;
  assign n67339 = pi18 ? n32 : n67338;
  assign n67340 = pi17 ? n32 : n67339;
  assign n67341 = pi16 ? n32 : n67340;
  assign n67342 = pi15 ? n67341 : n16913;
  assign n67343 = pi14 ? n67337 : n67342;
  assign n67344 = pi13 ? n67332 : n67343;
  assign n67345 = pi12 ? n67198 : n67344;
  assign n67346 = pi11 ? n67326 : n67345;
  assign n67347 = pi20 ? n2077 : ~n141;
  assign n67348 = pi19 ? n32 : n67347;
  assign n67349 = pi18 ? n32 : n67348;
  assign n67350 = pi17 ? n32 : n67349;
  assign n67351 = pi16 ? n32 : n67350;
  assign n67352 = pi15 ? n16832 : n67351;
  assign n67353 = pi15 ? n67100 : n17039;
  assign n67354 = pi14 ? n67352 : n67353;
  assign n67355 = pi15 ? n16392 : n16298;
  assign n67356 = pi19 ? n322 : n39565;
  assign n67357 = pi18 ? n32 : n67356;
  assign n67358 = pi17 ? n32 : n67357;
  assign n67359 = pi16 ? n32 : n67358;
  assign n67360 = pi19 ? n322 : ~n1265;
  assign n67361 = pi18 ? n32 : n67360;
  assign n67362 = pi17 ? n32 : n67361;
  assign n67363 = pi16 ? n32 : n67362;
  assign n67364 = pi15 ? n67359 : n67363;
  assign n67365 = pi14 ? n67355 : n67364;
  assign n67366 = pi13 ? n67354 : n67365;
  assign n67367 = pi19 ? n589 : ~n47180;
  assign n67368 = pi20 ? n220 : n1331;
  assign n67369 = pi19 ? n67368 : ~n67232;
  assign n67370 = pi18 ? n67367 : n67369;
  assign n67371 = pi17 ? n67370 : n15228;
  assign n67372 = pi16 ? n32 : n67371;
  assign n67373 = pi15 ? n15230 : n67372;
  assign n67374 = pi14 ? n64615 : n67373;
  assign n67375 = pi19 ? n32 : n57780;
  assign n67376 = pi18 ? n32 : n67375;
  assign n67377 = pi17 ? n32 : n67376;
  assign n67378 = pi16 ? n32 : n67377;
  assign n67379 = pi15 ? n67247 : n67378;
  assign n67380 = pi14 ? n67243 : n67379;
  assign n67381 = pi13 ? n67374 : n67380;
  assign n67382 = pi12 ? n67366 : n67381;
  assign n67383 = pi16 ? n32 : n66969;
  assign n67384 = pi15 ? n16105 : n67383;
  assign n67385 = pi18 ? n51851 : n20164;
  assign n67386 = pi17 ? n32 : n67385;
  assign n67387 = pi16 ? n32 : n67386;
  assign n67388 = pi15 ? n16105 : n67387;
  assign n67389 = pi14 ? n67384 : n67388;
  assign n67390 = pi19 ? n594 : ~n821;
  assign n67391 = pi18 ? n32 : n67390;
  assign n67392 = pi17 ? n32 : n67391;
  assign n67393 = pi16 ? n32 : n67392;
  assign n67394 = pi20 ? n1839 : ~n314;
  assign n67395 = pi19 ? n67394 : n16304;
  assign n67396 = pi18 ? n67395 : n32;
  assign n67397 = pi17 ? n67396 : n66984;
  assign n67398 = pi16 ? n32 : n67397;
  assign n67399 = pi15 ? n67393 : n67398;
  assign n67400 = pi19 ? n2848 : n3692;
  assign n67401 = pi18 ? n67400 : n32;
  assign n67402 = pi17 ? n67401 : n67268;
  assign n67403 = pi16 ? n32 : n67402;
  assign n67404 = pi15 ? n67403 : n67274;
  assign n67405 = pi14 ? n67399 : n67404;
  assign n67406 = pi13 ? n67389 : n67405;
  assign n67407 = pi17 ? n3553 : ~n8989;
  assign n67408 = pi16 ? n32 : n67407;
  assign n67409 = pi17 ? n3553 : ~n2616;
  assign n67410 = pi16 ? n32 : n67409;
  assign n67411 = pi15 ? n67408 : n67410;
  assign n67412 = pi18 ? n36119 : ~n25732;
  assign n67413 = pi17 ? n3855 : ~n67412;
  assign n67414 = pi16 ? n32 : n67413;
  assign n67415 = pi15 ? n67414 : n14580;
  assign n67416 = pi14 ? n67411 : n67415;
  assign n67417 = pi17 ? n1697 : ~n7931;
  assign n67418 = pi16 ? n32 : n67417;
  assign n67419 = pi19 ? n53582 : ~n32;
  assign n67420 = pi18 ? n32 : n67419;
  assign n67421 = pi17 ? n4037 : ~n67420;
  assign n67422 = pi16 ? n32 : n67421;
  assign n67423 = pi15 ? n67418 : n67422;
  assign n67424 = pi14 ? n67423 : n67306;
  assign n67425 = pi13 ? n67416 : n67424;
  assign n67426 = pi12 ? n67406 : n67425;
  assign n67427 = pi11 ? n67382 : n67426;
  assign n67428 = pi10 ? n67346 : n67427;
  assign n67429 = pi09 ? n67318 : n67428;
  assign n67430 = pi08 ? n67312 : n67429;
  assign n67431 = pi07 ? n67178 : n67430;
  assign n67432 = pi12 ? n32 : n26135;
  assign n67433 = pi11 ? n32 : n67432;
  assign n67434 = pi10 ? n32 : n67433;
  assign n67435 = pi14 ? n26097 : n67313;
  assign n67436 = pi15 ? n25904 : n26322;
  assign n67437 = pi14 ? n67436 : n52128;
  assign n67438 = pi13 ? n67435 : n67437;
  assign n67439 = pi15 ? n17216 : n25904;
  assign n67440 = pi14 ? n27057 : n67439;
  assign n67441 = pi13 ? n67440 : n32;
  assign n67442 = pi12 ? n67438 : n67441;
  assign n67443 = pi15 ? n25904 : n17367;
  assign n67444 = pi14 ? n38290 : n67443;
  assign n67445 = pi15 ? n25997 : n26201;
  assign n67446 = pi19 ? n32 : n21493;
  assign n67447 = pi18 ? n32 : n67446;
  assign n67448 = pi17 ? n32 : n67447;
  assign n67449 = pi16 ? n32 : n67448;
  assign n67450 = pi15 ? n16804 : n67449;
  assign n67451 = pi14 ? n67445 : n67450;
  assign n67452 = pi13 ? n67444 : n67451;
  assign n67453 = pi17 ? n32 : n52189;
  assign n67454 = pi16 ? n32 : n67453;
  assign n67455 = pi15 ? n67449 : n67454;
  assign n67456 = pi19 ? n507 : ~n804;
  assign n67457 = pi18 ? n32 : n67456;
  assign n67458 = pi17 ? n32 : n67457;
  assign n67459 = pi16 ? n32 : n67458;
  assign n67460 = pi20 ? n67 : n207;
  assign n67461 = pi19 ? n32 : ~n67460;
  assign n67462 = pi18 ? n32 : n67461;
  assign n67463 = pi17 ? n32 : n67462;
  assign n67464 = pi16 ? n32 : n67463;
  assign n67465 = pi15 ? n67459 : n67464;
  assign n67466 = pi14 ? n67455 : n67465;
  assign n67467 = pi19 ? n32 : ~n244;
  assign n67468 = pi18 ? n32 : n67467;
  assign n67469 = pi17 ? n32 : n67468;
  assign n67470 = pi16 ? n32 : n67469;
  assign n67471 = pi19 ? n20006 : ~n429;
  assign n67472 = pi18 ? n32 : n67471;
  assign n67473 = pi17 ? n32 : n67472;
  assign n67474 = pi16 ? n32 : n67473;
  assign n67475 = pi15 ? n67470 : n67474;
  assign n67476 = pi15 ? n16105 : n17066;
  assign n67477 = pi14 ? n67475 : n67476;
  assign n67478 = pi13 ? n67466 : n67477;
  assign n67479 = pi12 ? n67452 : n67478;
  assign n67480 = pi11 ? n67442 : n67479;
  assign n67481 = pi15 ? n17066 : n17188;
  assign n67482 = pi14 ? n67481 : n17039;
  assign n67483 = pi19 ? n322 : n19847;
  assign n67484 = pi18 ? n32 : n67483;
  assign n67485 = pi17 ? n32 : n67484;
  assign n67486 = pi16 ? n32 : n67485;
  assign n67487 = pi15 ? n67486 : n16606;
  assign n67488 = pi14 ? n67487 : n52242;
  assign n67489 = pi13 ? n67482 : n67488;
  assign n67490 = pi15 ? n37182 : n24367;
  assign n67491 = pi19 ? n32 : ~n3507;
  assign n67492 = pi18 ? n32 : n67491;
  assign n67493 = pi17 ? n32 : n67492;
  assign n67494 = pi16 ? n32 : n67493;
  assign n67495 = pi19 ? n531 : ~n39054;
  assign n67496 = pi19 ? n18728 : n4126;
  assign n67497 = pi18 ? n67495 : n67496;
  assign n67498 = pi18 ? n248 : n24697;
  assign n67499 = pi17 ? n67497 : n67498;
  assign n67500 = pi16 ? n32 : n67499;
  assign n67501 = pi15 ? n67494 : n67500;
  assign n67502 = pi14 ? n67490 : n67501;
  assign n67503 = pi18 ? n32 : n52163;
  assign n67504 = pi17 ? n32 : n67503;
  assign n67505 = pi16 ? n32 : n67504;
  assign n67506 = pi15 ? n67505 : n24640;
  assign n67507 = pi21 ? n631 : ~n124;
  assign n67508 = pi20 ? n67507 : ~n32;
  assign n67509 = pi19 ? n507 : ~n67508;
  assign n67510 = pi18 ? n32 : n67509;
  assign n67511 = pi17 ? n32 : n67510;
  assign n67512 = pi16 ? n32 : n67511;
  assign n67513 = pi15 ? n24367 : n67512;
  assign n67514 = pi14 ? n67506 : n67513;
  assign n67515 = pi13 ? n67502 : n67514;
  assign n67516 = pi12 ? n67489 : n67515;
  assign n67517 = pi20 ? n38686 : n32;
  assign n67518 = pi19 ? n507 : n67517;
  assign n67519 = pi18 ? n32 : n67518;
  assign n67520 = pi17 ? n32 : n67519;
  assign n67521 = pi16 ? n32 : n67520;
  assign n67522 = pi15 ? n40057 : n67521;
  assign n67523 = pi19 ? n32 : ~n6683;
  assign n67524 = pi18 ? n32 : n67523;
  assign n67525 = pi17 ? n32 : n67524;
  assign n67526 = pi16 ? n32 : n67525;
  assign n67527 = pi15 ? n24582 : n67526;
  assign n67528 = pi14 ? n67522 : n67527;
  assign n67529 = pi19 ? n1464 : ~n20022;
  assign n67530 = pi18 ? n32 : n67529;
  assign n67531 = pi17 ? n32 : n67530;
  assign n67532 = pi16 ? n32 : n67531;
  assign n67533 = pi20 ? n101 : ~n342;
  assign n67534 = pi19 ? n67533 : ~n32;
  assign n67535 = pi18 ? n67534 : ~n350;
  assign n67536 = pi19 ? n322 : n19892;
  assign n67537 = pi18 ? n32 : n67536;
  assign n67538 = pi17 ? n67535 : n67537;
  assign n67539 = pi16 ? n32 : n67538;
  assign n67540 = pi15 ? n67532 : n67539;
  assign n67541 = pi19 ? n67533 : ~n24218;
  assign n67542 = pi18 ? n67541 : n32;
  assign n67543 = pi17 ? n67542 : n53496;
  assign n67544 = pi16 ? n32 : n67543;
  assign n67545 = pi19 ? n221 : ~n1941;
  assign n67546 = pi18 ? n32 : n67545;
  assign n67547 = pi17 ? n50213 : n67546;
  assign n67548 = pi16 ? n32 : n67547;
  assign n67549 = pi15 ? n67544 : n67548;
  assign n67550 = pi14 ? n67540 : n67549;
  assign n67551 = pi13 ? n67528 : n67550;
  assign n67552 = pi19 ? n322 : n1941;
  assign n67553 = pi18 ? n32 : n67552;
  assign n67554 = pi17 ? n4034 : ~n67553;
  assign n67555 = pi16 ? n32 : n67554;
  assign n67556 = pi19 ? n2025 : ~n5626;
  assign n67557 = pi18 ? n32 : n67556;
  assign n67558 = pi17 ? n4034 : ~n67557;
  assign n67559 = pi16 ? n32 : n67558;
  assign n67560 = pi15 ? n67555 : n67559;
  assign n67561 = pi18 ? n23073 : ~n25244;
  assign n67562 = pi17 ? n38384 : ~n67561;
  assign n67563 = pi16 ? n32 : n67562;
  assign n67564 = pi15 ? n67563 : n14580;
  assign n67565 = pi14 ? n67560 : n67564;
  assign n67566 = pi19 ? n32 : ~n17194;
  assign n67567 = pi18 ? n67566 : ~n32;
  assign n67568 = pi17 ? n67567 : ~n2623;
  assign n67569 = pi16 ? n32 : n67568;
  assign n67570 = pi21 ? n1939 : ~n309;
  assign n67571 = pi20 ? n32 : n67570;
  assign n67572 = pi19 ? n67571 : ~n28686;
  assign n67573 = pi18 ? n67572 : n38402;
  assign n67574 = pi19 ? n38407 : ~n1105;
  assign n67575 = pi18 ? n38406 : n67574;
  assign n67576 = pi17 ? n67573 : n67575;
  assign n67577 = pi16 ? n32 : n67576;
  assign n67578 = pi15 ? n67569 : n67577;
  assign n67579 = pi18 ? n21138 : n32;
  assign n67580 = pi17 ? n67579 : n34844;
  assign n67581 = pi16 ? n32 : n67580;
  assign n67582 = pi19 ? n32 : ~n52205;
  assign n67583 = pi18 ? n67582 : ~n6059;
  assign n67584 = pi18 ? n32 : n65572;
  assign n67585 = pi17 ? n67583 : ~n67584;
  assign n67586 = pi16 ? n32 : n67585;
  assign n67587 = pi15 ? n67581 : n67586;
  assign n67588 = pi14 ? n67578 : n67587;
  assign n67589 = pi13 ? n67565 : n67588;
  assign n67590 = pi12 ? n67551 : n67589;
  assign n67591 = pi11 ? n67516 : n67590;
  assign n67592 = pi10 ? n67480 : n67591;
  assign n67593 = pi09 ? n67434 : n67592;
  assign n67594 = pi13 ? n67435 : n52226;
  assign n67595 = pi15 ? n32 : n26310;
  assign n67596 = pi15 ? n16850 : n25984;
  assign n67597 = pi14 ? n67595 : n67596;
  assign n67598 = pi14 ? n32 : n26034;
  assign n67599 = pi13 ? n67597 : n67598;
  assign n67600 = pi12 ? n67594 : n67599;
  assign n67601 = pi15 ? n25904 : n17121;
  assign n67602 = pi14 ? n38290 : n67601;
  assign n67603 = pi15 ? n25997 : n17061;
  assign n67604 = pi15 ? n25997 : n67449;
  assign n67605 = pi14 ? n67603 : n67604;
  assign n67606 = pi13 ? n67602 : n67605;
  assign n67607 = pi19 ? n32 : ~n1969;
  assign n67608 = pi18 ? n32 : n67607;
  assign n67609 = pi17 ? n32 : n67608;
  assign n67610 = pi16 ? n32 : n67609;
  assign n67611 = pi15 ? n16352 : n67610;
  assign n67612 = pi19 ? n507 : ~n1394;
  assign n67613 = pi18 ? n32 : n67612;
  assign n67614 = pi17 ? n32 : n67613;
  assign n67615 = pi16 ? n32 : n67614;
  assign n67616 = pi19 ? n32 : ~n2168;
  assign n67617 = pi18 ? n32 : n67616;
  assign n67618 = pi17 ? n32 : n67617;
  assign n67619 = pi16 ? n32 : n67618;
  assign n67620 = pi15 ? n67615 : n67619;
  assign n67621 = pi14 ? n67611 : n67620;
  assign n67622 = pi19 ? n32 : ~n14065;
  assign n67623 = pi18 ? n32 : n67622;
  assign n67624 = pi17 ? n32 : n67623;
  assign n67625 = pi16 ? n32 : n67624;
  assign n67626 = pi15 ? n67625 : n67474;
  assign n67627 = pi19 ? n32 : n59936;
  assign n67628 = pi18 ? n32 : n67627;
  assign n67629 = pi17 ? n32 : n67628;
  assign n67630 = pi16 ? n32 : n67629;
  assign n67631 = pi19 ? n32 : n21969;
  assign n67632 = pi18 ? n32 : n67631;
  assign n67633 = pi17 ? n32 : n67632;
  assign n67634 = pi16 ? n32 : n67633;
  assign n67635 = pi15 ? n67630 : n67634;
  assign n67636 = pi14 ? n67626 : n67635;
  assign n67637 = pi13 ? n67621 : n67636;
  assign n67638 = pi12 ? n67606 : n67637;
  assign n67639 = pi11 ? n67600 : n67638;
  assign n67640 = pi14 ? n17412 : n17090;
  assign n67641 = pi15 ? n67486 : n38447;
  assign n67642 = pi15 ? n27304 : n15633;
  assign n67643 = pi14 ? n67641 : n67642;
  assign n67644 = pi13 ? n67640 : n67643;
  assign n67645 = pi15 ? n24511 : n24237;
  assign n67646 = pi19 ? n750 : ~n39054;
  assign n67647 = pi18 ? n67646 : n67496;
  assign n67648 = pi18 ? n248 : n27525;
  assign n67649 = pi17 ? n67647 : n67648;
  assign n67650 = pi16 ? n32 : n67649;
  assign n67651 = pi15 ? n27528 : n67650;
  assign n67652 = pi14 ? n67645 : n67651;
  assign n67653 = pi19 ? n4342 : ~n766;
  assign n67654 = pi18 ? n32 : n67653;
  assign n67655 = pi17 ? n32 : n67654;
  assign n67656 = pi16 ? n32 : n67655;
  assign n67657 = pi15 ? n67656 : n64148;
  assign n67658 = pi20 ? n41008 : n32;
  assign n67659 = pi19 ? n32 : n67658;
  assign n67660 = pi18 ? n32 : n67659;
  assign n67661 = pi17 ? n32 : n67660;
  assign n67662 = pi16 ? n32 : n67661;
  assign n67663 = pi19 ? n507 : ~n54737;
  assign n67664 = pi18 ? n32 : n67663;
  assign n67665 = pi17 ? n32 : n67664;
  assign n67666 = pi16 ? n32 : n67665;
  assign n67667 = pi15 ? n67662 : n67666;
  assign n67668 = pi14 ? n67657 : n67667;
  assign n67669 = pi13 ? n67652 : n67668;
  assign n67670 = pi12 ? n67644 : n67669;
  assign n67671 = pi21 ? n1009 : ~n140;
  assign n67672 = pi20 ? n67671 : n32;
  assign n67673 = pi19 ? n507 : n67672;
  assign n67674 = pi18 ? n32 : n67673;
  assign n67675 = pi17 ? n32 : n67674;
  assign n67676 = pi16 ? n32 : n67675;
  assign n67677 = pi15 ? n40057 : n67676;
  assign n67678 = pi14 ? n67677 : n67527;
  assign n67679 = pi20 ? n32 : n10862;
  assign n67680 = pi19 ? n67679 : ~n32;
  assign n67681 = pi18 ? n67680 : ~n350;
  assign n67682 = pi17 ? n67681 : n67537;
  assign n67683 = pi16 ? n32 : n67682;
  assign n67684 = pi15 ? n67532 : n67683;
  assign n67685 = pi19 ? n67679 : ~n24218;
  assign n67686 = pi18 ? n67685 : n32;
  assign n67687 = pi17 ? n67686 : n53496;
  assign n67688 = pi16 ? n32 : n67687;
  assign n67689 = pi15 ? n67688 : n67548;
  assign n67690 = pi14 ? n67684 : n67689;
  assign n67691 = pi13 ? n67678 : n67690;
  assign n67692 = pi17 ? n4515 : ~n67553;
  assign n67693 = pi16 ? n32 : n67692;
  assign n67694 = pi19 ? n208 : ~n5626;
  assign n67695 = pi18 ? n32 : n67694;
  assign n67696 = pi17 ? n4515 : ~n67695;
  assign n67697 = pi16 ? n32 : n67696;
  assign n67698 = pi15 ? n67693 : n67697;
  assign n67699 = pi17 ? n38459 : ~n67561;
  assign n67700 = pi16 ? n32 : n67699;
  assign n67701 = pi15 ? n67700 : n14580;
  assign n67702 = pi14 ? n67698 : n67701;
  assign n67703 = pi19 ? n32 : ~n38468;
  assign n67704 = pi18 ? n67703 : ~n32;
  assign n67705 = pi17 ? n67704 : ~n2750;
  assign n67706 = pi16 ? n32 : n67705;
  assign n67707 = pi19 ? n507 : ~n28686;
  assign n67708 = pi18 ? n67707 : n38402;
  assign n67709 = pi17 ? n67708 : n67575;
  assign n67710 = pi16 ? n32 : n67709;
  assign n67711 = pi15 ? n67706 : n67710;
  assign n67712 = pi19 ? n32 : ~n30681;
  assign n67713 = pi18 ? n67712 : ~n6059;
  assign n67714 = pi17 ? n67713 : ~n67584;
  assign n67715 = pi16 ? n32 : n67714;
  assign n67716 = pi15 ? n34846 : n67715;
  assign n67717 = pi14 ? n67711 : n67716;
  assign n67718 = pi13 ? n67702 : n67717;
  assign n67719 = pi12 ? n67691 : n67718;
  assign n67720 = pi11 ? n67670 : n67719;
  assign n67721 = pi10 ? n67639 : n67720;
  assign n67722 = pi09 ? n67434 : n67721;
  assign n67723 = pi08 ? n67593 : n67722;
  assign n67724 = pi15 ? n26225 : n26183;
  assign n67725 = pi14 ? n32 : n67724;
  assign n67726 = pi13 ? n32 : n67725;
  assign n67727 = pi12 ? n32 : n67726;
  assign n67728 = pi11 ? n32 : n67727;
  assign n67729 = pi10 ? n32 : n67728;
  assign n67730 = pi14 ? n26226 : n17348;
  assign n67731 = pi13 ? n67730 : n52301;
  assign n67732 = pi15 ? n25904 : n26310;
  assign n67733 = pi14 ? n67732 : n26144;
  assign n67734 = pi13 ? n67733 : n32;
  assign n67735 = pi12 ? n67731 : n67734;
  assign n67736 = pi15 ? n17348 : n17431;
  assign n67737 = pi19 ? n32 : n61517;
  assign n67738 = pi18 ? n32 : n67737;
  assign n67739 = pi17 ? n32 : n67738;
  assign n67740 = pi16 ? n32 : n67739;
  assign n67741 = pi15 ? n67740 : n17056;
  assign n67742 = pi14 ? n67736 : n67741;
  assign n67743 = pi15 ? n26479 : n16352;
  assign n67744 = pi14 ? n26479 : n67743;
  assign n67745 = pi13 ? n67742 : n67744;
  assign n67746 = pi15 ? n54872 : n67330;
  assign n67747 = pi15 ? n67459 : n67454;
  assign n67748 = pi14 ? n67746 : n67747;
  assign n67749 = pi19 ? n32 : ~n1348;
  assign n67750 = pi18 ? n32 : n67749;
  assign n67751 = pi17 ? n32 : n67750;
  assign n67752 = pi16 ? n32 : n67751;
  assign n67753 = pi15 ? n67752 : n50513;
  assign n67754 = pi15 ? n25556 : n25814;
  assign n67755 = pi14 ? n67753 : n67754;
  assign n67756 = pi13 ? n67748 : n67755;
  assign n67757 = pi12 ? n67745 : n67756;
  assign n67758 = pi11 ? n67735 : n67757;
  assign n67759 = pi20 ? n9641 : ~n141;
  assign n67760 = pi19 ? n32 : n67759;
  assign n67761 = pi18 ? n32 : n67760;
  assign n67762 = pi17 ? n32 : n67761;
  assign n67763 = pi16 ? n32 : n67762;
  assign n67764 = pi15 ? n67763 : n16832;
  assign n67765 = pi14 ? n17412 : n67764;
  assign n67766 = pi20 ? n7007 : n32;
  assign n67767 = pi19 ? n322 : n67766;
  assign n67768 = pi18 ? n32 : n67767;
  assign n67769 = pi17 ? n32 : n67768;
  assign n67770 = pi16 ? n32 : n67769;
  assign n67771 = pi15 ? n67770 : n24874;
  assign n67772 = pi19 ? n32 : n20610;
  assign n67773 = pi18 ? n32 : n67772;
  assign n67774 = pi17 ? n32 : n67773;
  assign n67775 = pi16 ? n32 : n67774;
  assign n67776 = pi15 ? n67775 : n40231;
  assign n67777 = pi14 ? n67771 : n67776;
  assign n67778 = pi13 ? n67765 : n67777;
  assign n67779 = pi17 ? n52276 : n16450;
  assign n67780 = pi16 ? n32 : n67779;
  assign n67781 = pi15 ? n40313 : n67780;
  assign n67782 = pi20 ? n260 : n1385;
  assign n67783 = pi19 ? n507 : n67782;
  assign n67784 = pi18 ? n67783 : ~n618;
  assign n67785 = pi17 ? n67784 : n27526;
  assign n67786 = pi16 ? n32 : n67785;
  assign n67787 = pi18 ? n508 : ~n16389;
  assign n67788 = pi19 ? n4670 : ~n6042;
  assign n67789 = pi18 ? n28421 : ~n67788;
  assign n67790 = pi17 ? n67787 : ~n67789;
  assign n67791 = pi16 ? n32 : n67790;
  assign n67792 = pi15 ? n67786 : n67791;
  assign n67793 = pi14 ? n67781 : n67792;
  assign n67794 = pi19 ? n4342 : ~n60048;
  assign n67795 = pi18 ? n32 : n67794;
  assign n67796 = pi17 ? n32 : n67795;
  assign n67797 = pi16 ? n32 : n67796;
  assign n67798 = pi15 ? n67797 : n50341;
  assign n67799 = pi21 ? n140 : n242;
  assign n67800 = pi20 ? n67799 : ~n32;
  assign n67801 = pi19 ? n507 : ~n67800;
  assign n67802 = pi18 ? n32 : n67801;
  assign n67803 = pi17 ? n32 : n67802;
  assign n67804 = pi16 ? n32 : n67803;
  assign n67805 = pi15 ? n16101 : n67804;
  assign n67806 = pi14 ? n67798 : n67805;
  assign n67807 = pi13 ? n67793 : n67806;
  assign n67808 = pi12 ? n67778 : n67807;
  assign n67809 = pi20 ? n38925 : n32;
  assign n67810 = pi19 ? n32 : n67809;
  assign n67811 = pi18 ? n32 : n67810;
  assign n67812 = pi17 ? n32 : n67811;
  assign n67813 = pi16 ? n32 : n67812;
  assign n67814 = pi15 ? n67813 : n52178;
  assign n67815 = pi14 ? n67814 : n67527;
  assign n67816 = pi18 ? n2747 : ~n350;
  assign n67817 = pi17 ? n67816 : n37195;
  assign n67818 = pi16 ? n32 : n67817;
  assign n67819 = pi15 ? n37644 : n67818;
  assign n67820 = pi19 ? n1320 : ~n267;
  assign n67821 = pi18 ? n67820 : ~n237;
  assign n67822 = pi17 ? n67821 : n53496;
  assign n67823 = pi16 ? n32 : n67822;
  assign n67824 = pi17 ? n43398 : n35032;
  assign n67825 = pi16 ? n32 : n67824;
  assign n67826 = pi15 ? n67823 : n67825;
  assign n67827 = pi14 ? n67819 : n67826;
  assign n67828 = pi13 ? n67815 : n67827;
  assign n67829 = pi17 ? n4682 : ~n67553;
  assign n67830 = pi16 ? n32 : n67829;
  assign n67831 = pi19 ? n750 : ~n5626;
  assign n67832 = pi18 ? n32 : n67831;
  assign n67833 = pi17 ? n4682 : ~n67832;
  assign n67834 = pi16 ? n32 : n67833;
  assign n67835 = pi15 ? n67830 : n67834;
  assign n67836 = pi18 ? n702 : ~n38521;
  assign n67837 = pi18 ? n22159 : ~n25244;
  assign n67838 = pi17 ? n67836 : ~n67837;
  assign n67839 = pi16 ? n32 : n67838;
  assign n67840 = pi15 ? n67839 : n14580;
  assign n67841 = pi14 ? n67835 : n67840;
  assign n67842 = pi17 ? n58767 : ~n2750;
  assign n67843 = pi16 ? n32 : n67842;
  assign n67844 = pi20 ? n564 : ~n831;
  assign n67845 = pi19 ? n32 : n67844;
  assign n67846 = pi18 ? n67845 : n38541;
  assign n67847 = pi19 ? n38545 : ~n1105;
  assign n67848 = pi18 ? n38544 : n67847;
  assign n67849 = pi17 ? n67846 : n67848;
  assign n67850 = pi16 ? n32 : n67849;
  assign n67851 = pi15 ? n67843 : n67850;
  assign n67852 = pi18 ? n24271 : n32;
  assign n67853 = pi17 ? n67852 : n34844;
  assign n67854 = pi16 ? n32 : n67853;
  assign n67855 = pi18 ? n268 : n350;
  assign n67856 = pi18 ? n4671 : n65572;
  assign n67857 = pi17 ? n67855 : ~n67856;
  assign n67858 = pi16 ? n32 : n67857;
  assign n67859 = pi15 ? n67854 : n67858;
  assign n67860 = pi14 ? n67851 : n67859;
  assign n67861 = pi13 ? n67841 : n67860;
  assign n67862 = pi12 ? n67828 : n67861;
  assign n67863 = pi11 ? n67808 : n67862;
  assign n67864 = pi10 ? n67758 : n67863;
  assign n67865 = pi09 ? n67729 : n67864;
  assign n67866 = pi13 ? n67730 : n52406;
  assign n67867 = pi19 ? n32 : n26857;
  assign n67868 = pi18 ? n32 : n67867;
  assign n67869 = pi17 ? n32 : n67868;
  assign n67870 = pi16 ? n32 : n67869;
  assign n67871 = pi15 ? n25904 : n67870;
  assign n67872 = pi14 ? n67871 : n38489;
  assign n67873 = pi14 ? n26100 : n32;
  assign n67874 = pi13 ? n67872 : n67873;
  assign n67875 = pi12 ? n67866 : n67874;
  assign n67876 = pi19 ? n32 : n21817;
  assign n67877 = pi18 ? n32 : n67876;
  assign n67878 = pi17 ? n32 : n67877;
  assign n67879 = pi16 ? n32 : n67878;
  assign n67880 = pi15 ? n16824 : n67879;
  assign n67881 = pi14 ? n16824 : n67880;
  assign n67882 = pi13 ? n67742 : n67881;
  assign n67883 = pi19 ? n507 : ~n1969;
  assign n67884 = pi18 ? n32 : n67883;
  assign n67885 = pi17 ? n32 : n67884;
  assign n67886 = pi16 ? n32 : n67885;
  assign n67887 = pi15 ? n67886 : n67610;
  assign n67888 = pi14 ? n67746 : n67887;
  assign n67889 = pi15 ? n27528 : n50513;
  assign n67890 = pi15 ? n32 : n25814;
  assign n67891 = pi14 ? n67889 : n67890;
  assign n67892 = pi13 ? n67888 : n67891;
  assign n67893 = pi12 ? n67882 : n67892;
  assign n67894 = pi11 ? n67875 : n67893;
  assign n67895 = pi20 ? n10183 : ~n243;
  assign n67896 = pi19 ? n32 : n67895;
  assign n67897 = pi18 ? n32 : n67896;
  assign n67898 = pi17 ? n32 : n67897;
  assign n67899 = pi16 ? n32 : n67898;
  assign n67900 = pi15 ? n67899 : n25814;
  assign n67901 = pi14 ? n17178 : n67900;
  assign n67902 = pi21 ? n32 : ~n20130;
  assign n67903 = pi20 ? n67902 : ~n32;
  assign n67904 = pi19 ? n32 : ~n67903;
  assign n67905 = pi18 ? n32 : n67904;
  assign n67906 = pi17 ? n32 : n67905;
  assign n67907 = pi16 ? n32 : n67906;
  assign n67908 = pi15 ? n67775 : n67907;
  assign n67909 = pi14 ? n67771 : n67908;
  assign n67910 = pi13 ? n67901 : n67909;
  assign n67911 = pi21 ? n32 : n16091;
  assign n67912 = pi20 ? n67911 : ~n32;
  assign n67913 = pi19 ? n32 : ~n67912;
  assign n67914 = pi18 ? n32 : n67913;
  assign n67915 = pi17 ? n32 : n67914;
  assign n67916 = pi16 ? n32 : n67915;
  assign n67917 = pi15 ? n67916 : n24237;
  assign n67918 = pi20 ? n831 : n321;
  assign n67919 = pi19 ? n32 : n67918;
  assign n67920 = pi18 ? n67919 : ~n618;
  assign n67921 = pi18 ? n19232 : n27525;
  assign n67922 = pi17 ? n67920 : n67921;
  assign n67923 = pi16 ? n32 : n67922;
  assign n67924 = pi18 ? n1750 : ~n16389;
  assign n67925 = pi17 ? n67924 : ~n67789;
  assign n67926 = pi16 ? n32 : n67925;
  assign n67927 = pi15 ? n67923 : n67926;
  assign n67928 = pi14 ? n67917 : n67927;
  assign n67929 = pi13 ? n67928 : n67806;
  assign n67930 = pi12 ? n67910 : n67929;
  assign n67931 = pi18 ? n2622 : ~n350;
  assign n67932 = pi17 ? n67931 : n37195;
  assign n67933 = pi16 ? n32 : n67932;
  assign n67934 = pi15 ? n67532 : n67933;
  assign n67935 = pi20 ? n141 : ~n266;
  assign n67936 = pi19 ? n32 : n67935;
  assign n67937 = pi18 ? n67936 : ~n237;
  assign n67938 = pi17 ? n67937 : n53496;
  assign n67939 = pi16 ? n32 : n67938;
  assign n67940 = pi17 ? n43398 : n67546;
  assign n67941 = pi16 ? n32 : n67940;
  assign n67942 = pi15 ? n67939 : n67941;
  assign n67943 = pi14 ? n67934 : n67942;
  assign n67944 = pi13 ? n67815 : n67943;
  assign n67945 = pi17 ? n4822 : ~n67553;
  assign n67946 = pi16 ? n32 : n67945;
  assign n67947 = pi17 ? n4822 : ~n67832;
  assign n67948 = pi16 ? n32 : n67947;
  assign n67949 = pi15 ? n67946 : n67948;
  assign n67950 = pi18 ? n38575 : ~n25244;
  assign n67951 = pi17 ? n38573 : ~n67950;
  assign n67952 = pi16 ? n32 : n67951;
  assign n67953 = pi15 ? n67952 : n14580;
  assign n67954 = pi14 ? n67949 : n67953;
  assign n67955 = pi20 ? n175 : n260;
  assign n67956 = pi19 ? n32 : n67955;
  assign n67957 = pi18 ? n67956 : ~n19654;
  assign n67958 = pi19 ? n6057 : n1105;
  assign n67959 = pi18 ? n32 : n67958;
  assign n67960 = pi17 ? n67957 : ~n67959;
  assign n67961 = pi16 ? n32 : n67960;
  assign n67962 = pi17 ? n17883 : n24999;
  assign n67963 = pi16 ? n32 : n67962;
  assign n67964 = pi15 ? n67961 : n67963;
  assign n67965 = pi15 ? n34846 : n67858;
  assign n67966 = pi14 ? n67964 : n67965;
  assign n67967 = pi13 ? n67954 : n67966;
  assign n67968 = pi12 ? n67944 : n67967;
  assign n67969 = pi11 ? n67930 : n67968;
  assign n67970 = pi10 ? n67894 : n67969;
  assign n67971 = pi09 ? n67729 : n67970;
  assign n67972 = pi08 ? n67865 : n67971;
  assign n67973 = pi07 ? n67723 : n67972;
  assign n67974 = pi06 ? n67431 : n67973;
  assign n67975 = pi05 ? n66867 : n67974;
  assign n67976 = pi04 ? n65731 : n67975;
  assign n67977 = pi03 ? n63759 : n67976;
  assign n67978 = pi02 ? n60306 : n67977;
  assign n67979 = pi01 ? n32 : n67978;
  assign n67980 = pi14 ? n32 : n26269;
  assign n67981 = pi13 ? n32 : n67980;
  assign n67982 = pi12 ? n32 : n67981;
  assign n67983 = pi11 ? n32 : n67982;
  assign n67984 = pi10 ? n32 : n67983;
  assign n67985 = pi14 ? n26904 : n26231;
  assign n67986 = pi15 ? n16850 : n26400;
  assign n67987 = pi14 ? n67986 : n26235;
  assign n67988 = pi13 ? n67985 : n67987;
  assign n67989 = pi15 ? n17348 : n26225;
  assign n67990 = pi14 ? n67989 : n38616;
  assign n67991 = pi13 ? n67990 : n32;
  assign n67992 = pi12 ? n67988 : n67991;
  assign n67993 = pi14 ? n26235 : n26145;
  assign n67994 = pi14 ? n67187 : n52055;
  assign n67995 = pi13 ? n67993 : n67994;
  assign n67996 = pi15 ? n16804 : n26201;
  assign n67997 = pi14 ? n26323 : n67996;
  assign n67998 = pi19 ? n32 : n29270;
  assign n67999 = pi18 ? n32 : n67998;
  assign n68000 = pi17 ? n32 : n67999;
  assign n68001 = pi16 ? n32 : n68000;
  assign n68002 = pi18 ? n32 : n19245;
  assign n68003 = pi17 ? n32 : n68002;
  assign n68004 = pi16 ? n32 : n68003;
  assign n68005 = pi15 ? n68001 : n68004;
  assign n68006 = pi15 ? n32 : n66880;
  assign n68007 = pi14 ? n68005 : n68006;
  assign n68008 = pi13 ? n67997 : n68007;
  assign n68009 = pi12 ? n67995 : n68008;
  assign n68010 = pi11 ? n67992 : n68009;
  assign n68011 = pi20 ? n382 : ~n339;
  assign n68012 = pi19 ? n32 : n68011;
  assign n68013 = pi18 ? n32 : n68012;
  assign n68014 = pi17 ? n32 : n68013;
  assign n68015 = pi16 ? n32 : n68014;
  assign n68016 = pi15 ? n17121 : n68015;
  assign n68017 = pi20 ? n7377 : n481;
  assign n68018 = pi19 ? n32 : n68017;
  assign n68019 = pi18 ? n32 : n68018;
  assign n68020 = pi17 ? n32 : n68019;
  assign n68021 = pi16 ? n32 : n68020;
  assign n68022 = pi20 ? n518 : n481;
  assign n68023 = pi19 ? n32 : n68022;
  assign n68024 = pi18 ? n32 : n68023;
  assign n68025 = pi17 ? n32 : n68024;
  assign n68026 = pi16 ? n32 : n68025;
  assign n68027 = pi15 ? n68021 : n68026;
  assign n68028 = pi14 ? n68016 : n68027;
  assign n68029 = pi20 ? n53136 : ~n339;
  assign n68030 = pi19 ? n1464 : n68029;
  assign n68031 = pi18 ? n32 : n68030;
  assign n68032 = pi17 ? n32 : n68031;
  assign n68033 = pi16 ? n32 : n68032;
  assign n68034 = pi20 ? n1817 : ~n339;
  assign n68035 = pi19 ? n322 : n68034;
  assign n68036 = pi18 ? n32 : n68035;
  assign n68037 = pi17 ? n32 : n68036;
  assign n68038 = pi16 ? n32 : n68037;
  assign n68039 = pi15 ? n68033 : n68038;
  assign n68040 = pi20 ? n1076 : n141;
  assign n68041 = pi19 ? n507 : ~n68040;
  assign n68042 = pi18 ? n32 : n68041;
  assign n68043 = pi17 ? n32 : n68042;
  assign n68044 = pi16 ? n32 : n68043;
  assign n68045 = pi20 ? n17712 : ~n32;
  assign n68046 = pi19 ? n32 : ~n68045;
  assign n68047 = pi18 ? n32 : n68046;
  assign n68048 = pi17 ? n32 : n68047;
  assign n68049 = pi16 ? n32 : n68048;
  assign n68050 = pi15 ? n68044 : n68049;
  assign n68051 = pi14 ? n68039 : n68050;
  assign n68052 = pi13 ? n68028 : n68051;
  assign n68053 = pi19 ? n507 : ~n53777;
  assign n68054 = pi18 ? n32 : n68053;
  assign n68055 = pi17 ? n32 : n68054;
  assign n68056 = pi16 ? n32 : n68055;
  assign n68057 = pi17 ? n52508 : n15228;
  assign n68058 = pi16 ? n32 : n68057;
  assign n68059 = pi15 ? n68056 : n68058;
  assign n68060 = pi18 ? n17650 : n20565;
  assign n68061 = pi17 ? n52518 : n68060;
  assign n68062 = pi16 ? n32 : n68061;
  assign n68063 = pi19 ? n5694 : n176;
  assign n68064 = pi18 ? n940 : ~n68063;
  assign n68065 = pi17 ? n34891 : ~n68064;
  assign n68066 = pi16 ? n32 : n68065;
  assign n68067 = pi15 ? n68062 : n68066;
  assign n68068 = pi14 ? n68059 : n68067;
  assign n68069 = pi19 ? n349 : n321;
  assign n68070 = pi19 ? n5694 : n112;
  assign n68071 = pi18 ? n68069 : ~n68070;
  assign n68072 = pi17 ? n15401 : ~n68071;
  assign n68073 = pi16 ? n32 : n68072;
  assign n68074 = pi15 ? n68073 : n50341;
  assign n68075 = pi15 ? n16452 : n67804;
  assign n68076 = pi14 ? n68074 : n68075;
  assign n68077 = pi13 ? n68068 : n68076;
  assign n68078 = pi12 ? n68052 : n68077;
  assign n68079 = pi20 ? n27922 : n32;
  assign n68080 = pi19 ? n32 : n68079;
  assign n68081 = pi18 ? n32 : n68080;
  assign n68082 = pi17 ? n32 : n68081;
  assign n68083 = pi16 ? n32 : n68082;
  assign n68084 = pi15 ? n68083 : n52178;
  assign n68085 = pi19 ? n1464 : ~n6683;
  assign n68086 = pi18 ? n32 : n68085;
  assign n68087 = pi17 ? n32 : n68086;
  assign n68088 = pi16 ? n32 : n68087;
  assign n68089 = pi15 ? n24582 : n68088;
  assign n68090 = pi14 ? n68084 : n68089;
  assign n68091 = pi18 ? n41652 : ~n23440;
  assign n68092 = pi19 ? n4982 : ~n20022;
  assign n68093 = pi18 ? n12811 : n68092;
  assign n68094 = pi17 ? n68091 : n68093;
  assign n68095 = pi16 ? n32 : n68094;
  assign n68096 = pi20 ? n38783 : ~n321;
  assign n68097 = pi19 ? n32 : n68096;
  assign n68098 = pi19 ? n20006 : n1464;
  assign n68099 = pi18 ? n68097 : ~n68098;
  assign n68100 = pi19 ? n4721 : n19892;
  assign n68101 = pi18 ? n45507 : n68100;
  assign n68102 = pi17 ? n68099 : n68101;
  assign n68103 = pi16 ? n32 : n68102;
  assign n68104 = pi15 ? n68095 : n68103;
  assign n68105 = pi19 ? n32302 : n349;
  assign n68106 = pi18 ? n68097 : ~n68105;
  assign n68107 = pi19 ? n208 : n5614;
  assign n68108 = pi18 ? n17642 : n68107;
  assign n68109 = pi17 ? n68106 : n68108;
  assign n68110 = pi16 ? n32 : n68109;
  assign n68111 = pi17 ? n17951 : n14573;
  assign n68112 = pi16 ? n32 : n68111;
  assign n68113 = pi15 ? n68110 : n68112;
  assign n68114 = pi14 ? n68104 : n68113;
  assign n68115 = pi13 ? n68090 : n68114;
  assign n68116 = pi17 ? n6439 : ~n67553;
  assign n68117 = pi16 ? n32 : n68116;
  assign n68118 = pi17 ? n6439 : ~n9961;
  assign n68119 = pi16 ? n32 : n68118;
  assign n68120 = pi15 ? n68117 : n68119;
  assign n68121 = pi18 ? n684 : n52537;
  assign n68122 = pi18 ? n52539 : n25244;
  assign n68123 = pi17 ? n68121 : n68122;
  assign n68124 = pi16 ? n32 : n68123;
  assign n68125 = pi15 ? n68124 : n22923;
  assign n68126 = pi14 ? n68120 : n68125;
  assign n68127 = pi18 ? n11930 : ~n38663;
  assign n68128 = pi19 ? n38778 : n1105;
  assign n68129 = pi18 ? n38665 : n68128;
  assign n68130 = pi17 ? n68127 : ~n68129;
  assign n68131 = pi16 ? n32 : n68130;
  assign n68132 = pi20 ? n67 : n1331;
  assign n68133 = pi19 ? n32 : n68132;
  assign n68134 = pi18 ? n68133 : n9170;
  assign n68135 = pi17 ? n68134 : n25670;
  assign n68136 = pi16 ? n32 : n68135;
  assign n68137 = pi15 ? n68131 : n68136;
  assign n68138 = pi18 ? n36848 : n15844;
  assign n68139 = pi21 ? n206 : ~n12274;
  assign n68140 = pi20 ? n32 : n68139;
  assign n68141 = pi19 ? n68140 : n32;
  assign n68142 = pi18 ? n52258 : n68141;
  assign n68143 = pi17 ? n68138 : n68142;
  assign n68144 = pi16 ? n32 : n68143;
  assign n68145 = pi18 ? n11930 : n52561;
  assign n68146 = pi18 ? n5731 : n65572;
  assign n68147 = pi17 ? n68145 : ~n68146;
  assign n68148 = pi16 ? n32 : n68147;
  assign n68149 = pi15 ? n68144 : n68148;
  assign n68150 = pi14 ? n68137 : n68149;
  assign n68151 = pi13 ? n68126 : n68150;
  assign n68152 = pi12 ? n68115 : n68151;
  assign n68153 = pi11 ? n68078 : n68152;
  assign n68154 = pi10 ? n68010 : n68153;
  assign n68155 = pi09 ? n67984 : n68154;
  assign n68156 = pi13 ? n67985 : n52572;
  assign n68157 = pi14 ? n38491 : n26269;
  assign n68158 = pi13 ? n68157 : n52574;
  assign n68159 = pi12 ? n68156 : n68158;
  assign n68160 = pi15 ? n16850 : n16397;
  assign n68161 = pi14 ? n67187 : n68160;
  assign n68162 = pi13 ? n67993 : n68161;
  assign n68163 = pi15 ? n16736 : n16824;
  assign n68164 = pi15 ? n16824 : n17056;
  assign n68165 = pi14 ? n68163 : n68164;
  assign n68166 = pi13 ? n68165 : n68007;
  assign n68167 = pi12 ? n68162 : n68166;
  assign n68168 = pi11 ? n68159 : n68167;
  assign n68169 = pi20 ? n1076 : ~n339;
  assign n68170 = pi19 ? n1464 : n68169;
  assign n68171 = pi18 ? n32 : n68170;
  assign n68172 = pi17 ? n32 : n68171;
  assign n68173 = pi16 ? n32 : n68172;
  assign n68174 = pi15 ? n68173 : n68038;
  assign n68175 = pi14 ? n68174 : n68050;
  assign n68176 = pi13 ? n68028 : n68175;
  assign n68177 = pi15 ? n68056 : n36100;
  assign n68178 = pi17 ? n52598 : n68060;
  assign n68179 = pi16 ? n32 : n68178;
  assign n68180 = pi17 ? n1966 : ~n68064;
  assign n68181 = pi16 ? n32 : n68180;
  assign n68182 = pi15 ? n68179 : n68181;
  assign n68183 = pi14 ? n68177 : n68182;
  assign n68184 = pi20 ? n46830 : ~n32;
  assign n68185 = pi19 ? n507 : ~n68184;
  assign n68186 = pi18 ? n32 : n68185;
  assign n68187 = pi17 ? n32 : n68186;
  assign n68188 = pi16 ? n32 : n68187;
  assign n68189 = pi15 ? n16452 : n68188;
  assign n68190 = pi14 ? n68074 : n68189;
  assign n68191 = pi13 ? n68183 : n68190;
  assign n68192 = pi12 ? n68176 : n68191;
  assign n68193 = pi19 ? n507 : ~n40268;
  assign n68194 = pi18 ? n32 : n68193;
  assign n68195 = pi17 ? n32 : n68194;
  assign n68196 = pi16 ? n32 : n68195;
  assign n68197 = pi15 ? n68083 : n68196;
  assign n68198 = pi14 ? n68197 : n68089;
  assign n68199 = pi18 ? n863 : ~n23440;
  assign n68200 = pi17 ? n68199 : n68093;
  assign n68201 = pi16 ? n32 : n68200;
  assign n68202 = pi18 ? n16666 : ~n68098;
  assign n68203 = pi19 ? n4721 : n7488;
  assign n68204 = pi18 ? n45507 : n68203;
  assign n68205 = pi17 ? n68202 : n68204;
  assign n68206 = pi16 ? n32 : n68205;
  assign n68207 = pi15 ? n68201 : n68206;
  assign n68208 = pi20 ? n2140 : ~n206;
  assign n68209 = pi19 ? n68208 : n349;
  assign n68210 = pi18 ? n16666 : ~n68209;
  assign n68211 = pi17 ? n68210 : n68108;
  assign n68212 = pi16 ? n32 : n68211;
  assign n68213 = pi15 ? n68212 : n68112;
  assign n68214 = pi14 ? n68207 : n68213;
  assign n68215 = pi13 ? n68198 : n68214;
  assign n68216 = pi17 ? n4798 : ~n67553;
  assign n68217 = pi16 ? n32 : n68216;
  assign n68218 = pi17 ? n4798 : ~n9961;
  assign n68219 = pi16 ? n32 : n68218;
  assign n68220 = pi15 ? n68217 : n68219;
  assign n68221 = pi18 ? n366 : n52537;
  assign n68222 = pi17 ? n68221 : n68122;
  assign n68223 = pi16 ? n32 : n68222;
  assign n68224 = pi15 ? n68223 : n1109;
  assign n68225 = pi14 ? n68220 : n68224;
  assign n68226 = pi18 ? n863 : ~n38714;
  assign n68227 = pi19 ? n750 : n1105;
  assign n68228 = pi18 ? n38665 : n68227;
  assign n68229 = pi17 ? n68226 : ~n68228;
  assign n68230 = pi16 ? n32 : n68229;
  assign n68231 = pi15 ? n68230 : n66700;
  assign n68232 = pi20 ? n32 : n20507;
  assign n68233 = pi19 ? n68232 : n32;
  assign n68234 = pi18 ? n52258 : n68233;
  assign n68235 = pi17 ? n15845 : n68234;
  assign n68236 = pi16 ? n32 : n68235;
  assign n68237 = pi18 ? n858 : n52622;
  assign n68238 = pi17 ? n68237 : ~n68146;
  assign n68239 = pi16 ? n32 : n68238;
  assign n68240 = pi15 ? n68236 : n68239;
  assign n68241 = pi14 ? n68231 : n68240;
  assign n68242 = pi13 ? n68225 : n68241;
  assign n68243 = pi12 ? n68215 : n68242;
  assign n68244 = pi11 ? n68192 : n68243;
  assign n68245 = pi10 ? n68168 : n68244;
  assign n68246 = pi09 ? n67984 : n68245;
  assign n68247 = pi08 ? n68155 : n68246;
  assign n68248 = pi15 ? n32 : n26354;
  assign n68249 = pi14 ? n32 : n68248;
  assign n68250 = pi13 ? n32 : n68249;
  assign n68251 = pi12 ? n32 : n68250;
  assign n68252 = pi11 ? n32 : n68251;
  assign n68253 = pi10 ? n32 : n68252;
  assign n68254 = pi15 ? n26269 : n17531;
  assign n68255 = pi15 ? n17348 : n26272;
  assign n68256 = pi14 ? n68254 : n68255;
  assign n68257 = pi13 ? n68256 : n52642;
  assign n68258 = pi14 ? n32 : n26904;
  assign n68259 = pi13 ? n52487 : n68258;
  assign n68260 = pi12 ? n68257 : n68259;
  assign n68261 = pi15 ? n26272 : n16850;
  assign n68262 = pi15 ? n17061 : n16850;
  assign n68263 = pi14 ? n68261 : n68262;
  assign n68264 = pi15 ? n16850 : n17061;
  assign n68265 = pi14 ? n68264 : n68262;
  assign n68266 = pi13 ? n68263 : n68265;
  assign n68267 = pi20 ? n428 : ~n501;
  assign n68268 = pi19 ? n32 : n68267;
  assign n68269 = pi18 ? n32 : n68268;
  assign n68270 = pi17 ? n32 : n68269;
  assign n68271 = pi16 ? n32 : n68270;
  assign n68272 = pi15 ? n68271 : n16824;
  assign n68273 = pi14 ? n68272 : n27341;
  assign n68274 = pi15 ? n16804 : n40426;
  assign n68275 = pi15 ? n25904 : n66880;
  assign n68276 = pi14 ? n68274 : n68275;
  assign n68277 = pi13 ? n68273 : n68276;
  assign n68278 = pi12 ? n68266 : n68277;
  assign n68279 = pi11 ? n68260 : n68278;
  assign n68280 = pi20 ? n8630 : ~n1940;
  assign n68281 = pi19 ? n32 : n68280;
  assign n68282 = pi18 ? n32 : n68281;
  assign n68283 = pi17 ? n32 : n68282;
  assign n68284 = pi16 ? n32 : n68283;
  assign n68285 = pi15 ? n25997 : n68284;
  assign n68286 = pi20 ? n7377 : ~n243;
  assign n68287 = pi19 ? n32 : n68286;
  assign n68288 = pi18 ? n32 : n68287;
  assign n68289 = pi17 ? n32585 : n68288;
  assign n68290 = pi16 ? n32 : n68289;
  assign n68291 = pi15 ? n68290 : n68026;
  assign n68292 = pi14 ? n68285 : n68291;
  assign n68293 = pi19 ? n32 : n68169;
  assign n68294 = pi18 ? n32 : n68293;
  assign n68295 = pi17 ? n32 : n68294;
  assign n68296 = pi16 ? n32 : n68295;
  assign n68297 = pi19 ? n507 : n68034;
  assign n68298 = pi18 ? n32 : n68297;
  assign n68299 = pi17 ? n32 : n68298;
  assign n68300 = pi16 ? n32 : n68299;
  assign n68301 = pi15 ? n68296 : n68300;
  assign n68302 = pi20 ? n1076 : n339;
  assign n68303 = pi19 ? n507 : ~n68302;
  assign n68304 = pi18 ? n32 : n68303;
  assign n68305 = pi17 ? n32 : n68304;
  assign n68306 = pi16 ? n32 : n68305;
  assign n68307 = pi15 ? n68306 : n27388;
  assign n68308 = pi14 ? n68301 : n68307;
  assign n68309 = pi13 ? n68292 : n68308;
  assign n68310 = pi19 ? n507 : ~n3524;
  assign n68311 = pi18 ? n32 : n68310;
  assign n68312 = pi17 ? n32 : n68311;
  assign n68313 = pi16 ? n32 : n68312;
  assign n68314 = pi15 ? n68056 : n68313;
  assign n68315 = pi17 ? n52666 : n24872;
  assign n68316 = pi16 ? n32 : n68315;
  assign n68317 = pi18 ? n4281 : ~n32;
  assign n68318 = pi17 ? n68317 : ~n68064;
  assign n68319 = pi16 ? n32 : n68318;
  assign n68320 = pi15 ? n68316 : n68319;
  assign n68321 = pi14 ? n68314 : n68320;
  assign n68322 = pi20 ? n246 : n333;
  assign n68323 = pi19 ? n68322 : n5707;
  assign n68324 = pi18 ? n32 : n68323;
  assign n68325 = pi19 ? n6298 : n321;
  assign n68326 = pi18 ? n68325 : ~n68070;
  assign n68327 = pi17 ? n68324 : ~n68326;
  assign n68328 = pi16 ? n32 : n68327;
  assign n68329 = pi15 ? n68328 : n50341;
  assign n68330 = pi19 ? n594 : n19317;
  assign n68331 = pi18 ? n32 : n68330;
  assign n68332 = pi17 ? n32 : n68331;
  assign n68333 = pi16 ? n32 : n68332;
  assign n68334 = pi15 ? n16452 : n68333;
  assign n68335 = pi14 ? n68329 : n68334;
  assign n68336 = pi13 ? n68321 : n68335;
  assign n68337 = pi12 ? n68309 : n68336;
  assign n68338 = pi19 ? n857 : ~n40268;
  assign n68339 = pi18 ? n32 : n68338;
  assign n68340 = pi17 ? n32 : n68339;
  assign n68341 = pi16 ? n32 : n68340;
  assign n68342 = pi15 ? n24705 : n68341;
  assign n68343 = pi19 ? n594 : n52364;
  assign n68344 = pi18 ? n32 : n68343;
  assign n68345 = pi17 ? n32 : n68344;
  assign n68346 = pi16 ? n32 : n68345;
  assign n68347 = pi19 ? n322 : ~n502;
  assign n68348 = pi18 ? n32 : n68347;
  assign n68349 = pi17 ? n32 : n68348;
  assign n68350 = pi16 ? n32 : n68349;
  assign n68351 = pi15 ? n68346 : n68350;
  assign n68352 = pi14 ? n68342 : n68351;
  assign n68353 = pi18 ? n1379 : ~n23440;
  assign n68354 = pi22 ? n50 : ~n84;
  assign n68355 = pi21 ? n68354 : ~n32;
  assign n68356 = pi20 ? n68355 : ~n32;
  assign n68357 = pi19 ? n17918 : ~n68356;
  assign n68358 = pi18 ? n12811 : n68357;
  assign n68359 = pi17 ? n68353 : n68358;
  assign n68360 = pi16 ? n32 : n68359;
  assign n68361 = pi21 ? n13784 : n259;
  assign n68362 = pi20 ? n32 : n68361;
  assign n68363 = pi19 ? n32 : n68362;
  assign n68364 = pi18 ? n68363 : ~n32;
  assign n68365 = pi19 ? n343 : ~n6298;
  assign n68366 = pi21 ? n12274 : ~n32;
  assign n68367 = pi20 ? n68366 : ~n32;
  assign n68368 = pi19 ? n5694 : ~n68367;
  assign n68369 = pi18 ? n68365 : n68368;
  assign n68370 = pi17 ? n68364 : n68369;
  assign n68371 = pi16 ? n32 : n68370;
  assign n68372 = pi15 ? n68360 : n68371;
  assign n68373 = pi18 ? n68363 : ~n496;
  assign n68374 = pi19 ? n18396 : n32;
  assign n68375 = pi18 ? n68374 : n14567;
  assign n68376 = pi17 ? n68373 : n68375;
  assign n68377 = pi16 ? n32 : n68376;
  assign n68378 = pi17 ? n17849 : n14573;
  assign n68379 = pi16 ? n32 : n68378;
  assign n68380 = pi15 ? n68377 : n68379;
  assign n68381 = pi14 ? n68372 : n68380;
  assign n68382 = pi13 ? n68352 : n68381;
  assign n68383 = pi19 ? n1325 : ~n7502;
  assign n68384 = pi18 ? n32 : n68383;
  assign n68385 = pi17 ? n1971 : ~n68384;
  assign n68386 = pi16 ? n32 : n68385;
  assign n68387 = pi17 ? n1971 : ~n65547;
  assign n68388 = pi16 ? n32 : n68387;
  assign n68389 = pi15 ? n68386 : n68388;
  assign n68390 = pi18 ? n1819 : n52697;
  assign n68391 = pi18 ? n4965 : n27463;
  assign n68392 = pi17 ? n68390 : n68391;
  assign n68393 = pi16 ? n32 : n68392;
  assign n68394 = pi19 ? n5748 : ~n1105;
  assign n68395 = pi18 ? n38787 : n68394;
  assign n68396 = pi17 ? n17820 : n68395;
  assign n68397 = pi16 ? n32 : n68396;
  assign n68398 = pi15 ? n68393 : n68397;
  assign n68399 = pi14 ? n68389 : n68398;
  assign n68400 = pi18 ? n17819 : n28160;
  assign n68401 = pi19 ? n28686 : n39206;
  assign n68402 = pi19 ? n208 : n1105;
  assign n68403 = pi18 ? n68401 : ~n68402;
  assign n68404 = pi17 ? n68400 : n68403;
  assign n68405 = pi16 ? n32 : n68404;
  assign n68406 = pi17 ? n18292 : n27469;
  assign n68407 = pi16 ? n32 : n68406;
  assign n68408 = pi15 ? n68405 : n68407;
  assign n68409 = pi18 ? n28273 : n15844;
  assign n68410 = pi17 ? n68409 : n68234;
  assign n68411 = pi16 ? n32 : n68410;
  assign n68412 = pi18 ? n17819 : n52561;
  assign n68413 = pi18 ? n14153 : n65572;
  assign n68414 = pi17 ? n68412 : ~n68413;
  assign n68415 = pi16 ? n32 : n68414;
  assign n68416 = pi15 ? n68411 : n68415;
  assign n68417 = pi14 ? n68408 : n68416;
  assign n68418 = pi13 ? n68399 : n68417;
  assign n68419 = pi12 ? n68382 : n68418;
  assign n68420 = pi11 ? n68337 : n68419;
  assign n68421 = pi10 ? n68279 : n68420;
  assign n68422 = pi09 ? n68253 : n68421;
  assign n68423 = pi15 ? n26272 : n17152;
  assign n68424 = pi14 ? n68254 : n68423;
  assign n68425 = pi13 ? n68424 : n52739;
  assign n68426 = pi15 ? n17348 : n17531;
  assign n68427 = pi14 ? n68426 : n32;
  assign n68428 = pi13 ? n68427 : n68258;
  assign n68429 = pi12 ? n68425 : n68428;
  assign n68430 = pi15 ? n26183 : n16850;
  assign n68431 = pi14 ? n68430 : n68262;
  assign n68432 = pi13 ? n68431 : n68265;
  assign n68433 = pi14 ? n68274 : n68006;
  assign n68434 = pi13 ? n68273 : n68433;
  assign n68435 = pi12 ? n68432 : n68434;
  assign n68436 = pi11 ? n68429 : n68435;
  assign n68437 = pi20 ? n8630 : ~n339;
  assign n68438 = pi19 ? n32 : n68437;
  assign n68439 = pi18 ? n32 : n68438;
  assign n68440 = pi17 ? n32 : n68439;
  assign n68441 = pi16 ? n32 : n68440;
  assign n68442 = pi15 ? n26201 : n68441;
  assign n68443 = pi14 ? n68442 : n68291;
  assign n68444 = pi15 ? n68044 : n27388;
  assign n68445 = pi14 ? n68301 : n68444;
  assign n68446 = pi13 ? n68443 : n68445;
  assign n68447 = pi17 ? n17849 : n37996;
  assign n68448 = pi16 ? n32 : n68447;
  assign n68449 = pi15 ? n68056 : n68448;
  assign n68450 = pi17 ? n52749 : n24872;
  assign n68451 = pi16 ? n32 : n68450;
  assign n68452 = pi17 ? n1580 : ~n68064;
  assign n68453 = pi16 ? n32 : n68452;
  assign n68454 = pi15 ? n68451 : n68453;
  assign n68455 = pi14 ? n68449 : n68454;
  assign n68456 = pi18 ? n17848 : n68323;
  assign n68457 = pi17 ? n68456 : ~n68326;
  assign n68458 = pi16 ? n32 : n68457;
  assign n68459 = pi15 ? n68458 : n50341;
  assign n68460 = pi19 ? n1574 : n19317;
  assign n68461 = pi18 ? n32 : n68460;
  assign n68462 = pi17 ? n32 : n68461;
  assign n68463 = pi16 ? n32 : n68462;
  assign n68464 = pi15 ? n16452 : n68463;
  assign n68465 = pi14 ? n68459 : n68464;
  assign n68466 = pi13 ? n68455 : n68465;
  assign n68467 = pi12 ? n68446 : n68466;
  assign n68468 = pi19 ? n857 : n67517;
  assign n68469 = pi18 ? n32 : n68468;
  assign n68470 = pi17 ? n32 : n68469;
  assign n68471 = pi16 ? n32 : n68470;
  assign n68472 = pi15 ? n24705 : n68471;
  assign n68473 = pi19 ? n594 : ~n6683;
  assign n68474 = pi18 ? n32 : n68473;
  assign n68475 = pi17 ? n32 : n68474;
  assign n68476 = pi16 ? n32 : n68475;
  assign n68477 = pi19 ? n322 : ~n20022;
  assign n68478 = pi18 ? n32 : n68477;
  assign n68479 = pi17 ? n32 : n68478;
  assign n68480 = pi16 ? n32 : n68479;
  assign n68481 = pi15 ? n68476 : n68480;
  assign n68482 = pi14 ? n68472 : n68481;
  assign n68483 = pi18 ? n1841 : ~n23440;
  assign n68484 = pi19 ? n17918 : n6230;
  assign n68485 = pi18 ? n12811 : n68484;
  assign n68486 = pi17 ? n68483 : n68485;
  assign n68487 = pi16 ? n32 : n68486;
  assign n68488 = pi19 ? n5694 : n5614;
  assign n68489 = pi18 ? n68365 : n68488;
  assign n68490 = pi17 ? n1842 : n68489;
  assign n68491 = pi16 ? n32 : n68490;
  assign n68492 = pi15 ? n68487 : n68491;
  assign n68493 = pi17 ? n12700 : n68375;
  assign n68494 = pi16 ? n32 : n68493;
  assign n68495 = pi15 ? n68494 : n68379;
  assign n68496 = pi14 ? n68492 : n68495;
  assign n68497 = pi13 ? n68482 : n68496;
  assign n68498 = pi19 ? n1325 : ~n5626;
  assign n68499 = pi18 ? n32 : n68498;
  assign n68500 = pi17 ? n1322 : ~n68499;
  assign n68501 = pi16 ? n32 : n68500;
  assign n68502 = pi17 ? n1322 : ~n65547;
  assign n68503 = pi16 ? n32 : n68502;
  assign n68504 = pi15 ? n68501 : n68503;
  assign n68505 = pi18 ? n32 : n52697;
  assign n68506 = pi17 ? n68505 : n68391;
  assign n68507 = pi16 ? n32 : n68506;
  assign n68508 = pi17 ? n32 : n68395;
  assign n68509 = pi16 ? n32 : n68508;
  assign n68510 = pi15 ? n68507 : n68509;
  assign n68511 = pi14 ? n68504 : n68510;
  assign n68512 = pi18 ? n32 : n28160;
  assign n68513 = pi17 ? n68512 : n68403;
  assign n68514 = pi16 ? n32 : n68513;
  assign n68515 = pi15 ? n68514 : n22825;
  assign n68516 = pi18 ? n1575 : n15844;
  assign n68517 = pi17 ? n68516 : n68234;
  assign n68518 = pi16 ? n32 : n68517;
  assign n68519 = pi18 ? n32 : n52561;
  assign n68520 = pi18 ? n14153 : n35545;
  assign n68521 = pi17 ? n68519 : ~n68520;
  assign n68522 = pi16 ? n32 : n68521;
  assign n68523 = pi15 ? n68518 : n68522;
  assign n68524 = pi14 ? n68515 : n68523;
  assign n68525 = pi13 ? n68511 : n68524;
  assign n68526 = pi12 ? n68497 : n68525;
  assign n68527 = pi11 ? n68467 : n68526;
  assign n68528 = pi10 ? n68436 : n68527;
  assign n68529 = pi09 ? n68253 : n68528;
  assign n68530 = pi08 ? n68422 : n68529;
  assign n68531 = pi07 ? n68247 : n68530;
  assign n68532 = pi14 ? n32 : n26462;
  assign n68533 = pi13 ? n32 : n68532;
  assign n68534 = pi12 ? n32 : n68533;
  assign n68535 = pi11 ? n32 : n68534;
  assign n68536 = pi10 ? n32 : n68535;
  assign n68537 = pi15 ? n32 : n26462;
  assign n68538 = pi14 ? n68537 : n17421;
  assign n68539 = pi14 ? n26434 : n52805;
  assign n68540 = pi13 ? n68538 : n68539;
  assign n68541 = pi15 ? n38855 : n17531;
  assign n68542 = pi14 ? n68541 : n26904;
  assign n68543 = pi13 ? n68542 : n32;
  assign n68544 = pi12 ? n68540 : n68543;
  assign n68545 = pi20 ? n321 : n17509;
  assign n68546 = pi19 ? n32 : n68545;
  assign n68547 = pi18 ? n32 : n68546;
  assign n68548 = pi17 ? n32 : n68547;
  assign n68549 = pi16 ? n32 : n68548;
  assign n68550 = pi18 ? n32 : n56417;
  assign n68551 = pi17 ? n32 : n68550;
  assign n68552 = pi16 ? n32 : n68551;
  assign n68553 = pi15 ? n68549 : n68552;
  assign n68554 = pi15 ? n53119 : n17205;
  assign n68555 = pi14 ? n68553 : n68554;
  assign n68556 = pi15 ? n17205 : n53119;
  assign n68557 = pi15 ? n53119 : n26400;
  assign n68558 = pi14 ? n68556 : n68557;
  assign n68559 = pi13 ? n68555 : n68558;
  assign n68560 = pi20 ? n428 : ~n1839;
  assign n68561 = pi19 ? n32 : n68560;
  assign n68562 = pi18 ? n32 : n68561;
  assign n68563 = pi17 ? n32 : n68562;
  assign n68564 = pi16 ? n32 : n68563;
  assign n68565 = pi15 ? n26400 : n68564;
  assign n68566 = pi15 ? n26322 : n25984;
  assign n68567 = pi14 ? n68565 : n68566;
  assign n68568 = pi15 ? n16804 : n26479;
  assign n68569 = pi15 ? n52818 : n16452;
  assign n68570 = pi14 ? n68568 : n68569;
  assign n68571 = pi13 ? n68567 : n68570;
  assign n68572 = pi12 ? n68559 : n68571;
  assign n68573 = pi11 ? n68544 : n68572;
  assign n68574 = pi20 ? n7007 : n481;
  assign n68575 = pi19 ? n32 : n68574;
  assign n68576 = pi18 ? n32 : n68575;
  assign n68577 = pi17 ? n32 : n68576;
  assign n68578 = pi16 ? n32 : n68577;
  assign n68579 = pi15 ? n40478 : n68578;
  assign n68580 = pi14 ? n68285 : n68579;
  assign n68581 = pi21 ? n206 : n124;
  assign n68582 = pi20 ? n68581 : ~n339;
  assign n68583 = pi19 ? n32 : n68582;
  assign n68584 = pi18 ? n32 : n68583;
  assign n68585 = pi17 ? n32 : n68584;
  assign n68586 = pi16 ? n32 : n68585;
  assign n68587 = pi15 ? n25708 : n68586;
  assign n68588 = pi20 ? n16521 : ~n339;
  assign n68589 = pi19 ? n32 : n68588;
  assign n68590 = pi18 ? n32 : n68589;
  assign n68591 = pi17 ? n32 : n68590;
  assign n68592 = pi16 ? n32 : n68591;
  assign n68593 = pi15 ? n68592 : n16467;
  assign n68594 = pi14 ? n68587 : n68593;
  assign n68595 = pi13 ? n68580 : n68594;
  assign n68596 = pi19 ? n9037 : n4342;
  assign n68597 = pi18 ? n32 : n68596;
  assign n68598 = pi21 ? n174 : n35;
  assign n68599 = pi20 ? n68598 : ~n32;
  assign n68600 = pi19 ? n32 : ~n68599;
  assign n68601 = pi18 ? n16847 : n68600;
  assign n68602 = pi17 ? n68597 : n68601;
  assign n68603 = pi16 ? n32 : n68602;
  assign n68604 = pi17 ? n52850 : n14983;
  assign n68605 = pi16 ? n32 : n68604;
  assign n68606 = pi15 ? n68603 : n68605;
  assign n68607 = pi14 ? n68606 : n25572;
  assign n68608 = pi19 ? n507 : n25448;
  assign n68609 = pi18 ? n32 : n68608;
  assign n68610 = pi17 ? n32 : n68609;
  assign n68611 = pi16 ? n32 : n68610;
  assign n68612 = pi15 ? n37182 : n68611;
  assign n68613 = pi19 ? n1574 : ~n2317;
  assign n68614 = pi18 ? n32 : n68613;
  assign n68615 = pi17 ? n32 : n68614;
  assign n68616 = pi16 ? n32 : n68615;
  assign n68617 = pi15 ? n55295 : n68616;
  assign n68618 = pi14 ? n68612 : n68617;
  assign n68619 = pi13 ? n68607 : n68618;
  assign n68620 = pi12 ? n68595 : n68619;
  assign n68621 = pi17 ? n32 : n66683;
  assign n68622 = pi16 ? n32 : n68621;
  assign n68623 = pi15 ? n24640 : n68622;
  assign n68624 = pi19 ? n267 : n6049;
  assign n68625 = pi18 ? n32 : n68624;
  assign n68626 = pi20 ? n501 : n321;
  assign n68627 = pi20 ? n10889 : ~n206;
  assign n68628 = pi19 ? n68626 : n68627;
  assign n68629 = pi19 ? n349 : n7480;
  assign n68630 = pi18 ? n68628 : ~n68629;
  assign n68631 = pi17 ? n68625 : n68630;
  assign n68632 = pi16 ? n32 : n68631;
  assign n68633 = pi15 ? n16105 : n68632;
  assign n68634 = pi14 ? n68623 : n68633;
  assign n68635 = pi18 ? n322 : ~n63394;
  assign n68636 = pi17 ? n32149 : ~n68635;
  assign n68637 = pi16 ? n32 : n68636;
  assign n68638 = pi18 ? n1575 : n532;
  assign n68639 = pi19 ? n4982 : ~n813;
  assign n68640 = pi18 ? n322 : ~n68639;
  assign n68641 = pi17 ? n68638 : ~n68640;
  assign n68642 = pi16 ? n32 : n68641;
  assign n68643 = pi15 ? n68637 : n68642;
  assign n68644 = pi18 ? n32 : ~n32317;
  assign n68645 = pi18 ? n940 : n37658;
  assign n68646 = pi17 ? n68644 : n68645;
  assign n68647 = pi16 ? n32 : n68646;
  assign n68648 = pi19 ? n507 : n18665;
  assign n68649 = pi18 ? n32 : n68648;
  assign n68650 = pi19 ? n4721 : n7502;
  assign n68651 = pi18 ? n32 : n68650;
  assign n68652 = pi17 ? n68649 : n68651;
  assign n68653 = pi16 ? n32 : n68652;
  assign n68654 = pi15 ? n68647 : n68653;
  assign n68655 = pi14 ? n68643 : n68654;
  assign n68656 = pi13 ? n68634 : n68655;
  assign n68657 = pi19 ? n4721 : n2614;
  assign n68658 = pi18 ? n32 : n68657;
  assign n68659 = pi17 ? n1677 : ~n68658;
  assign n68660 = pi16 ? n32 : n68659;
  assign n68661 = pi20 ? n1611 : ~n321;
  assign n68662 = pi19 ? n68661 : n322;
  assign n68663 = pi18 ? n32 : n68662;
  assign n68664 = pi18 ? n46739 : ~n15515;
  assign n68665 = pi17 ? n68663 : ~n68664;
  assign n68666 = pi16 ? n32 : n68665;
  assign n68667 = pi15 ? n68660 : n68666;
  assign n68668 = pi19 ? n1844 : n507;
  assign n68669 = pi18 ? n32 : n68668;
  assign n68670 = pi19 ? n5356 : n1105;
  assign n68671 = pi18 ? n4380 : ~n68670;
  assign n68672 = pi17 ? n68669 : n68671;
  assign n68673 = pi16 ? n32 : n68672;
  assign n68674 = pi20 ? n16079 : ~n207;
  assign n68675 = pi19 ? n68674 : n32;
  assign n68676 = pi18 ? n32 : n68675;
  assign n68677 = pi19 ? n5694 : n1105;
  assign n68678 = pi18 ? n20164 : ~n68677;
  assign n68679 = pi17 ? n68676 : n68678;
  assign n68680 = pi16 ? n32 : n68679;
  assign n68681 = pi15 ? n68673 : n68680;
  assign n68682 = pi14 ? n68667 : n68681;
  assign n68683 = pi19 ? n9822 : n32;
  assign n68684 = pi18 ? n32 : n68683;
  assign n68685 = pi17 ? n57774 : n68684;
  assign n68686 = pi16 ? n32 : n68685;
  assign n68687 = pi17 ? n16317 : n33968;
  assign n68688 = pi16 ? n32 : n68687;
  assign n68689 = pi15 ? n68686 : n68688;
  assign n68690 = pi19 ? n51391 : ~n236;
  assign n68691 = pi18 ? n32 : n68690;
  assign n68692 = pi18 ? n32 : n6140;
  assign n68693 = pi17 ? n68691 : n68692;
  assign n68694 = pi16 ? n32 : n68693;
  assign n68695 = pi19 ? n15685 : ~n5694;
  assign n68696 = pi18 ? n32 : n68695;
  assign n68697 = pi17 ? n68696 : ~n7535;
  assign n68698 = pi16 ? n32 : n68697;
  assign n68699 = pi15 ? n68694 : n68698;
  assign n68700 = pi14 ? n68689 : n68699;
  assign n68701 = pi13 ? n68682 : n68700;
  assign n68702 = pi12 ? n68656 : n68701;
  assign n68703 = pi11 ? n68620 : n68702;
  assign n68704 = pi10 ? n68573 : n68703;
  assign n68705 = pi09 ? n68536 : n68704;
  assign n68706 = pi14 ? n68537 : n17619;
  assign n68707 = pi13 ? n68706 : n52901;
  assign n68708 = pi18 ? n32 : n56696;
  assign n68709 = pi17 ? n32 : n68708;
  assign n68710 = pi16 ? n32 : n68709;
  assign n68711 = pi15 ? n68710 : n32;
  assign n68712 = pi14 ? n68711 : n26904;
  assign n68713 = pi13 ? n68712 : n38814;
  assign n68714 = pi12 ? n68707 : n68713;
  assign n68715 = pi15 ? n53119 : n17152;
  assign n68716 = pi14 ? n68553 : n68715;
  assign n68717 = pi15 ? n17152 : n53119;
  assign n68718 = pi15 ? n53119 : n16850;
  assign n68719 = pi14 ? n68717 : n68718;
  assign n68720 = pi13 ? n68716 : n68719;
  assign n68721 = pi19 ? n32 : n24209;
  assign n68722 = pi18 ? n32 : n68721;
  assign n68723 = pi17 ? n32 : n68722;
  assign n68724 = pi16 ? n32 : n68723;
  assign n68725 = pi15 ? n16850 : n68724;
  assign n68726 = pi14 ? n68725 : n68566;
  assign n68727 = pi13 ? n68726 : n68570;
  assign n68728 = pi12 ? n68720 : n68727;
  assign n68729 = pi11 ? n68714 : n68728;
  assign n68730 = pi20 ? n1076 : ~n1940;
  assign n68731 = pi19 ? n32 : n68730;
  assign n68732 = pi18 ? n32 : n68731;
  assign n68733 = pi17 ? n32 : n68732;
  assign n68734 = pi16 ? n32 : n68733;
  assign n68735 = pi15 ? n26201 : n68734;
  assign n68736 = pi20 ? n14286 : ~n243;
  assign n68737 = pi19 ? n32 : n68736;
  assign n68738 = pi18 ? n32 : n68737;
  assign n68739 = pi17 ? n32 : n68738;
  assign n68740 = pi16 ? n32 : n68739;
  assign n68741 = pi15 ? n68740 : n68026;
  assign n68742 = pi14 ? n68735 : n68741;
  assign n68743 = pi20 ? n16521 : ~n141;
  assign n68744 = pi19 ? n32 : n68743;
  assign n68745 = pi18 ? n32 : n68744;
  assign n68746 = pi17 ? n32 : n68745;
  assign n68747 = pi16 ? n32 : n68746;
  assign n68748 = pi15 ? n68747 : n16467;
  assign n68749 = pi14 ? n68587 : n68748;
  assign n68750 = pi13 ? n68742 : n68749;
  assign n68751 = pi17 ? n52924 : n27526;
  assign n68752 = pi16 ? n32 : n68751;
  assign n68753 = pi15 ? n68603 : n68752;
  assign n68754 = pi17 ? n20280 : n24872;
  assign n68755 = pi16 ? n32 : n68754;
  assign n68756 = pi15 ? n68755 : n32;
  assign n68757 = pi14 ? n68753 : n68756;
  assign n68758 = pi19 ? n507 : n16294;
  assign n68759 = pi18 ? n32 : n68758;
  assign n68760 = pi17 ? n32 : n68759;
  assign n68761 = pi16 ? n32 : n68760;
  assign n68762 = pi15 ? n37182 : n68761;
  assign n68763 = pi15 ? n55295 : n24640;
  assign n68764 = pi14 ? n68762 : n68763;
  assign n68765 = pi13 ? n68757 : n68764;
  assign n68766 = pi12 ? n68750 : n68765;
  assign n68767 = pi15 ? n24247 : n68622;
  assign n68768 = pi20 ? n39175 : ~n2358;
  assign n68769 = pi20 ? n6050 : ~n2385;
  assign n68770 = pi19 ? n68768 : ~n68769;
  assign n68771 = pi18 ? n32 : n68770;
  assign n68772 = pi19 ? n349 : ~n7488;
  assign n68773 = pi18 ? n68628 : ~n68772;
  assign n68774 = pi17 ? n68771 : n68773;
  assign n68775 = pi16 ? n32 : n68774;
  assign n68776 = pi15 ? n16105 : n68775;
  assign n68777 = pi14 ? n68767 : n68776;
  assign n68778 = pi17 ? n2531 : ~n68640;
  assign n68779 = pi16 ? n32 : n68778;
  assign n68780 = pi15 ? n68637 : n68779;
  assign n68781 = pi17 ? n14154 : n68645;
  assign n68782 = pi16 ? n32 : n68781;
  assign n68783 = pi19 ? n28926 : ~n10410;
  assign n68784 = pi18 ? n32 : n68783;
  assign n68785 = pi17 ? n68784 : n38173;
  assign n68786 = pi16 ? n32 : n68785;
  assign n68787 = pi15 ? n68782 : n68786;
  assign n68788 = pi14 ? n68780 : n68787;
  assign n68789 = pi13 ? n68777 : n68788;
  assign n68790 = pi17 ? n2136 : ~n68658;
  assign n68791 = pi16 ? n32 : n68790;
  assign n68792 = pi20 ? n9628 : ~n321;
  assign n68793 = pi19 ? n68792 : n322;
  assign n68794 = pi18 ? n32 : n68793;
  assign n68795 = pi17 ? n68794 : ~n68664;
  assign n68796 = pi16 ? n32 : n68795;
  assign n68797 = pi15 ? n68791 : n68796;
  assign n68798 = pi17 ? n2954 : n68671;
  assign n68799 = pi16 ? n32 : n68798;
  assign n68800 = pi17 ? n21344 : n68678;
  assign n68801 = pi16 ? n32 : n68800;
  assign n68802 = pi15 ? n68799 : n68801;
  assign n68803 = pi14 ? n68797 : n68802;
  assign n68804 = pi17 ? n32 : n68684;
  assign n68805 = pi16 ? n32 : n68804;
  assign n68806 = pi17 ? n52948 : n33968;
  assign n68807 = pi16 ? n32 : n68806;
  assign n68808 = pi15 ? n68805 : n68807;
  assign n68809 = pi19 ? n28926 : ~n236;
  assign n68810 = pi18 ? n32 : n68809;
  assign n68811 = pi17 ? n68810 : n68692;
  assign n68812 = pi16 ? n32 : n68811;
  assign n68813 = pi19 ? n15983 : ~n5694;
  assign n68814 = pi18 ? n32 : n68813;
  assign n68815 = pi17 ? n68814 : ~n7535;
  assign n68816 = pi16 ? n32 : n68815;
  assign n68817 = pi15 ? n68812 : n68816;
  assign n68818 = pi14 ? n68808 : n68817;
  assign n68819 = pi13 ? n68803 : n68818;
  assign n68820 = pi12 ? n68789 : n68819;
  assign n68821 = pi11 ? n68766 : n68820;
  assign n68822 = pi10 ? n68729 : n68821;
  assign n68823 = pi09 ? n68536 : n68822;
  assign n68824 = pi08 ? n68705 : n68823;
  assign n68825 = pi14 ? n38967 : n38973;
  assign n68826 = pi13 ? n32 : n68825;
  assign n68827 = pi12 ? n32 : n68826;
  assign n68828 = pi11 ? n32 : n68827;
  assign n68829 = pi10 ? n32 : n68828;
  assign n68830 = pi15 ? n26951 : n38913;
  assign n68831 = pi14 ? n68830 : n17466;
  assign n68832 = pi15 ? n17348 : n26425;
  assign n68833 = pi14 ? n17465 : n68832;
  assign n68834 = pi13 ? n68831 : n68833;
  assign n68835 = pi15 ? n26462 : n32;
  assign n68836 = pi14 ? n68835 : n38938;
  assign n68837 = pi14 ? n38814 : n52973;
  assign n68838 = pi13 ? n68836 : n68837;
  assign n68839 = pi12 ? n68834 : n68838;
  assign n68840 = pi20 ? n321 : n20353;
  assign n68841 = pi19 ? n32 : n68840;
  assign n68842 = pi18 ? n32 : n68841;
  assign n68843 = pi17 ? n32 : n68842;
  assign n68844 = pi16 ? n32 : n68843;
  assign n68845 = pi15 ? n68844 : n68552;
  assign n68846 = pi15 ? n53963 : n26272;
  assign n68847 = pi14 ? n68845 : n68846;
  assign n68848 = pi15 ? n17348 : n53119;
  assign n68849 = pi15 ? n53119 : n17286;
  assign n68850 = pi14 ? n68848 : n68849;
  assign n68851 = pi13 ? n68847 : n68850;
  assign n68852 = pi15 ? n26400 : n68724;
  assign n68853 = pi14 ? n68852 : n26760;
  assign n68854 = pi20 ? n246 : n274;
  assign n68855 = pi19 ? n32 : n68854;
  assign n68856 = pi18 ? n32 : n68855;
  assign n68857 = pi17 ? n32 : n68856;
  assign n68858 = pi16 ? n32 : n68857;
  assign n68859 = pi15 ? n25904 : n68858;
  assign n68860 = pi14 ? n68568 : n68859;
  assign n68861 = pi13 ? n68853 : n68860;
  assign n68862 = pi12 ? n68851 : n68861;
  assign n68863 = pi11 ? n68839 : n68862;
  assign n68864 = pi19 ? n32 : n32856;
  assign n68865 = pi18 ? n32 : n68864;
  assign n68866 = pi17 ? n32 : n68865;
  assign n68867 = pi16 ? n32 : n68866;
  assign n68868 = pi15 ? n68867 : n39775;
  assign n68869 = pi14 ? n25997 : n68868;
  assign n68870 = pi15 ? n68747 : n16392;
  assign n68871 = pi14 ? n68587 : n68870;
  assign n68872 = pi13 ? n68869 : n68871;
  assign n68873 = pi20 ? n151 : n321;
  assign n68874 = pi19 ? n68873 : n4342;
  assign n68875 = pi18 ? n32 : n68874;
  assign n68876 = pi18 ? n16847 : n24054;
  assign n68877 = pi17 ? n68875 : n68876;
  assign n68878 = pi16 ? n32 : n68877;
  assign n68879 = pi19 ? n594 : n176;
  assign n68880 = pi18 ? n32 : n68879;
  assign n68881 = pi17 ? n68880 : n55195;
  assign n68882 = pi16 ? n32 : n68881;
  assign n68883 = pi15 ? n68878 : n68882;
  assign n68884 = pi21 ? n405 : ~n7659;
  assign n68885 = pi20 ? n68884 : n32;
  assign n68886 = pi19 ? n18330 : n68885;
  assign n68887 = pi18 ? n32 : n68886;
  assign n68888 = pi17 ? n68887 : n24872;
  assign n68889 = pi16 ? n32 : n68888;
  assign n68890 = pi17 ? n21541 : n16784;
  assign n68891 = pi16 ? n32 : n68890;
  assign n68892 = pi15 ? n68889 : n68891;
  assign n68893 = pi14 ? n68883 : n68892;
  assign n68894 = pi19 ? n32 : ~n60048;
  assign n68895 = pi18 ? n32 : n68894;
  assign n68896 = pi17 ? n32 : n68895;
  assign n68897 = pi16 ? n32 : n68896;
  assign n68898 = pi15 ? n68897 : n50949;
  assign n68899 = pi14 ? n68898 : n27453;
  assign n68900 = pi13 ? n68893 : n68899;
  assign n68901 = pi12 ? n68872 : n68900;
  assign n68902 = pi19 ? n857 : ~n7014;
  assign n68903 = pi18 ? n32 : n68902;
  assign n68904 = pi17 ? n32 : n68903;
  assign n68905 = pi16 ? n32 : n68904;
  assign n68906 = pi15 ? n68905 : n68622;
  assign n68907 = pi19 ? n14260 : ~n28957;
  assign n68908 = pi18 ? n32 : n68907;
  assign n68909 = pi19 ? n321 : n32302;
  assign n68910 = pi19 ? n349 : ~n6230;
  assign n68911 = pi18 ? n68909 : ~n68910;
  assign n68912 = pi17 ? n68908 : n68911;
  assign n68913 = pi16 ? n32 : n68912;
  assign n68914 = pi15 ? n23725 : n68913;
  assign n68915 = pi14 ? n68906 : n68914;
  assign n68916 = pi18 ? n322 : ~n35698;
  assign n68917 = pi17 ? n2531 : ~n68916;
  assign n68918 = pi16 ? n32 : n68917;
  assign n68919 = pi15 ? n68918 : n68779;
  assign n68920 = pi18 ? n940 : n38172;
  assign n68921 = pi17 ? n14154 : n68920;
  assign n68922 = pi16 ? n32 : n68921;
  assign n68923 = pi19 ? n1464 : ~n5626;
  assign n68924 = pi18 ? n17879 : n68923;
  assign n68925 = pi17 ? n2531 : ~n68924;
  assign n68926 = pi16 ? n32 : n68925;
  assign n68927 = pi15 ? n68922 : n68926;
  assign n68928 = pi14 ? n68919 : n68927;
  assign n68929 = pi13 ? n68915 : n68928;
  assign n68930 = pi17 ? n2319 : ~n68658;
  assign n68931 = pi16 ? n32 : n68930;
  assign n68932 = pi20 ? n428 : n915;
  assign n68933 = pi19 ? n68932 : n322;
  assign n68934 = pi18 ? n32 : n68933;
  assign n68935 = pi18 ? n46739 : ~n1541;
  assign n68936 = pi17 ? n68934 : ~n68935;
  assign n68937 = pi16 ? n32 : n68936;
  assign n68938 = pi15 ? n68931 : n68937;
  assign n68939 = pi20 ? n32 : ~n259;
  assign n68940 = pi19 ? n68939 : n19749;
  assign n68941 = pi18 ? n32 : n68940;
  assign n68942 = pi19 ? n5356 : ~n32;
  assign n68943 = pi18 ? n1819 : ~n68942;
  assign n68944 = pi17 ? n68941 : n68943;
  assign n68945 = pi16 ? n32 : n68944;
  assign n68946 = pi18 ? n20164 : ~n48270;
  assign n68947 = pi17 ? n13950 : n68946;
  assign n68948 = pi16 ? n32 : n68947;
  assign n68949 = pi15 ? n68945 : n68948;
  assign n68950 = pi14 ? n68938 : n68949;
  assign n68951 = pi20 ? n101 : n357;
  assign n68952 = pi19 ? n68951 : n32;
  assign n68953 = pi18 ? n32 : n68952;
  assign n68954 = pi17 ? n68953 : n68684;
  assign n68955 = pi16 ? n32 : n68954;
  assign n68956 = pi20 ? n101 : n2358;
  assign n68957 = pi19 ? n68956 : n18396;
  assign n68958 = pi18 ? n32 : n68957;
  assign n68959 = pi19 ? n5694 : n267;
  assign n68960 = pi20 ? n32 : n7448;
  assign n68961 = pi19 ? n68960 : n32;
  assign n68962 = pi18 ? n68959 : n68961;
  assign n68963 = pi17 ? n68958 : n68962;
  assign n68964 = pi16 ? n32 : n68963;
  assign n68965 = pi15 ? n68955 : n68964;
  assign n68966 = pi20 ? n101 : ~n260;
  assign n68967 = pi19 ? n68966 : ~n207;
  assign n68968 = pi18 ? n32 : n68967;
  assign n68969 = pi17 ? n68968 : n38114;
  assign n68970 = pi16 ? n32 : n68969;
  assign n68971 = pi19 ? n16915 : ~n5694;
  assign n68972 = pi18 ? n32 : n68971;
  assign n68973 = pi17 ? n68972 : ~n5779;
  assign n68974 = pi16 ? n32 : n68973;
  assign n68975 = pi15 ? n68970 : n68974;
  assign n68976 = pi14 ? n68965 : n68975;
  assign n68977 = pi13 ? n68950 : n68976;
  assign n68978 = pi12 ? n68929 : n68977;
  assign n68979 = pi11 ? n68901 : n68978;
  assign n68980 = pi10 ? n68863 : n68979;
  assign n68981 = pi09 ? n68829 : n68980;
  assign n68982 = pi13 ? n68831 : n39034;
  assign n68983 = pi14 ? n68835 : n32;
  assign n68984 = pi13 ? n68983 : n32;
  assign n68985 = pi12 ? n68982 : n68984;
  assign n68986 = pi20 ? n321 : n726;
  assign n68987 = pi19 ? n32 : n68986;
  assign n68988 = pi18 ? n32 : n68987;
  assign n68989 = pi17 ? n32 : n68988;
  assign n68990 = pi16 ? n32 : n68989;
  assign n68991 = pi16 ? n32 : n48276;
  assign n68992 = pi15 ? n68991 : n26272;
  assign n68993 = pi14 ? n68990 : n68992;
  assign n68994 = pi13 ? n68993 : n68850;
  assign n68995 = pi14 ? n68725 : n26760;
  assign n68996 = pi15 ? n25904 : n16452;
  assign n68997 = pi14 ? n68568 : n68996;
  assign n68998 = pi13 ? n68995 : n68997;
  assign n68999 = pi12 ? n68994 : n68998;
  assign n69000 = pi11 ? n68985 : n68999;
  assign n69001 = pi20 ? n749 : n481;
  assign n69002 = pi19 ? n32 : n69001;
  assign n69003 = pi18 ? n32 : n69002;
  assign n69004 = pi17 ? n32 : n69003;
  assign n69005 = pi16 ? n32 : n69004;
  assign n69006 = pi15 ? n68867 : n69005;
  assign n69007 = pi14 ? n25997 : n69006;
  assign n69008 = pi18 ? n32 : n28640;
  assign n69009 = pi17 ? n32 : n69008;
  assign n69010 = pi16 ? n32 : n69009;
  assign n69011 = pi19 ? n32 : n42365;
  assign n69012 = pi18 ? n32 : n69011;
  assign n69013 = pi17 ? n32 : n69012;
  assign n69014 = pi16 ? n32 : n69013;
  assign n69015 = pi15 ? n69010 : n69014;
  assign n69016 = pi21 ? n405 : n1392;
  assign n69017 = pi20 ? n69016 : n32;
  assign n69018 = pi19 ? n32 : n69017;
  assign n69019 = pi18 ? n32 : n69018;
  assign n69020 = pi17 ? n32 : n69019;
  assign n69021 = pi16 ? n32 : n69020;
  assign n69022 = pi15 ? n68747 : n69021;
  assign n69023 = pi14 ? n69015 : n69022;
  assign n69024 = pi13 ? n69007 : n69023;
  assign n69025 = pi17 ? n53130 : n68876;
  assign n69026 = pi16 ? n32 : n69025;
  assign n69027 = pi20 ? n32 : n55061;
  assign n69028 = pi19 ? n69027 : n4670;
  assign n69029 = pi18 ? n32 : n69028;
  assign n69030 = pi21 ? n405 : ~n13784;
  assign n69031 = pi20 ? n69030 : ~n32;
  assign n69032 = pi19 ? n32 : ~n69031;
  assign n69033 = pi18 ? n32 : n69032;
  assign n69034 = pi17 ? n69029 : n69033;
  assign n69035 = pi16 ? n32 : n69034;
  assign n69036 = pi15 ? n69026 : n69035;
  assign n69037 = pi21 ? n174 : n14513;
  assign n69038 = pi20 ? n32 : n69037;
  assign n69039 = pi19 ? n69038 : n18789;
  assign n69040 = pi18 ? n32 : n69039;
  assign n69041 = pi17 ? n69040 : n24872;
  assign n69042 = pi16 ? n32 : n69041;
  assign n69043 = pi19 ? n1818 : n16542;
  assign n69044 = pi18 ? n32 : n69043;
  assign n69045 = pi21 ? n405 : n51;
  assign n69046 = pi20 ? n69045 : n32;
  assign n69047 = pi19 ? n32 : n69046;
  assign n69048 = pi18 ? n32 : n69047;
  assign n69049 = pi17 ? n69044 : n69048;
  assign n69050 = pi16 ? n32 : n69049;
  assign n69051 = pi15 ? n69042 : n69050;
  assign n69052 = pi14 ? n69036 : n69051;
  assign n69053 = pi14 ? n68898 : n38638;
  assign n69054 = pi13 ? n69052 : n69053;
  assign n69055 = pi12 ? n69024 : n69054;
  assign n69056 = pi19 ? n507 : ~n7014;
  assign n69057 = pi18 ? n32 : n69056;
  assign n69058 = pi17 ? n32 : n69057;
  assign n69059 = pi16 ? n32 : n69058;
  assign n69060 = pi15 ? n69059 : n68622;
  assign n69061 = pi19 ? n208 : ~n28957;
  assign n69062 = pi18 ? n32 : n69061;
  assign n69063 = pi17 ? n69062 : n68911;
  assign n69064 = pi16 ? n32 : n69063;
  assign n69065 = pi15 ? n23725 : n69064;
  assign n69066 = pi14 ? n69060 : n69065;
  assign n69067 = pi17 ? n2299 : ~n68916;
  assign n69068 = pi16 ? n32 : n69067;
  assign n69069 = pi17 ? n2299 : ~n68640;
  assign n69070 = pi16 ? n32 : n69069;
  assign n69071 = pi15 ? n69068 : n69070;
  assign n69072 = pi18 ? n32 : n68923;
  assign n69073 = pi17 ? n2531 : ~n69072;
  assign n69074 = pi16 ? n32 : n69073;
  assign n69075 = pi15 ? n68922 : n69074;
  assign n69076 = pi14 ? n69071 : n69075;
  assign n69077 = pi13 ? n69066 : n69076;
  assign n69078 = pi17 ? n2653 : ~n68658;
  assign n69079 = pi16 ? n32 : n69078;
  assign n69080 = pi19 ? n267 : n322;
  assign n69081 = pi18 ? n32 : n69080;
  assign n69082 = pi17 ? n69081 : ~n68935;
  assign n69083 = pi16 ? n32 : n69082;
  assign n69084 = pi15 ? n69079 : n69083;
  assign n69085 = pi19 ? n1818 : n3495;
  assign n69086 = pi18 ? n32 : n69085;
  assign n69087 = pi18 ? n32 : ~n68942;
  assign n69088 = pi17 ? n69086 : n69087;
  assign n69089 = pi16 ? n32 : n69088;
  assign n69090 = pi17 ? n32 : n68946;
  assign n69091 = pi16 ? n32 : n69090;
  assign n69092 = pi15 ? n69089 : n69091;
  assign n69093 = pi14 ? n69084 : n69092;
  assign n69094 = pi20 ? n321 : n175;
  assign n69095 = pi19 ? n69094 : n32;
  assign n69096 = pi18 ? n32 : n69095;
  assign n69097 = pi17 ? n32 : n69096;
  assign n69098 = pi16 ? n32 : n69097;
  assign n69099 = pi19 ? n322 : n41419;
  assign n69100 = pi18 ? n32 : n69099;
  assign n69101 = pi17 ? n69100 : n68962;
  assign n69102 = pi16 ? n32 : n69101;
  assign n69103 = pi15 ? n69098 : n69102;
  assign n69104 = pi19 ? n507 : ~n207;
  assign n69105 = pi18 ? n32 : n69104;
  assign n69106 = pi18 ? n268 : n25116;
  assign n69107 = pi17 ? n69105 : n69106;
  assign n69108 = pi16 ? n32 : n69107;
  assign n69109 = pi19 ? n6057 : ~n5694;
  assign n69110 = pi18 ? n32 : n69109;
  assign n69111 = pi17 ? n69110 : ~n5779;
  assign n69112 = pi16 ? n32 : n69111;
  assign n69113 = pi15 ? n69108 : n69112;
  assign n69114 = pi14 ? n69103 : n69113;
  assign n69115 = pi13 ? n69093 : n69114;
  assign n69116 = pi12 ? n69077 : n69115;
  assign n69117 = pi11 ? n69055 : n69116;
  assign n69118 = pi10 ? n69000 : n69117;
  assign n69119 = pi09 ? n68829 : n69118;
  assign n69120 = pi08 ? n68981 : n69119;
  assign n69121 = pi07 ? n68824 : n69120;
  assign n69122 = pi06 ? n68531 : n69121;
  assign n69123 = pi14 ? n32 : n17488;
  assign n69124 = pi13 ? n32 : n69123;
  assign n69125 = pi12 ? n32 : n69124;
  assign n69126 = pi11 ? n32 : n69125;
  assign n69127 = pi10 ? n32 : n69126;
  assign n69128 = pi15 ? n17316 : n17607;
  assign n69129 = pi15 ? n17316 : n17193;
  assign n69130 = pi14 ? n69128 : n69129;
  assign n69131 = pi13 ? n69130 : n17278;
  assign n69132 = pi14 ? n32 : n39083;
  assign n69133 = pi13 ? n27102 : n69132;
  assign n69134 = pi12 ? n69131 : n69133;
  assign n69135 = pi17 ? n32 : n47671;
  assign n69136 = pi16 ? n32 : n69135;
  assign n69137 = pi15 ? n15847 : n69136;
  assign n69138 = pi15 ? n68991 : n26269;
  assign n69139 = pi14 ? n69137 : n69138;
  assign n69140 = pi20 ? n428 : n1817;
  assign n69141 = pi19 ? n32 : n69140;
  assign n69142 = pi18 ? n32 : n69141;
  assign n69143 = pi17 ? n32 : n69142;
  assign n69144 = pi16 ? n32 : n69143;
  assign n69145 = pi15 ? n69144 : n26269;
  assign n69146 = pi14 ? n16852 : n69145;
  assign n69147 = pi13 ? n69139 : n69146;
  assign n69148 = pi15 ? n16736 : n68724;
  assign n69149 = pi14 ? n69148 : n67185;
  assign n69150 = pi15 ? n16452 : n66880;
  assign n69151 = pi14 ? n68568 : n69150;
  assign n69152 = pi13 ? n69149 : n69151;
  assign n69153 = pi12 ? n69147 : n69152;
  assign n69154 = pi11 ? n69134 : n69153;
  assign n69155 = pi19 ? n322 : n21486;
  assign n69156 = pi18 ? n32 : n69155;
  assign n69157 = pi17 ? n32 : n69156;
  assign n69158 = pi16 ? n32 : n69157;
  assign n69159 = pi19 ? n322 : n8622;
  assign n69160 = pi18 ? n32 : n69159;
  assign n69161 = pi17 ? n32 : n69160;
  assign n69162 = pi16 ? n32 : n69161;
  assign n69163 = pi15 ? n69158 : n69162;
  assign n69164 = pi20 ? n207 : n481;
  assign n69165 = pi19 ? n32 : n69164;
  assign n69166 = pi18 ? n32 : n69165;
  assign n69167 = pi17 ? n32 : n69166;
  assign n69168 = pi16 ? n32 : n69167;
  assign n69169 = pi15 ? n69168 : n15531;
  assign n69170 = pi14 ? n69163 : n69169;
  assign n69171 = pi15 ? n16984 : n15847;
  assign n69172 = pi20 ? n382 : n141;
  assign n69173 = pi19 ? n322 : ~n69172;
  assign n69174 = pi18 ? n32 : n69173;
  assign n69175 = pi17 ? n32 : n69174;
  assign n69176 = pi16 ? n32 : n69175;
  assign n69177 = pi18 ? n32 : n9745;
  assign n69178 = pi19 ? n5356 : n6298;
  assign n69179 = pi18 ? n32 : ~n69178;
  assign n69180 = pi17 ? n69177 : n69179;
  assign n69181 = pi16 ? n32 : n69180;
  assign n69182 = pi15 ? n69176 : n69181;
  assign n69183 = pi14 ? n69171 : n69182;
  assign n69184 = pi13 ? n69170 : n69183;
  assign n69185 = pi15 ? n32 : n27528;
  assign n69186 = pi17 ? n21926 : n15228;
  assign n69187 = pi16 ? n32 : n69186;
  assign n69188 = pi20 ? n7939 : ~n175;
  assign n69189 = pi19 ? n69188 : ~n507;
  assign n69190 = pi19 ? n1612 : n112;
  assign n69191 = pi18 ? n69189 : ~n69190;
  assign n69192 = pi17 ? n22085 : ~n69191;
  assign n69193 = pi16 ? n32 : n69192;
  assign n69194 = pi15 ? n69187 : n69193;
  assign n69195 = pi14 ? n69185 : n69194;
  assign n69196 = pi15 ? n50949 : n24700;
  assign n69197 = pi15 ? n24247 : n22817;
  assign n69198 = pi14 ? n69196 : n69197;
  assign n69199 = pi13 ? n69195 : n69198;
  assign n69200 = pi12 ? n69184 : n69199;
  assign n69201 = pi15 ? n66408 : n24247;
  assign n69202 = pi19 ? n1818 : n321;
  assign n69203 = pi18 ? n32 : n69202;
  assign n69204 = pi19 ? n28686 : ~n1490;
  assign n69205 = pi18 ? n69204 : ~n34250;
  assign n69206 = pi17 ? n69203 : n69205;
  assign n69207 = pi16 ? n32 : n69206;
  assign n69208 = pi18 ? n32 : n59923;
  assign n69209 = pi17 ? n69208 : ~n2724;
  assign n69210 = pi16 ? n32 : n69209;
  assign n69211 = pi15 ? n69207 : n69210;
  assign n69212 = pi14 ? n69201 : n69211;
  assign n69213 = pi19 ? n267 : ~n32;
  assign n69214 = pi18 ? n32 : n69213;
  assign n69215 = pi17 ? n69214 : ~n8472;
  assign n69216 = pi16 ? n32 : n69215;
  assign n69217 = pi17 ? n69214 : ~n7931;
  assign n69218 = pi16 ? n32 : n69217;
  assign n69219 = pi15 ? n69216 : n69218;
  assign n69220 = pi17 ? n48428 : ~n2750;
  assign n69221 = pi16 ? n32 : n69220;
  assign n69222 = pi19 ? n1508 : ~n5626;
  assign n69223 = pi18 ? n32 : n69222;
  assign n69224 = pi17 ? n2292 : ~n69223;
  assign n69225 = pi16 ? n32 : n69224;
  assign n69226 = pi15 ? n69221 : n69225;
  assign n69227 = pi14 ? n69219 : n69226;
  assign n69228 = pi13 ? n69212 : n69227;
  assign n69229 = pi19 ? n4982 : n617;
  assign n69230 = pi18 ? n32 : n69229;
  assign n69231 = pi17 ? n2292 : ~n69230;
  assign n69232 = pi16 ? n32 : n69231;
  assign n69233 = pi19 ? n267 : n23895;
  assign n69234 = pi18 ? n69233 : n6145;
  assign n69235 = pi17 ? n15845 : n69234;
  assign n69236 = pi16 ? n32 : n69235;
  assign n69237 = pi15 ? n69232 : n69236;
  assign n69238 = pi18 ? n16847 : n20912;
  assign n69239 = pi17 ? n19886 : n69238;
  assign n69240 = pi16 ? n32 : n69239;
  assign n69241 = pi15 ? n22817 : n69240;
  assign n69242 = pi14 ? n69237 : n69241;
  assign n69243 = pi17 ? n20011 : n32;
  assign n69244 = pi16 ? n32 : n69243;
  assign n69245 = pi15 ? n69244 : n648;
  assign n69246 = pi19 ? n32 : ~n11899;
  assign n69247 = pi18 ? n32 : n69246;
  assign n69248 = pi19 ? n34031 : n28179;
  assign n69249 = pi19 ? n6308 : n32;
  assign n69250 = pi18 ? n69248 : ~n69249;
  assign n69251 = pi17 ? n69247 : ~n69250;
  assign n69252 = pi16 ? n32 : n69251;
  assign n69253 = pi19 ? n519 : n25120;
  assign n69254 = pi18 ? n32 : n69253;
  assign n69255 = pi18 ? n350 : ~n46010;
  assign n69256 = pi17 ? n69254 : n69255;
  assign n69257 = pi16 ? n32 : n69256;
  assign n69258 = pi15 ? n69252 : n69257;
  assign n69259 = pi14 ? n69245 : n69258;
  assign n69260 = pi13 ? n69242 : n69259;
  assign n69261 = pi12 ? n69228 : n69260;
  assign n69262 = pi11 ? n69200 : n69261;
  assign n69263 = pi10 ? n69154 : n69262;
  assign n69264 = pi09 ? n69127 : n69263;
  assign n69265 = pi15 ? n17278 : n17316;
  assign n69266 = pi14 ? n69265 : n53212;
  assign n69267 = pi13 ? n69130 : n69266;
  assign n69268 = pi14 ? n32 : n17279;
  assign n69269 = pi13 ? n27102 : n69268;
  assign n69270 = pi12 ? n69267 : n69269;
  assign n69271 = pi20 ? n321 : n111;
  assign n69272 = pi19 ? n32 : n69271;
  assign n69273 = pi18 ? n32 : n69272;
  assign n69274 = pi17 ? n32 : n69273;
  assign n69275 = pi16 ? n32 : n69274;
  assign n69276 = pi20 ? n321 : ~n17134;
  assign n69277 = pi19 ? n32 : n69276;
  assign n69278 = pi18 ? n32 : n69277;
  assign n69279 = pi17 ? n32 : n69278;
  assign n69280 = pi16 ? n32 : n69279;
  assign n69281 = pi15 ? n69275 : n69280;
  assign n69282 = pi14 ? n69281 : n69138;
  assign n69283 = pi13 ? n69282 : n69146;
  assign n69284 = pi12 ? n69283 : n69152;
  assign n69285 = pi11 ? n69270 : n69284;
  assign n69286 = pi15 ? n66910 : n69181;
  assign n69287 = pi14 ? n69171 : n69286;
  assign n69288 = pi13 ? n69170 : n69287;
  assign n69289 = pi15 ? n16377 : n27528;
  assign n69290 = pi19 ? n69188 : ~n857;
  assign n69291 = pi18 ? n69290 : ~n69190;
  assign n69292 = pi17 ? n32 : ~n69291;
  assign n69293 = pi16 ? n32 : n69292;
  assign n69294 = pi15 ? n69187 : n69293;
  assign n69295 = pi14 ? n69289 : n69294;
  assign n69296 = pi13 ? n69295 : n69198;
  assign n69297 = pi12 ? n69288 : n69296;
  assign n69298 = pi19 ? n1464 : n321;
  assign n69299 = pi18 ? n32 : n69298;
  assign n69300 = pi19 ? n18377 : ~n54803;
  assign n69301 = pi19 ? n12572 : ~n32;
  assign n69302 = pi18 ? n69300 : ~n69301;
  assign n69303 = pi17 ? n69299 : n69302;
  assign n69304 = pi16 ? n32 : n69303;
  assign n69305 = pi17 ? n2519 : ~n2724;
  assign n69306 = pi16 ? n32 : n69305;
  assign n69307 = pi15 ? n69304 : n69306;
  assign n69308 = pi14 ? n69201 : n69307;
  assign n69309 = pi17 ? n2750 : ~n6236;
  assign n69310 = pi16 ? n32 : n69309;
  assign n69311 = pi17 ? n2750 : ~n7931;
  assign n69312 = pi16 ? n32 : n69311;
  assign n69313 = pi15 ? n69310 : n69312;
  assign n69314 = pi17 ? n2748 : ~n69223;
  assign n69315 = pi16 ? n32 : n69314;
  assign n69316 = pi15 ? n69221 : n69315;
  assign n69317 = pi14 ? n69313 : n69316;
  assign n69318 = pi13 ? n69308 : n69317;
  assign n69319 = pi17 ? n2748 : ~n69230;
  assign n69320 = pi16 ? n32 : n69319;
  assign n69321 = pi15 ? n69320 : n69236;
  assign n69322 = pi19 ? n1320 : n32;
  assign n69323 = pi18 ? n32 : n69322;
  assign n69324 = pi17 ? n32 : n69323;
  assign n69325 = pi16 ? n32 : n69324;
  assign n69326 = pi17 ? n32 : n69238;
  assign n69327 = pi16 ? n32 : n69326;
  assign n69328 = pi15 ? n69325 : n69327;
  assign n69329 = pi14 ? n69321 : n69328;
  assign n69330 = pi17 ? n40575 : n21317;
  assign n69331 = pi16 ? n32 : n69330;
  assign n69332 = pi15 ? n69331 : n648;
  assign n69333 = pi19 ? n1574 : ~n11899;
  assign n69334 = pi18 ? n32 : n69333;
  assign n69335 = pi17 ? n69334 : ~n69250;
  assign n69336 = pi16 ? n32 : n69335;
  assign n69337 = pi19 ? n32 : n25120;
  assign n69338 = pi18 ? n32 : n69337;
  assign n69339 = pi18 ? n350 : ~n22872;
  assign n69340 = pi17 ? n69338 : n69339;
  assign n69341 = pi16 ? n32 : n69340;
  assign n69342 = pi15 ? n69336 : n69341;
  assign n69343 = pi14 ? n69332 : n69342;
  assign n69344 = pi13 ? n69329 : n69343;
  assign n69345 = pi12 ? n69318 : n69344;
  assign n69346 = pi11 ? n69297 : n69345;
  assign n69347 = pi10 ? n69285 : n69346;
  assign n69348 = pi09 ? n69127 : n69347;
  assign n69349 = pi08 ? n69264 : n69348;
  assign n69350 = pi14 ? n32 : n17465;
  assign n69351 = pi14 ? n32 : n39155;
  assign n69352 = pi13 ? n69350 : n69351;
  assign n69353 = pi12 ? n17465 : n69352;
  assign n69354 = pi15 ? n69275 : n69136;
  assign n69355 = pi14 ? n69354 : n69138;
  assign n69356 = pi15 ? n16850 : n53119;
  assign n69357 = pi15 ? n26269 : n32;
  assign n69358 = pi14 ? n69356 : n69357;
  assign n69359 = pi13 ? n69355 : n69358;
  assign n69360 = pi15 ? n68564 : n68724;
  assign n69361 = pi14 ? n69360 : n67185;
  assign n69362 = pi15 ? n24874 : n67449;
  assign n69363 = pi14 ? n26322 : n69362;
  assign n69364 = pi13 ? n69361 : n69363;
  assign n69365 = pi12 ? n69359 : n69364;
  assign n69366 = pi11 ? n69353 : n69365;
  assign n69367 = pi19 ? n322 : n8035;
  assign n69368 = pi18 ? n32 : n69367;
  assign n69369 = pi17 ? n32 : n69368;
  assign n69370 = pi16 ? n32 : n69369;
  assign n69371 = pi15 ? n69158 : n69370;
  assign n69372 = pi15 ? n69005 : n69010;
  assign n69373 = pi14 ? n69371 : n69372;
  assign n69374 = pi15 ? n69014 : n16485;
  assign n69375 = pi19 ? n4964 : n349;
  assign n69376 = pi18 ? n32 : ~n69375;
  assign n69377 = pi17 ? n8193 : n69376;
  assign n69378 = pi16 ? n32 : n69377;
  assign n69379 = pi15 ? n66910 : n69378;
  assign n69380 = pi14 ? n69374 : n69379;
  assign n69381 = pi13 ? n69373 : n69380;
  assign n69382 = pi20 ? n65551 : n32;
  assign n69383 = pi19 ? n32 : n69382;
  assign n69384 = pi18 ? n32 : n69383;
  assign n69385 = pi17 ? n32 : n69384;
  assign n69386 = pi16 ? n32 : n69385;
  assign n69387 = pi15 ? n69386 : n27528;
  assign n69388 = pi19 ? n18489 : ~n343;
  assign n69389 = pi18 ? n32 : n69388;
  assign n69390 = pi17 ? n53261 : n69389;
  assign n69391 = pi16 ? n32 : n69390;
  assign n69392 = pi15 ? n69391 : n22540;
  assign n69393 = pi14 ? n69387 : n69392;
  assign n69394 = pi19 ? n857 : n247;
  assign n69395 = pi18 ? n32 : n69394;
  assign n69396 = pi17 ? n32 : n69395;
  assign n69397 = pi16 ? n32 : n69396;
  assign n69398 = pi19 ? n857 : ~n343;
  assign n69399 = pi18 ? n32 : n69398;
  assign n69400 = pi17 ? n32 : n69399;
  assign n69401 = pi16 ? n32 : n69400;
  assign n69402 = pi15 ? n69397 : n69401;
  assign n69403 = pi15 ? n15362 : n69325;
  assign n69404 = pi14 ? n69402 : n69403;
  assign n69405 = pi13 ? n69393 : n69404;
  assign n69406 = pi12 ? n69381 : n69405;
  assign n69407 = pi19 ? n4518 : ~n2848;
  assign n69408 = pi18 ? n32 : n69407;
  assign n69409 = pi17 ? n32 : n69408;
  assign n69410 = pi16 ? n32 : n69409;
  assign n69411 = pi15 ? n69410 : n15244;
  assign n69412 = pi19 ? n32 : n18502;
  assign n69413 = pi18 ? n32 : n69412;
  assign n69414 = pi19 ? n29444 : n342;
  assign n69415 = pi19 ? n12572 : ~n5614;
  assign n69416 = pi18 ? n69414 : n69415;
  assign n69417 = pi17 ? n69413 : ~n69416;
  assign n69418 = pi16 ? n32 : n69417;
  assign n69419 = pi17 ? n2736 : ~n2724;
  assign n69420 = pi16 ? n32 : n69419;
  assign n69421 = pi15 ? n69418 : n69420;
  assign n69422 = pi14 ? n69411 : n69421;
  assign n69423 = pi19 ? n1574 : n617;
  assign n69424 = pi18 ? n32 : n69423;
  assign n69425 = pi17 ? n69424 : ~n6236;
  assign n69426 = pi16 ? n32 : n69425;
  assign n69427 = pi17 ? n69424 : ~n35572;
  assign n69428 = pi16 ? n32 : n69427;
  assign n69429 = pi15 ? n69426 : n69428;
  assign n69430 = pi18 ? n32 : n1886;
  assign n69431 = pi17 ? n69430 : ~n2750;
  assign n69432 = pi16 ? n32 : n69431;
  assign n69433 = pi17 ? n2750 : ~n68658;
  assign n69434 = pi16 ? n32 : n69433;
  assign n69435 = pi15 ? n69432 : n69434;
  assign n69436 = pi14 ? n69429 : n69435;
  assign n69437 = pi13 ? n69422 : n69436;
  assign n69438 = pi19 ? n4982 : n1105;
  assign n69439 = pi18 ? n32 : n69438;
  assign n69440 = pi17 ? n2855 : ~n69439;
  assign n69441 = pi16 ? n32 : n69440;
  assign n69442 = pi20 ? n357 : ~n9491;
  assign n69443 = pi19 ? n69442 : n36184;
  assign n69444 = pi20 ? n14286 : n342;
  assign n69445 = pi19 ? n69444 : n32;
  assign n69446 = pi18 ? n69443 : n69445;
  assign n69447 = pi17 ? n15964 : n69446;
  assign n69448 = pi16 ? n32 : n69447;
  assign n69449 = pi15 ? n69441 : n69448;
  assign n69450 = pi17 ? n23572 : n69238;
  assign n69451 = pi16 ? n32 : n69450;
  assign n69452 = pi15 ? n22437 : n69451;
  assign n69453 = pi14 ? n69449 : n69452;
  assign n69454 = pi17 ? n23572 : n14392;
  assign n69455 = pi16 ? n32 : n69454;
  assign n69456 = pi15 ? n69455 : n648;
  assign n69457 = pi20 ? n10878 : ~n6303;
  assign n69458 = pi19 ? n32 : n69457;
  assign n69459 = pi18 ? n32 : n69458;
  assign n69460 = pi19 ? n45418 : ~n32;
  assign n69461 = pi18 ? n53303 : n69460;
  assign n69462 = pi17 ? n69459 : ~n69461;
  assign n69463 = pi16 ? n32 : n69462;
  assign n69464 = pi19 ? n32 : n34502;
  assign n69465 = pi18 ? n32 : n69464;
  assign n69466 = pi17 ? n69465 : n69339;
  assign n69467 = pi16 ? n32 : n69466;
  assign n69468 = pi15 ? n69463 : n69467;
  assign n69469 = pi14 ? n69456 : n69468;
  assign n69470 = pi13 ? n69453 : n69469;
  assign n69471 = pi12 ? n69437 : n69470;
  assign n69472 = pi11 ? n69406 : n69471;
  assign n69473 = pi10 ? n69366 : n69472;
  assign n69474 = pi09 ? n17493 : n69473;
  assign n69475 = pi19 ? n18489 : ~n2303;
  assign n69476 = pi18 ? n32 : n69475;
  assign n69477 = pi17 ? n26423 : n69476;
  assign n69478 = pi16 ? n32 : n69477;
  assign n69479 = pi15 ? n69478 : n22540;
  assign n69480 = pi14 ? n69387 : n69479;
  assign n69481 = pi19 ? n1785 : n247;
  assign n69482 = pi18 ? n32 : n69481;
  assign n69483 = pi17 ? n32 : n69482;
  assign n69484 = pi16 ? n32 : n69483;
  assign n69485 = pi19 ? n1785 : ~n589;
  assign n69486 = pi18 ? n32 : n69485;
  assign n69487 = pi17 ? n32 : n69486;
  assign n69488 = pi16 ? n32 : n69487;
  assign n69489 = pi15 ? n69484 : n69488;
  assign n69490 = pi19 ? n519 : n161;
  assign n69491 = pi18 ? n32 : n69490;
  assign n69492 = pi17 ? n32 : n69491;
  assign n69493 = pi16 ? n32 : n69492;
  assign n69494 = pi15 ? n15362 : n69493;
  assign n69495 = pi14 ? n69489 : n69494;
  assign n69496 = pi13 ? n69480 : n69495;
  assign n69497 = pi12 ? n69381 : n69496;
  assign n69498 = pi20 ? n243 : ~n266;
  assign n69499 = pi19 ? n32 : n69498;
  assign n69500 = pi18 ? n32 : n69499;
  assign n69501 = pi17 ? n69500 : ~n69416;
  assign n69502 = pi16 ? n32 : n69501;
  assign n69503 = pi17 ? n2616 : ~n2724;
  assign n69504 = pi16 ? n32 : n69503;
  assign n69505 = pi15 ? n69502 : n69504;
  assign n69506 = pi14 ? n69411 : n69505;
  assign n69507 = pi17 ? n2736 : ~n6236;
  assign n69508 = pi16 ? n32 : n69507;
  assign n69509 = pi17 ? n2736 : ~n35572;
  assign n69510 = pi16 ? n32 : n69509;
  assign n69511 = pi15 ? n69508 : n69510;
  assign n69512 = pi17 ? n3067 : ~n2616;
  assign n69513 = pi16 ? n32 : n69512;
  assign n69514 = pi17 ? n4245 : ~n68658;
  assign n69515 = pi16 ? n32 : n69514;
  assign n69516 = pi15 ? n69513 : n69515;
  assign n69517 = pi14 ? n69511 : n69516;
  assign n69518 = pi13 ? n69506 : n69517;
  assign n69519 = pi17 ? n4245 : ~n69439;
  assign n69520 = pi16 ? n32 : n69519;
  assign n69521 = pi19 ? n267 : n36184;
  assign n69522 = pi18 ? n69521 : n69445;
  assign n69523 = pi17 ? n32 : n69522;
  assign n69524 = pi16 ? n32 : n69523;
  assign n69525 = pi15 ? n69520 : n69524;
  assign n69526 = pi19 ? n1369 : n32;
  assign n69527 = pi18 ? n16847 : n69526;
  assign n69528 = pi17 ? n32 : n69527;
  assign n69529 = pi16 ? n32 : n69528;
  assign n69530 = pi15 ? n22437 : n69529;
  assign n69531 = pi14 ? n69525 : n69530;
  assign n69532 = pi15 ? n22958 : n14973;
  assign n69533 = pi20 ? n175 : ~n1091;
  assign n69534 = pi19 ? n32 : n69533;
  assign n69535 = pi18 ? n32 : n69534;
  assign n69536 = pi20 ? n175 : ~n1685;
  assign n69537 = pi19 ? n69536 : ~n32;
  assign n69538 = pi18 ? n53349 : n69537;
  assign n69539 = pi17 ? n69535 : ~n69538;
  assign n69540 = pi16 ? n32 : n69539;
  assign n69541 = pi19 ? n32 : n68873;
  assign n69542 = pi18 ? n32 : n69541;
  assign n69543 = pi17 ? n69542 : n69339;
  assign n69544 = pi16 ? n32 : n69543;
  assign n69545 = pi15 ? n69540 : n69544;
  assign n69546 = pi14 ? n69532 : n69545;
  assign n69547 = pi13 ? n69531 : n69546;
  assign n69548 = pi12 ? n69518 : n69547;
  assign n69549 = pi11 ? n69497 : n69548;
  assign n69550 = pi10 ? n69366 : n69549;
  assign n69551 = pi09 ? n17493 : n69550;
  assign n69552 = pi08 ? n69474 : n69551;
  assign n69553 = pi07 ? n69349 : n69552;
  assign n69554 = pi13 ? n32 : n69132;
  assign n69555 = pi12 ? n32 : n69554;
  assign n69556 = pi15 ? n69275 : n68991;
  assign n69557 = pi18 ? n32 : n22885;
  assign n69558 = pi17 ? n32 : n69557;
  assign n69559 = pi16 ? n32 : n69558;
  assign n69560 = pi15 ? n69559 : n16392;
  assign n69561 = pi14 ? n69556 : n69560;
  assign n69562 = pi13 ? n69561 : n69358;
  assign n69563 = pi20 ? n175 : ~n11048;
  assign n69564 = pi19 ? n32 : n69563;
  assign n69565 = pi18 ? n32 : n69564;
  assign n69566 = pi17 ? n32 : n69565;
  assign n69567 = pi16 ? n32 : n69566;
  assign n69568 = pi15 ? n32 : n69567;
  assign n69569 = pi14 ? n68564 : n69568;
  assign n69570 = pi15 ? n38750 : n68858;
  assign n69571 = pi15 ? n16237 : n25997;
  assign n69572 = pi14 ? n69570 : n69571;
  assign n69573 = pi13 ? n69569 : n69572;
  assign n69574 = pi12 ? n69562 : n69573;
  assign n69575 = pi11 ? n69555 : n69574;
  assign n69576 = pi19 ? n322 : n21493;
  assign n69577 = pi18 ? n32 : n69576;
  assign n69578 = pi17 ? n32 : n69577;
  assign n69579 = pi16 ? n32 : n69578;
  assign n69580 = pi19 ? n322 : n39771;
  assign n69581 = pi18 ? n248 : n69580;
  assign n69582 = pi17 ? n32 : n69581;
  assign n69583 = pi16 ? n32 : n69582;
  assign n69584 = pi15 ? n69579 : n69583;
  assign n69585 = pi20 ? n266 : ~n243;
  assign n69586 = pi19 ? n32 : n69585;
  assign n69587 = pi18 ? n248 : n69586;
  assign n69588 = pi17 ? n32 : n69587;
  assign n69589 = pi16 ? n32 : n69588;
  assign n69590 = pi19 ? n32 : n7840;
  assign n69591 = pi18 ? n32 : n69590;
  assign n69592 = pi17 ? n32 : n69591;
  assign n69593 = pi16 ? n32 : n69592;
  assign n69594 = pi15 ? n69589 : n69593;
  assign n69595 = pi14 ? n69584 : n69594;
  assign n69596 = pi20 ? n501 : ~n339;
  assign n69597 = pi19 ? n322 : n69596;
  assign n69598 = pi18 ? n32 : n69597;
  assign n69599 = pi17 ? n32 : n69598;
  assign n69600 = pi16 ? n32 : n69599;
  assign n69601 = pi19 ? n1757 : n16828;
  assign n69602 = pi18 ? n53382 : n69601;
  assign n69603 = pi17 ? n4319 : n69602;
  assign n69604 = pi16 ? n32 : n69603;
  assign n69605 = pi15 ? n69600 : n69604;
  assign n69606 = pi19 ? n208 : ~n9340;
  assign n69607 = pi18 ? n32 : ~n69606;
  assign n69608 = pi17 ? n53392 : ~n69607;
  assign n69609 = pi16 ? n32 : n69608;
  assign n69610 = pi18 ? n350 : ~n14567;
  assign n69611 = pi17 ? n32 : ~n69610;
  assign n69612 = pi16 ? n32 : n69611;
  assign n69613 = pi15 ? n69609 : n69612;
  assign n69614 = pi14 ? n69605 : n69613;
  assign n69615 = pi13 ? n69595 : n69614;
  assign n69616 = pi21 ? n405 : ~n10182;
  assign n69617 = pi20 ? n69616 : n32;
  assign n69618 = pi19 ? n9007 : n69617;
  assign n69619 = pi18 ? n32 : n69618;
  assign n69620 = pi17 ? n32 : n69619;
  assign n69621 = pi16 ? n32 : n69620;
  assign n69622 = pi20 ? n18255 : n32;
  assign n69623 = pi19 ? n462 : n69622;
  assign n69624 = pi18 ? n32 : n69623;
  assign n69625 = pi17 ? n32 : n69624;
  assign n69626 = pi16 ? n32 : n69625;
  assign n69627 = pi15 ? n69621 : n69626;
  assign n69628 = pi21 ? n405 : ~n51;
  assign n69629 = pi20 ? n69628 : ~n32;
  assign n69630 = pi19 ? n11374 : ~n69629;
  assign n69631 = pi18 ? n32 : n69630;
  assign n69632 = pi17 ? n32 : n69631;
  assign n69633 = pi16 ? n32 : n69632;
  assign n69634 = pi15 ? n69633 : n16452;
  assign n69635 = pi14 ? n69627 : n69634;
  assign n69636 = pi15 ? n16298 : n55403;
  assign n69637 = pi19 ? n1325 : ~n813;
  assign n69638 = pi18 ? n32 : n69637;
  assign n69639 = pi17 ? n32 : n69638;
  assign n69640 = pi16 ? n32 : n69639;
  assign n69641 = pi19 ? n519 : n7693;
  assign n69642 = pi18 ? n32 : n69641;
  assign n69643 = pi17 ? n32 : n69642;
  assign n69644 = pi16 ? n32 : n69643;
  assign n69645 = pi15 ? n69640 : n69644;
  assign n69646 = pi14 ? n69636 : n69645;
  assign n69647 = pi13 ? n69635 : n69646;
  assign n69648 = pi12 ? n69615 : n69647;
  assign n69649 = pi19 ? n1165 : ~n9368;
  assign n69650 = pi18 ? n32 : n69649;
  assign n69651 = pi17 ? n32 : n69650;
  assign n69652 = pi16 ? n32 : n69651;
  assign n69653 = pi19 ? n594 : n7488;
  assign n69654 = pi18 ? n863 : n69653;
  assign n69655 = pi17 ? n32 : n69654;
  assign n69656 = pi16 ? n32 : n69655;
  assign n69657 = pi15 ? n69652 : n69656;
  assign n69658 = pi19 ? n857 : ~n5614;
  assign n69659 = pi18 ? n32 : n69658;
  assign n69660 = pi17 ? n7039 : ~n69659;
  assign n69661 = pi16 ? n32 : n69660;
  assign n69662 = pi19 ? n1325 : n236;
  assign n69663 = pi18 ? n32 : n69662;
  assign n69664 = pi17 ? n7039 : ~n69663;
  assign n69665 = pi16 ? n32 : n69664;
  assign n69666 = pi15 ? n69661 : n69665;
  assign n69667 = pi14 ? n69657 : n69666;
  assign n69668 = pi19 ? n32 : n13793;
  assign n69669 = pi18 ? n32 : n69668;
  assign n69670 = pi17 ? n69669 : ~n3201;
  assign n69671 = pi16 ? n32 : n69670;
  assign n69672 = pi19 ? n267 : n2614;
  assign n69673 = pi18 ? n32 : n69672;
  assign n69674 = pi17 ? n69669 : ~n69673;
  assign n69675 = pi16 ? n32 : n69674;
  assign n69676 = pi15 ? n69671 : n69675;
  assign n69677 = pi19 ? n208 : n2614;
  assign n69678 = pi18 ? n32 : n69677;
  assign n69679 = pi17 ? n64060 : ~n69678;
  assign n69680 = pi16 ? n32 : n69679;
  assign n69681 = pi17 ? n2733 : ~n7515;
  assign n69682 = pi16 ? n32 : n69681;
  assign n69683 = pi15 ? n69680 : n69682;
  assign n69684 = pi14 ? n69676 : n69683;
  assign n69685 = pi13 ? n69667 : n69684;
  assign n69686 = pi17 ? n2733 : ~n69439;
  assign n69687 = pi16 ? n32 : n69686;
  assign n69688 = pi15 ? n69687 : n22540;
  assign n69689 = pi18 ? n9012 : n14964;
  assign n69690 = pi17 ? n32 : n69689;
  assign n69691 = pi16 ? n32 : n69690;
  assign n69692 = pi20 ? n321 : n10878;
  assign n69693 = pi19 ? n69692 : n32;
  assign n69694 = pi18 ? n32 : n69693;
  assign n69695 = pi17 ? n32 : n69694;
  assign n69696 = pi16 ? n32 : n69695;
  assign n69697 = pi15 ? n69691 : n69696;
  assign n69698 = pi14 ? n69688 : n69697;
  assign n69699 = pi20 ? n32 : n22331;
  assign n69700 = pi19 ? n69699 : n32;
  assign n69701 = pi18 ? n32 : n69700;
  assign n69702 = pi17 ? n16982 : n69701;
  assign n69703 = pi16 ? n32 : n69702;
  assign n69704 = pi17 ? n48231 : n26670;
  assign n69705 = pi16 ? n32 : n69704;
  assign n69706 = pi15 ? n69703 : n69705;
  assign n69707 = pi18 ? n4343 : ~n24476;
  assign n69708 = pi17 ? n17346 : n69707;
  assign n69709 = pi16 ? n32 : n69708;
  assign n69710 = pi20 ? n32 : n406;
  assign n69711 = pi19 ? n32 : n69710;
  assign n69712 = pi18 ? n32 : n69711;
  assign n69713 = pi18 ? n20729 : ~n22872;
  assign n69714 = pi17 ? n69712 : n69713;
  assign n69715 = pi16 ? n32 : n69714;
  assign n69716 = pi15 ? n69709 : n69715;
  assign n69717 = pi14 ? n69706 : n69716;
  assign n69718 = pi13 ? n69698 : n69717;
  assign n69719 = pi12 ? n69685 : n69718;
  assign n69720 = pi11 ? n69648 : n69719;
  assign n69721 = pi10 ? n69575 : n69720;
  assign n69722 = pi09 ? n17493 : n69721;
  assign n69723 = pi13 ? n32 : n69268;
  assign n69724 = pi12 ? n32 : n69723;
  assign n69725 = pi15 ? n15847 : n68991;
  assign n69726 = pi14 ? n69725 : n69560;
  assign n69727 = pi13 ? n69726 : n69358;
  assign n69728 = pi15 ? n67449 : n25997;
  assign n69729 = pi14 ? n69570 : n69728;
  assign n69730 = pi13 ? n69569 : n69729;
  assign n69731 = pi12 ? n69727 : n69730;
  assign n69732 = pi11 ? n69724 : n69731;
  assign n69733 = pi19 ? n322 : n6420;
  assign n69734 = pi18 ? n32 : n69733;
  assign n69735 = pi17 ? n32 : n69734;
  assign n69736 = pi16 ? n32 : n69735;
  assign n69737 = pi20 ? n1475 : n481;
  assign n69738 = pi19 ? n322 : n69737;
  assign n69739 = pi18 ? n248 : n69738;
  assign n69740 = pi17 ? n32 : n69739;
  assign n69741 = pi16 ? n32 : n69740;
  assign n69742 = pi15 ? n69736 : n69741;
  assign n69743 = pi18 ? n19232 : n69586;
  assign n69744 = pi17 ? n32 : n69743;
  assign n69745 = pi16 ? n32 : n69744;
  assign n69746 = pi20 ? n53469 : ~n339;
  assign n69747 = pi19 ? n32 : n69746;
  assign n69748 = pi18 ? n32 : n69747;
  assign n69749 = pi17 ? n32 : n69748;
  assign n69750 = pi16 ? n32 : n69749;
  assign n69751 = pi15 ? n69745 : n69750;
  assign n69752 = pi14 ? n69742 : n69751;
  assign n69753 = pi19 ? n322 : n12854;
  assign n69754 = pi18 ? n32 : n69753;
  assign n69755 = pi17 ? n32 : n69754;
  assign n69756 = pi16 ? n32 : n69755;
  assign n69757 = pi20 ? n9628 : ~n141;
  assign n69758 = pi19 ? n1757 : n69757;
  assign n69759 = pi18 ? n53480 : n69758;
  assign n69760 = pi17 ? n53478 : n69759;
  assign n69761 = pi16 ? n32 : n69760;
  assign n69762 = pi15 ? n69756 : n69761;
  assign n69763 = pi20 ? n220 : n141;
  assign n69764 = pi19 ? n208 : ~n69763;
  assign n69765 = pi18 ? n32 : ~n69764;
  assign n69766 = pi17 ? n53487 : ~n69765;
  assign n69767 = pi16 ? n32 : n69766;
  assign n69768 = pi15 ? n69767 : n69612;
  assign n69769 = pi14 ? n69762 : n69768;
  assign n69770 = pi13 ? n69752 : n69769;
  assign n69771 = pi18 ? n19774 : n69623;
  assign n69772 = pi17 ? n32 : n69771;
  assign n69773 = pi16 ? n32 : n69772;
  assign n69774 = pi15 ? n69621 : n69773;
  assign n69775 = pi14 ? n69774 : n69634;
  assign n69776 = pi13 ? n69775 : n69646;
  assign n69777 = pi12 ? n69770 : n69776;
  assign n69778 = pi17 ? n2963 : ~n69659;
  assign n69779 = pi16 ? n32 : n69778;
  assign n69780 = pi17 ? n2963 : ~n69663;
  assign n69781 = pi16 ? n32 : n69780;
  assign n69782 = pi15 ? n69779 : n69781;
  assign n69783 = pi14 ? n69657 : n69782;
  assign n69784 = pi17 ? n2726 : ~n69673;
  assign n69785 = pi16 ? n32 : n69784;
  assign n69786 = pi15 ? n9403 : n69785;
  assign n69787 = pi17 ? n3050 : ~n67290;
  assign n69788 = pi16 ? n32 : n69787;
  assign n69789 = pi15 ? n69680 : n69788;
  assign n69790 = pi14 ? n69786 : n69789;
  assign n69791 = pi13 ? n69783 : n69790;
  assign n69792 = pi17 ? n3050 : ~n69439;
  assign n69793 = pi16 ? n32 : n69792;
  assign n69794 = pi15 ? n69793 : n32;
  assign n69795 = pi14 ? n69794 : n69697;
  assign n69796 = pi17 ? n23052 : n14788;
  assign n69797 = pi16 ? n32 : n69796;
  assign n69798 = pi15 ? n22958 : n69797;
  assign n69799 = pi17 ? n32 : n69707;
  assign n69800 = pi16 ? n32 : n69799;
  assign n69801 = pi18 ? n32 : n18331;
  assign n69802 = pi21 ? n9485 : n32;
  assign n69803 = pi20 ? n32 : n69802;
  assign n69804 = pi19 ? n69803 : n32;
  assign n69805 = pi18 ? n69804 : ~n5372;
  assign n69806 = pi17 ? n69801 : n69805;
  assign n69807 = pi16 ? n32 : n69806;
  assign n69808 = pi15 ? n69800 : n69807;
  assign n69809 = pi14 ? n69798 : n69808;
  assign n69810 = pi13 ? n69795 : n69809;
  assign n69811 = pi12 ? n69791 : n69810;
  assign n69812 = pi11 ? n69777 : n69811;
  assign n69813 = pi10 ? n69732 : n69812;
  assign n69814 = pi09 ? n17493 : n69813;
  assign n69815 = pi08 ? n69722 : n69814;
  assign n69816 = pi15 ? n16397 : n17286;
  assign n69817 = pi15 ? n26269 : n17039;
  assign n69818 = pi14 ? n69816 : n69817;
  assign n69819 = pi13 ? n69726 : n69818;
  assign n69820 = pi15 ? n68564 : n26400;
  assign n69821 = pi20 ? n342 : ~n11048;
  assign n69822 = pi19 ? n32 : n69821;
  assign n69823 = pi18 ? n32 : n69822;
  assign n69824 = pi17 ? n32 : n69823;
  assign n69825 = pi16 ? n32 : n69824;
  assign n69826 = pi15 ? n32 : n69825;
  assign n69827 = pi14 ? n69820 : n69826;
  assign n69828 = pi20 ? n1385 : n274;
  assign n69829 = pi19 ? n32 : n69828;
  assign n69830 = pi18 ? n32 : n69829;
  assign n69831 = pi17 ? n32 : n69830;
  assign n69832 = pi16 ? n32 : n69831;
  assign n69833 = pi15 ? n25904 : n69832;
  assign n69834 = pi15 ? n67449 : n26201;
  assign n69835 = pi14 ? n69833 : n69834;
  assign n69836 = pi13 ? n69827 : n69835;
  assign n69837 = pi12 ? n69819 : n69836;
  assign n69838 = pi11 ? n69724 : n69837;
  assign n69839 = pi18 ? n32 : n69738;
  assign n69840 = pi17 ? n32 : n69839;
  assign n69841 = pi16 ? n32 : n69840;
  assign n69842 = pi15 ? n53132 : n69841;
  assign n69843 = pi19 ? n32 : n7829;
  assign n69844 = pi18 ? n32 : n69843;
  assign n69845 = pi17 ? n32 : n69844;
  assign n69846 = pi16 ? n32 : n69845;
  assign n69847 = pi15 ? n69846 : n69750;
  assign n69848 = pi14 ? n69842 : n69847;
  assign n69849 = pi19 ? n322 : n55659;
  assign n69850 = pi18 ? n32 : n69849;
  assign n69851 = pi17 ? n32 : n69850;
  assign n69852 = pi16 ? n32 : n69851;
  assign n69853 = pi19 ? n1248 : n18502;
  assign n69854 = pi19 ? n349 : ~n69757;
  assign n69855 = pi18 ? n69853 : ~n69854;
  assign n69856 = pi17 ? n4111 : n69855;
  assign n69857 = pi16 ? n32 : n69856;
  assign n69858 = pi15 ? n69852 : n69857;
  assign n69859 = pi21 ? n405 : ~n2076;
  assign n69860 = pi20 ? n69859 : ~n32;
  assign n69861 = pi19 ? n208 : ~n69860;
  assign n69862 = pi18 ? n32 : ~n69861;
  assign n69863 = pi17 ? n32 : ~n69862;
  assign n69864 = pi16 ? n32 : n69863;
  assign n69865 = pi19 ? n208 : ~n8645;
  assign n69866 = pi18 ? n350 : ~n69865;
  assign n69867 = pi17 ? n32 : ~n69866;
  assign n69868 = pi16 ? n32 : n69867;
  assign n69869 = pi15 ? n69864 : n69868;
  assign n69870 = pi14 ? n69858 : n69869;
  assign n69871 = pi13 ? n69848 : n69870;
  assign n69872 = pi19 ? n42008 : n32;
  assign n69873 = pi21 ? n405 : ~n8275;
  assign n69874 = pi20 ? n69873 : n32;
  assign n69875 = pi19 ? n9007 : n69874;
  assign n69876 = pi18 ? n69872 : n69875;
  assign n69877 = pi17 ? n32 : n69876;
  assign n69878 = pi16 ? n32 : n69877;
  assign n69879 = pi19 ? n32 : n61101;
  assign n69880 = pi18 ? n32 : n69879;
  assign n69881 = pi17 ? n32 : n69880;
  assign n69882 = pi16 ? n32 : n69881;
  assign n69883 = pi15 ? n69878 : n69882;
  assign n69884 = pi19 ? n32 : ~n8645;
  assign n69885 = pi18 ? n32 : n69884;
  assign n69886 = pi17 ? n32 : n69885;
  assign n69887 = pi16 ? n32 : n69886;
  assign n69888 = pi15 ? n69887 : n16101;
  assign n69889 = pi14 ? n69883 : n69888;
  assign n69890 = pi15 ? n24237 : n55403;
  assign n69891 = pi15 ? n15080 : n37654;
  assign n69892 = pi14 ? n69890 : n69891;
  assign n69893 = pi13 ? n69889 : n69892;
  assign n69894 = pi12 ? n69871 : n69893;
  assign n69895 = pi19 ? n322 : ~n9368;
  assign n69896 = pi18 ? n32 : n69895;
  assign n69897 = pi17 ? n32 : n69896;
  assign n69898 = pi16 ? n32 : n69897;
  assign n69899 = pi19 ? n32 : n18489;
  assign n69900 = pi19 ? n17842 : n7488;
  assign n69901 = pi18 ? n69899 : n69900;
  assign n69902 = pi17 ? n23052 : n69901;
  assign n69903 = pi16 ? n32 : n69902;
  assign n69904 = pi15 ? n69898 : n69903;
  assign n69905 = pi19 ? n519 : ~n5614;
  assign n69906 = pi18 ? n32 : n69905;
  assign n69907 = pi17 ? n3164 : ~n69906;
  assign n69908 = pi16 ? n32 : n69907;
  assign n69909 = pi18 ? n32 : n11386;
  assign n69910 = pi17 ? n4128 : ~n69909;
  assign n69911 = pi16 ? n32 : n69910;
  assign n69912 = pi15 ? n69908 : n69911;
  assign n69913 = pi14 ? n69904 : n69912;
  assign n69914 = pi17 ? n4128 : ~n2736;
  assign n69915 = pi16 ? n32 : n69914;
  assign n69916 = pi19 ? n32 : n53174;
  assign n69917 = pi18 ? n32 : n69916;
  assign n69918 = pi17 ? n69917 : ~n69673;
  assign n69919 = pi16 ? n32 : n69918;
  assign n69920 = pi15 ? n69915 : n69919;
  assign n69921 = pi17 ? n69917 : ~n69678;
  assign n69922 = pi16 ? n32 : n69921;
  assign n69923 = pi19 ? n14786 : n1105;
  assign n69924 = pi18 ? n32 : n69923;
  assign n69925 = pi17 ? n3164 : ~n69924;
  assign n69926 = pi16 ? n32 : n69925;
  assign n69927 = pi15 ? n69922 : n69926;
  assign n69928 = pi14 ? n69920 : n69927;
  assign n69929 = pi13 ? n69913 : n69928;
  assign n69930 = pi20 ? n32 : ~n974;
  assign n69931 = pi19 ? n69930 : n1105;
  assign n69932 = pi18 ? n32 : n69931;
  assign n69933 = pi17 ? n3164 : ~n69932;
  assign n69934 = pi16 ? n32 : n69933;
  assign n69935 = pi15 ? n69934 : n32;
  assign n69936 = pi20 ? n246 : n175;
  assign n69937 = pi19 ? n69936 : n32;
  assign n69938 = pi18 ? n22305 : n69937;
  assign n69939 = pi17 ? n32 : n69938;
  assign n69940 = pi16 ? n32 : n69939;
  assign n69941 = pi20 ? n321 : n18624;
  assign n69942 = pi19 ? n69941 : n32;
  assign n69943 = pi18 ? n32 : n69942;
  assign n69944 = pi17 ? n2954 : n69943;
  assign n69945 = pi16 ? n32 : n69944;
  assign n69946 = pi15 ? n69940 : n69945;
  assign n69947 = pi14 ? n69935 : n69946;
  assign n69948 = pi15 ? n14790 : n21686;
  assign n69949 = pi19 ? n18478 : ~n32;
  assign n69950 = pi18 ? n4343 : ~n69949;
  assign n69951 = pi17 ? n2954 : n69950;
  assign n69952 = pi16 ? n32 : n69951;
  assign n69953 = pi18 ? n69949 : n5372;
  assign n69954 = pi17 ? n3728 : ~n69953;
  assign n69955 = pi16 ? n32 : n69954;
  assign n69956 = pi15 ? n69952 : n69955;
  assign n69957 = pi14 ? n69948 : n69956;
  assign n69958 = pi13 ? n69947 : n69957;
  assign n69959 = pi12 ? n69929 : n69958;
  assign n69960 = pi11 ? n69894 : n69959;
  assign n69961 = pi10 ? n69838 : n69960;
  assign n69962 = pi09 ? n17493 : n69961;
  assign n69963 = pi20 ? n653 : ~n243;
  assign n69964 = pi19 ? n32 : n69963;
  assign n69965 = pi18 ? n32 : n69964;
  assign n69966 = pi17 ? n32 : n69965;
  assign n69967 = pi16 ? n32 : n69966;
  assign n69968 = pi15 ? n69967 : n69750;
  assign n69969 = pi14 ? n69842 : n69968;
  assign n69970 = pi19 ? n322 : n13074;
  assign n69971 = pi18 ? n32 : n69970;
  assign n69972 = pi17 ? n32 : n69971;
  assign n69973 = pi16 ? n32 : n69972;
  assign n69974 = pi15 ? n69973 : n69857;
  assign n69975 = pi21 ? n100 : ~n2076;
  assign n69976 = pi20 ? n69975 : ~n32;
  assign n69977 = pi19 ? n208 : ~n69976;
  assign n69978 = pi18 ? n32 : ~n69977;
  assign n69979 = pi17 ? n32 : ~n69978;
  assign n69980 = pi16 ? n32 : n69979;
  assign n69981 = pi15 ? n69980 : n69868;
  assign n69982 = pi14 ? n69974 : n69981;
  assign n69983 = pi13 ? n69969 : n69982;
  assign n69984 = pi18 ? n53618 : n69875;
  assign n69985 = pi17 ? n32 : n69984;
  assign n69986 = pi16 ? n32 : n69985;
  assign n69987 = pi20 ? n27539 : n32;
  assign n69988 = pi19 ? n32 : n69987;
  assign n69989 = pi18 ? n32 : n69988;
  assign n69990 = pi17 ? n32 : n69989;
  assign n69991 = pi16 ? n32 : n69990;
  assign n69992 = pi15 ? n69986 : n69991;
  assign n69993 = pi15 ? n69887 : n16298;
  assign n69994 = pi14 ? n69992 : n69993;
  assign n69995 = pi19 ? n507 : n8064;
  assign n69996 = pi18 ? n32 : n69995;
  assign n69997 = pi17 ? n32 : n69996;
  assign n69998 = pi16 ? n32 : n69997;
  assign n69999 = pi15 ? n24237 : n69998;
  assign n70000 = pi19 ? n519 : ~n9368;
  assign n70001 = pi18 ? n32 : n70000;
  assign n70002 = pi17 ? n32 : n70001;
  assign n70003 = pi16 ? n32 : n70002;
  assign n70004 = pi19 ? n1165 : n7693;
  assign n70005 = pi18 ? n32 : n70004;
  assign n70006 = pi17 ? n32 : n70005;
  assign n70007 = pi16 ? n32 : n70006;
  assign n70008 = pi15 ? n70003 : n70007;
  assign n70009 = pi14 ? n69999 : n70008;
  assign n70010 = pi13 ? n69994 : n70009;
  assign n70011 = pi12 ? n69983 : n70010;
  assign n70012 = pi19 ? n1320 : ~n1812;
  assign n70013 = pi18 ? n32 : n70012;
  assign n70014 = pi17 ? n32 : n70013;
  assign n70015 = pi16 ? n32 : n70014;
  assign n70016 = pi15 ? n70015 : n69903;
  assign n70017 = pi17 ? n3728 : ~n69909;
  assign n70018 = pi16 ? n32 : n70017;
  assign n70019 = pi15 ? n53580 : n70018;
  assign n70020 = pi14 ? n70016 : n70019;
  assign n70021 = pi21 ? n206 : n66;
  assign n70022 = pi20 ? n32 : n70021;
  assign n70023 = pi19 ? n70022 : n2614;
  assign n70024 = pi18 ? n32 : n70023;
  assign n70025 = pi17 ? n2954 : ~n70024;
  assign n70026 = pi16 ? n32 : n70025;
  assign n70027 = pi15 ? n9954 : n70026;
  assign n70028 = pi19 ? n14589 : n2614;
  assign n70029 = pi18 ? n32 : n70028;
  assign n70030 = pi17 ? n2954 : ~n70029;
  assign n70031 = pi16 ? n32 : n70030;
  assign n70032 = pi17 ? n2954 : ~n69924;
  assign n70033 = pi16 ? n32 : n70032;
  assign n70034 = pi15 ? n70031 : n70033;
  assign n70035 = pi14 ? n70027 : n70034;
  assign n70036 = pi13 ? n70020 : n70035;
  assign n70037 = pi20 ? n32 : ~n52847;
  assign n70038 = pi19 ? n70037 : ~n32;
  assign n70039 = pi18 ? n32 : n70038;
  assign n70040 = pi17 ? n2954 : ~n70039;
  assign n70041 = pi16 ? n32 : n70040;
  assign n70042 = pi15 ? n70041 : n21543;
  assign n70043 = pi20 ? n10644 : ~n266;
  assign n70044 = pi19 ? n5694 : ~n70043;
  assign n70045 = pi18 ? n70044 : n69937;
  assign n70046 = pi17 ? n32 : n70045;
  assign n70047 = pi16 ? n32 : n70046;
  assign n70048 = pi17 ? n32 : n69943;
  assign n70049 = pi16 ? n32 : n70048;
  assign n70050 = pi15 ? n70047 : n70049;
  assign n70051 = pi14 ? n70042 : n70050;
  assign n70052 = pi17 ? n32 : n69950;
  assign n70053 = pi16 ? n32 : n70052;
  assign n70054 = pi17 ? n32 : ~n69953;
  assign n70055 = pi16 ? n32 : n70054;
  assign n70056 = pi15 ? n70053 : n70055;
  assign n70057 = pi14 ? n69948 : n70056;
  assign n70058 = pi13 ? n70051 : n70057;
  assign n70059 = pi12 ? n70036 : n70058;
  assign n70060 = pi11 ? n70011 : n70059;
  assign n70061 = pi10 ? n69838 : n70060;
  assign n70062 = pi09 ? n17493 : n70061;
  assign n70063 = pi08 ? n69962 : n70062;
  assign n70064 = pi07 ? n69815 : n70063;
  assign n70065 = pi06 ? n69553 : n70064;
  assign n70066 = pi05 ? n69122 : n70065;
  assign n70067 = pi15 ? n17278 : n16392;
  assign n70068 = pi14 ? n17443 : n70067;
  assign n70069 = pi13 ? n32 : n70068;
  assign n70070 = pi12 ? n32 : n70069;
  assign n70071 = pi15 ? n32 : n69559;
  assign n70072 = pi15 ? n68991 : n16397;
  assign n70073 = pi14 ? n70071 : n70072;
  assign n70074 = pi15 ? n17286 : n68564;
  assign n70075 = pi14 ? n26904 : n70074;
  assign n70076 = pi13 ? n70073 : n70075;
  assign n70077 = pi15 ? n68564 : n25948;
  assign n70078 = pi20 ? n321 : n7487;
  assign n70079 = pi19 ? n32 : n70078;
  assign n70080 = pi18 ? n32 : n70079;
  assign n70081 = pi17 ? n32 : n70080;
  assign n70082 = pi16 ? n32 : n70081;
  assign n70083 = pi15 ? n16804 : n70082;
  assign n70084 = pi14 ? n70077 : n70083;
  assign n70085 = pi19 ? n32 : n39001;
  assign n70086 = pi18 ? n32 : n70085;
  assign n70087 = pi17 ? n32 : n70086;
  assign n70088 = pi16 ? n32 : n70087;
  assign n70089 = pi15 ? n70088 : n53803;
  assign n70090 = pi20 ? n6621 : n1940;
  assign n70091 = pi19 ? n322 : ~n70090;
  assign n70092 = pi18 ? n32 : n70091;
  assign n70093 = pi17 ? n32 : n70092;
  assign n70094 = pi16 ? n32 : n70093;
  assign n70095 = pi15 ? n69579 : n70094;
  assign n70096 = pi14 ? n70089 : n70095;
  assign n70097 = pi13 ? n70084 : n70096;
  assign n70098 = pi12 ? n70076 : n70097;
  assign n70099 = pi11 ? n70070 : n70098;
  assign n70100 = pi19 ? n32 : ~n6619;
  assign n70101 = pi18 ? n32 : n70100;
  assign n70102 = pi17 ? n32 : n70101;
  assign n70103 = pi16 ? n32 : n70102;
  assign n70104 = pi15 ? n70103 : n69967;
  assign n70105 = pi20 ? n2385 : n243;
  assign n70106 = pi19 ? n267 : ~n70105;
  assign n70107 = pi18 ? n32 : n70106;
  assign n70108 = pi17 ? n32 : n70107;
  assign n70109 = pi16 ? n32 : n70108;
  assign n70110 = pi15 ? n70109 : n66344;
  assign n70111 = pi14 ? n70104 : n70110;
  assign n70112 = pi19 ? n322 : n59251;
  assign n70113 = pi18 ? n23440 : n70112;
  assign n70114 = pi17 ? n32 : n70113;
  assign n70115 = pi16 ? n32 : n70114;
  assign n70116 = pi19 ? n68626 : n5694;
  assign n70117 = pi19 ? n322 : ~n10158;
  assign n70118 = pi18 ? n70116 : n70117;
  assign n70119 = pi17 ? n32 : n70118;
  assign n70120 = pi16 ? n32 : n70119;
  assign n70121 = pi15 ? n70115 : n70120;
  assign n70122 = pi21 ? n100 : n9326;
  assign n70123 = pi20 ? n70122 : ~n32;
  assign n70124 = pi19 ? n267 : ~n70123;
  assign n70125 = pi18 ? n32 : n70124;
  assign n70126 = pi17 ? n32 : n70125;
  assign n70127 = pi16 ? n32 : n70126;
  assign n70128 = pi15 ? n70127 : n23981;
  assign n70129 = pi14 ? n70121 : n70128;
  assign n70130 = pi13 ? n70111 : n70129;
  assign n70131 = pi20 ? n64109 : n32;
  assign n70132 = pi19 ? n322 : n70131;
  assign n70133 = pi18 ? n32 : n70132;
  assign n70134 = pi17 ? n32 : n70133;
  assign n70135 = pi16 ? n32 : n70134;
  assign n70136 = pi19 ? n322 : ~n9646;
  assign n70137 = pi18 ? n6867 : n70136;
  assign n70138 = pi17 ? n32 : n70137;
  assign n70139 = pi16 ? n32 : n70138;
  assign n70140 = pi15 ? n70135 : n70139;
  assign n70141 = pi14 ? n70140 : n25301;
  assign n70142 = pi19 ? n1320 : ~n288;
  assign n70143 = pi18 ? n32 : n70142;
  assign n70144 = pi17 ? n32 : n70143;
  assign n70145 = pi16 ? n32 : n70144;
  assign n70146 = pi15 ? n24237 : n70145;
  assign n70147 = pi20 ? n32 : n7205;
  assign n70148 = pi19 ? n70147 : ~n6887;
  assign n70149 = pi18 ? n32 : n70148;
  assign n70150 = pi17 ? n32 : n70149;
  assign n70151 = pi16 ? n32 : n70150;
  assign n70152 = pi15 ? n35889 : n70151;
  assign n70153 = pi14 ? n70146 : n70152;
  assign n70154 = pi13 ? n70141 : n70153;
  assign n70155 = pi12 ? n70130 : n70154;
  assign n70156 = pi20 ? n32 : n58757;
  assign n70157 = pi19 ? n70156 : ~n1812;
  assign n70158 = pi18 ? n32 : n70157;
  assign n70159 = pi17 ? n32 : n70158;
  assign n70160 = pi16 ? n32 : n70159;
  assign n70161 = pi19 ? n617 : n349;
  assign n70162 = pi21 ? n34 : ~n32;
  assign n70163 = pi20 ? n70162 : ~n32;
  assign n70164 = pi19 ? n1165 : n70163;
  assign n70165 = pi18 ? n70161 : ~n70164;
  assign n70166 = pi17 ? n3569 : n70165;
  assign n70167 = pi16 ? n32 : n70166;
  assign n70168 = pi15 ? n70160 : n70167;
  assign n70169 = pi20 ? n32 : ~n18256;
  assign n70170 = pi19 ? n70169 : ~n32;
  assign n70171 = pi18 ? n618 : ~n70170;
  assign n70172 = pi17 ? n3569 : n70171;
  assign n70173 = pi16 ? n32 : n70172;
  assign n70174 = pi18 ? n31385 : ~n3200;
  assign n70175 = pi17 ? n32 : n70174;
  assign n70176 = pi16 ? n32 : n70175;
  assign n70177 = pi15 ? n70173 : n70176;
  assign n70178 = pi14 ? n70168 : n70177;
  assign n70179 = pi19 ? n5688 : n32;
  assign n70180 = pi19 ? n22558 : n236;
  assign n70181 = pi18 ? n70179 : n70180;
  assign n70182 = pi17 ? n32 : ~n70181;
  assign n70183 = pi16 ? n32 : n70182;
  assign n70184 = pi19 ? n30659 : n2614;
  assign n70185 = pi18 ? n70179 : n70184;
  assign n70186 = pi17 ? n32 : ~n70185;
  assign n70187 = pi16 ? n32 : n70186;
  assign n70188 = pi15 ? n70183 : n70187;
  assign n70189 = pi19 ? n267 : n1105;
  assign n70190 = pi18 ? n350 : ~n70189;
  assign n70191 = pi17 ? n32 : n70190;
  assign n70192 = pi16 ? n32 : n70191;
  assign n70193 = pi21 ? n32 : ~n30090;
  assign n70194 = pi20 ? n32 : n70193;
  assign n70195 = pi19 ? n70194 : ~n32;
  assign n70196 = pi18 ? n3350 : ~n70195;
  assign n70197 = pi17 ? n32 : n70196;
  assign n70198 = pi16 ? n32 : n70197;
  assign n70199 = pi15 ? n70192 : n70198;
  assign n70200 = pi14 ? n70188 : n70199;
  assign n70201 = pi13 ? n70178 : n70200;
  assign n70202 = pi18 ? n19629 : n33739;
  assign n70203 = pi17 ? n32 : n70202;
  assign n70204 = pi16 ? n32 : n70203;
  assign n70205 = pi15 ? n70204 : n24543;
  assign n70206 = pi18 ? n32478 : n22431;
  assign n70207 = pi17 ? n32 : n70206;
  assign n70208 = pi16 ? n32 : n70207;
  assign n70209 = pi18 ? n4343 : n5502;
  assign n70210 = pi17 ? n32 : n70209;
  assign n70211 = pi16 ? n32 : n70210;
  assign n70212 = pi15 ? n70208 : n70211;
  assign n70213 = pi14 ? n70205 : n70212;
  assign n70214 = pi18 ? n9170 : n32;
  assign n70215 = pi17 ? n32 : n70214;
  assign n70216 = pi16 ? n32 : n70215;
  assign n70217 = pi15 ? n70216 : n60798;
  assign n70218 = pi20 ? n52702 : ~n32;
  assign n70219 = pi19 ? n70218 : ~n32;
  assign n70220 = pi18 ? n70219 : ~n323;
  assign n70221 = pi17 ? n32 : n70220;
  assign n70222 = pi16 ? n32 : n70221;
  assign n70223 = pi15 ? n70222 : n10250;
  assign n70224 = pi14 ? n70217 : n70223;
  assign n70225 = pi13 ? n70213 : n70224;
  assign n70226 = pi12 ? n70201 : n70225;
  assign n70227 = pi11 ? n70155 : n70226;
  assign n70228 = pi10 ? n70099 : n70227;
  assign n70229 = pi09 ? n17493 : n70228;
  assign n70230 = pi19 ? n32 : n40908;
  assign n70231 = pi18 ? n32 : n70230;
  assign n70232 = pi17 ? n32 : n70231;
  assign n70233 = pi16 ? n32 : n70232;
  assign n70234 = pi15 ? n17278 : n70233;
  assign n70235 = pi14 ? n17443 : n70234;
  assign n70236 = pi13 ? n32 : n70235;
  assign n70237 = pi12 ? n32 : n70236;
  assign n70238 = pi15 ? n17188 : n69559;
  assign n70239 = pi20 ? n342 : n726;
  assign n70240 = pi19 ? n32 : n70239;
  assign n70241 = pi18 ? n32 : n70240;
  assign n70242 = pi17 ? n32 : n70241;
  assign n70243 = pi16 ? n32 : n70242;
  assign n70244 = pi15 ? n70243 : n16397;
  assign n70245 = pi14 ? n70238 : n70244;
  assign n70246 = pi13 ? n70245 : n70075;
  assign n70247 = pi20 ? n206 : ~n1940;
  assign n70248 = pi19 ? n32 : n70247;
  assign n70249 = pi18 ? n32 : n70248;
  assign n70250 = pi17 ? n32 : n70249;
  assign n70251 = pi16 ? n32 : n70250;
  assign n70252 = pi15 ? n70088 : n70251;
  assign n70253 = pi20 ? n6621 : n339;
  assign n70254 = pi19 ? n322 : ~n70253;
  assign n70255 = pi18 ? n32 : n70254;
  assign n70256 = pi17 ? n32 : n70255;
  assign n70257 = pi16 ? n32 : n70256;
  assign n70258 = pi15 ? n69579 : n70257;
  assign n70259 = pi14 ? n70252 : n70258;
  assign n70260 = pi13 ? n70084 : n70259;
  assign n70261 = pi12 ? n70246 : n70260;
  assign n70262 = pi11 ? n70237 : n70261;
  assign n70263 = pi15 ? n70103 : n69846;
  assign n70264 = pi19 ? n32 : n20768;
  assign n70265 = pi18 ? n32 : n70264;
  assign n70266 = pi17 ? n32 : n70265;
  assign n70267 = pi16 ? n32 : n70266;
  assign n70268 = pi15 ? n70109 : n70267;
  assign n70269 = pi14 ? n70263 : n70268;
  assign n70270 = pi19 ? n321 : n5694;
  assign n70271 = pi19 ? n322 : ~n10394;
  assign n70272 = pi18 ? n70270 : n70271;
  assign n70273 = pi17 ? n32 : n70272;
  assign n70274 = pi16 ? n32 : n70273;
  assign n70275 = pi15 ? n70115 : n70274;
  assign n70276 = pi14 ? n70275 : n70128;
  assign n70277 = pi13 ? n70269 : n70276;
  assign n70278 = pi18 ? n6867 : n53686;
  assign n70279 = pi17 ? n32 : n70278;
  assign n70280 = pi16 ? n32 : n70279;
  assign n70281 = pi15 ? n70135 : n70280;
  assign n70282 = pi15 ? n25301 : n16105;
  assign n70283 = pi14 ? n70281 : n70282;
  assign n70284 = pi19 ? n32 : ~n54655;
  assign n70285 = pi18 ? n32 : n70284;
  assign n70286 = pi17 ? n32 : n70285;
  assign n70287 = pi16 ? n32 : n70286;
  assign n70288 = pi15 ? n70287 : n70145;
  assign n70289 = pi19 ? n322 : ~n6693;
  assign n70290 = pi18 ? n32 : n70289;
  assign n70291 = pi17 ? n32 : n70290;
  assign n70292 = pi16 ? n32 : n70291;
  assign n70293 = pi15 ? n49496 : n70292;
  assign n70294 = pi14 ? n70288 : n70293;
  assign n70295 = pi13 ? n70283 : n70294;
  assign n70296 = pi12 ? n70277 : n70295;
  assign n70297 = pi19 ? n322 : n617;
  assign n70298 = pi18 ? n30839 : ~n70297;
  assign n70299 = pi17 ? n32 : n70298;
  assign n70300 = pi16 ? n32 : n70299;
  assign n70301 = pi15 ? n24443 : n70300;
  assign n70302 = pi18 ? n237 : ~n37093;
  assign n70303 = pi17 ? n32 : n70302;
  assign n70304 = pi16 ? n32 : n70303;
  assign n70305 = pi15 ? n70304 : n70176;
  assign n70306 = pi14 ? n70301 : n70305;
  assign n70307 = pi19 ? n15993 : ~n32;
  assign n70308 = pi19 ? n1508 : n236;
  assign n70309 = pi18 ? n70307 : ~n70308;
  assign n70310 = pi17 ? n32 : n70309;
  assign n70311 = pi16 ? n32 : n70310;
  assign n70312 = pi19 ? n4982 : n2614;
  assign n70313 = pi18 ? n35564 : ~n70312;
  assign n70314 = pi17 ? n32 : n70313;
  assign n70315 = pi16 ? n32 : n70314;
  assign n70316 = pi15 ? n70311 : n70315;
  assign n70317 = pi18 ? n350 : ~n47144;
  assign n70318 = pi17 ? n32 : n70317;
  assign n70319 = pi16 ? n32 : n70318;
  assign n70320 = pi15 ? n70192 : n70319;
  assign n70321 = pi14 ? n70316 : n70320;
  assign n70322 = pi13 ? n70306 : n70321;
  assign n70323 = pi15 ? n33742 : n24543;
  assign n70324 = pi18 ? n5749 : n22431;
  assign n70325 = pi17 ? n32 : n70324;
  assign n70326 = pi16 ? n32 : n70325;
  assign n70327 = pi18 ? n4671 : n5502;
  assign n70328 = pi17 ? n32 : n70327;
  assign n70329 = pi16 ? n32 : n70328;
  assign n70330 = pi15 ? n70326 : n70329;
  assign n70331 = pi14 ? n70323 : n70330;
  assign n70332 = pi15 ? n32 : n60798;
  assign n70333 = pi14 ? n70332 : n10490;
  assign n70334 = pi13 ? n70331 : n70333;
  assign n70335 = pi12 ? n70322 : n70334;
  assign n70336 = pi11 ? n70296 : n70335;
  assign n70337 = pi10 ? n70262 : n70336;
  assign n70338 = pi09 ? n17493 : n70337;
  assign n70339 = pi08 ? n70229 : n70338;
  assign n70340 = pi14 ? n26904 : n68557;
  assign n70341 = pi13 ? n70245 : n70340;
  assign n70342 = pi15 ? n26400 : n26479;
  assign n70343 = pi20 ? n246 : n7487;
  assign n70344 = pi19 ? n32 : n70343;
  assign n70345 = pi18 ? n32 : n70344;
  assign n70346 = pi17 ? n32 : n70345;
  assign n70347 = pi16 ? n32 : n70346;
  assign n70348 = pi15 ? n17061 : n70347;
  assign n70349 = pi14 ? n70342 : n70348;
  assign n70350 = pi20 ? n6621 : n274;
  assign n70351 = pi19 ? n32 : n70350;
  assign n70352 = pi18 ? n32 : n70351;
  assign n70353 = pi17 ? n32 : n70352;
  assign n70354 = pi16 ? n32 : n70353;
  assign n70355 = pi20 ? n11107 : ~n1940;
  assign n70356 = pi19 ? n32 : n70355;
  assign n70357 = pi18 ? n32 : n70356;
  assign n70358 = pi17 ? n32 : n70357;
  assign n70359 = pi16 ? n32 : n70358;
  assign n70360 = pi15 ? n70354 : n70359;
  assign n70361 = pi20 ? n1324 : ~n1940;
  assign n70362 = pi19 ? n322 : n70361;
  assign n70363 = pi18 ? n32 : n70362;
  assign n70364 = pi17 ? n32 : n70363;
  assign n70365 = pi16 ? n32 : n70364;
  assign n70366 = pi19 ? n322 : ~n8818;
  assign n70367 = pi18 ? n32 : n70366;
  assign n70368 = pi17 ? n32 : n70367;
  assign n70369 = pi16 ? n32 : n70368;
  assign n70370 = pi15 ? n70365 : n70369;
  assign n70371 = pi14 ? n70360 : n70370;
  assign n70372 = pi13 ? n70349 : n70371;
  assign n70373 = pi12 ? n70341 : n70372;
  assign n70374 = pi11 ? n70237 : n70373;
  assign n70375 = pi18 ? n32 : n69586;
  assign n70376 = pi17 ? n32 : n70375;
  assign n70377 = pi16 ? n32 : n70376;
  assign n70378 = pi15 ? n55261 : n70377;
  assign n70379 = pi20 ? n4279 : n243;
  assign n70380 = pi19 ? n267 : ~n70379;
  assign n70381 = pi18 ? n32 : n70380;
  assign n70382 = pi17 ? n32 : n70381;
  assign n70383 = pi16 ? n32 : n70382;
  assign n70384 = pi19 ? n32 : n59251;
  assign n70385 = pi18 ? n32 : n70384;
  assign n70386 = pi17 ? n32 : n70385;
  assign n70387 = pi16 ? n32 : n70386;
  assign n70388 = pi15 ? n70383 : n70387;
  assign n70389 = pi14 ? n70378 : n70388;
  assign n70390 = pi20 ? n40685 : n141;
  assign n70391 = pi19 ? n322 : ~n70390;
  assign n70392 = pi18 ? n23440 : n70391;
  assign n70393 = pi17 ? n32 : n70392;
  assign n70394 = pi16 ? n32 : n70393;
  assign n70395 = pi20 ? n14286 : n321;
  assign n70396 = pi19 ? n70395 : n5694;
  assign n70397 = pi19 ? n322 : ~n45479;
  assign n70398 = pi18 ? n70396 : n70397;
  assign n70399 = pi17 ? n32 : n70398;
  assign n70400 = pi16 ? n32 : n70399;
  assign n70401 = pi15 ? n70394 : n70400;
  assign n70402 = pi19 ? n916 : n58730;
  assign n70403 = pi18 ? n32 : n70402;
  assign n70404 = pi17 ? n32 : n70403;
  assign n70405 = pi16 ? n32 : n70404;
  assign n70406 = pi20 ? n40382 : n32;
  assign n70407 = pi19 ? n32 : n70406;
  assign n70408 = pi18 ? n32 : n70407;
  assign n70409 = pi17 ? n32 : n70408;
  assign n70410 = pi16 ? n32 : n70409;
  assign n70411 = pi15 ? n70405 : n70410;
  assign n70412 = pi14 ? n70401 : n70411;
  assign n70413 = pi13 ? n70389 : n70412;
  assign n70414 = pi19 ? n9169 : n176;
  assign n70415 = pi20 ? n38783 : ~n32;
  assign n70416 = pi19 ? n322 : ~n70415;
  assign n70417 = pi18 ? n70414 : n70416;
  assign n70418 = pi17 ? n32 : n70417;
  assign n70419 = pi16 ? n32 : n70418;
  assign n70420 = pi20 ? n14968 : n7487;
  assign n70421 = pi20 ? n246 : n1331;
  assign n70422 = pi19 ? n70420 : n70421;
  assign n70423 = pi21 ? n16175 : ~n206;
  assign n70424 = pi20 ? n70423 : n32;
  assign n70425 = pi19 ? n322 : n70424;
  assign n70426 = pi18 ? n70422 : n70425;
  assign n70427 = pi17 ? n32 : n70426;
  assign n70428 = pi16 ? n32 : n70427;
  assign n70429 = pi15 ? n70419 : n70428;
  assign n70430 = pi15 ? n53986 : n32;
  assign n70431 = pi14 ? n70429 : n70430;
  assign n70432 = pi21 ? n10445 : n259;
  assign n70433 = pi20 ? n70432 : ~n32;
  assign n70434 = pi19 ? n32 : ~n70433;
  assign n70435 = pi18 ? n32 : n70434;
  assign n70436 = pi17 ? n32 : n70435;
  assign n70437 = pi16 ? n32 : n70436;
  assign n70438 = pi19 ? n507 : n10662;
  assign n70439 = pi18 ? n32 : n70438;
  assign n70440 = pi17 ? n32 : n70439;
  assign n70441 = pi16 ? n32 : n70440;
  assign n70442 = pi15 ? n70437 : n70441;
  assign n70443 = pi19 ? n322 : n29950;
  assign n70444 = pi18 ? n32 : n70443;
  assign n70445 = pi17 ? n32 : n70444;
  assign n70446 = pi16 ? n32 : n70445;
  assign n70447 = pi15 ? n70446 : n37274;
  assign n70448 = pi14 ? n70442 : n70447;
  assign n70449 = pi13 ? n70431 : n70448;
  assign n70450 = pi12 ? n70413 : n70449;
  assign n70451 = pi19 ? n6298 : n349;
  assign n70452 = pi18 ? n70451 : ~n323;
  assign n70453 = pi17 ? n32 : n70452;
  assign n70454 = pi16 ? n32 : n70453;
  assign n70455 = pi15 ? n33970 : n70454;
  assign n70456 = pi19 ? n31100 : n236;
  assign n70457 = pi18 ? n53778 : ~n70456;
  assign n70458 = pi17 ? n32 : n70457;
  assign n70459 = pi16 ? n32 : n70458;
  assign n70460 = pi21 ? n7107 : ~n259;
  assign n70461 = pi20 ? n32 : n70460;
  assign n70462 = pi19 ? n70461 : n236;
  assign n70463 = pi18 ? n430 : ~n70462;
  assign n70464 = pi17 ? n32 : n70463;
  assign n70465 = pi16 ? n32 : n70464;
  assign n70466 = pi15 ? n70459 : n70465;
  assign n70467 = pi14 ? n70455 : n70466;
  assign n70468 = pi19 ? n17194 : n617;
  assign n70469 = pi18 ? n48270 : ~n70468;
  assign n70470 = pi17 ? n32 : n70469;
  assign n70471 = pi16 ? n32 : n70470;
  assign n70472 = pi19 ? n4867 : ~n32;
  assign n70473 = pi18 ? n48270 : ~n70472;
  assign n70474 = pi17 ? n32 : n70473;
  assign n70475 = pi16 ? n32 : n70474;
  assign n70476 = pi15 ? n70471 : n70475;
  assign n70477 = pi18 ? n344 : ~n63633;
  assign n70478 = pi17 ? n32 : n70477;
  assign n70479 = pi16 ? n32 : n70478;
  assign n70480 = pi15 ? n53852 : n70479;
  assign n70481 = pi14 ? n70476 : n70480;
  assign n70482 = pi13 ? n70467 : n70481;
  assign n70483 = pi18 ? n4671 : n24667;
  assign n70484 = pi17 ? n32 : n70483;
  assign n70485 = pi16 ? n32 : n70484;
  assign n70486 = pi15 ? n70485 : n55015;
  assign n70487 = pi21 ? n7478 : ~n206;
  assign n70488 = pi20 ? n32 : n70487;
  assign n70489 = pi19 ? n70488 : n32;
  assign n70490 = pi18 ? n13945 : n70489;
  assign n70491 = pi17 ? n32 : n70490;
  assign n70492 = pi16 ? n32 : n70491;
  assign n70493 = pi15 ? n70492 : n20836;
  assign n70494 = pi14 ? n70486 : n70493;
  assign n70495 = pi19 ? n13939 : n1757;
  assign n70496 = pi20 ? n206 : n9367;
  assign n70497 = pi19 ? n70496 : ~n32;
  assign n70498 = pi18 ? n70495 : ~n70497;
  assign n70499 = pi17 ? n32 : n70498;
  assign n70500 = pi16 ? n32 : n70499;
  assign n70501 = pi15 ? n32 : n70500;
  assign n70502 = pi19 ? n340 : ~n462;
  assign n70503 = pi19 ? n1868 : ~n32;
  assign n70504 = pi18 ? n70502 : ~n70503;
  assign n70505 = pi17 ? n32 : n70504;
  assign n70506 = pi16 ? n32 : n70505;
  assign n70507 = pi15 ? n10725 : n70506;
  assign n70508 = pi14 ? n70501 : n70507;
  assign n70509 = pi13 ? n70494 : n70508;
  assign n70510 = pi12 ? n70482 : n70509;
  assign n70511 = pi11 ? n70450 : n70510;
  assign n70512 = pi10 ? n70374 : n70511;
  assign n70513 = pi09 ? n17493 : n70512;
  assign n70514 = pi20 ? n342 : ~n16253;
  assign n70515 = pi19 ? n32 : n70514;
  assign n70516 = pi18 ? n32 : n70515;
  assign n70517 = pi17 ? n32 : n70516;
  assign n70518 = pi16 ? n32 : n70517;
  assign n70519 = pi15 ? n17278 : n70518;
  assign n70520 = pi14 ? n17443 : n70519;
  assign n70521 = pi13 ? n32 : n70520;
  assign n70522 = pi12 ? n32 : n70521;
  assign n70523 = pi15 ? n32 : n26515;
  assign n70524 = pi15 ? n16875 : n16397;
  assign n70525 = pi14 ? n70523 : n70524;
  assign n70526 = pi15 ? n16736 : n26400;
  assign n70527 = pi14 ? n26904 : n70526;
  assign n70528 = pi13 ? n70525 : n70527;
  assign n70529 = pi12 ? n70528 : n70372;
  assign n70530 = pi11 ? n70522 : n70529;
  assign n70531 = pi21 ? n1939 : n206;
  assign n70532 = pi20 ? n70531 : ~n141;
  assign n70533 = pi19 ? n32 : n70532;
  assign n70534 = pi18 ? n32 : n70533;
  assign n70535 = pi17 ? n32 : n70534;
  assign n70536 = pi16 ? n32 : n70535;
  assign n70537 = pi15 ? n70383 : n70536;
  assign n70538 = pi14 ? n70378 : n70537;
  assign n70539 = pi20 ? n7839 : n141;
  assign n70540 = pi19 ? n322 : ~n70539;
  assign n70541 = pi18 ? n23440 : n70540;
  assign n70542 = pi17 ? n32 : n70541;
  assign n70543 = pi16 ? n32 : n70542;
  assign n70544 = pi19 ? n322 : ~n12801;
  assign n70545 = pi18 ? n46739 : n70544;
  assign n70546 = pi17 ? n32 : n70545;
  assign n70547 = pi16 ? n32 : n70546;
  assign n70548 = pi15 ? n70543 : n70547;
  assign n70549 = pi20 ? n29452 : n32;
  assign n70550 = pi19 ? n32 : n70549;
  assign n70551 = pi18 ? n32 : n70550;
  assign n70552 = pi17 ? n32 : n70551;
  assign n70553 = pi16 ? n32 : n70552;
  assign n70554 = pi15 ? n70405 : n70553;
  assign n70555 = pi14 ? n70548 : n70554;
  assign n70556 = pi13 ? n70538 : n70555;
  assign n70557 = pi19 ? n17713 : n4670;
  assign n70558 = pi20 ? n38586 : ~n32;
  assign n70559 = pi19 ? n322 : ~n70558;
  assign n70560 = pi18 ? n70557 : n70559;
  assign n70561 = pi17 ? n32 : n70560;
  assign n70562 = pi16 ? n32 : n70561;
  assign n70563 = pi19 ? n322 : n247;
  assign n70564 = pi18 ? n32 : n70563;
  assign n70565 = pi17 ? n32 : n70564;
  assign n70566 = pi16 ? n32 : n70565;
  assign n70567 = pi15 ? n70562 : n70566;
  assign n70568 = pi15 ? n24289 : n24256;
  assign n70569 = pi14 ? n70567 : n70568;
  assign n70570 = pi19 ? n507 : n16304;
  assign n70571 = pi18 ? n32 : n70570;
  assign n70572 = pi17 ? n32 : n70571;
  assign n70573 = pi16 ? n32 : n70572;
  assign n70574 = pi15 ? n70287 : n70573;
  assign n70575 = pi14 ? n70574 : n70447;
  assign n70576 = pi13 ? n70569 : n70575;
  assign n70577 = pi12 ? n70556 : n70576;
  assign n70578 = pi19 ? n42677 : n32;
  assign n70579 = pi18 ? n32 : n70578;
  assign n70580 = pi17 ? n32 : n70579;
  assign n70581 = pi16 ? n32 : n70580;
  assign n70582 = pi19 ? n2297 : n349;
  assign n70583 = pi18 ? n70582 : ~n2291;
  assign n70584 = pi17 ? n32 : n70583;
  assign n70585 = pi16 ? n32 : n70584;
  assign n70586 = pi15 ? n70581 : n70585;
  assign n70587 = pi20 ? n32 : ~n7839;
  assign n70588 = pi19 ? n70587 : n236;
  assign n70589 = pi18 ? n532 : ~n70588;
  assign n70590 = pi17 ? n32 : n70589;
  assign n70591 = pi16 ? n32 : n70590;
  assign n70592 = pi18 ? n532 : ~n1465;
  assign n70593 = pi17 ? n32 : n70592;
  assign n70594 = pi16 ? n32 : n70593;
  assign n70595 = pi15 ? n70591 : n70594;
  assign n70596 = pi14 ? n70586 : n70595;
  assign n70597 = pi20 ? n32 : ~n10889;
  assign n70598 = pi19 ? n70597 : n617;
  assign n70599 = pi18 ? n48270 : ~n70598;
  assign n70600 = pi17 ? n32 : n70599;
  assign n70601 = pi16 ? n32 : n70600;
  assign n70602 = pi18 ? n48270 : ~n7278;
  assign n70603 = pi17 ? n32 : n70602;
  assign n70604 = pi16 ? n32 : n70603;
  assign n70605 = pi15 ? n70601 : n70604;
  assign n70606 = pi18 ? n2424 : ~n63633;
  assign n70607 = pi17 ? n32 : n70606;
  assign n70608 = pi16 ? n32 : n70607;
  assign n70609 = pi15 ? n10721 : n70608;
  assign n70610 = pi14 ? n70605 : n70609;
  assign n70611 = pi13 ? n70596 : n70610;
  assign n70612 = pi20 ? n32 : ~n44237;
  assign n70613 = pi19 ? n70612 : n32;
  assign n70614 = pi18 ? n32 : n70613;
  assign n70615 = pi17 ? n32 : n70614;
  assign n70616 = pi16 ? n32 : n70615;
  assign n70617 = pi15 ? n54196 : n70616;
  assign n70618 = pi15 ? n21801 : n20836;
  assign n70619 = pi14 ? n70617 : n70618;
  assign n70620 = pi18 ? n34485 : ~n70497;
  assign n70621 = pi17 ? n32 : n70620;
  assign n70622 = pi16 ? n32 : n70621;
  assign n70623 = pi15 ? n32 : n70622;
  assign n70624 = pi19 ? n14781 : n53946;
  assign n70625 = pi18 ? n70624 : ~n70503;
  assign n70626 = pi17 ? n32 : n70625;
  assign n70627 = pi16 ? n32 : n70626;
  assign n70628 = pi15 ? n10963 : n70627;
  assign n70629 = pi14 ? n70623 : n70628;
  assign n70630 = pi13 ? n70619 : n70629;
  assign n70631 = pi12 ? n70611 : n70630;
  assign n70632 = pi11 ? n70577 : n70631;
  assign n70633 = pi10 ? n70530 : n70632;
  assign n70634 = pi09 ? n17493 : n70633;
  assign n70635 = pi08 ? n70513 : n70634;
  assign n70636 = pi07 ? n70339 : n70635;
  assign n70637 = pi20 ? n342 : n9000;
  assign n70638 = pi19 ? n32 : n70637;
  assign n70639 = pi18 ? n32 : n70638;
  assign n70640 = pi17 ? n32 : n70639;
  assign n70641 = pi16 ? n32 : n70640;
  assign n70642 = pi15 ? n70641 : n70518;
  assign n70643 = pi14 ? n17443 : n70642;
  assign n70644 = pi13 ? n32 : n70643;
  assign n70645 = pi12 ? n32 : n70644;
  assign n70646 = pi15 ? n17465 : n26515;
  assign n70647 = pi18 ? n32 : n35345;
  assign n70648 = pi17 ? n32 : n70647;
  assign n70649 = pi16 ? n32 : n70648;
  assign n70650 = pi15 ? n70649 : n16397;
  assign n70651 = pi14 ? n70646 : n70650;
  assign n70652 = pi19 ? n32 : n6281;
  assign n70653 = pi18 ? n32 : n70652;
  assign n70654 = pi17 ? n32 : n70653;
  assign n70655 = pi16 ? n32 : n70654;
  assign n70656 = pi15 ? n16452 : n70655;
  assign n70657 = pi19 ? n32 : ~n8202;
  assign n70658 = pi18 ? n32 : n70657;
  assign n70659 = pi17 ? n32 : n70658;
  assign n70660 = pi16 ? n32 : n70659;
  assign n70661 = pi15 ? n70660 : n26400;
  assign n70662 = pi14 ? n70656 : n70661;
  assign n70663 = pi13 ? n70651 : n70662;
  assign n70664 = pi20 ? n175 : n6229;
  assign n70665 = pi19 ? n32 : n70664;
  assign n70666 = pi18 ? n32 : n70665;
  assign n70667 = pi17 ? n32 : n70666;
  assign n70668 = pi16 ? n32 : n70667;
  assign n70669 = pi15 ? n70668 : n16352;
  assign n70670 = pi19 ? n32 : n23301;
  assign n70671 = pi18 ? n32 : n70670;
  assign n70672 = pi17 ? n32 : n70671;
  assign n70673 = pi16 ? n32 : n70672;
  assign n70674 = pi15 ? n70673 : n25984;
  assign n70675 = pi14 ? n70669 : n70674;
  assign n70676 = pi19 ? n32 : ~n8230;
  assign n70677 = pi18 ? n32 : n70676;
  assign n70678 = pi17 ? n32 : n70677;
  assign n70679 = pi16 ? n32 : n70678;
  assign n70680 = pi19 ? n32 : n70361;
  assign n70681 = pi18 ? n32 : n70680;
  assign n70682 = pi17 ? n32 : n70681;
  assign n70683 = pi16 ? n32 : n70682;
  assign n70684 = pi15 ? n70679 : n70683;
  assign n70685 = pi15 ? n38071 : n51565;
  assign n70686 = pi14 ? n70684 : n70685;
  assign n70687 = pi13 ? n70675 : n70686;
  assign n70688 = pi12 ? n70663 : n70687;
  assign n70689 = pi11 ? n70645 : n70688;
  assign n70690 = pi19 ? n322 : n31395;
  assign n70691 = pi18 ? n32 : n70690;
  assign n70692 = pi17 ? n32 : n70691;
  assign n70693 = pi16 ? n32 : n70692;
  assign n70694 = pi15 ? n53814 : n70693;
  assign n70695 = pi15 ? n24504 : n70536;
  assign n70696 = pi14 ? n70694 : n70695;
  assign n70697 = pi21 ? n405 : ~n14158;
  assign n70698 = pi20 ? n70697 : ~n32;
  assign n70699 = pi19 ? n21349 : ~n70698;
  assign n70700 = pi18 ? n32 : n70699;
  assign n70701 = pi17 ? n32 : n70700;
  assign n70702 = pi16 ? n32 : n70701;
  assign n70703 = pi15 ? n70702 : n25846;
  assign n70704 = pi19 ? n9007 : n50732;
  assign n70705 = pi18 ? n16389 : n70704;
  assign n70706 = pi17 ? n32 : n70705;
  assign n70707 = pi16 ? n32 : n70706;
  assign n70708 = pi19 ? n5371 : n70558;
  assign n70709 = pi18 ? n15844 : ~n70708;
  assign n70710 = pi17 ? n32 : n70709;
  assign n70711 = pi16 ? n32 : n70710;
  assign n70712 = pi15 ? n70707 : n70711;
  assign n70713 = pi14 ? n70703 : n70712;
  assign n70714 = pi13 ? n70696 : n70713;
  assign n70715 = pi20 ? n70531 : ~n32;
  assign n70716 = pi19 ? n208 : ~n70715;
  assign n70717 = pi18 ? n6399 : n70716;
  assign n70718 = pi17 ? n32 : n70717;
  assign n70719 = pi16 ? n32 : n70718;
  assign n70720 = pi15 ? n70719 : n54016;
  assign n70721 = pi15 ? n32 : n24247;
  assign n70722 = pi14 ? n70720 : n70721;
  assign n70723 = pi15 ? n39247 : n36109;
  assign n70724 = pi19 ? n1476 : ~n1941;
  assign n70725 = pi18 ? n32 : n70724;
  assign n70726 = pi17 ? n32 : n70725;
  assign n70727 = pi16 ? n32 : n70726;
  assign n70728 = pi15 ? n25466 : n70727;
  assign n70729 = pi14 ? n70723 : n70728;
  assign n70730 = pi13 ? n70722 : n70729;
  assign n70731 = pi12 ? n70714 : n70730;
  assign n70732 = pi19 ? n654 : ~n32;
  assign n70733 = pi18 ? n1712 : ~n70732;
  assign n70734 = pi17 ? n32 : n70733;
  assign n70735 = pi16 ? n32 : n70734;
  assign n70736 = pi19 ? n9220 : ~n32;
  assign n70737 = pi20 ? n32 : ~n7377;
  assign n70738 = pi19 ? n70737 : ~n32;
  assign n70739 = pi18 ? n70736 : ~n70738;
  assign n70740 = pi17 ? n32 : n70739;
  assign n70741 = pi16 ? n32 : n70740;
  assign n70742 = pi15 ? n70735 : n70741;
  assign n70743 = pi21 ? n174 : n124;
  assign n70744 = pi20 ? n32 : n70743;
  assign n70745 = pi19 ? n70744 : n236;
  assign n70746 = pi18 ? n1465 : ~n70745;
  assign n70747 = pi17 ? n32 : n70746;
  assign n70748 = pi16 ? n32 : n70747;
  assign n70749 = pi19 ? n6355 : n617;
  assign n70750 = pi18 ? n69213 : ~n70749;
  assign n70751 = pi17 ? n32 : n70750;
  assign n70752 = pi16 ? n32 : n70751;
  assign n70753 = pi15 ? n70748 : n70752;
  assign n70754 = pi14 ? n70742 : n70753;
  assign n70755 = pi21 ? n174 : n27422;
  assign n70756 = pi20 ? n321 : ~n70755;
  assign n70757 = pi19 ? n70756 : ~n32;
  assign n70758 = pi18 ? n697 : ~n70757;
  assign n70759 = pi17 ? n32 : n70758;
  assign n70760 = pi16 ? n32 : n70759;
  assign n70761 = pi20 ? n321 : n7861;
  assign n70762 = pi19 ? n70761 : ~n32;
  assign n70763 = pi18 ? n697 : ~n70762;
  assign n70764 = pi17 ? n32 : n70763;
  assign n70765 = pi16 ? n32 : n70764;
  assign n70766 = pi15 ? n70760 : n70765;
  assign n70767 = pi20 ? n321 : ~n16309;
  assign n70768 = pi19 ? n70767 : ~n32;
  assign n70769 = pi18 ? n8086 : ~n70768;
  assign n70770 = pi17 ? n32 : n70769;
  assign n70771 = pi16 ? n32 : n70770;
  assign n70772 = pi18 ? n20020 : n35411;
  assign n70773 = pi17 ? n32 : n70772;
  assign n70774 = pi16 ? n32 : n70773;
  assign n70775 = pi15 ? n70771 : n70774;
  assign n70776 = pi14 ? n70766 : n70775;
  assign n70777 = pi13 ? n70754 : n70776;
  assign n70778 = pi15 ? n14798 : n21389;
  assign n70779 = pi18 ? n20172 : n2278;
  assign n70780 = pi17 ? n32 : n70779;
  assign n70781 = pi16 ? n32 : n70780;
  assign n70782 = pi18 ? n8106 : n5158;
  assign n70783 = pi17 ? n32 : n70782;
  assign n70784 = pi16 ? n32 : n70783;
  assign n70785 = pi15 ? n70781 : n70784;
  assign n70786 = pi14 ? n70778 : n70785;
  assign n70787 = pi18 ? n1326 : ~n54044;
  assign n70788 = pi17 ? n32 : n70787;
  assign n70789 = pi16 ? n32 : n70788;
  assign n70790 = pi15 ? n33290 : n70789;
  assign n70791 = pi19 ? n857 : ~n247;
  assign n70792 = pi18 ? n70791 : ~n323;
  assign n70793 = pi17 ? n32 : n70792;
  assign n70794 = pi16 ? n32 : n70793;
  assign n70795 = pi15 ? n70794 : n32219;
  assign n70796 = pi14 ? n70790 : n70795;
  assign n70797 = pi13 ? n70786 : n70796;
  assign n70798 = pi12 ? n70777 : n70797;
  assign n70799 = pi11 ? n70731 : n70798;
  assign n70800 = pi10 ? n70689 : n70799;
  assign n70801 = pi09 ? n17493 : n70800;
  assign n70802 = pi15 ? n68991 : n70518;
  assign n70803 = pi14 ? n17443 : n70802;
  assign n70804 = pi13 ? n32 : n70803;
  assign n70805 = pi12 ? n32 : n70804;
  assign n70806 = pi11 ? n70805 : n70688;
  assign n70807 = pi20 ? n7939 : ~n141;
  assign n70808 = pi19 ? n32 : n70807;
  assign n70809 = pi18 ? n32 : n70808;
  assign n70810 = pi17 ? n32 : n70809;
  assign n70811 = pi16 ? n32 : n70810;
  assign n70812 = pi15 ? n24504 : n70811;
  assign n70813 = pi14 ? n70694 : n70812;
  assign n70814 = pi21 ? n1939 : ~n14158;
  assign n70815 = pi20 ? n70814 : ~n32;
  assign n70816 = pi19 ? n21349 : ~n70815;
  assign n70817 = pi18 ? n32 : n70816;
  assign n70818 = pi17 ? n32 : n70817;
  assign n70819 = pi16 ? n32 : n70818;
  assign n70820 = pi15 ? n70819 : n25846;
  assign n70821 = pi21 ? n1939 : n2076;
  assign n70822 = pi20 ? n70821 : n32;
  assign n70823 = pi19 ? n9007 : n70822;
  assign n70824 = pi18 ? n16389 : n70823;
  assign n70825 = pi17 ? n32 : n70824;
  assign n70826 = pi16 ? n32 : n70825;
  assign n70827 = pi15 ? n70826 : n70711;
  assign n70828 = pi14 ? n70820 : n70827;
  assign n70829 = pi13 ? n70813 : n70828;
  assign n70830 = pi18 ? n14970 : n70716;
  assign n70831 = pi17 ? n32 : n70830;
  assign n70832 = pi16 ? n32 : n70831;
  assign n70833 = pi15 ? n70832 : n54016;
  assign n70834 = pi14 ? n70833 : n70721;
  assign n70835 = pi19 ? n244 : ~n236;
  assign n70836 = pi18 ? n32 : n70835;
  assign n70837 = pi17 ? n32 : n70836;
  assign n70838 = pi16 ? n32 : n70837;
  assign n70839 = pi15 ? n70727 : n70838;
  assign n70840 = pi14 ? n70723 : n70839;
  assign n70841 = pi13 ? n70834 : n70840;
  assign n70842 = pi12 ? n70829 : n70841;
  assign n70843 = pi19 ? n4721 : ~n53;
  assign n70844 = pi18 ? n4428 : ~n70843;
  assign n70845 = pi17 ? n32 : n70844;
  assign n70846 = pi16 ? n32 : n70845;
  assign n70847 = pi15 ? n70735 : n70846;
  assign n70848 = pi19 ? n44258 : n2614;
  assign n70849 = pi18 ? n1465 : ~n70848;
  assign n70850 = pi17 ? n32 : n70849;
  assign n70851 = pi16 ? n32 : n70850;
  assign n70852 = pi22 ? n65 : ~n84;
  assign n70853 = pi21 ? n206 : ~n70852;
  assign n70854 = pi20 ? n32 : ~n70853;
  assign n70855 = pi19 ? n70854 : ~n32;
  assign n70856 = pi18 ? n702 : ~n70855;
  assign n70857 = pi17 ? n32 : n70856;
  assign n70858 = pi16 ? n32 : n70857;
  assign n70859 = pi15 ? n70851 : n70858;
  assign n70860 = pi14 ? n70847 : n70859;
  assign n70861 = pi21 ? n174 : ~n7478;
  assign n70862 = pi20 ? n321 : ~n70861;
  assign n70863 = pi19 ? n70862 : ~n32;
  assign n70864 = pi18 ? n697 : ~n70863;
  assign n70865 = pi17 ? n32 : n70864;
  assign n70866 = pi16 ? n32 : n70865;
  assign n70867 = pi21 ? n206 : ~n14792;
  assign n70868 = pi20 ? n321 : n70867;
  assign n70869 = pi19 ? n70868 : ~n32;
  assign n70870 = pi18 ? n697 : ~n70869;
  assign n70871 = pi17 ? n32 : n70870;
  assign n70872 = pi16 ? n32 : n70871;
  assign n70873 = pi15 ? n70866 : n70872;
  assign n70874 = pi18 ? n8086 : ~n22486;
  assign n70875 = pi17 ? n32 : n70874;
  assign n70876 = pi16 ? n32 : n70875;
  assign n70877 = pi15 ? n70876 : n35414;
  assign n70878 = pi14 ? n70873 : n70877;
  assign n70879 = pi13 ? n70860 : n70878;
  assign n70880 = pi15 ? n14790 : n21389;
  assign n70881 = pi15 ? n29701 : n32;
  assign n70882 = pi14 ? n70880 : n70881;
  assign n70883 = pi18 ? n17118 : n22779;
  assign n70884 = pi17 ? n32 : n70883;
  assign n70885 = pi16 ? n32 : n70884;
  assign n70886 = pi15 ? n70885 : n11423;
  assign n70887 = pi18 ? n36557 : ~n605;
  assign n70888 = pi17 ? n32 : n70887;
  assign n70889 = pi16 ? n32 : n70888;
  assign n70890 = pi15 ? n70889 : n12098;
  assign n70891 = pi14 ? n70886 : n70890;
  assign n70892 = pi13 ? n70882 : n70891;
  assign n70893 = pi12 ? n70879 : n70892;
  assign n70894 = pi11 ? n70842 : n70893;
  assign n70895 = pi10 ? n70806 : n70894;
  assign n70896 = pi09 ? n17493 : n70895;
  assign n70897 = pi08 ? n70801 : n70896;
  assign n70898 = pi15 ? n69144 : n16736;
  assign n70899 = pi14 ? n26515 : n70898;
  assign n70900 = pi20 ? n1324 : n1817;
  assign n70901 = pi19 ? n32 : n70900;
  assign n70902 = pi18 ? n32 : n70901;
  assign n70903 = pi17 ? n32 : n70902;
  assign n70904 = pi16 ? n32 : n70903;
  assign n70905 = pi15 ? n70655 : n70904;
  assign n70906 = pi19 ? n32 : ~n9846;
  assign n70907 = pi18 ? n32 : n70906;
  assign n70908 = pi17 ? n32 : n70907;
  assign n70909 = pi16 ? n32 : n70908;
  assign n70910 = pi15 ? n70909 : n26400;
  assign n70911 = pi14 ? n70905 : n70910;
  assign n70912 = pi13 ? n70899 : n70911;
  assign n70913 = pi20 ? n1324 : ~n11048;
  assign n70914 = pi19 ? n32 : n70913;
  assign n70915 = pi18 ? n32 : n70914;
  assign n70916 = pi17 ? n32 : n70915;
  assign n70917 = pi16 ? n32 : n70916;
  assign n70918 = pi15 ? n70917 : n25984;
  assign n70919 = pi14 ? n70669 : n70918;
  assign n70920 = pi19 ? n32 : ~n7823;
  assign n70921 = pi18 ? n32 : n70920;
  assign n70922 = pi17 ? n32 : n70921;
  assign n70923 = pi16 ? n32 : n70922;
  assign n70924 = pi15 ? n70923 : n70683;
  assign n70925 = pi14 ? n70924 : n70685;
  assign n70926 = pi13 ? n70919 : n70925;
  assign n70927 = pi12 ? n70912 : n70926;
  assign n70928 = pi11 ? n70805 : n70927;
  assign n70929 = pi20 ? n18624 : ~n339;
  assign n70930 = pi19 ? n322 : n70929;
  assign n70931 = pi18 ? n32 : n70930;
  assign n70932 = pi17 ? n32 : n70931;
  assign n70933 = pi16 ? n32 : n70932;
  assign n70934 = pi19 ? n322 : n23227;
  assign n70935 = pi18 ? n32 : n70934;
  assign n70936 = pi17 ? n32 : n70935;
  assign n70937 = pi16 ? n32 : n70936;
  assign n70938 = pi15 ? n70933 : n70937;
  assign n70939 = pi20 ? n18256 : n32;
  assign n70940 = pi19 ? n32 : n70939;
  assign n70941 = pi18 ? n32 : n70940;
  assign n70942 = pi17 ? n32 : n70941;
  assign n70943 = pi16 ? n32 : n70942;
  assign n70944 = pi19 ? n358 : ~n2297;
  assign n70945 = pi18 ? n32 : n70944;
  assign n70946 = pi17 ? n32 : n70945;
  assign n70947 = pi16 ? n32 : n70946;
  assign n70948 = pi15 ? n70943 : n70947;
  assign n70949 = pi14 ? n70938 : n70948;
  assign n70950 = pi19 ? n21349 : ~n11561;
  assign n70951 = pi18 ? n32 : n70950;
  assign n70952 = pi17 ? n32 : n70951;
  assign n70953 = pi16 ? n32 : n70952;
  assign n70954 = pi15 ? n70953 : n54174;
  assign n70955 = pi20 ? n915 : ~n207;
  assign n70956 = pi20 ? n35409 : n32;
  assign n70957 = pi19 ? n70955 : n70956;
  assign n70958 = pi18 ? n16834 : n70957;
  assign n70959 = pi17 ? n32 : n70958;
  assign n70960 = pi16 ? n32 : n70959;
  assign n70961 = pi19 ? n594 : ~n54219;
  assign n70962 = pi21 ? n1939 : n10445;
  assign n70963 = pi20 ? n70962 : ~n32;
  assign n70964 = pi19 ? n5371 : n70963;
  assign n70965 = pi18 ? n70961 : ~n70964;
  assign n70966 = pi17 ? n32 : n70965;
  assign n70967 = pi16 ? n32 : n70966;
  assign n70968 = pi15 ? n70960 : n70967;
  assign n70969 = pi14 ? n70954 : n70968;
  assign n70970 = pi13 ? n70949 : n70969;
  assign n70971 = pi20 ? n17712 : n342;
  assign n70972 = pi19 ? n32 : n70971;
  assign n70973 = pi19 ? n14260 : ~n10890;
  assign n70974 = pi18 ? n70972 : n70973;
  assign n70975 = pi17 ? n32 : n70974;
  assign n70976 = pi16 ? n32 : n70975;
  assign n70977 = pi15 ? n70976 : n36109;
  assign n70978 = pi15 ? n23484 : n24511;
  assign n70979 = pi14 ? n70977 : n70978;
  assign n70980 = pi19 ? n11972 : ~n1941;
  assign n70981 = pi18 ? n32 : n70980;
  assign n70982 = pi17 ? n32 : n70981;
  assign n70983 = pi16 ? n32 : n70982;
  assign n70984 = pi19 ? n1150 : ~n236;
  assign n70985 = pi18 ? n32 : n70984;
  assign n70986 = pi17 ? n32 : n70985;
  assign n70987 = pi16 ? n32 : n70986;
  assign n70988 = pi15 ? n70983 : n70987;
  assign n70989 = pi14 ? n70723 : n70988;
  assign n70990 = pi13 ? n70979 : n70989;
  assign n70991 = pi12 ? n70970 : n70990;
  assign n70992 = pi18 ? n6235 : ~n70732;
  assign n70993 = pi17 ? n32 : n70992;
  assign n70994 = pi16 ? n32 : n70993;
  assign n70995 = pi19 ? n4721 : n10447;
  assign n70996 = pi18 ? n6235 : ~n70995;
  assign n70997 = pi17 ? n32 : n70996;
  assign n70998 = pi16 ? n32 : n70997;
  assign n70999 = pi15 ? n70994 : n70998;
  assign n71000 = pi19 ? n221 : n2614;
  assign n71001 = pi18 ? n1750 : ~n71000;
  assign n71002 = pi17 ? n32 : n71001;
  assign n71003 = pi16 ? n32 : n71002;
  assign n71004 = pi20 ? n32 : ~n20507;
  assign n71005 = pi19 ? n71004 : ~n32;
  assign n71006 = pi18 ? n1750 : ~n71005;
  assign n71007 = pi17 ? n32 : n71006;
  assign n71008 = pi16 ? n32 : n71007;
  assign n71009 = pi15 ? n71003 : n71008;
  assign n71010 = pi14 ? n70999 : n71009;
  assign n71011 = pi20 ? n321 : ~n13084;
  assign n71012 = pi19 ? n71011 : ~n32;
  assign n71013 = pi18 ? n697 : ~n71012;
  assign n71014 = pi17 ? n32 : n71013;
  assign n71015 = pi16 ? n32 : n71014;
  assign n71016 = pi21 ? n405 : n10445;
  assign n71017 = pi20 ? n321 : n71016;
  assign n71018 = pi19 ? n71017 : ~n32;
  assign n71019 = pi18 ? n697 : ~n71018;
  assign n71020 = pi17 ? n32 : n71019;
  assign n71021 = pi16 ? n32 : n71020;
  assign n71022 = pi15 ? n71015 : n71021;
  assign n71023 = pi18 ? n702 : ~n47074;
  assign n71024 = pi17 ? n32 : n71023;
  assign n71025 = pi16 ? n32 : n71024;
  assign n71026 = pi18 ? n20172 : n23091;
  assign n71027 = pi17 ? n32 : n71026;
  assign n71028 = pi16 ? n32 : n71027;
  assign n71029 = pi15 ? n71025 : n71028;
  assign n71030 = pi14 ? n71022 : n71029;
  assign n71031 = pi13 ? n71010 : n71030;
  assign n71032 = pi15 ? n14790 : n21464;
  assign n71033 = pi14 ? n71032 : n33991;
  assign n71034 = pi20 ? n220 : ~n2385;
  assign n71035 = pi19 ? n32 : n71034;
  assign n71036 = pi20 ? n314 : n1839;
  assign n71037 = pi19 ? n71036 : ~n32;
  assign n71038 = pi18 ? n71035 : ~n71037;
  assign n71039 = pi17 ? n32 : n71038;
  assign n71040 = pi16 ? n32 : n71039;
  assign n71041 = pi18 ? n962 : ~n323;
  assign n71042 = pi17 ? n32 : n71041;
  assign n71043 = pi16 ? n32 : n71042;
  assign n71044 = pi15 ? n71040 : n71043;
  assign n71045 = pi18 ? n496 : ~n605;
  assign n71046 = pi17 ? n32 : n71045;
  assign n71047 = pi16 ? n32 : n71046;
  assign n71048 = pi18 ? n8819 : ~n418;
  assign n71049 = pi17 ? n32 : n71048;
  assign n71050 = pi16 ? n32 : n71049;
  assign n71051 = pi15 ? n71047 : n71050;
  assign n71052 = pi14 ? n71044 : n71051;
  assign n71053 = pi13 ? n71033 : n71052;
  assign n71054 = pi12 ? n71031 : n71053;
  assign n71055 = pi11 ? n70991 : n71054;
  assign n71056 = pi10 ? n70928 : n71055;
  assign n71057 = pi09 ? n17493 : n71056;
  assign n71058 = pi15 ? n38071 : n67775;
  assign n71059 = pi14 ? n70924 : n71058;
  assign n71060 = pi13 ? n70919 : n71059;
  assign n71061 = pi12 ? n70912 : n71060;
  assign n71062 = pi11 ? n70805 : n71061;
  assign n71063 = pi20 ? n25513 : ~n243;
  assign n71064 = pi19 ? n322 : n71063;
  assign n71065 = pi18 ? n32 : n71064;
  assign n71066 = pi17 ? n32 : n71065;
  assign n71067 = pi16 ? n32 : n71066;
  assign n71068 = pi20 ? n19604 : ~n243;
  assign n71069 = pi19 ? n322 : n71068;
  assign n71070 = pi18 ? n32 : n71069;
  assign n71071 = pi17 ? n32 : n71070;
  assign n71072 = pi16 ? n32 : n71071;
  assign n71073 = pi15 ? n71067 : n71072;
  assign n71074 = pi20 ? n16008 : ~n141;
  assign n71075 = pi19 ? n32 : n71074;
  assign n71076 = pi18 ? n32 : n71075;
  assign n71077 = pi17 ? n32 : n71076;
  assign n71078 = pi16 ? n32 : n71077;
  assign n71079 = pi18 ? n16962 : n70944;
  assign n71080 = pi17 ? n32 : n71079;
  assign n71081 = pi16 ? n32 : n71080;
  assign n71082 = pi15 ? n71078 : n71081;
  assign n71083 = pi14 ? n71073 : n71082;
  assign n71084 = pi19 ? n21349 : ~n11108;
  assign n71085 = pi18 ? n32 : n71084;
  assign n71086 = pi17 ? n32 : n71085;
  assign n71087 = pi16 ? n32 : n71086;
  assign n71088 = pi19 ? n322 : n70822;
  assign n71089 = pi18 ? n32 : n71088;
  assign n71090 = pi17 ? n32 : n71089;
  assign n71091 = pi16 ? n32 : n71090;
  assign n71092 = pi15 ? n71087 : n71091;
  assign n71093 = pi21 ? n51 : n14158;
  assign n71094 = pi20 ? n71093 : n32;
  assign n71095 = pi19 ? n4391 : ~n71094;
  assign n71096 = pi18 ? n16389 : ~n71095;
  assign n71097 = pi17 ? n32 : n71096;
  assign n71098 = pi16 ? n32 : n71097;
  assign n71099 = pi20 ? n1939 : ~n32;
  assign n71100 = pi19 ? n5371 : n71099;
  assign n71101 = pi18 ? n15844 : ~n71100;
  assign n71102 = pi17 ? n32 : n71101;
  assign n71103 = pi16 ? n32 : n71102;
  assign n71104 = pi15 ? n71098 : n71103;
  assign n71105 = pi14 ? n71092 : n71104;
  assign n71106 = pi13 ? n71083 : n71105;
  assign n71107 = pi19 ? n208 : ~n39789;
  assign n71108 = pi18 ? n46659 : n71107;
  assign n71109 = pi17 ? n32 : n71108;
  assign n71110 = pi16 ? n32 : n71109;
  assign n71111 = pi15 ? n71110 : n36109;
  assign n71112 = pi19 ? n32 : ~n6652;
  assign n71113 = pi18 ? n32 : n71112;
  assign n71114 = pi17 ? n32 : n71113;
  assign n71115 = pi16 ? n32 : n71114;
  assign n71116 = pi15 ? n71115 : n24511;
  assign n71117 = pi14 ? n71111 : n71116;
  assign n71118 = pi19 ? n322 : n7693;
  assign n71119 = pi18 ? n32 : n71118;
  assign n71120 = pi17 ? n32 : n71119;
  assign n71121 = pi16 ? n32 : n71120;
  assign n71122 = pi15 ? n71121 : n39808;
  assign n71123 = pi15 ? n14575 : n70987;
  assign n71124 = pi14 ? n71122 : n71123;
  assign n71125 = pi13 ? n71117 : n71124;
  assign n71126 = pi12 ? n71106 : n71125;
  assign n71127 = pi19 ? n17859 : ~n53;
  assign n71128 = pi18 ? n697 : ~n71127;
  assign n71129 = pi17 ? n32 : n71128;
  assign n71130 = pi16 ? n32 : n71129;
  assign n71131 = pi19 ? n4721 : n1941;
  assign n71132 = pi18 ? n697 : ~n71131;
  assign n71133 = pi17 ? n32 : n71132;
  assign n71134 = pi16 ? n32 : n71133;
  assign n71135 = pi15 ? n71130 : n71134;
  assign n71136 = pi18 ? n697 : ~n8975;
  assign n71137 = pi17 ? n32 : n71136;
  assign n71138 = pi16 ? n32 : n71137;
  assign n71139 = pi18 ? n697 : ~n71005;
  assign n71140 = pi17 ? n32 : n71139;
  assign n71141 = pi16 ? n32 : n71140;
  assign n71142 = pi15 ? n71138 : n71141;
  assign n71143 = pi14 ? n71135 : n71142;
  assign n71144 = pi20 ? n321 : ~n10644;
  assign n71145 = pi19 ? n71144 : ~n32;
  assign n71146 = pi18 ? n697 : ~n71145;
  assign n71147 = pi17 ? n32 : n71146;
  assign n71148 = pi16 ? n32 : n71147;
  assign n71149 = pi21 ? n405 : n6898;
  assign n71150 = pi20 ? n321 : n71149;
  assign n71151 = pi19 ? n71150 : ~n32;
  assign n71152 = pi18 ? n697 : ~n71151;
  assign n71153 = pi17 ? n32 : n71152;
  assign n71154 = pi16 ? n32 : n71153;
  assign n71155 = pi15 ? n71148 : n71154;
  assign n71156 = pi20 ? n321 : ~n18158;
  assign n71157 = pi19 ? n71156 : ~n32;
  assign n71158 = pi18 ? n496 : ~n71157;
  assign n71159 = pi17 ? n32 : n71158;
  assign n71160 = pi16 ? n32 : n71159;
  assign n71161 = pi15 ? n71160 : n22437;
  assign n71162 = pi14 ? n71155 : n71161;
  assign n71163 = pi13 ? n71143 : n71162;
  assign n71164 = pi14 ? n23534 : n62112;
  assign n71165 = pi20 ? n1324 : ~n2385;
  assign n71166 = pi19 ? n32 : n71165;
  assign n71167 = pi19 ? n8212 : ~n32;
  assign n71168 = pi18 ? n71166 : ~n71167;
  assign n71169 = pi17 ? n32 : n71168;
  assign n71170 = pi16 ? n32 : n71169;
  assign n71171 = pi15 ? n71170 : n11856;
  assign n71172 = pi15 ? n11860 : n20883;
  assign n71173 = pi14 ? n71171 : n71172;
  assign n71174 = pi13 ? n71164 : n71173;
  assign n71175 = pi12 ? n71163 : n71174;
  assign n71176 = pi11 ? n71126 : n71175;
  assign n71177 = pi10 ? n71062 : n71176;
  assign n71178 = pi09 ? n17493 : n71177;
  assign n71179 = pi08 ? n71057 : n71178;
  assign n71180 = pi07 ? n70897 : n71179;
  assign n71181 = pi06 ? n70636 : n71180;
  assign n71182 = pi20 ? n321 : ~n9000;
  assign n71183 = pi19 ? n32 : ~n71182;
  assign n71184 = pi18 ? n32 : n71183;
  assign n71185 = pi17 ? n32 : n71184;
  assign n71186 = pi16 ? n32 : n71185;
  assign n71187 = pi15 ? n24247 : n71186;
  assign n71188 = pi15 ? n25708 : n70518;
  assign n71189 = pi14 ? n71187 : n71188;
  assign n71190 = pi13 ? n32 : n71189;
  assign n71191 = pi12 ? n32 : n71190;
  assign n71192 = pi20 ? n175 : n726;
  assign n71193 = pi19 ? n32 : n71192;
  assign n71194 = pi18 ? n32 : n71193;
  assign n71195 = pi17 ? n32 : n71194;
  assign n71196 = pi16 ? n32 : n71195;
  assign n71197 = pi15 ? n71196 : n70243;
  assign n71198 = pi15 ? n17039 : n16850;
  assign n71199 = pi14 ? n71197 : n71198;
  assign n71200 = pi15 ? n17286 : n53119;
  assign n71201 = pi20 ? n220 : ~n1839;
  assign n71202 = pi19 ? n32 : n71201;
  assign n71203 = pi18 ? n32 : n71202;
  assign n71204 = pi17 ? n32 : n71203;
  assign n71205 = pi16 ? n32 : n71204;
  assign n71206 = pi15 ? n70909 : n71205;
  assign n71207 = pi14 ? n71200 : n71206;
  assign n71208 = pi13 ? n71199 : n71207;
  assign n71209 = pi20 ? n14286 : ~n11048;
  assign n71210 = pi19 ? n32 : n71209;
  assign n71211 = pi18 ? n32 : n71210;
  assign n71212 = pi17 ? n32 : n71211;
  assign n71213 = pi16 ? n32 : n71212;
  assign n71214 = pi15 ? n71213 : n55787;
  assign n71215 = pi19 ? n32 : ~n12657;
  assign n71216 = pi18 ? n32 : n71215;
  assign n71217 = pi17 ? n32 : n71216;
  assign n71218 = pi16 ? n32 : n71217;
  assign n71219 = pi19 ? n32 : ~n23396;
  assign n71220 = pi18 ? n32 : n71219;
  assign n71221 = pi17 ? n32 : n71220;
  assign n71222 = pi16 ? n32 : n71221;
  assign n71223 = pi15 ? n71218 : n71222;
  assign n71224 = pi14 ? n71214 : n71223;
  assign n71225 = pi20 ? n39764 : n1940;
  assign n71226 = pi19 ? n32 : ~n71225;
  assign n71227 = pi18 ? n32 : n71226;
  assign n71228 = pi17 ? n32 : n71227;
  assign n71229 = pi16 ? n32 : n71228;
  assign n71230 = pi15 ? n70923 : n71229;
  assign n71231 = pi15 ? n39775 : n15403;
  assign n71232 = pi14 ? n71230 : n71231;
  assign n71233 = pi13 ? n71224 : n71232;
  assign n71234 = pi12 ? n71208 : n71233;
  assign n71235 = pi11 ? n71191 : n71234;
  assign n71236 = pi19 ? n531 : ~n22901;
  assign n71237 = pi18 ? n32 : n71236;
  assign n71238 = pi17 ? n32 : n71237;
  assign n71239 = pi16 ? n32 : n71238;
  assign n71240 = pi19 ? n5694 : n21042;
  assign n71241 = pi18 ? n32 : n71240;
  assign n71242 = pi17 ? n32 : n71241;
  assign n71243 = pi16 ? n32 : n71242;
  assign n71244 = pi15 ? n71239 : n71243;
  assign n71245 = pi20 ? n7229 : ~n141;
  assign n71246 = pi19 ? n32 : n71245;
  assign n71247 = pi18 ? n32 : n71246;
  assign n71248 = pi17 ? n32 : n71247;
  assign n71249 = pi16 ? n32 : n71248;
  assign n71250 = pi15 ? n71249 : n54320;
  assign n71251 = pi14 ? n71244 : n71250;
  assign n71252 = pi20 ? n321 : n915;
  assign n71253 = pi19 ? n71252 : ~n65785;
  assign n71254 = pi18 ? n54334 : n71253;
  assign n71255 = pi17 ? n32 : n71254;
  assign n71256 = pi16 ? n32 : n71255;
  assign n71257 = pi21 ? n1939 : ~n9326;
  assign n71258 = pi20 ? n71257 : n32;
  assign n71259 = pi19 ? n267 : n71258;
  assign n71260 = pi18 ? n54334 : n71259;
  assign n71261 = pi17 ? n32 : n71260;
  assign n71262 = pi16 ? n32 : n71261;
  assign n71263 = pi15 ? n71256 : n71262;
  assign n71264 = pi21 ? n51 : ~n100;
  assign n71265 = pi20 ? n71264 : n32;
  assign n71266 = pi19 ? n34188 : ~n71265;
  assign n71267 = pi18 ? n32 : ~n71266;
  assign n71268 = pi17 ? n32 : n71267;
  assign n71269 = pi16 ? n32 : n71268;
  assign n71270 = pi20 ? n342 : ~n357;
  assign n71271 = pi21 ? n51 : ~n1939;
  assign n71272 = pi20 ? n71271 : n32;
  assign n71273 = pi19 ? n71270 : ~n71272;
  assign n71274 = pi18 ? n32 : ~n71273;
  assign n71275 = pi17 ? n32 : n71274;
  assign n71276 = pi16 ? n32 : n71275;
  assign n71277 = pi15 ? n71269 : n71276;
  assign n71278 = pi14 ? n71263 : n71277;
  assign n71279 = pi13 ? n71251 : n71278;
  assign n71280 = pi21 ? n1939 : ~n124;
  assign n71281 = pi20 ? n71280 : ~n32;
  assign n71282 = pi19 ? n507 : ~n71281;
  assign n71283 = pi18 ? n32 : n71282;
  assign n71284 = pi17 ? n32 : n71283;
  assign n71285 = pi16 ? n32 : n71284;
  assign n71286 = pi15 ? n71285 : n24511;
  assign n71287 = pi14 ? n54434 : n71286;
  assign n71288 = pi15 ? n71121 : n14575;
  assign n71289 = pi19 ? n20006 : n358;
  assign n71290 = pi18 ? n32 : n71289;
  assign n71291 = pi17 ? n32 : n71290;
  assign n71292 = pi16 ? n32 : n71291;
  assign n71293 = pi15 ? n25466 : n71292;
  assign n71294 = pi14 ? n71288 : n71293;
  assign n71295 = pi13 ? n71287 : n71294;
  assign n71296 = pi12 ? n71279 : n71295;
  assign n71297 = pi19 ? n21137 : n1941;
  assign n71298 = pi18 ? n590 : ~n71297;
  assign n71299 = pi17 ? n32 : n71298;
  assign n71300 = pi16 ? n32 : n71299;
  assign n71301 = pi19 ? n9007 : n1941;
  assign n71302 = pi18 ? n4392 : ~n71301;
  assign n71303 = pi17 ? n32 : n71302;
  assign n71304 = pi16 ? n32 : n71303;
  assign n71305 = pi15 ? n71300 : n71304;
  assign n71306 = pi20 ? n32 : ~n7007;
  assign n71307 = pi19 ? n71306 : n236;
  assign n71308 = pi18 ? n7368 : ~n71307;
  assign n71309 = pi17 ? n32 : n71308;
  assign n71310 = pi16 ? n32 : n71309;
  assign n71311 = pi20 ? n32 : n20501;
  assign n71312 = pi19 ? n71311 : ~n32;
  assign n71313 = pi18 ? n940 : ~n71312;
  assign n71314 = pi17 ? n32 : n71313;
  assign n71315 = pi16 ? n32 : n71314;
  assign n71316 = pi15 ? n71310 : n71315;
  assign n71317 = pi14 ? n71305 : n71316;
  assign n71318 = pi18 ? n16847 : ~n508;
  assign n71319 = pi17 ? n32 : n71318;
  assign n71320 = pi16 ? n32 : n71319;
  assign n71321 = pi20 ? n342 : ~n17654;
  assign n71322 = pi19 ? n71321 : ~n32;
  assign n71323 = pi18 ? n4722 : ~n71322;
  assign n71324 = pi17 ? n32 : n71323;
  assign n71325 = pi16 ? n32 : n71324;
  assign n71326 = pi15 ? n71320 : n71325;
  assign n71327 = pi20 ? n518 : ~n18158;
  assign n71328 = pi19 ? n71327 : ~n32;
  assign n71329 = pi18 ? n684 : ~n71328;
  assign n71330 = pi17 ? n32 : n71329;
  assign n71331 = pi16 ? n32 : n71330;
  assign n71332 = pi19 ? n32 : n18396;
  assign n71333 = pi18 ? n71332 : n25185;
  assign n71334 = pi17 ? n32 : n71333;
  assign n71335 = pi16 ? n32 : n71334;
  assign n71336 = pi15 ? n71331 : n71335;
  assign n71337 = pi14 ? n71326 : n71336;
  assign n71338 = pi13 ? n71317 : n71337;
  assign n71339 = pi15 ? n22376 : n14397;
  assign n71340 = pi19 ? n52399 : n32;
  assign n71341 = pi18 ? n17118 : n71340;
  assign n71342 = pi17 ? n32 : n71341;
  assign n71343 = pi16 ? n32 : n71342;
  assign n71344 = pi20 ? n266 : ~n1839;
  assign n71345 = pi19 ? n71344 : n32;
  assign n71346 = pi18 ? n16981 : n71345;
  assign n71347 = pi17 ? n32 : n71346;
  assign n71348 = pi16 ? n32 : n71347;
  assign n71349 = pi15 ? n71343 : n71348;
  assign n71350 = pi14 ? n71339 : n71349;
  assign n71351 = pi18 ? n47419 : ~n1914;
  assign n71352 = pi17 ? n32 : n71351;
  assign n71353 = pi16 ? n32 : n71352;
  assign n71354 = pi15 ? n71353 : n12091;
  assign n71355 = pi18 ? n42416 : ~n605;
  assign n71356 = pi17 ? n32 : n71355;
  assign n71357 = pi16 ? n32 : n71356;
  assign n71358 = pi18 ? n268 : ~n418;
  assign n71359 = pi17 ? n32 : n71358;
  assign n71360 = pi16 ? n32 : n71359;
  assign n71361 = pi15 ? n71357 : n71360;
  assign n71362 = pi14 ? n71354 : n71361;
  assign n71363 = pi13 ? n71350 : n71362;
  assign n71364 = pi12 ? n71338 : n71363;
  assign n71365 = pi11 ? n71296 : n71364;
  assign n71366 = pi10 ? n71235 : n71365;
  assign n71367 = pi09 ? n17493 : n71366;
  assign n71368 = pi15 ? n16485 : n70518;
  assign n71369 = pi14 ? n71187 : n71368;
  assign n71370 = pi13 ? n40837 : n71369;
  assign n71371 = pi12 ? n32 : n71370;
  assign n71372 = pi15 ? n16587 : n55787;
  assign n71373 = pi19 ? n32 : ~n12666;
  assign n71374 = pi18 ? n32 : n71373;
  assign n71375 = pi17 ? n32 : n71374;
  assign n71376 = pi16 ? n32 : n71375;
  assign n71377 = pi15 ? n71218 : n71376;
  assign n71378 = pi14 ? n71372 : n71377;
  assign n71379 = pi19 ? n32 : ~n8247;
  assign n71380 = pi18 ? n32 : n71379;
  assign n71381 = pi17 ? n32 : n71380;
  assign n71382 = pi16 ? n32 : n71381;
  assign n71383 = pi15 ? n70923 : n71382;
  assign n71384 = pi20 ? n339 : n481;
  assign n71385 = pi19 ? n32 : n71384;
  assign n71386 = pi18 ? n32 : n71385;
  assign n71387 = pi17 ? n32 : n71386;
  assign n71388 = pi16 ? n32 : n71387;
  assign n71389 = pi15 ? n15847 : n71388;
  assign n71390 = pi14 ? n71383 : n71389;
  assign n71391 = pi13 ? n71378 : n71390;
  assign n71392 = pi12 ? n71208 : n71391;
  assign n71393 = pi11 ? n71371 : n71392;
  assign n71394 = pi19 ? n5694 : n7405;
  assign n71395 = pi18 ? n32 : n71394;
  assign n71396 = pi17 ? n32 : n71395;
  assign n71397 = pi16 ? n32 : n71396;
  assign n71398 = pi15 ? n71239 : n71397;
  assign n71399 = pi19 ? n68 : n27066;
  assign n71400 = pi18 ? n32 : n71399;
  assign n71401 = pi17 ? n32 : n71400;
  assign n71402 = pi16 ? n32 : n71401;
  assign n71403 = pi15 ? n71402 : n54320;
  assign n71404 = pi14 ? n71398 : n71403;
  assign n71405 = pi21 ? n51 : ~n405;
  assign n71406 = pi20 ? n71405 : n32;
  assign n71407 = pi19 ? n34188 : ~n71406;
  assign n71408 = pi18 ? n32 : ~n71407;
  assign n71409 = pi17 ? n32 : n71408;
  assign n71410 = pi16 ? n32 : n71409;
  assign n71411 = pi19 ? n71270 : ~n3495;
  assign n71412 = pi18 ? n32 : ~n71411;
  assign n71413 = pi17 ? n32 : n71412;
  assign n71414 = pi16 ? n32 : n71413;
  assign n71415 = pi15 ? n71410 : n71414;
  assign n71416 = pi14 ? n71263 : n71415;
  assign n71417 = pi13 ? n71404 : n71416;
  assign n71418 = pi19 ? n507 : ~n11123;
  assign n71419 = pi18 ? n32 : n71418;
  assign n71420 = pi17 ? n32 : n71419;
  assign n71421 = pi16 ? n32 : n71420;
  assign n71422 = pi15 ? n71421 : n24511;
  assign n71423 = pi14 ? n54347 : n71422;
  assign n71424 = pi21 ? n7410 : n206;
  assign n71425 = pi20 ? n32 : ~n71424;
  assign n71426 = pi19 ? n71425 : n53;
  assign n71427 = pi18 ? n32 : n71426;
  assign n71428 = pi17 ? n32 : n71427;
  assign n71429 = pi16 ? n32 : n71428;
  assign n71430 = pi15 ? n25466 : n71429;
  assign n71431 = pi14 ? n71288 : n71430;
  assign n71432 = pi13 ? n71423 : n71431;
  assign n71433 = pi12 ? n71417 : n71432;
  assign n71434 = pi19 ? n275 : n1941;
  assign n71435 = pi18 ? n684 : ~n71434;
  assign n71436 = pi17 ? n32 : n71435;
  assign n71437 = pi16 ? n32 : n71436;
  assign n71438 = pi19 ? n9007 : n236;
  assign n71439 = pi18 ? n1741 : ~n71438;
  assign n71440 = pi17 ? n32 : n71439;
  assign n71441 = pi16 ? n32 : n71440;
  assign n71442 = pi15 ? n71437 : n71441;
  assign n71443 = pi19 ? n5730 : n1105;
  assign n71444 = pi18 ? n209 : ~n71443;
  assign n71445 = pi17 ? n32 : n71444;
  assign n71446 = pi16 ? n32 : n71445;
  assign n71447 = pi21 ? n174 : n12274;
  assign n71448 = pi20 ? n32 : n71447;
  assign n71449 = pi19 ? n71448 : ~n32;
  assign n71450 = pi18 ? n940 : ~n71449;
  assign n71451 = pi17 ? n32 : n71450;
  assign n71452 = pi16 ? n32 : n71451;
  assign n71453 = pi15 ? n71446 : n71452;
  assign n71454 = pi14 ? n71442 : n71453;
  assign n71455 = pi20 ? n342 : ~n26934;
  assign n71456 = pi19 ? n71455 : ~n32;
  assign n71457 = pi18 ? n4722 : ~n71456;
  assign n71458 = pi17 ? n32 : n71457;
  assign n71459 = pi16 ? n32 : n71458;
  assign n71460 = pi15 ? n71320 : n71459;
  assign n71461 = pi18 ? n880 : ~n71157;
  assign n71462 = pi17 ? n32 : n71461;
  assign n71463 = pi16 ? n32 : n71462;
  assign n71464 = pi18 ? n4380 : n25116;
  assign n71465 = pi17 ? n32 : n71464;
  assign n71466 = pi16 ? n32 : n71465;
  assign n71467 = pi15 ? n71463 : n71466;
  assign n71468 = pi14 ? n71460 : n71467;
  assign n71469 = pi13 ? n71454 : n71468;
  assign n71470 = pi20 ? n32 : n31747;
  assign n71471 = pi19 ? n71470 : n32;
  assign n71472 = pi18 ? n32 : n71471;
  assign n71473 = pi17 ? n32 : n71472;
  assign n71474 = pi16 ? n32 : n71473;
  assign n71475 = pi20 ? n11560 : ~n1839;
  assign n71476 = pi19 ? n71475 : n32;
  assign n71477 = pi18 ? n32 : n71476;
  assign n71478 = pi17 ? n32 : n71477;
  assign n71479 = pi16 ? n32 : n71478;
  assign n71480 = pi15 ? n71474 : n71479;
  assign n71481 = pi14 ? n27189 : n71480;
  assign n71482 = pi18 ? n209 : ~n1914;
  assign n71483 = pi17 ? n32 : n71482;
  assign n71484 = pi16 ? n32 : n71483;
  assign n71485 = pi20 ? n101 : n1940;
  assign n71486 = pi19 ? n71485 : ~n32;
  assign n71487 = pi18 ? n209 : ~n71486;
  assign n71488 = pi17 ? n32 : n71487;
  assign n71489 = pi16 ? n32 : n71488;
  assign n71490 = pi15 ? n71484 : n71489;
  assign n71491 = pi18 ? n222 : ~n605;
  assign n71492 = pi17 ? n32 : n71491;
  assign n71493 = pi16 ? n32 : n71492;
  assign n71494 = pi18 ? n268 : ~n3786;
  assign n71495 = pi17 ? n32 : n71494;
  assign n71496 = pi16 ? n32 : n71495;
  assign n71497 = pi15 ? n71493 : n71496;
  assign n71498 = pi14 ? n71490 : n71497;
  assign n71499 = pi13 ? n71481 : n71498;
  assign n71500 = pi12 ? n71469 : n71499;
  assign n71501 = pi11 ? n71433 : n71500;
  assign n71502 = pi10 ? n71393 : n71501;
  assign n71503 = pi09 ? n17493 : n71502;
  assign n71504 = pi08 ? n71367 : n71503;
  assign n71505 = pi20 ? n246 : ~n9000;
  assign n71506 = pi19 ? n32 : ~n71505;
  assign n71507 = pi18 ? n32 : n71506;
  assign n71508 = pi17 ? n32 : n71507;
  assign n71509 = pi16 ? n32 : n71508;
  assign n71510 = pi15 ? n24247 : n71509;
  assign n71511 = pi20 ? n32 : ~n16253;
  assign n71512 = pi19 ? n32 : n71511;
  assign n71513 = pi18 ? n32 : n71512;
  assign n71514 = pi17 ? n32 : n71513;
  assign n71515 = pi16 ? n32 : n71514;
  assign n71516 = pi15 ? n16485 : n71515;
  assign n71517 = pi14 ? n71510 : n71516;
  assign n71518 = pi13 ? n36490 : n71517;
  assign n71519 = pi12 ? n32 : n71518;
  assign n71520 = pi15 ? n26515 : n68991;
  assign n71521 = pi14 ? n71520 : n16851;
  assign n71522 = pi19 ? n32 : ~n8212;
  assign n71523 = pi18 ? n32 : n71522;
  assign n71524 = pi17 ? n32 : n71523;
  assign n71525 = pi16 ? n32 : n71524;
  assign n71526 = pi20 ? n10644 : ~n1839;
  assign n71527 = pi19 ? n32 : n71526;
  assign n71528 = pi18 ? n32 : n71527;
  assign n71529 = pi17 ? n32 : n71528;
  assign n71530 = pi16 ? n32 : n71529;
  assign n71531 = pi15 ? n71525 : n71530;
  assign n71532 = pi14 ? n53119 : n71531;
  assign n71533 = pi13 ? n71521 : n71532;
  assign n71534 = pi15 ? n54872 : n26009;
  assign n71535 = pi14 ? n71534 : n71377;
  assign n71536 = pi19 ? n32 : ~n8803;
  assign n71537 = pi18 ? n32 : n71536;
  assign n71538 = pi17 ? n32 : n71537;
  assign n71539 = pi16 ? n32 : n71538;
  assign n71540 = pi15 ? n71539 : n54472;
  assign n71541 = pi20 ? n220 : n481;
  assign n71542 = pi19 ? n32 : n71541;
  assign n71543 = pi18 ? n32 : n71542;
  assign n71544 = pi17 ? n32 : n71543;
  assign n71545 = pi16 ? n32 : n71544;
  assign n71546 = pi15 ? n24874 : n71545;
  assign n71547 = pi14 ? n71540 : n71546;
  assign n71548 = pi13 ? n71535 : n71547;
  assign n71549 = pi12 ? n71533 : n71548;
  assign n71550 = pi11 ? n71519 : n71549;
  assign n71551 = pi19 ? n531 : n21154;
  assign n71552 = pi18 ? n32 : n71551;
  assign n71553 = pi17 ? n32 : n71552;
  assign n71554 = pi16 ? n32 : n71553;
  assign n71555 = pi15 ? n71554 : n71397;
  assign n71556 = pi19 ? n236 : n11108;
  assign n71557 = pi18 ? n32 : ~n71556;
  assign n71558 = pi17 ? n32 : n71557;
  assign n71559 = pi16 ? n32 : n71558;
  assign n71560 = pi19 ? n142 : ~n236;
  assign n71561 = pi18 ? n32 : n71560;
  assign n71562 = pi17 ? n32 : n71561;
  assign n71563 = pi16 ? n32 : n71562;
  assign n71564 = pi15 ? n71559 : n71563;
  assign n71565 = pi14 ? n71555 : n71564;
  assign n71566 = pi21 ? n140 : ~n2076;
  assign n71567 = pi20 ? n71566 : ~n32;
  assign n71568 = pi19 ? n4964 : ~n71567;
  assign n71569 = pi18 ? n863 : n71568;
  assign n71570 = pi17 ? n32 : n71569;
  assign n71571 = pi16 ? n32 : n71570;
  assign n71572 = pi19 ? n267 : n19847;
  assign n71573 = pi18 ? n863 : n71572;
  assign n71574 = pi17 ? n32 : n71573;
  assign n71575 = pi16 ? n32 : n71574;
  assign n71576 = pi15 ? n71571 : n71575;
  assign n71577 = pi19 ? n4964 : n429;
  assign n71578 = pi18 ? n32 : ~n71577;
  assign n71579 = pi17 ? n32 : n71578;
  assign n71580 = pi16 ? n32 : n71579;
  assign n71581 = pi15 ? n71580 : n12784;
  assign n71582 = pi14 ? n71576 : n71581;
  assign n71583 = pi13 ? n71565 : n71582;
  assign n71584 = pi15 ? n32 : n24813;
  assign n71585 = pi19 ? n507 : ~n10890;
  assign n71586 = pi18 ? n32 : n71585;
  assign n71587 = pi17 ? n32 : n71586;
  assign n71588 = pi16 ? n32 : n71587;
  assign n71589 = pi15 ? n71588 : n24504;
  assign n71590 = pi14 ? n71584 : n71589;
  assign n71591 = pi15 ? n39520 : n14580;
  assign n71592 = pi21 ? n35 : ~n9326;
  assign n71593 = pi20 ? n339 : ~n71592;
  assign n71594 = pi19 ? n71593 : ~n7502;
  assign n71595 = pi18 ? n1012 : ~n71594;
  assign n71596 = pi17 ? n32 : n71595;
  assign n71597 = pi16 ? n32 : n71596;
  assign n71598 = pi15 ? n22825 : n71597;
  assign n71599 = pi14 ? n71591 : n71598;
  assign n71600 = pi13 ? n71590 : n71599;
  assign n71601 = pi12 ? n71583 : n71600;
  assign n71602 = pi19 ? n221 : n1941;
  assign n71603 = pi18 ? n940 : ~n71602;
  assign n71604 = pi17 ? n32 : n71603;
  assign n71605 = pi16 ? n32 : n71604;
  assign n71606 = pi19 ? n662 : n236;
  assign n71607 = pi18 ? n940 : ~n71606;
  assign n71608 = pi17 ? n32 : n71607;
  assign n71609 = pi16 ? n32 : n71608;
  assign n71610 = pi15 ? n71605 : n71609;
  assign n71611 = pi21 ? n85 : ~n32;
  assign n71612 = pi20 ? n32 : ~n71611;
  assign n71613 = pi19 ? n71612 : n1105;
  assign n71614 = pi18 ? n751 : ~n71613;
  assign n71615 = pi17 ? n32 : n71614;
  assign n71616 = pi16 ? n32 : n71615;
  assign n71617 = pi19 ? n14661 : ~n32;
  assign n71618 = pi18 ? n751 : ~n71617;
  assign n71619 = pi17 ? n32 : n71618;
  assign n71620 = pi16 ? n32 : n71619;
  assign n71621 = pi15 ? n71616 : n71620;
  assign n71622 = pi14 ? n71610 : n71621;
  assign n71623 = pi21 ? n140 : ~n7107;
  assign n71624 = pi20 ? n32 : n71623;
  assign n71625 = pi19 ? n71624 : ~n32;
  assign n71626 = pi18 ? n268 : ~n71625;
  assign n71627 = pi17 ? n32 : n71626;
  assign n71628 = pi16 ? n32 : n71627;
  assign n71629 = pi20 ? n342 : ~n27235;
  assign n71630 = pi19 ? n71629 : ~n32;
  assign n71631 = pi18 ? n4127 : ~n71630;
  assign n71632 = pi17 ? n32 : n71631;
  assign n71633 = pi16 ? n32 : n71632;
  assign n71634 = pi15 ? n71628 : n71633;
  assign n71635 = pi18 ? n940 : ~n23200;
  assign n71636 = pi17 ? n32 : n71635;
  assign n71637 = pi16 ? n32 : n71636;
  assign n71638 = pi18 ? n4380 : n21683;
  assign n71639 = pi17 ? n32 : n71638;
  assign n71640 = pi16 ? n32 : n71639;
  assign n71641 = pi15 ? n71637 : n71640;
  assign n71642 = pi14 ? n71634 : n71641;
  assign n71643 = pi13 ? n71622 : n71642;
  assign n71644 = pi18 ? n1819 : n14165;
  assign n71645 = pi17 ? n32 : n71644;
  assign n71646 = pi16 ? n32 : n71645;
  assign n71647 = pi18 ? n1592 : n32474;
  assign n71648 = pi17 ? n32 : n71647;
  assign n71649 = pi16 ? n32 : n71648;
  assign n71650 = pi15 ? n71646 : n71649;
  assign n71651 = pi14 ? n27172 : n71650;
  assign n71652 = pi15 ? n12781 : n12538;
  assign n71653 = pi15 ? n12542 : n12791;
  assign n71654 = pi14 ? n71652 : n71653;
  assign n71655 = pi13 ? n71651 : n71654;
  assign n71656 = pi12 ? n71643 : n71655;
  assign n71657 = pi11 ? n71601 : n71656;
  assign n71658 = pi10 ? n71550 : n71657;
  assign n71659 = pi09 ? n17493 : n71658;
  assign n71660 = pi19 ? n32 : ~n40989;
  assign n71661 = pi18 ? n32 : n71660;
  assign n71662 = pi17 ? n32 : n71661;
  assign n71663 = pi16 ? n32 : n71662;
  assign n71664 = pi15 ? n24247 : n71663;
  assign n71665 = pi15 ? n16485 : n26951;
  assign n71666 = pi14 ? n71664 : n71665;
  assign n71667 = pi13 ? n36490 : n71666;
  assign n71668 = pi12 ? n32 : n71667;
  assign n71669 = pi15 ? n54872 : n32;
  assign n71670 = pi19 ? n32 : ~n1476;
  assign n71671 = pi18 ? n32 : n71670;
  assign n71672 = pi17 ? n32 : n71671;
  assign n71673 = pi16 ? n32 : n71672;
  assign n71674 = pi15 ? n71218 : n71673;
  assign n71675 = pi14 ? n71669 : n71674;
  assign n71676 = pi13 ? n71675 : n71547;
  assign n71677 = pi12 ? n71533 : n71676;
  assign n71678 = pi11 ? n71668 : n71677;
  assign n71679 = pi15 ? n71559 : n23484;
  assign n71680 = pi14 ? n71555 : n71679;
  assign n71681 = pi19 ? n2025 : ~n32;
  assign n71682 = pi18 ? n32 : ~n71681;
  assign n71683 = pi17 ? n32 : n71682;
  assign n71684 = pi16 ? n32 : n71683;
  assign n71685 = pi15 ? n71580 : n71684;
  assign n71686 = pi14 ? n71576 : n71685;
  assign n71687 = pi13 ? n71680 : n71686;
  assign n71688 = pi15 ? n32 : n40057;
  assign n71689 = pi19 ? n462 : ~n6693;
  assign n71690 = pi18 ? n32 : n71689;
  assign n71691 = pi17 ? n32 : n71690;
  assign n71692 = pi16 ? n32 : n71691;
  assign n71693 = pi15 ? n71588 : n71692;
  assign n71694 = pi14 ? n71688 : n71693;
  assign n71695 = pi19 ? n2359 : ~n813;
  assign n71696 = pi18 ? n32 : n71695;
  assign n71697 = pi17 ? n32 : n71696;
  assign n71698 = pi16 ? n32 : n71697;
  assign n71699 = pi15 ? n71698 : n14580;
  assign n71700 = pi20 ? n339 : ~n53890;
  assign n71701 = pi19 ? n71700 : ~n7502;
  assign n71702 = pi18 ? n1575 : ~n71701;
  assign n71703 = pi17 ? n32 : n71702;
  assign n71704 = pi16 ? n32 : n71703;
  assign n71705 = pi15 ? n22825 : n71704;
  assign n71706 = pi14 ? n71699 : n71705;
  assign n71707 = pi13 ? n71694 : n71706;
  assign n71708 = pi12 ? n71687 : n71707;
  assign n71709 = pi19 ? n9220 : n1941;
  assign n71710 = pi18 ? n940 : ~n71709;
  assign n71711 = pi17 ? n32 : n71710;
  assign n71712 = pi16 ? n32 : n71711;
  assign n71713 = pi19 ? n462 : n617;
  assign n71714 = pi18 ? n940 : ~n71713;
  assign n71715 = pi17 ? n32 : n71714;
  assign n71716 = pi16 ? n32 : n71715;
  assign n71717 = pi15 ? n71712 : n71716;
  assign n71718 = pi19 ? n572 : n1105;
  assign n71719 = pi18 ? n940 : ~n71718;
  assign n71720 = pi17 ? n32 : n71719;
  assign n71721 = pi16 ? n32 : n71720;
  assign n71722 = pi19 ? n1145 : ~n32;
  assign n71723 = pi18 ? n940 : ~n71722;
  assign n71724 = pi17 ? n32 : n71723;
  assign n71725 = pi16 ? n32 : n71724;
  assign n71726 = pi15 ? n71721 : n71725;
  assign n71727 = pi14 ? n71717 : n71726;
  assign n71728 = pi18 ? n32 : ~n47421;
  assign n71729 = pi17 ? n32 : n71728;
  assign n71730 = pi16 ? n32 : n71729;
  assign n71731 = pi21 ? n313 : n100;
  assign n71732 = pi20 ? n342 : n71731;
  assign n71733 = pi19 ? n71732 : ~n32;
  assign n71734 = pi18 ? n863 : ~n71733;
  assign n71735 = pi17 ? n32 : n71734;
  assign n71736 = pi16 ? n32 : n71735;
  assign n71737 = pi15 ? n71730 : n71736;
  assign n71738 = pi18 ? n863 : ~n23200;
  assign n71739 = pi17 ? n32 : n71738;
  assign n71740 = pi16 ? n32 : n71739;
  assign n71741 = pi15 ? n71740 : n21686;
  assign n71742 = pi14 ? n71737 : n71741;
  assign n71743 = pi13 ? n71727 : n71742;
  assign n71744 = pi15 ? n22006 : n14156;
  assign n71745 = pi20 ? n206 : n439;
  assign n71746 = pi19 ? n71745 : n32;
  assign n71747 = pi18 ? n863 : n71746;
  assign n71748 = pi17 ? n32 : n71747;
  assign n71749 = pi16 ? n32 : n71748;
  assign n71750 = pi15 ? n14168 : n71749;
  assign n71751 = pi14 ? n71744 : n71750;
  assign n71752 = pi13 ? n71751 : n12793;
  assign n71753 = pi12 ? n71743 : n71752;
  assign n71754 = pi11 ? n71708 : n71753;
  assign n71755 = pi10 ? n71678 : n71754;
  assign n71756 = pi09 ? n17493 : n71755;
  assign n71757 = pi08 ? n71659 : n71756;
  assign n71758 = pi07 ? n71504 : n71757;
  assign n71759 = pi19 ? n507 : n13906;
  assign n71760 = pi18 ? n32 : n71759;
  assign n71761 = pi17 ? n32 : n71760;
  assign n71762 = pi16 ? n32 : n71761;
  assign n71763 = pi15 ? n17278 : n71762;
  assign n71764 = pi15 ? n65606 : n26951;
  assign n71765 = pi14 ? n71763 : n71764;
  assign n71766 = pi13 ? n32 : n71765;
  assign n71767 = pi12 ? n32 : n71766;
  assign n71768 = pi20 ? n321 : ~n564;
  assign n71769 = pi19 ? n32 : ~n71768;
  assign n71770 = pi18 ? n32 : n71769;
  assign n71771 = pi17 ? n32 : n71770;
  assign n71772 = pi16 ? n32 : n71771;
  assign n71773 = pi15 ? n71772 : n24247;
  assign n71774 = pi14 ? n68991 : n71773;
  assign n71775 = pi20 ? n9641 : ~n518;
  assign n71776 = pi19 ? n507 : n71775;
  assign n71777 = pi18 ? n32 : n71776;
  assign n71778 = pi17 ? n32 : n71777;
  assign n71779 = pi16 ? n32 : n71778;
  assign n71780 = pi20 ? n1324 : ~n518;
  assign n71781 = pi19 ? n1818 : n71780;
  assign n71782 = pi18 ? n32 : n71781;
  assign n71783 = pi17 ? n32 : n71782;
  assign n71784 = pi16 ? n32 : n71783;
  assign n71785 = pi15 ? n71779 : n71784;
  assign n71786 = pi19 ? n1818 : ~n8212;
  assign n71787 = pi18 ? n32 : n71786;
  assign n71788 = pi17 ? n32 : n71787;
  assign n71789 = pi16 ? n32 : n71788;
  assign n71790 = pi20 ? n1817 : n1475;
  assign n71791 = pi19 ? n32 : ~n71790;
  assign n71792 = pi18 ? n32 : n71791;
  assign n71793 = pi17 ? n32 : n71792;
  assign n71794 = pi16 ? n32 : n71793;
  assign n71795 = pi15 ? n71789 : n71794;
  assign n71796 = pi14 ? n71785 : n71795;
  assign n71797 = pi13 ? n71774 : n71796;
  assign n71798 = pi19 ? n322 : ~n12657;
  assign n71799 = pi18 ? n32 : n71798;
  assign n71800 = pi17 ? n32 : n71799;
  assign n71801 = pi16 ? n32 : n71800;
  assign n71802 = pi15 ? n16546 : n71801;
  assign n71803 = pi20 ? n9641 : n1475;
  assign n71804 = pi19 ? n322 : ~n71803;
  assign n71805 = pi18 ? n32 : n71804;
  assign n71806 = pi17 ? n32 : n71805;
  assign n71807 = pi16 ? n32 : n71806;
  assign n71808 = pi15 ? n71807 : n16352;
  assign n71809 = pi14 ? n71802 : n71808;
  assign n71810 = pi15 ? n54636 : n24700;
  assign n71811 = pi19 ? n507 : ~n12957;
  assign n71812 = pi18 ? n32 : n71811;
  assign n71813 = pi17 ? n32 : n71812;
  assign n71814 = pi16 ? n32 : n71813;
  assign n71815 = pi19 ? n32 : ~n33595;
  assign n71816 = pi18 ? n32 : n71815;
  assign n71817 = pi17 ? n32 : n71816;
  assign n71818 = pi16 ? n32 : n71817;
  assign n71819 = pi15 ? n71814 : n71818;
  assign n71820 = pi14 ? n71810 : n71819;
  assign n71821 = pi13 ? n71809 : n71820;
  assign n71822 = pi12 ? n71797 : n71821;
  assign n71823 = pi11 ? n71767 : n71822;
  assign n71824 = pi19 ? n5741 : n68169;
  assign n71825 = pi18 ? n32 : n71824;
  assign n71826 = pi17 ? n32 : n71825;
  assign n71827 = pi16 ? n32 : n71826;
  assign n71828 = pi20 ? n47301 : n32;
  assign n71829 = pi19 ? n236 : n71828;
  assign n71830 = pi18 ? n32 : n71829;
  assign n71831 = pi17 ? n32 : n71830;
  assign n71832 = pi16 ? n32 : n71831;
  assign n71833 = pi15 ? n71827 : n71832;
  assign n71834 = pi20 ? n915 : ~n321;
  assign n71835 = pi20 ? n18540 : ~n32;
  assign n71836 = pi19 ? n71834 : ~n71835;
  assign n71837 = pi18 ? n32 : n71836;
  assign n71838 = pi17 ? n32 : n71837;
  assign n71839 = pi16 ? n32 : n71838;
  assign n71840 = pi18 ? n1575 : n20172;
  assign n71841 = pi17 ? n32 : n71840;
  assign n71842 = pi16 ? n32 : n71841;
  assign n71843 = pi15 ? n71839 : n71842;
  assign n71844 = pi14 ? n71833 : n71843;
  assign n71845 = pi21 ? n259 : n2076;
  assign n71846 = pi20 ? n71845 : n32;
  assign n71847 = pi19 ? n62288 : n71846;
  assign n71848 = pi18 ? n936 : n71847;
  assign n71849 = pi17 ? n32 : n71848;
  assign n71850 = pi16 ? n32 : n71849;
  assign n71851 = pi21 ? n1392 : ~n100;
  assign n71852 = pi20 ? n71851 : n32;
  assign n71853 = pi19 ? n4721 : n71852;
  assign n71854 = pi18 ? n32 : n71853;
  assign n71855 = pi17 ? n32 : n71854;
  assign n71856 = pi16 ? n32 : n71855;
  assign n71857 = pi15 ? n71850 : n71856;
  assign n71858 = pi20 ? n12882 : ~n32;
  assign n71859 = pi19 ? n62288 : n71858;
  assign n71860 = pi18 ? n32 : ~n71859;
  assign n71861 = pi17 ? n32 : n71860;
  assign n71862 = pi16 ? n32 : n71861;
  assign n71863 = pi20 ? n260 : ~n342;
  assign n71864 = pi19 ? n71863 : ~n32;
  assign n71865 = pi18 ? n936 : ~n71864;
  assign n71866 = pi17 ? n32 : n71865;
  assign n71867 = pi16 ? n32 : n71866;
  assign n71868 = pi15 ? n71862 : n71867;
  assign n71869 = pi14 ? n71857 : n71868;
  assign n71870 = pi13 ? n71844 : n71869;
  assign n71871 = pi19 ? n221 : n9724;
  assign n71872 = pi18 ? n32 : n71871;
  assign n71873 = pi17 ? n32 : n71872;
  assign n71874 = pi16 ? n32 : n71873;
  assign n71875 = pi15 ? n52178 : n71874;
  assign n71876 = pi19 ? n4982 : ~n10890;
  assign n71877 = pi18 ? n32 : n71876;
  assign n71878 = pi17 ? n32 : n71877;
  assign n71879 = pi16 ? n32 : n71878;
  assign n71880 = pi19 ? n4721 : n7693;
  assign n71881 = pi18 ? n32 : n71880;
  assign n71882 = pi17 ? n32 : n71881;
  assign n71883 = pi16 ? n32 : n71882;
  assign n71884 = pi15 ? n71879 : n71883;
  assign n71885 = pi14 ? n71875 : n71884;
  assign n71886 = pi19 ? n42677 : ~n813;
  assign n71887 = pi18 ? n32 : n71886;
  assign n71888 = pi17 ? n32 : n71887;
  assign n71889 = pi16 ? n32 : n71888;
  assign n71890 = pi19 ? n47981 : ~n236;
  assign n71891 = pi18 ? n32 : n71890;
  assign n71892 = pi17 ? n32 : n71891;
  assign n71893 = pi16 ? n32 : n71892;
  assign n71894 = pi15 ? n71889 : n71893;
  assign n71895 = pi19 ? n617 : ~n1941;
  assign n71896 = pi18 ? n32 : n71895;
  assign n71897 = pi17 ? n32 : n71896;
  assign n71898 = pi16 ? n32 : n71897;
  assign n71899 = pi15 ? n71898 : n24179;
  assign n71900 = pi14 ? n71894 : n71899;
  assign n71901 = pi13 ? n71885 : n71900;
  assign n71902 = pi12 ? n71870 : n71901;
  assign n71903 = pi19 ? n8388 : ~n617;
  assign n71904 = pi18 ? n863 : n71903;
  assign n71905 = pi17 ? n32 : n71904;
  assign n71906 = pi16 ? n32 : n71905;
  assign n71907 = pi19 ? n36510 : ~n1105;
  assign n71908 = pi18 ? n863 : n71907;
  assign n71909 = pi17 ? n32 : n71908;
  assign n71910 = pi16 ? n32 : n71909;
  assign n71911 = pi15 ? n71906 : n71910;
  assign n71912 = pi20 ? n321 : ~n12884;
  assign n71913 = pi19 ? n71912 : ~n1105;
  assign n71914 = pi18 ? n32 : n71913;
  assign n71915 = pi17 ? n32 : n71914;
  assign n71916 = pi16 ? n32 : n71915;
  assign n71917 = pi20 ? n220 : n13084;
  assign n71918 = pi19 ? n71917 : n32;
  assign n71919 = pi18 ? n32 : n71918;
  assign n71920 = pi17 ? n32 : n71919;
  assign n71921 = pi16 ? n32 : n71920;
  assign n71922 = pi15 ? n71916 : n71921;
  assign n71923 = pi14 ? n71911 : n71922;
  assign n71924 = pi19 ? n30681 : n32;
  assign n71925 = pi18 ? n32 : n71924;
  assign n71926 = pi17 ? n32 : n71925;
  assign n71927 = pi16 ? n32 : n71926;
  assign n71928 = pi19 ? n51660 : n32;
  assign n71929 = pi18 ? n32 : n71928;
  assign n71930 = pi17 ? n32 : n71929;
  assign n71931 = pi16 ? n32 : n71930;
  assign n71932 = pi15 ? n71927 : n71931;
  assign n71933 = pi20 ? n207 : ~n7852;
  assign n71934 = pi19 ? n71933 : ~n32;
  assign n71935 = pi18 ? n32 : ~n71934;
  assign n71936 = pi17 ? n32 : n71935;
  assign n71937 = pi16 ? n32 : n71936;
  assign n71938 = pi20 ? n820 : ~n623;
  assign n71939 = pi19 ? n71938 : ~n32;
  assign n71940 = pi18 ? n32 : ~n71939;
  assign n71941 = pi17 ? n32 : n71940;
  assign n71942 = pi16 ? n32 : n71941;
  assign n71943 = pi15 ? n71937 : n71942;
  assign n71944 = pi14 ? n71932 : n71943;
  assign n71945 = pi13 ? n71923 : n71944;
  assign n71946 = pi20 ? n246 : n6229;
  assign n71947 = pi19 ? n71946 : n32;
  assign n71948 = pi18 ? n32 : n71947;
  assign n71949 = pi17 ? n32 : n71948;
  assign n71950 = pi16 ? n32 : n71949;
  assign n71951 = pi19 ? n68854 : n32;
  assign n71952 = pi18 ? n32 : n71951;
  assign n71953 = pi17 ? n32 : n71952;
  assign n71954 = pi16 ? n32 : n71953;
  assign n71955 = pi15 ? n71950 : n71954;
  assign n71956 = pi20 ? n405 : n439;
  assign n71957 = pi19 ? n71956 : n32;
  assign n71958 = pi18 ? n32 : n71957;
  assign n71959 = pi17 ? n32 : n71958;
  assign n71960 = pi16 ? n32 : n71959;
  assign n71961 = pi15 ? n71960 : n13066;
  assign n71962 = pi14 ? n71955 : n71961;
  assign n71963 = pi20 ? n21111 : ~n207;
  assign n71964 = pi19 ? n71963 : n32;
  assign n71965 = pi18 ? n32 : n71964;
  assign n71966 = pi17 ? n32 : n71965;
  assign n71967 = pi16 ? n32 : n71966;
  assign n71968 = pi15 ? n71967 : n13380;
  assign n71969 = pi18 ? n32 : n31340;
  assign n71970 = pi17 ? n32 : n71969;
  assign n71971 = pi16 ? n32 : n71970;
  assign n71972 = pi15 ? n71971 : n13089;
  assign n71973 = pi14 ? n71968 : n71972;
  assign n71974 = pi13 ? n71962 : n71973;
  assign n71975 = pi12 ? n71945 : n71974;
  assign n71976 = pi11 ? n71902 : n71975;
  assign n71977 = pi10 ? n71823 : n71976;
  assign n71978 = pi09 ? n32 : n71977;
  assign n71979 = pi15 ? n65606 : n71515;
  assign n71980 = pi14 ? n71763 : n71979;
  assign n71981 = pi13 ? n32 : n71980;
  assign n71982 = pi12 ? n32 : n71981;
  assign n71983 = pi15 ? n68991 : n70243;
  assign n71984 = pi14 ? n71983 : n71773;
  assign n71985 = pi20 ? n1817 : n749;
  assign n71986 = pi19 ? n32 : ~n71985;
  assign n71987 = pi18 ? n32 : n71986;
  assign n71988 = pi17 ? n32 : n71987;
  assign n71989 = pi16 ? n32 : n71988;
  assign n71990 = pi15 ? n71789 : n71989;
  assign n71991 = pi14 ? n71785 : n71990;
  assign n71992 = pi13 ? n71984 : n71991;
  assign n71993 = pi15 ? n54472 : n24700;
  assign n71994 = pi14 ? n71993 : n71819;
  assign n71995 = pi13 ? n71809 : n71994;
  assign n71996 = pi12 ? n71992 : n71995;
  assign n71997 = pi11 ? n71982 : n71996;
  assign n71998 = pi19 ? n2614 : ~n11561;
  assign n71999 = pi18 ? n32 : n71998;
  assign n72000 = pi17 ? n32 : n71999;
  assign n72001 = pi16 ? n32 : n72000;
  assign n72002 = pi15 ? n71827 : n72001;
  assign n72003 = pi20 ? n15961 : ~n321;
  assign n72004 = pi19 ? n72003 : ~n71835;
  assign n72005 = pi18 ? n32 : n72004;
  assign n72006 = pi17 ? n32 : n72005;
  assign n72007 = pi16 ? n32 : n72006;
  assign n72008 = pi19 ? n37 : n358;
  assign n72009 = pi18 ? n32 : n72008;
  assign n72010 = pi17 ? n32 : n72009;
  assign n72011 = pi16 ? n32 : n72010;
  assign n72012 = pi15 ? n72007 : n72011;
  assign n72013 = pi14 ? n72002 : n72012;
  assign n72014 = pi19 ? n62288 : ~n22911;
  assign n72015 = pi18 ? n32 : n72014;
  assign n72016 = pi17 ? n32 : n72015;
  assign n72017 = pi16 ? n32 : n72016;
  assign n72018 = pi20 ? n36 : ~n246;
  assign n72019 = pi20 ? n41915 : n32;
  assign n72020 = pi19 ? n72018 : n72019;
  assign n72021 = pi18 ? n32 : n72020;
  assign n72022 = pi17 ? n32 : n72021;
  assign n72023 = pi16 ? n32 : n72022;
  assign n72024 = pi15 ? n72017 : n72023;
  assign n72025 = pi20 ? n1377 : n220;
  assign n72026 = pi19 ? n72025 : ~n67800;
  assign n72027 = pi18 ? n32 : n72026;
  assign n72028 = pi17 ? n32 : n72027;
  assign n72029 = pi16 ? n32 : n72028;
  assign n72030 = pi19 ? n342 : n358;
  assign n72031 = pi18 ? n32 : n72030;
  assign n72032 = pi17 ? n32 : n72031;
  assign n72033 = pi16 ? n32 : n72032;
  assign n72034 = pi15 ? n72029 : n72033;
  assign n72035 = pi14 ? n72024 : n72034;
  assign n72036 = pi13 ? n72013 : n72035;
  assign n72037 = pi15 ? n24742 : n71874;
  assign n72038 = pi19 ? n4982 : n19136;
  assign n72039 = pi18 ? n32 : n72038;
  assign n72040 = pi17 ? n32 : n72039;
  assign n72041 = pi16 ? n32 : n72040;
  assign n72042 = pi18 ? n32 : n68203;
  assign n72043 = pi17 ? n32 : n72042;
  assign n72044 = pi16 ? n32 : n72043;
  assign n72045 = pi15 ? n72041 : n72044;
  assign n72046 = pi14 ? n72037 : n72045;
  assign n72047 = pi20 ? n36 : ~n428;
  assign n72048 = pi19 ? n72047 : ~n1941;
  assign n72049 = pi18 ? n32 : n72048;
  assign n72050 = pi17 ? n32 : n72049;
  assign n72051 = pi16 ? n32 : n72050;
  assign n72052 = pi15 ? n13309 : n72051;
  assign n72053 = pi14 ? n71894 : n72052;
  assign n72054 = pi13 ? n72046 : n72053;
  assign n72055 = pi12 ? n72036 : n72054;
  assign n72056 = pi20 ? n15930 : ~n32;
  assign n72057 = pi19 ? n72056 : ~n617;
  assign n72058 = pi18 ? n32 : n72057;
  assign n72059 = pi17 ? n32 : n72058;
  assign n72060 = pi16 ? n32 : n72059;
  assign n72061 = pi19 ? n71144 : ~n1105;
  assign n72062 = pi18 ? n32 : n72061;
  assign n72063 = pi17 ? n32 : n72062;
  assign n72064 = pi16 ? n32 : n72063;
  assign n72065 = pi15 ? n72060 : n72064;
  assign n72066 = pi19 ? n39206 : ~n1105;
  assign n72067 = pi18 ? n32 : n72066;
  assign n72068 = pi17 ? n32 : n72067;
  assign n72069 = pi16 ? n32 : n72068;
  assign n72070 = pi19 ? n46114 : n32;
  assign n72071 = pi18 ? n32 : n72070;
  assign n72072 = pi17 ? n32 : n72071;
  assign n72073 = pi16 ? n32 : n72072;
  assign n72074 = pi15 ? n72069 : n72073;
  assign n72075 = pi14 ? n72065 : n72074;
  assign n72076 = pi19 ? n34907 : n32;
  assign n72077 = pi18 ? n32 : n72076;
  assign n72078 = pi17 ? n32 : n72077;
  assign n72079 = pi16 ? n32 : n72078;
  assign n72080 = pi15 ? n71927 : n72079;
  assign n72081 = pi15 ? n22006 : n14152;
  assign n72082 = pi14 ? n72080 : n72081;
  assign n72083 = pi13 ? n72075 : n72082;
  assign n72084 = pi20 ? n246 : ~n6899;
  assign n72085 = pi19 ? n72084 : n32;
  assign n72086 = pi18 ? n32 : n72085;
  assign n72087 = pi17 ? n32 : n72086;
  assign n72088 = pi16 ? n32 : n72087;
  assign n72089 = pi20 ? n246 : ~n820;
  assign n72090 = pi19 ? n72089 : n32;
  assign n72091 = pi18 ? n32 : n72090;
  assign n72092 = pi17 ? n32 : n72091;
  assign n72093 = pi16 ? n32 : n72092;
  assign n72094 = pi15 ? n72088 : n72093;
  assign n72095 = pi20 ? n62438 : ~n17159;
  assign n72096 = pi19 ? n72095 : n32;
  assign n72097 = pi18 ? n32 : n72096;
  assign n72098 = pi17 ? n32 : n72097;
  assign n72099 = pi16 ? n32 : n72098;
  assign n72100 = pi15 ? n72099 : n13369;
  assign n72101 = pi14 ? n72094 : n72100;
  assign n72102 = pi15 ? n32730 : n13380;
  assign n72103 = pi14 ? n72102 : n13393;
  assign n72104 = pi13 ? n72101 : n72103;
  assign n72105 = pi12 ? n72083 : n72104;
  assign n72106 = pi11 ? n72055 : n72105;
  assign n72107 = pi10 ? n71997 : n72106;
  assign n72108 = pi09 ? n32 : n72107;
  assign n72109 = pi08 ? n71978 : n72108;
  assign n72110 = pi15 ? n65467 : n71515;
  assign n72111 = pi14 ? n71763 : n72110;
  assign n72112 = pi13 ? n32 : n72111;
  assign n72113 = pi12 ? n32 : n72112;
  assign n72114 = pi19 ? n507 : n53115;
  assign n72115 = pi18 ? n32 : n72114;
  assign n72116 = pi17 ? n32 : n72115;
  assign n72117 = pi16 ? n32 : n72116;
  assign n72118 = pi15 ? n72117 : n53119;
  assign n72119 = pi19 ? n32 : ~n13486;
  assign n72120 = pi18 ? n32 : n72119;
  assign n72121 = pi17 ? n32 : n72120;
  assign n72122 = pi16 ? n32 : n72121;
  assign n72123 = pi20 ? n1368 : n749;
  assign n72124 = pi19 ? n32 : ~n72123;
  assign n72125 = pi18 ? n32 : n72124;
  assign n72126 = pi17 ? n32 : n72125;
  assign n72127 = pi16 ? n32 : n72126;
  assign n72128 = pi15 ? n72122 : n72127;
  assign n72129 = pi14 ? n72118 : n72128;
  assign n72130 = pi13 ? n71984 : n72129;
  assign n72131 = pi15 ? n17039 : n71801;
  assign n72132 = pi20 ? n1324 : ~n749;
  assign n72133 = pi19 ? n32 : n72132;
  assign n72134 = pi18 ? n32 : n72133;
  assign n72135 = pi17 ? n32 : n72134;
  assign n72136 = pi16 ? n32 : n72135;
  assign n72137 = pi15 ? n71807 : n72136;
  assign n72138 = pi14 ? n72131 : n72137;
  assign n72139 = pi19 ? n6398 : ~n11546;
  assign n72140 = pi18 ? n32 : n72139;
  assign n72141 = pi17 ? n32 : n72140;
  assign n72142 = pi16 ? n32 : n72141;
  assign n72143 = pi15 ? n54885 : n72142;
  assign n72144 = pi19 ? n2092 : ~n12957;
  assign n72145 = pi18 ? n32 : n72144;
  assign n72146 = pi17 ? n32 : n72145;
  assign n72147 = pi16 ? n32 : n72146;
  assign n72148 = pi20 ? n14286 : n243;
  assign n72149 = pi19 ? n32 : ~n72148;
  assign n72150 = pi18 ? n32 : n72149;
  assign n72151 = pi17 ? n32 : n72150;
  assign n72152 = pi16 ? n32 : n72151;
  assign n72153 = pi15 ? n72147 : n72152;
  assign n72154 = pi14 ? n72143 : n72153;
  assign n72155 = pi13 ? n72138 : n72154;
  assign n72156 = pi12 ? n72130 : n72155;
  assign n72157 = pi11 ? n72113 : n72156;
  assign n72158 = pi19 ? n12578 : n25700;
  assign n72159 = pi18 ? n32 : n72158;
  assign n72160 = pi17 ? n32 : n72159;
  assign n72161 = pi16 ? n32 : n72160;
  assign n72162 = pi19 ? n343 : ~n54797;
  assign n72163 = pi18 ? n32 : n72162;
  assign n72164 = pi17 ? n32 : n72163;
  assign n72165 = pi16 ? n32 : n72164;
  assign n72166 = pi15 ? n72161 : n72165;
  assign n72167 = pi20 ? n16369 : ~n1385;
  assign n72168 = pi19 ? n72167 : ~n589;
  assign n72169 = pi18 ? n32 : n72168;
  assign n72170 = pi17 ? n32 : n72169;
  assign n72171 = pi16 ? n32 : n72170;
  assign n72172 = pi19 ? n52453 : n16969;
  assign n72173 = pi18 ? n32 : n72172;
  assign n72174 = pi17 ? n32 : n72173;
  assign n72175 = pi16 ? n32 : n72174;
  assign n72176 = pi15 ? n72171 : n72175;
  assign n72177 = pi14 ? n72166 : n72176;
  assign n72178 = pi21 ? n259 : n100;
  assign n72179 = pi20 ? n72178 : ~n32;
  assign n72180 = pi19 ? n34159 : ~n72179;
  assign n72181 = pi18 ? n32 : n72180;
  assign n72182 = pi17 ? n32 : n72181;
  assign n72183 = pi16 ? n32 : n72182;
  assign n72184 = pi20 ? n9628 : n7939;
  assign n72185 = pi19 ? n72184 : n15806;
  assign n72186 = pi18 ? n32 : n72185;
  assign n72187 = pi17 ? n32 : n72186;
  assign n72188 = pi16 ? n32 : n72187;
  assign n72189 = pi15 ? n72183 : n72188;
  assign n72190 = pi20 ? n18129 : n354;
  assign n72191 = pi21 ? n1392 : ~n85;
  assign n72192 = pi20 ? n72191 : ~n32;
  assign n72193 = pi19 ? n72190 : ~n72192;
  assign n72194 = pi18 ? n32 : n72193;
  assign n72195 = pi17 ? n32 : n72194;
  assign n72196 = pi16 ? n32 : n72195;
  assign n72197 = pi15 ? n72196 : n32;
  assign n72198 = pi14 ? n72189 : n72197;
  assign n72199 = pi13 ? n72177 : n72198;
  assign n72200 = pi21 ? n2076 : n259;
  assign n72201 = pi20 ? n72200 : ~n32;
  assign n72202 = pi19 ? n32 : ~n72201;
  assign n72203 = pi18 ? n32 : n72202;
  assign n72204 = pi17 ? n32 : n72203;
  assign n72205 = pi16 ? n32 : n72204;
  assign n72206 = pi19 ? n208 : n10662;
  assign n72207 = pi18 ? n32 : n72206;
  assign n72208 = pi17 ? n32 : n72207;
  assign n72209 = pi16 ? n32 : n72208;
  assign n72210 = pi15 ? n72205 : n72209;
  assign n72211 = pi19 ? n531 : ~n6900;
  assign n72212 = pi18 ? n32 : n72211;
  assign n72213 = pi17 ? n32 : n72212;
  assign n72214 = pi16 ? n32 : n72213;
  assign n72215 = pi19 ? n67266 : n5614;
  assign n72216 = pi18 ? n32 : n72215;
  assign n72217 = pi17 ? n32 : n72216;
  assign n72218 = pi16 ? n32 : n72217;
  assign n72219 = pi15 ? n72214 : n72218;
  assign n72220 = pi14 ? n72210 : n72219;
  assign n72221 = pi19 ? n4982 : ~n1941;
  assign n72222 = pi18 ? n32 : n72221;
  assign n72223 = pi17 ? n32 : n72222;
  assign n72224 = pi16 ? n32 : n72223;
  assign n72225 = pi15 ? n71889 : n72224;
  assign n72226 = pi20 ? n9628 : ~n56542;
  assign n72227 = pi19 ? n72226 : ~n617;
  assign n72228 = pi18 ? n32 : n72227;
  assign n72229 = pi17 ? n32 : n72228;
  assign n72230 = pi16 ? n32 : n72229;
  assign n72231 = pi20 ? n653 : n339;
  assign n72232 = pi19 ? n72231 : ~n617;
  assign n72233 = pi18 ? n32 : n72232;
  assign n72234 = pi17 ? n32 : n72233;
  assign n72235 = pi16 ? n32 : n72234;
  assign n72236 = pi15 ? n72230 : n72235;
  assign n72237 = pi14 ? n72225 : n72236;
  assign n72238 = pi13 ? n72220 : n72237;
  assign n72239 = pi12 ? n72199 : n72238;
  assign n72240 = pi19 ? n10148 : ~n1105;
  assign n72241 = pi18 ? n32 : n72240;
  assign n72242 = pi17 ? n32 : n72241;
  assign n72243 = pi16 ? n32 : n72242;
  assign n72244 = pi19 ? n44571 : n32;
  assign n72245 = pi18 ? n32 : n72244;
  assign n72246 = pi17 ? n32 : n72245;
  assign n72247 = pi16 ? n32 : n72246;
  assign n72248 = pi15 ? n72243 : n72247;
  assign n72249 = pi20 ? n321 : ~n7229;
  assign n72250 = pi19 ? n72249 : n32;
  assign n72251 = pi18 ? n32 : n72250;
  assign n72252 = pi17 ? n32 : n72251;
  assign n72253 = pi16 ? n32 : n72252;
  assign n72254 = pi20 ? n321 : n13171;
  assign n72255 = pi19 ? n72254 : n32;
  assign n72256 = pi18 ? n32 : n72255;
  assign n72257 = pi17 ? n32 : n72256;
  assign n72258 = pi16 ? n32 : n72257;
  assign n72259 = pi15 ? n72253 : n72258;
  assign n72260 = pi14 ? n72248 : n72259;
  assign n72261 = pi18 ? n32 : n64943;
  assign n72262 = pi17 ? n32 : n72261;
  assign n72263 = pi16 ? n32 : n72262;
  assign n72264 = pi20 ? n3523 : n20353;
  assign n72265 = pi19 ? n72264 : n32;
  assign n72266 = pi18 ? n32 : n72265;
  assign n72267 = pi17 ? n32 : n72266;
  assign n72268 = pi16 ? n32 : n72267;
  assign n72269 = pi15 ? n72263 : n72268;
  assign n72270 = pi20 ? n974 : n1685;
  assign n72271 = pi19 ? n72270 : n32;
  assign n72272 = pi18 ? n32 : n72271;
  assign n72273 = pi17 ? n32 : n72272;
  assign n72274 = pi16 ? n32 : n72273;
  assign n72275 = pi15 ? n72274 : n21033;
  assign n72276 = pi14 ? n72269 : n72275;
  assign n72277 = pi13 ? n72260 : n72276;
  assign n72278 = pi18 ? n32 : n21808;
  assign n72279 = pi17 ? n32 : n72278;
  assign n72280 = pi16 ? n32 : n72279;
  assign n72281 = pi19 ? n52220 : n32;
  assign n72282 = pi18 ? n32 : n72281;
  assign n72283 = pi17 ? n32 : n72282;
  assign n72284 = pi16 ? n32 : n72283;
  assign n72285 = pi15 ? n72280 : n72284;
  assign n72286 = pi20 ? n13792 : ~n207;
  assign n72287 = pi19 ? n72286 : n32;
  assign n72288 = pi18 ? n32 : n72287;
  assign n72289 = pi17 ? n32 : n72288;
  assign n72290 = pi16 ? n32 : n72289;
  assign n72291 = pi15 ? n72290 : n13671;
  assign n72292 = pi14 ? n72285 : n72291;
  assign n72293 = pi13 ? n72292 : n13686;
  assign n72294 = pi12 ? n72277 : n72293;
  assign n72295 = pi11 ? n72239 : n72294;
  assign n72296 = pi10 ? n72157 : n72295;
  assign n72297 = pi09 ? n32 : n72296;
  assign n72298 = pi19 ? n507 : n70637;
  assign n72299 = pi18 ? n32 : n72298;
  assign n72300 = pi17 ? n32 : n72299;
  assign n72301 = pi16 ? n32 : n72300;
  assign n72302 = pi15 ? n17278 : n72301;
  assign n72303 = pi14 ? n72302 : n72110;
  assign n72304 = pi13 ? n32 : n72303;
  assign n72305 = pi12 ? n32 : n72304;
  assign n72306 = pi15 ? n68991 : n16884;
  assign n72307 = pi14 ? n72306 : n71773;
  assign n72308 = pi15 ? n72117 : n68564;
  assign n72309 = pi19 ? n32 : ~n12425;
  assign n72310 = pi18 ? n32 : n72309;
  assign n72311 = pi17 ? n32 : n72310;
  assign n72312 = pi16 ? n32 : n72311;
  assign n72313 = pi19 ? n32 : ~n9597;
  assign n72314 = pi18 ? n32 : n72313;
  assign n72315 = pi17 ? n32 : n72314;
  assign n72316 = pi16 ? n32 : n72315;
  assign n72317 = pi15 ? n72312 : n72316;
  assign n72318 = pi14 ? n72308 : n72317;
  assign n72319 = pi13 ? n72307 : n72318;
  assign n72320 = pi20 ? n55121 : ~n6229;
  assign n72321 = pi19 ? n322 : ~n72320;
  assign n72322 = pi18 ? n32 : n72321;
  assign n72323 = pi17 ? n32 : n72322;
  assign n72324 = pi16 ? n32 : n72323;
  assign n72325 = pi15 ? n17039 : n72324;
  assign n72326 = pi19 ? n322 : ~n1868;
  assign n72327 = pi18 ? n32 : n72326;
  assign n72328 = pi17 ? n32 : n72327;
  assign n72329 = pi16 ? n32 : n72328;
  assign n72330 = pi20 ? n55121 : ~n243;
  assign n72331 = pi19 ? n32 : n72330;
  assign n72332 = pi18 ? n32 : n72331;
  assign n72333 = pi17 ? n32 : n72332;
  assign n72334 = pi16 ? n32 : n72333;
  assign n72335 = pi15 ? n72329 : n72334;
  assign n72336 = pi14 ? n72325 : n72335;
  assign n72337 = pi15 ? n54472 : n27528;
  assign n72338 = pi19 ? n32 : ~n12957;
  assign n72339 = pi18 ? n32 : n72338;
  assign n72340 = pi17 ? n32 : n72339;
  assign n72341 = pi16 ? n32 : n72340;
  assign n72342 = pi15 ? n72341 : n54636;
  assign n72343 = pi14 ? n72337 : n72342;
  assign n72344 = pi13 ? n72336 : n72343;
  assign n72345 = pi12 ? n72319 : n72344;
  assign n72346 = pi11 ? n72305 : n72345;
  assign n72347 = pi19 ? n343 : ~n11108;
  assign n72348 = pi18 ? n32 : n72347;
  assign n72349 = pi17 ? n32 : n72348;
  assign n72350 = pi16 ? n32 : n72349;
  assign n72351 = pi15 ? n72161 : n72350;
  assign n72352 = pi20 ? n151 : ~n1385;
  assign n72353 = pi19 ? n72352 : ~n589;
  assign n72354 = pi18 ? n32 : n72353;
  assign n72355 = pi17 ? n32 : n72354;
  assign n72356 = pi16 ? n32 : n72355;
  assign n72357 = pi20 ? n151 : n2140;
  assign n72358 = pi19 ? n72357 : n16969;
  assign n72359 = pi18 ? n32 : n72358;
  assign n72360 = pi17 ? n32 : n72359;
  assign n72361 = pi16 ? n32 : n72360;
  assign n72362 = pi15 ? n72356 : n72361;
  assign n72363 = pi14 ? n72351 : n72362;
  assign n72364 = pi20 ? n342 : ~n354;
  assign n72365 = pi19 ? n72364 : ~n72179;
  assign n72366 = pi18 ? n32 : n72365;
  assign n72367 = pi17 ? n32 : n72366;
  assign n72368 = pi16 ? n32 : n72367;
  assign n72369 = pi20 ? n1319 : n50285;
  assign n72370 = pi19 ? n72369 : n10632;
  assign n72371 = pi18 ? n32 : n72370;
  assign n72372 = pi17 ? n32 : n72371;
  assign n72373 = pi16 ? n32 : n72372;
  assign n72374 = pi15 ? n72368 : n72373;
  assign n72375 = pi20 ? n14286 : ~n9013;
  assign n72376 = pi21 ? n309 : n85;
  assign n72377 = pi20 ? n72376 : n32;
  assign n72378 = pi19 ? n72375 : n72377;
  assign n72379 = pi18 ? n32 : n72378;
  assign n72380 = pi17 ? n32 : n72379;
  assign n72381 = pi16 ? n32 : n72380;
  assign n72382 = pi19 ? n472 : n5635;
  assign n72383 = pi18 ? n32 : n72382;
  assign n72384 = pi17 ? n32 : n72383;
  assign n72385 = pi16 ? n32 : n72384;
  assign n72386 = pi15 ? n72381 : n72385;
  assign n72387 = pi14 ? n72374 : n72386;
  assign n72388 = pi13 ? n72363 : n72387;
  assign n72389 = pi15 ? n24511 : n72209;
  assign n72390 = pi14 ? n72389 : n72219;
  assign n72391 = pi20 ? n32 : n12882;
  assign n72392 = pi19 ? n72391 : ~n813;
  assign n72393 = pi18 ? n32 : n72392;
  assign n72394 = pi17 ? n32 : n72393;
  assign n72395 = pi16 ? n32 : n72394;
  assign n72396 = pi19 ? n727 : ~n236;
  assign n72397 = pi18 ? n32 : n72396;
  assign n72398 = pi17 ? n32 : n72397;
  assign n72399 = pi16 ? n32 : n72398;
  assign n72400 = pi15 ? n72395 : n72399;
  assign n72401 = pi20 ? n1319 : ~n18762;
  assign n72402 = pi19 ? n72401 : ~n617;
  assign n72403 = pi18 ? n32 : n72402;
  assign n72404 = pi17 ? n32 : n72403;
  assign n72405 = pi16 ? n32 : n72404;
  assign n72406 = pi19 ? n53777 : ~n617;
  assign n72407 = pi18 ? n32 : n72406;
  assign n72408 = pi17 ? n32 : n72407;
  assign n72409 = pi16 ? n32 : n72408;
  assign n72410 = pi15 ? n72405 : n72409;
  assign n72411 = pi14 ? n72400 : n72410;
  assign n72412 = pi13 ? n72390 : n72411;
  assign n72413 = pi12 ? n72388 : n72412;
  assign n72414 = pi15 ? n13900 : n72247;
  assign n72415 = pi21 ? n124 : ~n51;
  assign n72416 = pi20 ? n342 : ~n72415;
  assign n72417 = pi19 ? n72416 : n32;
  assign n72418 = pi18 ? n32 : n72417;
  assign n72419 = pi17 ? n32 : n72418;
  assign n72420 = pi16 ? n32 : n72419;
  assign n72421 = pi20 ? n342 : ~n16079;
  assign n72422 = pi19 ? n72421 : n32;
  assign n72423 = pi18 ? n32 : n72422;
  assign n72424 = pi17 ? n32 : n72423;
  assign n72425 = pi16 ? n32 : n72424;
  assign n72426 = pi15 ? n72420 : n72425;
  assign n72427 = pi14 ? n72414 : n72426;
  assign n72428 = pi18 ? n32 : n68374;
  assign n72429 = pi17 ? n32 : n72428;
  assign n72430 = pi16 ? n32 : n72429;
  assign n72431 = pi15 ? n72430 : n27328;
  assign n72432 = pi20 ? n428 : ~n2358;
  assign n72433 = pi19 ? n72432 : n32;
  assign n72434 = pi18 ? n32 : n72433;
  assign n72435 = pi17 ? n32 : n72434;
  assign n72436 = pi16 ? n32 : n72435;
  assign n72437 = pi15 ? n72436 : n21033;
  assign n72438 = pi14 ? n72431 : n72437;
  assign n72439 = pi13 ? n72427 : n72438;
  assign n72440 = pi12 ? n72439 : n13955;
  assign n72441 = pi11 ? n72413 : n72440;
  assign n72442 = pi10 ? n72346 : n72441;
  assign n72443 = pi09 ? n32 : n72442;
  assign n72444 = pi08 ? n72297 : n72443;
  assign n72445 = pi07 ? n72109 : n72444;
  assign n72446 = pi06 ? n71758 : n72445;
  assign n72447 = pi05 ? n71181 : n72446;
  assign n72448 = pi04 ? n70066 : n72447;
  assign n72449 = pi13 ? n32 : n51514;
  assign n72450 = pi12 ? n32 : n72449;
  assign n72451 = pi11 ? n32 : n72450;
  assign n72452 = pi10 ? n32 : n72451;
  assign n72453 = pi21 ? n1009 : n1939;
  assign n72454 = pi20 ? n32 : ~n72453;
  assign n72455 = pi19 ? n32 : n72454;
  assign n72456 = pi18 ? n32 : n72455;
  assign n72457 = pi17 ? n32 : n72456;
  assign n72458 = pi16 ? n32 : n72457;
  assign n72459 = pi15 ? n32 : n72458;
  assign n72460 = pi14 ? n17278 : n72459;
  assign n72461 = pi13 ? n32 : n72460;
  assign n72462 = pi12 ? n32 : n72461;
  assign n72463 = pi14 ? n72306 : n38744;
  assign n72464 = pi19 ? n142 : n7795;
  assign n72465 = pi18 ? n32 : n72464;
  assign n72466 = pi17 ? n32 : n72465;
  assign n72467 = pi16 ? n32 : n72466;
  assign n72468 = pi15 ? n53119 : n72467;
  assign n72469 = pi19 ? n275 : ~n7813;
  assign n72470 = pi18 ? n32 : n72469;
  assign n72471 = pi17 ? n32 : n72470;
  assign n72472 = pi16 ? n32 : n72471;
  assign n72473 = pi15 ? n72312 : n72472;
  assign n72474 = pi14 ? n72468 : n72473;
  assign n72475 = pi13 ? n72463 : n72474;
  assign n72476 = pi20 ? n14514 : ~n11048;
  assign n72477 = pi19 ? n4126 : n72476;
  assign n72478 = pi18 ? n32 : n72477;
  assign n72479 = pi17 ? n32 : n72478;
  assign n72480 = pi16 ? n32 : n72479;
  assign n72481 = pi15 ? n17039 : n72480;
  assign n72482 = pi20 ? n14286 : ~n749;
  assign n72483 = pi19 ? n32 : n72482;
  assign n72484 = pi18 ? n32 : n72483;
  assign n72485 = pi17 ? n32 : n72484;
  assign n72486 = pi16 ? n32 : n72485;
  assign n72487 = pi19 ? n4126 : ~n54632;
  assign n72488 = pi18 ? n32 : n72487;
  assign n72489 = pi17 ? n32 : n72488;
  assign n72490 = pi16 ? n32 : n72489;
  assign n72491 = pi15 ? n72486 : n72490;
  assign n72492 = pi14 ? n72481 : n72491;
  assign n72493 = pi19 ? n2386 : ~n13543;
  assign n72494 = pi18 ? n32 : n72493;
  assign n72495 = pi17 ? n32 : n72494;
  assign n72496 = pi16 ? n32 : n72495;
  assign n72497 = pi15 ? n72496 : n15230;
  assign n72498 = pi20 ? n518 : ~n481;
  assign n72499 = pi19 ? n32 : ~n72498;
  assign n72500 = pi18 ? n32 : n72499;
  assign n72501 = pi17 ? n32 : n72500;
  assign n72502 = pi16 ? n32 : n72501;
  assign n72503 = pi15 ? n72502 : n27213;
  assign n72504 = pi14 ? n72497 : n72503;
  assign n72505 = pi13 ? n72492 : n72504;
  assign n72506 = pi12 ? n72475 : n72505;
  assign n72507 = pi11 ? n72462 : n72506;
  assign n72508 = pi19 ? n6622 : n19852;
  assign n72509 = pi18 ? n32 : n72508;
  assign n72510 = pi17 ? n32 : n72509;
  assign n72511 = pi16 ? n32 : n72510;
  assign n72512 = pi19 ? n267 : n3692;
  assign n72513 = pi18 ? n32 : n72512;
  assign n72514 = pi17 ? n32 : n72513;
  assign n72515 = pi16 ? n32 : n72514;
  assign n72516 = pi15 ? n72511 : n72515;
  assign n72517 = pi19 ? n267 : ~n12008;
  assign n72518 = pi18 ? n32 : n72517;
  assign n72519 = pi17 ? n32 : n72518;
  assign n72520 = pi16 ? n32 : n72519;
  assign n72521 = pi15 ? n25584 : n72520;
  assign n72522 = pi14 ? n72516 : n72521;
  assign n72523 = pi15 ? n50949 : n22540;
  assign n72524 = pi19 ? n1348 : ~n58758;
  assign n72525 = pi18 ? n32 : n72524;
  assign n72526 = pi17 ? n32 : n72525;
  assign n72527 = pi16 ? n32 : n72526;
  assign n72528 = pi19 ? n32 : n54724;
  assign n72529 = pi18 ? n32 : n72528;
  assign n72530 = pi17 ? n32 : n72529;
  assign n72531 = pi16 ? n32 : n72530;
  assign n72532 = pi15 ? n72527 : n72531;
  assign n72533 = pi14 ? n72523 : n72532;
  assign n72534 = pi13 ? n72522 : n72533;
  assign n72535 = pi19 ? n267 : ~n40268;
  assign n72536 = pi18 ? n32 : n72535;
  assign n72537 = pi17 ? n32 : n72536;
  assign n72538 = pi16 ? n32 : n72537;
  assign n72539 = pi19 ? n322 : n6230;
  assign n72540 = pi18 ? n32 : n72539;
  assign n72541 = pi17 ? n32 : n72540;
  assign n72542 = pi16 ? n32 : n72541;
  assign n72543 = pi15 ? n72538 : n72542;
  assign n72544 = pi19 ? n261 : ~n821;
  assign n72545 = pi18 ? n32 : n72544;
  assign n72546 = pi17 ? n32 : n72545;
  assign n72547 = pi16 ? n32 : n72546;
  assign n72548 = pi15 ? n72547 : n24838;
  assign n72549 = pi14 ? n72543 : n72548;
  assign n72550 = pi15 ? n14138 : n55015;
  assign n72551 = pi20 ? n101 : n266;
  assign n72552 = pi19 ? n72551 : ~n617;
  assign n72553 = pi18 ? n32 : n72552;
  assign n72554 = pi17 ? n32 : n72553;
  assign n72555 = pi16 ? n32 : n72554;
  assign n72556 = pi19 ? n916 : ~n1105;
  assign n72557 = pi18 ? n32 : n72556;
  assign n72558 = pi17 ? n32 : n72557;
  assign n72559 = pi16 ? n32 : n72558;
  assign n72560 = pi15 ? n72555 : n72559;
  assign n72561 = pi14 ? n72550 : n72560;
  assign n72562 = pi13 ? n72549 : n72561;
  assign n72563 = pi12 ? n72534 : n72562;
  assign n72564 = pi19 ? n804 : n32;
  assign n72565 = pi18 ? n32 : n72564;
  assign n72566 = pi17 ? n32 : n72565;
  assign n72567 = pi16 ? n32 : n72566;
  assign n72568 = pi15 ? n72567 : n21853;
  assign n72569 = pi21 ? n309 : n51;
  assign n72570 = pi20 ? n32 : n72569;
  assign n72571 = pi19 ? n72570 : n32;
  assign n72572 = pi18 ? n32 : n72571;
  assign n72573 = pi17 ? n32 : n72572;
  assign n72574 = pi16 ? n32 : n72573;
  assign n72575 = pi20 ? n32 : ~n9491;
  assign n72576 = pi19 ? n72575 : n32;
  assign n72577 = pi18 ? n32 : n72576;
  assign n72578 = pi17 ? n32 : n72577;
  assign n72579 = pi16 ? n32 : n72578;
  assign n72580 = pi15 ? n72574 : n72579;
  assign n72581 = pi14 ? n72568 : n72580;
  assign n72582 = pi15 ? n32 : n14164;
  assign n72583 = pi14 ? n53575 : n72582;
  assign n72584 = pi13 ? n72581 : n72583;
  assign n72585 = pi12 ? n72584 : n32;
  assign n72586 = pi11 ? n72563 : n72585;
  assign n72587 = pi10 ? n72507 : n72586;
  assign n72588 = pi09 ? n72452 : n72587;
  assign n72589 = pi14 ? n72306 : n17364;
  assign n72590 = pi20 ? n175 : ~n1839;
  assign n72591 = pi19 ? n32 : n72590;
  assign n72592 = pi18 ? n32 : n72591;
  assign n72593 = pi17 ? n32 : n72592;
  assign n72594 = pi16 ? n32 : n72593;
  assign n72595 = pi15 ? n53119 : n72594;
  assign n72596 = pi15 ? n71222 : n72472;
  assign n72597 = pi14 ? n72595 : n72596;
  assign n72598 = pi13 ? n72589 : n72597;
  assign n72599 = pi20 ? n1385 : ~n11048;
  assign n72600 = pi19 ? n4126 : n72599;
  assign n72601 = pi18 ? n32 : n72600;
  assign n72602 = pi17 ? n32 : n72601;
  assign n72603 = pi16 ? n32 : n72602;
  assign n72604 = pi15 ? n16392 : n72603;
  assign n72605 = pi20 ? n151 : ~n749;
  assign n72606 = pi19 ? n126 : n72605;
  assign n72607 = pi18 ? n32 : n72606;
  assign n72608 = pi17 ? n32 : n72607;
  assign n72609 = pi16 ? n32 : n72608;
  assign n72610 = pi15 ? n72609 : n72490;
  assign n72611 = pi14 ? n72604 : n72610;
  assign n72612 = pi19 ? n55055 : ~n343;
  assign n72613 = pi18 ? n32 : n72612;
  assign n72614 = pi17 ? n32 : n72613;
  assign n72615 = pi16 ? n32 : n72614;
  assign n72616 = pi15 ? n72496 : n72615;
  assign n72617 = pi14 ? n72616 : n72503;
  assign n72618 = pi13 ? n72611 : n72617;
  assign n72619 = pi12 ? n72598 : n72618;
  assign n72620 = pi11 ? n72462 : n72619;
  assign n72621 = pi19 ? n267 : n19852;
  assign n72622 = pi18 ? n32 : n72621;
  assign n72623 = pi17 ? n32 : n72622;
  assign n72624 = pi16 ? n32 : n72623;
  assign n72625 = pi15 ? n72624 : n72515;
  assign n72626 = pi19 ? n1440 : ~n12008;
  assign n72627 = pi18 ? n32 : n72626;
  assign n72628 = pi17 ? n32 : n72627;
  assign n72629 = pi16 ? n32 : n72628;
  assign n72630 = pi15 ? n24582 : n72629;
  assign n72631 = pi14 ? n72625 : n72630;
  assign n72632 = pi20 ? n32 : n17134;
  assign n72633 = pi19 ? n72632 : n32;
  assign n72634 = pi18 ? n32 : n72633;
  assign n72635 = pi17 ? n32 : n72634;
  assign n72636 = pi16 ? n32 : n72635;
  assign n72637 = pi15 ? n50949 : n72636;
  assign n72638 = pi19 ? n340 : ~n58758;
  assign n72639 = pi18 ? n32 : n72638;
  assign n72640 = pi17 ? n32 : n72639;
  assign n72641 = pi16 ? n32 : n72640;
  assign n72642 = pi19 ? n32 : n29950;
  assign n72643 = pi18 ? n32 : n72642;
  assign n72644 = pi17 ? n32 : n72643;
  assign n72645 = pi16 ? n32 : n72644;
  assign n72646 = pi15 ? n72641 : n72645;
  assign n72647 = pi14 ? n72637 : n72646;
  assign n72648 = pi13 ? n72631 : n72647;
  assign n72649 = pi15 ? n40281 : n22437;
  assign n72650 = pi19 ? n267 : ~n617;
  assign n72651 = pi18 ? n32 : n72650;
  assign n72652 = pi17 ? n32 : n72651;
  assign n72653 = pi16 ? n32 : n72652;
  assign n72654 = pi19 ? n72391 : n32;
  assign n72655 = pi18 ? n32 : n72654;
  assign n72656 = pi17 ? n32 : n72655;
  assign n72657 = pi16 ? n32 : n72656;
  assign n72658 = pi15 ? n72653 : n72657;
  assign n72659 = pi14 ? n72649 : n72658;
  assign n72660 = pi13 ? n72549 : n72659;
  assign n72661 = pi12 ? n72648 : n72660;
  assign n72662 = pi15 ? n14373 : n21853;
  assign n72663 = pi18 ? n32 : n22554;
  assign n72664 = pi17 ? n32 : n72663;
  assign n72665 = pi16 ? n32 : n72664;
  assign n72666 = pi15 ? n648 : n72665;
  assign n72667 = pi14 ? n72662 : n72666;
  assign n72668 = pi15 ? n32 : n14405;
  assign n72669 = pi14 ? n53575 : n72668;
  assign n72670 = pi13 ? n72667 : n72669;
  assign n72671 = pi12 ? n72670 : n32;
  assign n72672 = pi11 ? n72661 : n72671;
  assign n72673 = pi10 ? n72620 : n72672;
  assign n72674 = pi09 ? n72452 : n72673;
  assign n72675 = pi08 ? n72588 : n72674;
  assign n72676 = pi15 ? n32 : n17193;
  assign n72677 = pi14 ? n17278 : n72676;
  assign n72678 = pi13 ? n32 : n72677;
  assign n72679 = pi12 ? n32 : n72678;
  assign n72680 = pi15 ? n17363 : n26269;
  assign n72681 = pi14 ? n72306 : n72680;
  assign n72682 = pi19 ? n6398 : n7795;
  assign n72683 = pi18 ? n32 : n72682;
  assign n72684 = pi17 ? n32 : n72683;
  assign n72685 = pi16 ? n32 : n72684;
  assign n72686 = pi15 ? n53963 : n72685;
  assign n72687 = pi19 ? n32 : ~n7813;
  assign n72688 = pi18 ? n32 : n72687;
  assign n72689 = pi17 ? n32 : n72688;
  assign n72690 = pi16 ? n32 : n72689;
  assign n72691 = pi15 ? n71673 : n72690;
  assign n72692 = pi14 ? n72686 : n72691;
  assign n72693 = pi13 ? n72681 : n72692;
  assign n72694 = pi20 ? n246 : ~n1475;
  assign n72695 = pi19 ? n507 : n72694;
  assign n72696 = pi18 ? n32 : n72695;
  assign n72697 = pi17 ? n32 : n72696;
  assign n72698 = pi16 ? n32 : n72697;
  assign n72699 = pi15 ? n25988 : n72698;
  assign n72700 = pi20 ? n1319 : ~n749;
  assign n72701 = pi19 ? n32 : n72700;
  assign n72702 = pi18 ? n32 : n72701;
  assign n72703 = pi17 ? n32 : n72702;
  assign n72704 = pi16 ? n32 : n72703;
  assign n72705 = pi19 ? n507 : ~n54632;
  assign n72706 = pi18 ? n32 : n72705;
  assign n72707 = pi17 ? n32 : n72706;
  assign n72708 = pi16 ? n32 : n72707;
  assign n72709 = pi15 ? n72704 : n72708;
  assign n72710 = pi14 ? n72699 : n72709;
  assign n72711 = pi19 ? n1165 : ~n1265;
  assign n72712 = pi18 ? n32 : n72711;
  assign n72713 = pi17 ? n32 : n72712;
  assign n72714 = pi16 ? n32 : n72713;
  assign n72715 = pi20 ? n32 : n39935;
  assign n72716 = pi19 ? n72715 : ~n12435;
  assign n72717 = pi18 ? n32 : n72716;
  assign n72718 = pi17 ? n32 : n72717;
  assign n72719 = pi16 ? n32 : n72718;
  assign n72720 = pi15 ? n72714 : n72719;
  assign n72721 = pi19 ? n32 : ~n15051;
  assign n72722 = pi18 ? n32 : n72721;
  assign n72723 = pi17 ? n32 : n72722;
  assign n72724 = pi16 ? n32 : n72723;
  assign n72725 = pi19 ? n1818 : ~n53777;
  assign n72726 = pi18 ? n32 : n72725;
  assign n72727 = pi17 ? n32 : n72726;
  assign n72728 = pi16 ? n32 : n72727;
  assign n72729 = pi15 ? n72724 : n72728;
  assign n72730 = pi14 ? n72720 : n72729;
  assign n72731 = pi13 ? n72710 : n72730;
  assign n72732 = pi12 ? n72693 : n72731;
  assign n72733 = pi11 ? n72679 : n72732;
  assign n72734 = pi21 ? n7659 : ~n174;
  assign n72735 = pi20 ? n32 : n72734;
  assign n72736 = pi22 ? n34 : n84;
  assign n72737 = pi21 ? n32 : n72736;
  assign n72738 = pi20 ? n72737 : n32;
  assign n72739 = pi19 ? n72735 : n72738;
  assign n72740 = pi18 ? n32 : n72739;
  assign n72741 = pi17 ? n32 : n72740;
  assign n72742 = pi16 ? n32 : n72741;
  assign n72743 = pi21 ? n242 : n173;
  assign n72744 = pi20 ? n32 : n72743;
  assign n72745 = pi19 ? n72744 : n10645;
  assign n72746 = pi18 ? n32 : n72745;
  assign n72747 = pi17 ? n32 : n72746;
  assign n72748 = pi16 ? n32 : n72747;
  assign n72749 = pi15 ? n72742 : n72748;
  assign n72750 = pi19 ? n857 : n7661;
  assign n72751 = pi18 ? n32 : n72750;
  assign n72752 = pi17 ? n32 : n72751;
  assign n72753 = pi16 ? n32 : n72752;
  assign n72754 = pi19 ? n9220 : ~n589;
  assign n72755 = pi18 ? n32 : n72754;
  assign n72756 = pi17 ? n32 : n72755;
  assign n72757 = pi16 ? n32 : n72756;
  assign n72758 = pi15 ? n72753 : n72757;
  assign n72759 = pi14 ? n72749 : n72758;
  assign n72760 = pi19 ? n18741 : n152;
  assign n72761 = pi18 ? n32 : n72760;
  assign n72762 = pi17 ? n32 : n72761;
  assign n72763 = pi16 ? n32 : n72762;
  assign n72764 = pi19 ? n519 : n3495;
  assign n72765 = pi18 ? n32 : n72764;
  assign n72766 = pi17 ? n32 : n72765;
  assign n72767 = pi16 ? n32 : n72766;
  assign n72768 = pi15 ? n72763 : n72767;
  assign n72769 = pi19 ? n4518 : ~n589;
  assign n72770 = pi18 ? n32 : n72769;
  assign n72771 = pi17 ? n32 : n72770;
  assign n72772 = pi16 ? n32 : n72771;
  assign n72773 = pi15 ? n72772 : n23484;
  assign n72774 = pi14 ? n72768 : n72773;
  assign n72775 = pi13 ? n72759 : n72774;
  assign n72776 = pi19 ? n1325 : n5614;
  assign n72777 = pi18 ? n32 : n72776;
  assign n72778 = pi17 ? n32 : n72777;
  assign n72779 = pi16 ? n32 : n72778;
  assign n72780 = pi19 ? n25184 : n19892;
  assign n72781 = pi18 ? n32 : n72780;
  assign n72782 = pi17 ? n32 : n72781;
  assign n72783 = pi16 ? n32 : n72782;
  assign n72784 = pi15 ? n72779 : n72783;
  assign n72785 = pi19 ? n19582 : ~n1941;
  assign n72786 = pi18 ? n32 : n72785;
  assign n72787 = pi17 ? n32 : n72786;
  assign n72788 = pi16 ? n32 : n72787;
  assign n72789 = pi15 ? n24167 : n72788;
  assign n72790 = pi14 ? n72784 : n72789;
  assign n72791 = pi19 ? n792 : n32;
  assign n72792 = pi18 ? n32 : n72791;
  assign n72793 = pi17 ? n32 : n72792;
  assign n72794 = pi16 ? n32 : n72793;
  assign n72795 = pi15 ? n72794 : n37312;
  assign n72796 = pi19 ? n47981 : ~n617;
  assign n72797 = pi18 ? n32 : n72796;
  assign n72798 = pi17 ? n32 : n72797;
  assign n72799 = pi16 ? n32 : n72798;
  assign n72800 = pi21 ? n66 : n405;
  assign n72801 = pi20 ? n32 : n72800;
  assign n72802 = pi19 ? n72801 : n32;
  assign n72803 = pi18 ? n32 : n72802;
  assign n72804 = pi17 ? n32 : n72803;
  assign n72805 = pi16 ? n32 : n72804;
  assign n72806 = pi15 ? n72799 : n72805;
  assign n72807 = pi14 ? n72795 : n72806;
  assign n72808 = pi13 ? n72790 : n72807;
  assign n72809 = pi12 ? n72775 : n72808;
  assign n72810 = pi15 ? n22437 : n26498;
  assign n72811 = pi15 ? n26672 : n32;
  assign n72812 = pi14 ? n72810 : n72811;
  assign n72813 = pi14 ? n659 : n21131;
  assign n72814 = pi13 ? n72812 : n72813;
  assign n72815 = pi12 ? n72814 : n32;
  assign n72816 = pi11 ? n72809 : n72815;
  assign n72817 = pi10 ? n72733 : n72816;
  assign n72818 = pi09 ? n72452 : n72817;
  assign n72819 = pi15 ? n16850 : n26269;
  assign n72820 = pi14 ? n72306 : n72819;
  assign n72821 = pi20 ? n3523 : ~n1839;
  assign n72822 = pi19 ? n6398 : n72821;
  assign n72823 = pi18 ? n32 : n72822;
  assign n72824 = pi17 ? n32 : n72823;
  assign n72825 = pi16 ? n32 : n72824;
  assign n72826 = pi15 ? n53963 : n72825;
  assign n72827 = pi19 ? n472 : ~n1476;
  assign n72828 = pi18 ? n32 : n72827;
  assign n72829 = pi17 ? n32 : n72828;
  assign n72830 = pi16 ? n32 : n72829;
  assign n72831 = pi15 ? n72830 : n72690;
  assign n72832 = pi14 ? n72826 : n72831;
  assign n72833 = pi13 ? n72820 : n72832;
  assign n72834 = pi20 ? n1817 : n6229;
  assign n72835 = pi19 ? n32 : n72834;
  assign n72836 = pi18 ? n32 : n72835;
  assign n72837 = pi17 ? n32 : n72836;
  assign n72838 = pi16 ? n32 : n72837;
  assign n72839 = pi15 ? n72838 : n72698;
  assign n72840 = pi20 ? n8661 : n243;
  assign n72841 = pi19 ? n507 : ~n72840;
  assign n72842 = pi18 ? n32 : n72841;
  assign n72843 = pi17 ? n32 : n72842;
  assign n72844 = pi16 ? n32 : n72843;
  assign n72845 = pi15 ? n72704 : n72844;
  assign n72846 = pi14 ? n72839 : n72845;
  assign n72847 = pi19 ? n507 : ~n14065;
  assign n72848 = pi18 ? n32 : n72847;
  assign n72849 = pi17 ? n32 : n72848;
  assign n72850 = pi16 ? n32 : n72849;
  assign n72851 = pi15 ? n15230 : n72850;
  assign n72852 = pi19 ? n32 : ~n14496;
  assign n72853 = pi18 ? n32 : n72852;
  assign n72854 = pi17 ? n32 : n72853;
  assign n72855 = pi16 ? n32 : n72854;
  assign n72856 = pi18 ? n32 : n44698;
  assign n72857 = pi17 ? n32 : n72856;
  assign n72858 = pi16 ? n32 : n72857;
  assign n72859 = pi15 ? n72855 : n72858;
  assign n72860 = pi14 ? n72851 : n72859;
  assign n72861 = pi13 ? n72846 : n72860;
  assign n72862 = pi12 ? n72833 : n72861;
  assign n72863 = pi11 ? n72679 : n72862;
  assign n72864 = pi19 ? n55204 : n152;
  assign n72865 = pi18 ? n32 : n72864;
  assign n72866 = pi17 ? n32 : n72865;
  assign n72867 = pi16 ? n32 : n72866;
  assign n72868 = pi19 ? n792 : n13085;
  assign n72869 = pi18 ? n32 : n72868;
  assign n72870 = pi17 ? n32 : n72869;
  assign n72871 = pi16 ? n32 : n72870;
  assign n72872 = pi15 ? n72867 : n72871;
  assign n72873 = pi21 ? n206 : ~n34;
  assign n72874 = pi20 ? n72873 : n32;
  assign n72875 = pi19 ? n857 : n72874;
  assign n72876 = pi18 ? n32 : n72875;
  assign n72877 = pi17 ? n32 : n72876;
  assign n72878 = pi16 ? n32 : n72877;
  assign n72879 = pi20 ? n23122 : ~n32;
  assign n72880 = pi19 ? n67679 : ~n72879;
  assign n72881 = pi18 ? n32 : n72880;
  assign n72882 = pi17 ? n32 : n72881;
  assign n72883 = pi16 ? n32 : n72882;
  assign n72884 = pi15 ? n72878 : n72883;
  assign n72885 = pi14 ? n72872 : n72884;
  assign n72886 = pi21 ? n14399 : ~n66;
  assign n72887 = pi20 ? n32 : n72886;
  assign n72888 = pi19 ? n72887 : n9169;
  assign n72889 = pi18 ? n32 : n72888;
  assign n72890 = pi17 ? n32 : n72889;
  assign n72891 = pi16 ? n32 : n72890;
  assign n72892 = pi19 ? n2141 : n19317;
  assign n72893 = pi18 ? n32 : n72892;
  assign n72894 = pi17 ? n32 : n72893;
  assign n72895 = pi16 ? n32 : n72894;
  assign n72896 = pi15 ? n72891 : n72895;
  assign n72897 = pi15 ? n72772 : n25888;
  assign n72898 = pi14 ? n72896 : n72897;
  assign n72899 = pi13 ? n72885 : n72898;
  assign n72900 = pi19 ? n54584 : n7488;
  assign n72901 = pi18 ? n32 : n72900;
  assign n72902 = pi17 ? n32 : n72901;
  assign n72903 = pi16 ? n32 : n72902;
  assign n72904 = pi15 ? n72903 : n72783;
  assign n72905 = pi19 ? n14602 : ~n1941;
  assign n72906 = pi18 ? n32 : n72905;
  assign n72907 = pi17 ? n32 : n72906;
  assign n72908 = pi16 ? n32 : n72907;
  assign n72909 = pi19 ? n14937 : ~n2614;
  assign n72910 = pi18 ? n32 : n72909;
  assign n72911 = pi17 ? n32 : n72910;
  assign n72912 = pi16 ? n32 : n72911;
  assign n72913 = pi15 ? n72908 : n72912;
  assign n72914 = pi14 ? n72904 : n72913;
  assign n72915 = pi15 ? n54026 : n37429;
  assign n72916 = pi21 ? n100 : ~n66;
  assign n72917 = pi20 ? n32 : n72916;
  assign n72918 = pi19 ? n72917 : ~n617;
  assign n72919 = pi18 ? n32 : n72918;
  assign n72920 = pi17 ? n32 : n72919;
  assign n72921 = pi16 ? n32 : n72920;
  assign n72922 = pi15 ? n72921 : n54026;
  assign n72923 = pi14 ? n72915 : n72922;
  assign n72924 = pi13 ? n72914 : n72923;
  assign n72925 = pi12 ? n72899 : n72924;
  assign n72926 = pi20 ? n32 : n39764;
  assign n72927 = pi19 ? n72926 : n32;
  assign n72928 = pi18 ? n32 : n72927;
  assign n72929 = pi17 ? n32 : n72928;
  assign n72930 = pi16 ? n32 : n72929;
  assign n72931 = pi15 ? n72930 : n14790;
  assign n72932 = pi14 ? n72931 : n14799;
  assign n72933 = pi13 ? n72932 : n32;
  assign n72934 = pi12 ? n72933 : n32;
  assign n72935 = pi11 ? n72925 : n72934;
  assign n72936 = pi10 ? n72863 : n72935;
  assign n72937 = pi09 ? n72452 : n72936;
  assign n72938 = pi08 ? n72818 : n72937;
  assign n72939 = pi07 ? n72675 : n72938;
  assign n72940 = pi14 ? n25818 : n32;
  assign n72941 = pi13 ? n72940 : n32;
  assign n72942 = pi14 ? n15848 : n32;
  assign n72943 = pi19 ? n32 : n13622;
  assign n72944 = pi18 ? n32 : n72943;
  assign n72945 = pi17 ? n32 : n72944;
  assign n72946 = pi16 ? n32 : n72945;
  assign n72947 = pi15 ? n32 : n72946;
  assign n72948 = pi14 ? n40412 : n72947;
  assign n72949 = pi13 ? n72942 : n72948;
  assign n72950 = pi12 ? n72941 : n72949;
  assign n72951 = pi15 ? n69136 : n17363;
  assign n72952 = pi19 ? n32 : ~n13529;
  assign n72953 = pi18 ? n32 : n72952;
  assign n72954 = pi17 ? n32 : n72953;
  assign n72955 = pi16 ? n32 : n72954;
  assign n72956 = pi15 ? n25763 : n72955;
  assign n72957 = pi14 ? n72951 : n72956;
  assign n72958 = pi20 ? n266 : ~n518;
  assign n72959 = pi19 ? n32 : n72958;
  assign n72960 = pi18 ? n32 : n72959;
  assign n72961 = pi17 ? n32 : n72960;
  assign n72962 = pi16 ? n32 : n72961;
  assign n72963 = pi19 ? n507 : n17752;
  assign n72964 = pi18 ? n32 : n72963;
  assign n72965 = pi17 ? n32 : n72964;
  assign n72966 = pi16 ? n32 : n72965;
  assign n72967 = pi15 ? n72962 : n72966;
  assign n72968 = pi19 ? n507 : n70078;
  assign n72969 = pi18 ? n32 : n72968;
  assign n72970 = pi17 ? n32 : n72969;
  assign n72971 = pi16 ? n32 : n72970;
  assign n72972 = pi19 ? n32 : n48082;
  assign n72973 = pi18 ? n32 : n72972;
  assign n72974 = pi17 ? n32 : n72973;
  assign n72975 = pi16 ? n32 : n72974;
  assign n72976 = pi15 ? n72971 : n72975;
  assign n72977 = pi14 ? n72967 : n72976;
  assign n72978 = pi13 ? n72957 : n72977;
  assign n72979 = pi19 ? n519 : ~n1476;
  assign n72980 = pi18 ? n32 : n72979;
  assign n72981 = pi17 ? n32 : n72980;
  assign n72982 = pi16 ? n32 : n72981;
  assign n72983 = pi15 ? n17216 : n72982;
  assign n72984 = pi19 ? n519 : n41918;
  assign n72985 = pi18 ? n32 : n72984;
  assign n72986 = pi17 ? n32 : n72985;
  assign n72987 = pi16 ? n32 : n72986;
  assign n72988 = pi19 ? n507 : ~n55276;
  assign n72989 = pi18 ? n32 : n72988;
  assign n72990 = pi17 ? n32 : n72989;
  assign n72991 = pi16 ? n32 : n72990;
  assign n72992 = pi15 ? n72987 : n72991;
  assign n72993 = pi14 ? n72983 : n72992;
  assign n72994 = pi19 ? n32 : ~n340;
  assign n72995 = pi18 ? n32 : n72994;
  assign n72996 = pi17 ? n32 : n72995;
  assign n72997 = pi16 ? n32 : n72996;
  assign n72998 = pi19 ? n519 : ~n14065;
  assign n72999 = pi18 ? n32 : n72998;
  assign n73000 = pi17 ? n32 : n72999;
  assign n73001 = pi16 ? n32 : n73000;
  assign n73002 = pi15 ? n72997 : n73001;
  assign n73003 = pi19 ? n507 : n21042;
  assign n73004 = pi18 ? n32 : n73003;
  assign n73005 = pi17 ? n32 : n73004;
  assign n73006 = pi16 ? n32 : n73005;
  assign n73007 = pi15 ? n73006 : n16392;
  assign n73008 = pi14 ? n73002 : n73007;
  assign n73009 = pi13 ? n72993 : n73008;
  assign n73010 = pi12 ? n72978 : n73009;
  assign n73011 = pi11 ? n72950 : n73010;
  assign n73012 = pi19 ? n6398 : ~n4406;
  assign n73013 = pi18 ? n32 : n73012;
  assign n73014 = pi17 ? n32 : n73013;
  assign n73015 = pi16 ? n32 : n73014;
  assign n73016 = pi19 ? n1165 : n39565;
  assign n73017 = pi18 ? n32 : n73016;
  assign n73018 = pi17 ? n32 : n73017;
  assign n73019 = pi16 ? n32 : n73018;
  assign n73020 = pi15 ? n73015 : n73019;
  assign n73021 = pi19 ? n1165 : n176;
  assign n73022 = pi18 ? n32 : n73021;
  assign n73023 = pi17 ? n32 : n73022;
  assign n73024 = pi16 ? n32 : n73023;
  assign n73025 = pi15 ? n73024 : n73015;
  assign n73026 = pi14 ? n73020 : n73025;
  assign n73027 = pi19 ? n14969 : n3692;
  assign n73028 = pi18 ? n32 : n73027;
  assign n73029 = pi17 ? n32 : n73028;
  assign n73030 = pi16 ? n32 : n73029;
  assign n73031 = pi15 ? n73030 : n72895;
  assign n73032 = pi19 ? n55229 : ~n589;
  assign n73033 = pi18 ? n32 : n73032;
  assign n73034 = pi17 ? n32 : n73033;
  assign n73035 = pi16 ? n32 : n73034;
  assign n73036 = pi19 ? n14786 : ~n236;
  assign n73037 = pi18 ? n32 : n73036;
  assign n73038 = pi17 ? n32 : n73037;
  assign n73039 = pi16 ? n32 : n73038;
  assign n73040 = pi15 ? n73035 : n73039;
  assign n73041 = pi14 ? n73031 : n73040;
  assign n73042 = pi13 ? n73026 : n73041;
  assign n73043 = pi19 ? n53174 : ~n1812;
  assign n73044 = pi18 ? n32 : n73043;
  assign n73045 = pi17 ? n32 : n73044;
  assign n73046 = pi16 ? n32 : n73045;
  assign n73047 = pi19 ? n40454 : ~n1812;
  assign n73048 = pi18 ? n32 : n73047;
  assign n73049 = pi17 ? n32 : n73048;
  assign n73050 = pi16 ? n32 : n73049;
  assign n73051 = pi15 ? n73046 : n73050;
  assign n73052 = pi19 ? n1840 : n5626;
  assign n73053 = pi18 ? n32 : n73052;
  assign n73054 = pi17 ? n32 : n73053;
  assign n73055 = pi16 ? n32 : n73054;
  assign n73056 = pi15 ? n14941 : n73055;
  assign n73057 = pi14 ? n73051 : n73056;
  assign n73058 = pi15 ? n39582 : n14958;
  assign n73059 = pi14 ? n15119 : n73058;
  assign n73060 = pi13 ? n73057 : n73059;
  assign n73061 = pi12 ? n73042 : n73060;
  assign n73062 = pi14 ? n22637 : n14975;
  assign n73063 = pi13 ? n73062 : n32;
  assign n73064 = pi12 ? n73063 : n32;
  assign n73065 = pi11 ? n73061 : n73064;
  assign n73066 = pi10 ? n73011 : n73065;
  assign n73067 = pi09 ? n72452 : n73066;
  assign n73068 = pi14 ? n17279 : n72947;
  assign n73069 = pi13 ? n72942 : n73068;
  assign n73070 = pi12 ? n72941 : n73069;
  assign n73071 = pi15 ? n16832 : n72955;
  assign n73072 = pi14 ? n72951 : n73071;
  assign n73073 = pi19 ? n519 : n70078;
  assign n73074 = pi18 ? n32 : n73073;
  assign n73075 = pi17 ? n32 : n73074;
  assign n73076 = pi16 ? n32 : n73075;
  assign n73077 = pi19 ? n6398 : n48082;
  assign n73078 = pi18 ? n32 : n73077;
  assign n73079 = pi17 ? n32 : n73078;
  assign n73080 = pi16 ? n32 : n73079;
  assign n73081 = pi15 ? n73076 : n73080;
  assign n73082 = pi14 ? n72967 : n73081;
  assign n73083 = pi13 ? n73072 : n73082;
  assign n73084 = pi19 ? n519 : n38221;
  assign n73085 = pi18 ? n32 : n73084;
  assign n73086 = pi17 ? n32 : n73085;
  assign n73087 = pi16 ? n32 : n73086;
  assign n73088 = pi19 ? n11183 : ~n55331;
  assign n73089 = pi18 ? n32 : n73088;
  assign n73090 = pi17 ? n32 : n73089;
  assign n73091 = pi16 ? n32 : n73090;
  assign n73092 = pi15 ? n73087 : n73091;
  assign n73093 = pi14 ? n72983 : n73092;
  assign n73094 = pi15 ? n67470 : n73001;
  assign n73095 = pi19 ? n507 : n7642;
  assign n73096 = pi18 ? n32 : n73095;
  assign n73097 = pi17 ? n32 : n73096;
  assign n73098 = pi16 ? n32 : n73097;
  assign n73099 = pi15 ? n73098 : n16392;
  assign n73100 = pi14 ? n73094 : n73099;
  assign n73101 = pi13 ? n73093 : n73100;
  assign n73102 = pi12 ? n73083 : n73101;
  assign n73103 = pi11 ? n73070 : n73102;
  assign n73104 = pi20 ? n63326 : ~n32;
  assign n73105 = pi19 ? n6398 : ~n73104;
  assign n73106 = pi18 ? n32 : n73105;
  assign n73107 = pi17 ? n32 : n73106;
  assign n73108 = pi16 ? n32 : n73107;
  assign n73109 = pi15 ? n73108 : n37468;
  assign n73110 = pi15 ? n22817 : n73015;
  assign n73111 = pi14 ? n73109 : n73110;
  assign n73112 = pi19 ? n6398 : n3692;
  assign n73113 = pi18 ? n32 : n73112;
  assign n73114 = pi17 ? n32 : n73113;
  assign n73115 = pi16 ? n32 : n73114;
  assign n73116 = pi15 ? n73115 : n55403;
  assign n73117 = pi19 ? n2141 : ~n57152;
  assign n73118 = pi18 ? n32 : n73117;
  assign n73119 = pi17 ? n32 : n73118;
  assign n73120 = pi16 ? n32 : n73119;
  assign n73121 = pi19 ? n6398 : ~n20022;
  assign n73122 = pi18 ? n32 : n73121;
  assign n73123 = pi17 ? n32 : n73122;
  assign n73124 = pi16 ? n32 : n73123;
  assign n73125 = pi15 ? n73120 : n73124;
  assign n73126 = pi14 ? n73116 : n73125;
  assign n73127 = pi13 ? n73111 : n73126;
  assign n73128 = pi19 ? n1840 : ~n1812;
  assign n73129 = pi18 ? n32 : n73128;
  assign n73130 = pi17 ? n32 : n73129;
  assign n73131 = pi16 ? n32 : n73130;
  assign n73132 = pi15 ? n73131 : n15248;
  assign n73133 = pi19 ? n975 : ~n1941;
  assign n73134 = pi18 ? n32 : n73133;
  assign n73135 = pi17 ? n32 : n73134;
  assign n73136 = pi16 ? n32 : n73135;
  assign n73137 = pi19 ? n975 : n5626;
  assign n73138 = pi18 ? n32 : n73137;
  assign n73139 = pi17 ? n32 : n73138;
  assign n73140 = pi16 ? n32 : n73139;
  assign n73141 = pi15 ? n73136 : n73140;
  assign n73142 = pi14 ? n73132 : n73141;
  assign n73143 = pi14 ? n15120 : n22252;
  assign n73144 = pi13 ? n73142 : n73143;
  assign n73145 = pi12 ? n73127 : n73144;
  assign n73146 = pi11 ? n73145 : n15130;
  assign n73147 = pi10 ? n73103 : n73146;
  assign n73148 = pi09 ? n72452 : n73147;
  assign n73149 = pi08 ? n73067 : n73148;
  assign n73150 = pi15 ? n15927 : n32;
  assign n73151 = pi14 ? n73150 : n32;
  assign n73152 = pi13 ? n73151 : n32;
  assign n73153 = pi14 ? n15848 : n22205;
  assign n73154 = pi13 ? n73153 : n73068;
  assign n73155 = pi12 ? n73152 : n73154;
  assign n73156 = pi15 ? n68990 : n16850;
  assign n73157 = pi19 ? n594 : ~n13529;
  assign n73158 = pi18 ? n32 : n73157;
  assign n73159 = pi17 ? n32 : n73158;
  assign n73160 = pi16 ? n32 : n73159;
  assign n73161 = pi15 ? n16832 : n73160;
  assign n73162 = pi14 ? n73156 : n73161;
  assign n73163 = pi18 ? n32 : n28126;
  assign n73164 = pi17 ? n32 : n73163;
  assign n73165 = pi16 ? n32 : n73164;
  assign n73166 = pi15 ? n72962 : n73165;
  assign n73167 = pi15 ? n15847 : n51565;
  assign n73168 = pi14 ? n73166 : n73167;
  assign n73169 = pi13 ? n73162 : n73168;
  assign n73170 = pi15 ? n17216 : n71673;
  assign n73171 = pi19 ? n472 : n9007;
  assign n73172 = pi18 ? n32 : n73171;
  assign n73173 = pi17 ? n32 : n73172;
  assign n73174 = pi16 ? n32 : n73173;
  assign n73175 = pi15 ? n73174 : n55390;
  assign n73176 = pi14 ? n73170 : n73175;
  assign n73177 = pi19 ? n507 : ~n244;
  assign n73178 = pi18 ? n32 : n73177;
  assign n73179 = pi17 ? n32 : n73178;
  assign n73180 = pi16 ? n32 : n73179;
  assign n73181 = pi15 ? n67470 : n73180;
  assign n73182 = pi19 ? n1320 : n4670;
  assign n73183 = pi18 ? n32 : n73182;
  assign n73184 = pi17 ? n32 : n73183;
  assign n73185 = pi16 ? n32 : n73184;
  assign n73186 = pi15 ? n73185 : n17039;
  assign n73187 = pi14 ? n73181 : n73186;
  assign n73188 = pi13 ? n73176 : n73187;
  assign n73189 = pi12 ? n73169 : n73188;
  assign n73190 = pi11 ? n73155 : n73189;
  assign n73191 = pi19 ? n507 : n70131;
  assign n73192 = pi18 ? n32 : n73191;
  assign n73193 = pi17 ? n32 : n73192;
  assign n73194 = pi16 ? n32 : n73193;
  assign n73195 = pi15 ? n50638 : n73194;
  assign n73196 = pi14 ? n73195 : n24563;
  assign n73197 = pi19 ? n1785 : n3495;
  assign n73198 = pi18 ? n32 : n73197;
  assign n73199 = pi17 ? n32 : n73198;
  assign n73200 = pi16 ? n32 : n73199;
  assign n73201 = pi15 ? n25050 : n73200;
  assign n73202 = pi15 ? n15244 : n26717;
  assign n73203 = pi14 ? n73201 : n73202;
  assign n73204 = pi13 ? n73196 : n73203;
  assign n73205 = pi19 ? n857 : ~n1812;
  assign n73206 = pi18 ? n32 : n73205;
  assign n73207 = pi17 ? n32 : n73206;
  assign n73208 = pi16 ? n32 : n73207;
  assign n73209 = pi15 ? n73208 : n22817;
  assign n73210 = pi15 ? n15518 : n15386;
  assign n73211 = pi14 ? n73209 : n73210;
  assign n73212 = pi14 ? n15119 : n22205;
  assign n73213 = pi13 ? n73211 : n73212;
  assign n73214 = pi12 ? n73204 : n73213;
  assign n73215 = pi11 ? n73214 : n15270;
  assign n73216 = pi10 ? n73190 : n73215;
  assign n73217 = pi09 ? n72452 : n73216;
  assign n73218 = pi15 ? n24237 : n15847;
  assign n73219 = pi14 ? n73218 : n32;
  assign n73220 = pi15 ? n17188 : n72946;
  assign n73221 = pi14 ? n17279 : n73220;
  assign n73222 = pi13 ? n73219 : n73221;
  assign n73223 = pi12 ? n73152 : n73222;
  assign n73224 = pi19 ? n1785 : n16828;
  assign n73225 = pi18 ? n32 : n73224;
  assign n73226 = pi17 ? n32 : n73225;
  assign n73227 = pi16 ? n32 : n73226;
  assign n73228 = pi20 ? n749 : ~n1817;
  assign n73229 = pi19 ? n2141 : ~n73228;
  assign n73230 = pi18 ? n32 : n73229;
  assign n73231 = pi17 ? n32 : n73230;
  assign n73232 = pi16 ? n32 : n73231;
  assign n73233 = pi15 ? n73227 : n73232;
  assign n73234 = pi14 ? n73156 : n73233;
  assign n73235 = pi20 ? n274 : ~n518;
  assign n73236 = pi19 ? n32 : n73235;
  assign n73237 = pi18 ? n32 : n73236;
  assign n73238 = pi17 ? n32 : n73237;
  assign n73239 = pi16 ? n32 : n73238;
  assign n73240 = pi15 ? n73239 : n73165;
  assign n73241 = pi19 ? n32 : n20884;
  assign n73242 = pi18 ? n32 : n73241;
  assign n73243 = pi17 ? n32 : n73242;
  assign n73244 = pi16 ? n32 : n73243;
  assign n73245 = pi15 ? n15847 : n73244;
  assign n73246 = pi14 ? n73240 : n73245;
  assign n73247 = pi13 ? n73234 : n73246;
  assign n73248 = pi19 ? n32 : n34319;
  assign n73249 = pi18 ? n32 : n73248;
  assign n73250 = pi17 ? n32 : n73249;
  assign n73251 = pi16 ? n32 : n73250;
  assign n73252 = pi19 ? n32 : ~n12680;
  assign n73253 = pi18 ? n32 : n73252;
  assign n73254 = pi17 ? n32 : n73253;
  assign n73255 = pi16 ? n32 : n73254;
  assign n73256 = pi15 ? n73251 : n73255;
  assign n73257 = pi14 ? n73170 : n73256;
  assign n73258 = pi15 ? n67470 : n15487;
  assign n73259 = pi19 ? n2141 : n4670;
  assign n73260 = pi18 ? n32 : n73259;
  assign n73261 = pi17 ? n32 : n73260;
  assign n73262 = pi16 ? n32 : n73261;
  assign n73263 = pi19 ? n1785 : n4491;
  assign n73264 = pi18 ? n32 : n73263;
  assign n73265 = pi17 ? n32 : n73264;
  assign n73266 = pi16 ? n32 : n73265;
  assign n73267 = pi15 ? n73262 : n73266;
  assign n73268 = pi14 ? n73258 : n73267;
  assign n73269 = pi13 ? n73257 : n73268;
  assign n73270 = pi12 ? n73247 : n73269;
  assign n73271 = pi11 ? n73223 : n73270;
  assign n73272 = pi19 ? n594 : n70131;
  assign n73273 = pi18 ? n32 : n73272;
  assign n73274 = pi17 ? n32 : n73273;
  assign n73275 = pi16 ? n32 : n73274;
  assign n73276 = pi15 ? n50638 : n73275;
  assign n73277 = pi15 ? n15263 : n16606;
  assign n73278 = pi14 ? n73276 : n73277;
  assign n73279 = pi15 ? n25050 : n24237;
  assign n73280 = pi14 ? n73279 : n27586;
  assign n73281 = pi13 ? n73278 : n73280;
  assign n73282 = pi19 ? n1785 : ~n1812;
  assign n73283 = pi18 ? n32 : n73282;
  assign n73284 = pi17 ? n32 : n73283;
  assign n73285 = pi16 ? n32 : n73284;
  assign n73286 = pi15 ? n73285 : n15263;
  assign n73287 = pi14 ? n73286 : n15387;
  assign n73288 = pi13 ? n73287 : n15391;
  assign n73289 = pi12 ? n73281 : n73288;
  assign n73290 = pi11 ? n73289 : n32;
  assign n73291 = pi10 ? n73271 : n73290;
  assign n73292 = pi09 ? n72452 : n73291;
  assign n73293 = pi08 ? n73217 : n73292;
  assign n73294 = pi07 ? n73149 : n73293;
  assign n73295 = pi06 ? n72939 : n73294;
  assign n73296 = pi14 ? n15847 : n32;
  assign n73297 = pi15 ? n17278 : n15927;
  assign n73298 = pi15 ? n16485 : n17193;
  assign n73299 = pi14 ? n73297 : n73298;
  assign n73300 = pi13 ? n73296 : n73299;
  assign n73301 = pi12 ? n32 : n73300;
  assign n73302 = pi20 ? n2385 : n726;
  assign n73303 = pi19 ? n32 : n73302;
  assign n73304 = pi18 ? n32 : n73303;
  assign n73305 = pi17 ? n32 : n73304;
  assign n73306 = pi16 ? n32 : n73305;
  assign n73307 = pi15 ? n73306 : n70267;
  assign n73308 = pi19 ? n32 : ~n9816;
  assign n73309 = pi18 ? n32 : n73308;
  assign n73310 = pi17 ? n32 : n73309;
  assign n73311 = pi16 ? n32 : n73310;
  assign n73312 = pi20 ? n357 : n1445;
  assign n73313 = pi19 ? n32 : n73312;
  assign n73314 = pi18 ? n32 : n73313;
  assign n73315 = pi17 ? n32 : n73314;
  assign n73316 = pi16 ? n32 : n73315;
  assign n73317 = pi15 ? n73311 : n73316;
  assign n73318 = pi14 ? n73307 : n73317;
  assign n73319 = pi20 ? n321 : n6229;
  assign n73320 = pi19 ? n594 : n73319;
  assign n73321 = pi18 ? n32 : n73320;
  assign n73322 = pi17 ? n32 : n73321;
  assign n73323 = pi16 ? n32 : n73322;
  assign n73324 = pi15 ? n53963 : n73323;
  assign n73325 = pi15 ? n55440 : n16824;
  assign n73326 = pi14 ? n73324 : n73325;
  assign n73327 = pi13 ? n73318 : n73326;
  assign n73328 = pi15 ? n16824 : n40567;
  assign n73329 = pi18 ? n32 : n36731;
  assign n73330 = pi17 ? n32 : n73329;
  assign n73331 = pi16 ? n32 : n73330;
  assign n73332 = pi15 ? n73331 : n66489;
  assign n73333 = pi14 ? n73328 : n73332;
  assign n73334 = pi19 ? n594 : ~n22704;
  assign n73335 = pi18 ? n32 : n73334;
  assign n73336 = pi17 ? n32 : n73335;
  assign n73337 = pi16 ? n32 : n73336;
  assign n73338 = pi15 ? n73337 : n55510;
  assign n73339 = pi19 ? n32 : n53064;
  assign n73340 = pi18 ? n32 : n73339;
  assign n73341 = pi17 ? n32 : n73340;
  assign n73342 = pi16 ? n32 : n73341;
  assign n73343 = pi15 ? n15847 : n73342;
  assign n73344 = pi14 ? n73338 : n73343;
  assign n73345 = pi13 ? n73333 : n73344;
  assign n73346 = pi12 ? n73327 : n73345;
  assign n73347 = pi11 ? n73301 : n73346;
  assign n73348 = pi15 ? n52315 : n55514;
  assign n73349 = pi19 ? n32 : ~n50852;
  assign n73350 = pi18 ? n32 : n73349;
  assign n73351 = pi17 ? n32 : n73350;
  assign n73352 = pi16 ? n32 : n73351;
  assign n73353 = pi15 ? n16606 : n73352;
  assign n73354 = pi14 ? n73348 : n73353;
  assign n73355 = pi15 ? n24528 : n16105;
  assign n73356 = pi15 ? n15834 : n15511;
  assign n73357 = pi14 ? n73355 : n73356;
  assign n73358 = pi13 ? n73354 : n73357;
  assign n73359 = pi15 ? n27631 : n32;
  assign n73360 = pi14 ? n73359 : n15520;
  assign n73361 = pi13 ? n73360 : n32;
  assign n73362 = pi12 ? n73358 : n73361;
  assign n73363 = pi11 ? n73362 : n32;
  assign n73364 = pi10 ? n73347 : n73363;
  assign n73365 = pi09 ? n32 : n73364;
  assign n73366 = pi20 ? n17287 : n32;
  assign n73367 = pi19 ? n32 : n73366;
  assign n73368 = pi18 ? n32 : n73367;
  assign n73369 = pi17 ? n32 : n73368;
  assign n73370 = pi16 ? n32 : n73369;
  assign n73371 = pi15 ? n15847 : n73370;
  assign n73372 = pi14 ? n73371 : n62899;
  assign n73373 = pi13 ? n73372 : n73299;
  assign n73374 = pi12 ? n32 : n73373;
  assign n73375 = pi20 ? n357 : ~n518;
  assign n73376 = pi19 ? n32 : n73375;
  assign n73377 = pi18 ? n32 : n73376;
  assign n73378 = pi17 ? n32 : n73377;
  assign n73379 = pi16 ? n32 : n73378;
  assign n73380 = pi15 ? n23484 : n73379;
  assign n73381 = pi14 ? n73307 : n73380;
  assign n73382 = pi15 ? n53963 : n15847;
  assign n73383 = pi19 ? n32 : n12885;
  assign n73384 = pi18 ? n32 : n73383;
  assign n73385 = pi17 ? n32 : n73384;
  assign n73386 = pi16 ? n32 : n73385;
  assign n73387 = pi15 ? n73386 : n16824;
  assign n73388 = pi14 ? n73382 : n73387;
  assign n73389 = pi13 ? n73381 : n73388;
  assign n73390 = pi15 ? n16824 : n15501;
  assign n73391 = pi19 ? n1574 : n32090;
  assign n73392 = pi18 ? n32 : n73391;
  assign n73393 = pi17 ? n32 : n73392;
  assign n73394 = pi16 ? n32 : n73393;
  assign n73395 = pi15 ? n73394 : n38065;
  assign n73396 = pi14 ? n73390 : n73395;
  assign n73397 = pi19 ? n32 : ~n22704;
  assign n73398 = pi18 ? n32 : n73397;
  assign n73399 = pi17 ? n32 : n73398;
  assign n73400 = pi16 ? n32 : n73399;
  assign n73401 = pi15 ? n73400 : n15507;
  assign n73402 = pi14 ? n73401 : n15847;
  assign n73403 = pi13 ? n73396 : n73402;
  assign n73404 = pi12 ? n73389 : n73403;
  assign n73405 = pi11 ? n73374 : n73404;
  assign n73406 = pi15 ? n52315 : n16105;
  assign n73407 = pi20 ? n55560 : n32;
  assign n73408 = pi19 ? n32 : n73407;
  assign n73409 = pi18 ? n32 : n73408;
  assign n73410 = pi17 ? n32 : n73409;
  assign n73411 = pi16 ? n32 : n73410;
  assign n73412 = pi15 ? n16452 : n73411;
  assign n73413 = pi14 ? n73406 : n73412;
  assign n73414 = pi15 ? n24274 : n15834;
  assign n73415 = pi14 ? n73414 : n15656;
  assign n73416 = pi13 ? n73413 : n73415;
  assign n73417 = pi14 ? n32 : n15666;
  assign n73418 = pi13 ? n73417 : n32;
  assign n73419 = pi12 ? n73416 : n73418;
  assign n73420 = pi11 ? n73419 : n32;
  assign n73421 = pi10 ? n73405 : n73420;
  assign n73422 = pi09 ? n32 : n73421;
  assign n73423 = pi08 ? n73365 : n73422;
  assign n73424 = pi15 ? n17278 : n16485;
  assign n73425 = pi15 ? n16485 : n17278;
  assign n73426 = pi14 ? n73424 : n73425;
  assign n73427 = pi13 ? n73296 : n73426;
  assign n73428 = pi12 ? n32 : n73427;
  assign n73429 = pi20 ? n17134 : ~n141;
  assign n73430 = pi19 ? n32 : n73429;
  assign n73431 = pi18 ? n32 : n73430;
  assign n73432 = pi17 ? n32 : n73431;
  assign n73433 = pi16 ? n32 : n73432;
  assign n73434 = pi15 ? n68991 : n73433;
  assign n73435 = pi15 ? n24274 : n72962;
  assign n73436 = pi14 ? n73434 : n73435;
  assign n73437 = pi20 ? n501 : ~n518;
  assign n73438 = pi19 ? n32 : n73437;
  assign n73439 = pi18 ? n32 : n73438;
  assign n73440 = pi17 ? n32 : n73439;
  assign n73441 = pi16 ? n32 : n73440;
  assign n73442 = pi15 ? n73441 : n15847;
  assign n73443 = pi20 ? n448 : n6229;
  assign n73444 = pi19 ? n32 : n73443;
  assign n73445 = pi18 ? n32 : n73444;
  assign n73446 = pi17 ? n32 : n73445;
  assign n73447 = pi16 ? n32 : n73446;
  assign n73448 = pi20 ? n339 : ~n1475;
  assign n73449 = pi19 ? n32 : n73448;
  assign n73450 = pi18 ? n32 : n73449;
  assign n73451 = pi17 ? n32 : n73450;
  assign n73452 = pi16 ? n32 : n73451;
  assign n73453 = pi15 ? n73447 : n73452;
  assign n73454 = pi14 ? n73442 : n73453;
  assign n73455 = pi13 ? n73436 : n73454;
  assign n73456 = pi20 ? n501 : ~n749;
  assign n73457 = pi19 ? n32 : n73456;
  assign n73458 = pi18 ? n32 : n73457;
  assign n73459 = pi17 ? n32 : n73458;
  assign n73460 = pi16 ? n32 : n73459;
  assign n73461 = pi21 ? n9485 : ~n206;
  assign n73462 = pi20 ? n73461 : n32;
  assign n73463 = pi19 ? n32 : n73462;
  assign n73464 = pi18 ? n32 : n73463;
  assign n73465 = pi17 ? n32 : n73464;
  assign n73466 = pi16 ? n32 : n73465;
  assign n73467 = pi15 ? n73460 : n73466;
  assign n73468 = pi21 ? n10445 : n32;
  assign n73469 = pi20 ? n73468 : ~n207;
  assign n73470 = pi19 ? n32 : n73469;
  assign n73471 = pi18 ? n32 : n73470;
  assign n73472 = pi17 ? n32 : n73471;
  assign n73473 = pi16 ? n32 : n73472;
  assign n73474 = pi19 ? n32 : n45341;
  assign n73475 = pi18 ? n32 : n73474;
  assign n73476 = pi17 ? n32 : n73475;
  assign n73477 = pi16 ? n32 : n73476;
  assign n73478 = pi15 ? n73473 : n73477;
  assign n73479 = pi14 ? n73467 : n73478;
  assign n73480 = pi21 ? n14792 : ~n32;
  assign n73481 = pi20 ? n73480 : ~n339;
  assign n73482 = pi19 ? n32 : n73481;
  assign n73483 = pi18 ? n32 : n73482;
  assign n73484 = pi17 ? n32 : n73483;
  assign n73485 = pi16 ? n32 : n73484;
  assign n73486 = pi15 ? n73485 : n15655;
  assign n73487 = pi20 ? n38586 : n32;
  assign n73488 = pi19 ? n32 : n73487;
  assign n73489 = pi18 ? n32 : n73488;
  assign n73490 = pi17 ? n32 : n73489;
  assign n73491 = pi16 ? n32 : n73490;
  assign n73492 = pi20 ? n13426 : n32;
  assign n73493 = pi19 ? n32 : n73492;
  assign n73494 = pi18 ? n32 : n73493;
  assign n73495 = pi17 ? n32 : n73494;
  assign n73496 = pi16 ? n32 : n73495;
  assign n73497 = pi15 ? n73491 : n73496;
  assign n73498 = pi14 ? n73486 : n73497;
  assign n73499 = pi13 ? n73479 : n73498;
  assign n73500 = pi12 ? n73455 : n73499;
  assign n73501 = pi11 ? n73428 : n73500;
  assign n73502 = pi21 ? n1009 : n174;
  assign n73503 = pi20 ? n73502 : n32;
  assign n73504 = pi19 ? n32 : n73503;
  assign n73505 = pi18 ? n32 : n73504;
  assign n73506 = pi17 ? n32 : n73505;
  assign n73507 = pi16 ? n32 : n73506;
  assign n73508 = pi20 ? n73468 : n32;
  assign n73509 = pi19 ? n32 : n73508;
  assign n73510 = pi18 ? n32 : n73509;
  assign n73511 = pi17 ? n32 : n73510;
  assign n73512 = pi16 ? n32 : n73511;
  assign n73513 = pi15 ? n73507 : n73512;
  assign n73514 = pi15 ? n16101 : n55727;
  assign n73515 = pi14 ? n73513 : n73514;
  assign n73516 = pi21 ? n50 : n32;
  assign n73517 = pi20 ? n73516 : n32;
  assign n73518 = pi19 ? n32 : n73517;
  assign n73519 = pi18 ? n32 : n73518;
  assign n73520 = pi17 ? n32 : n73519;
  assign n73521 = pi16 ? n32 : n73520;
  assign n73522 = pi15 ? n32 : n73521;
  assign n73523 = pi14 ? n73522 : n15837;
  assign n73524 = pi13 ? n73515 : n73523;
  assign n73525 = pi12 ? n73524 : n32;
  assign n73526 = pi11 ? n73525 : n32;
  assign n73527 = pi10 ? n73501 : n73526;
  assign n73528 = pi09 ? n32 : n73527;
  assign n73529 = pi15 ? n53963 : n16832;
  assign n73530 = pi15 ? n32 : n72962;
  assign n73531 = pi14 ? n73529 : n73530;
  assign n73532 = pi15 ? n73460 : n15847;
  assign n73533 = pi15 ? n73447 : n15766;
  assign n73534 = pi14 ? n73532 : n73533;
  assign n73535 = pi13 ? n73531 : n73534;
  assign n73536 = pi19 ? n32 : n6029;
  assign n73537 = pi18 ? n32 : n73536;
  assign n73538 = pi17 ? n32 : n73537;
  assign n73539 = pi16 ? n32 : n73538;
  assign n73540 = pi15 ? n73539 : n53895;
  assign n73541 = pi19 ? n32 : n45235;
  assign n73542 = pi18 ? n32 : n73541;
  assign n73543 = pi17 ? n32 : n73542;
  assign n73544 = pi16 ? n32 : n73543;
  assign n73545 = pi15 ? n73473 : n73544;
  assign n73546 = pi14 ? n73540 : n73545;
  assign n73547 = pi20 ? n11589 : n32;
  assign n73548 = pi19 ? n32 : n73547;
  assign n73549 = pi18 ? n32 : n73548;
  assign n73550 = pi17 ? n32 : n73549;
  assign n73551 = pi16 ? n32 : n73550;
  assign n73552 = pi15 ? n73551 : n15836;
  assign n73553 = pi21 ? n242 : ~n174;
  assign n73554 = pi20 ? n73553 : n32;
  assign n73555 = pi19 ? n32 : n73554;
  assign n73556 = pi18 ? n32 : n73555;
  assign n73557 = pi17 ? n32 : n73556;
  assign n73558 = pi16 ? n32 : n73557;
  assign n73559 = pi15 ? n73558 : n16105;
  assign n73560 = pi14 ? n73552 : n73559;
  assign n73561 = pi13 ? n73546 : n73560;
  assign n73562 = pi12 ? n73535 : n73561;
  assign n73563 = pi11 ? n73428 : n73562;
  assign n73564 = pi21 ? n48999 : n32;
  assign n73565 = pi20 ? n73564 : n32;
  assign n73566 = pi19 ? n32 : n73565;
  assign n73567 = pi18 ? n32 : n73566;
  assign n73568 = pi17 ? n32 : n73567;
  assign n73569 = pi16 ? n32 : n73568;
  assign n73570 = pi15 ? n32 : n73569;
  assign n73571 = pi19 ? n32 : n31748;
  assign n73572 = pi18 ? n32 : n73571;
  assign n73573 = pi17 ? n32 : n73572;
  assign n73574 = pi16 ? n32 : n73573;
  assign n73575 = pi15 ? n73574 : n16108;
  assign n73576 = pi14 ? n73570 : n73575;
  assign n73577 = pi15 ? n15836 : n15700;
  assign n73578 = pi14 ? n73577 : n15968;
  assign n73579 = pi13 ? n73576 : n73578;
  assign n73580 = pi12 ? n73579 : n32;
  assign n73581 = pi11 ? n73580 : n32;
  assign n73582 = pi10 ? n73563 : n73581;
  assign n73583 = pi09 ? n32 : n73582;
  assign n73584 = pi08 ? n73528 : n73583;
  assign n73585 = pi07 ? n73423 : n73584;
  assign n73586 = pi15 ? n17278 : n25713;
  assign n73587 = pi20 ? n266 : ~n10066;
  assign n73588 = pi19 ? n32 : n73587;
  assign n73589 = pi18 ? n32 : n73588;
  assign n73590 = pi17 ? n32 : n73589;
  assign n73591 = pi16 ? n32 : n73590;
  assign n73592 = pi20 ? n653 : n9000;
  assign n73593 = pi19 ? n32 : n73592;
  assign n73594 = pi18 ? n32 : n73593;
  assign n73595 = pi17 ? n32 : n73594;
  assign n73596 = pi16 ? n32 : n73595;
  assign n73597 = pi15 ? n73591 : n73596;
  assign n73598 = pi14 ? n73586 : n73597;
  assign n73599 = pi13 ? n73296 : n73598;
  assign n73600 = pi12 ? n32 : n73599;
  assign n73601 = pi20 ? n321 : n1685;
  assign n73602 = pi19 ? n32 : n73601;
  assign n73603 = pi18 ? n32 : n73602;
  assign n73604 = pi17 ? n32 : n73603;
  assign n73605 = pi16 ? n32 : n73604;
  assign n73606 = pi20 ? n12244 : ~n518;
  assign n73607 = pi19 ? n32 : n73606;
  assign n73608 = pi18 ? n32 : n73607;
  assign n73609 = pi17 ? n32 : n73608;
  assign n73610 = pi16 ? n32 : n73609;
  assign n73611 = pi15 ? n73605 : n73610;
  assign n73612 = pi14 ? n38744 : n73611;
  assign n73613 = pi20 ? n274 : ~n749;
  assign n73614 = pi19 ? n32 : n73613;
  assign n73615 = pi18 ? n32 : n73614;
  assign n73616 = pi17 ? n32 : n73615;
  assign n73617 = pi16 ? n32 : n73616;
  assign n73618 = pi15 ? n73617 : n32;
  assign n73619 = pi20 ? n749 : ~n11048;
  assign n73620 = pi19 ? n32 : n73619;
  assign n73621 = pi18 ? n32 : n73620;
  assign n73622 = pi17 ? n32 : n73621;
  assign n73623 = pi16 ? n32 : n73622;
  assign n73624 = pi20 ? n1940 : ~n749;
  assign n73625 = pi19 ? n32 : n73624;
  assign n73626 = pi18 ? n32 : n73625;
  assign n73627 = pi17 ? n32 : n73626;
  assign n73628 = pi16 ? n32 : n73627;
  assign n73629 = pi15 ? n73623 : n73628;
  assign n73630 = pi14 ? n73618 : n73629;
  assign n73631 = pi13 ? n73612 : n73630;
  assign n73632 = pi20 ? n11589 : ~n207;
  assign n73633 = pi19 ? n32 : n73632;
  assign n73634 = pi18 ? n32 : n73633;
  assign n73635 = pi17 ? n32 : n73634;
  assign n73636 = pi16 ? n32 : n73635;
  assign n73637 = pi15 ? n55571 : n73636;
  assign n73638 = pi21 ? n48999 : n206;
  assign n73639 = pi20 ? n73638 : ~n207;
  assign n73640 = pi19 ? n32 : n73639;
  assign n73641 = pi18 ? n32 : n73640;
  assign n73642 = pi17 ? n32 : n73641;
  assign n73643 = pi16 ? n32 : n73642;
  assign n73644 = pi20 ? n16079 : ~n339;
  assign n73645 = pi19 ? n32 : n73644;
  assign n73646 = pi18 ? n32 : n73645;
  assign n73647 = pi17 ? n32 : n73646;
  assign n73648 = pi16 ? n32 : n73647;
  assign n73649 = pi15 ? n73643 : n73648;
  assign n73650 = pi14 ? n73637 : n73649;
  assign n73651 = pi21 ? n35 : n1009;
  assign n73652 = pi20 ? n73651 : n32;
  assign n73653 = pi19 ? n32 : n73652;
  assign n73654 = pi18 ? n32 : n73653;
  assign n73655 = pi17 ? n32 : n73654;
  assign n73656 = pi16 ? n32 : n73655;
  assign n73657 = pi15 ? n55727 : n73656;
  assign n73658 = pi15 ? n15935 : n16108;
  assign n73659 = pi14 ? n73657 : n73658;
  assign n73660 = pi13 ? n73650 : n73659;
  assign n73661 = pi12 ? n73631 : n73660;
  assign n73662 = pi11 ? n73600 : n73661;
  assign n73663 = pi15 ? n16319 : n16204;
  assign n73664 = pi15 ? n16377 : n16108;
  assign n73665 = pi14 ? n73663 : n73664;
  assign n73666 = pi14 ? n16218 : n16110;
  assign n73667 = pi13 ? n73665 : n73666;
  assign n73668 = pi12 ? n73667 : n32;
  assign n73669 = pi11 ? n73668 : n32;
  assign n73670 = pi10 ? n73662 : n73669;
  assign n73671 = pi09 ? n32 : n73670;
  assign n73672 = pi20 ? n749 : ~n141;
  assign n73673 = pi19 ? n32 : n73672;
  assign n73674 = pi18 ? n32 : n73673;
  assign n73675 = pi17 ? n32 : n73674;
  assign n73676 = pi16 ? n32 : n73675;
  assign n73677 = pi15 ? n17278 : n73676;
  assign n73678 = pi20 ? n1331 : n220;
  assign n73679 = pi19 ? n32 : n73678;
  assign n73680 = pi18 ? n32 : n73679;
  assign n73681 = pi17 ? n32 : n73680;
  assign n73682 = pi16 ? n32 : n73681;
  assign n73683 = pi15 ? n73682 : n17278;
  assign n73684 = pi14 ? n73677 : n73683;
  assign n73685 = pi13 ? n73296 : n73684;
  assign n73686 = pi12 ? n32 : n73685;
  assign n73687 = pi20 ? n12244 : ~n1839;
  assign n73688 = pi19 ? n32 : n73687;
  assign n73689 = pi18 ? n32 : n73688;
  assign n73690 = pi17 ? n32 : n73689;
  assign n73691 = pi16 ? n32 : n73690;
  assign n73692 = pi15 ? n73605 : n73691;
  assign n73693 = pi14 ? n38744 : n73692;
  assign n73694 = pi15 ? n16049 : n55715;
  assign n73695 = pi14 ? n27376 : n73694;
  assign n73696 = pi13 ? n73693 : n73695;
  assign n73697 = pi15 ? n15847 : n16286;
  assign n73698 = pi19 ? n32 : n21415;
  assign n73699 = pi18 ? n32 : n73698;
  assign n73700 = pi17 ? n32 : n73699;
  assign n73701 = pi16 ? n32 : n73700;
  assign n73702 = pi15 ? n73701 : n25763;
  assign n73703 = pi14 ? n73697 : n73702;
  assign n73704 = pi21 ? n1939 : n1009;
  assign n73705 = pi20 ? n73704 : n32;
  assign n73706 = pi19 ? n32 : n73705;
  assign n73707 = pi18 ? n32 : n73706;
  assign n73708 = pi17 ? n32 : n73707;
  assign n73709 = pi16 ? n32 : n73708;
  assign n73710 = pi15 ? n55727 : n73709;
  assign n73711 = pi14 ? n73710 : n25818;
  assign n73712 = pi13 ? n73703 : n73711;
  assign n73713 = pi12 ? n73696 : n73712;
  assign n73714 = pi11 ? n73686 : n73713;
  assign n73715 = pi15 ? n15700 : n16204;
  assign n73716 = pi14 ? n73715 : n16378;
  assign n73717 = pi13 ? n73716 : n16219;
  assign n73718 = pi12 ? n73717 : n32;
  assign n73719 = pi11 ? n73718 : n32;
  assign n73720 = pi10 ? n73714 : n73719;
  assign n73721 = pi09 ? n32 : n73720;
  assign n73722 = pi08 ? n73671 : n73721;
  assign n73723 = pi14 ? n73424 : n17278;
  assign n73724 = pi13 ? n73296 : n73723;
  assign n73725 = pi12 ? n32 : n73724;
  assign n73726 = pi20 ? n321 : n1445;
  assign n73727 = pi19 ? n32 : n73726;
  assign n73728 = pi18 ? n32 : n73727;
  assign n73729 = pi17 ? n32 : n73728;
  assign n73730 = pi16 ? n32 : n73729;
  assign n73731 = pi19 ? n32 : n34129;
  assign n73732 = pi18 ? n32 : n73731;
  assign n73733 = pi17 ? n32 : n73732;
  assign n73734 = pi16 ? n32 : n73733;
  assign n73735 = pi15 ? n73730 : n73734;
  assign n73736 = pi14 ? n72819 : n73735;
  assign n73737 = pi20 ? n749 : ~n1475;
  assign n73738 = pi19 ? n32 : n73737;
  assign n73739 = pi18 ? n32 : n73738;
  assign n73740 = pi17 ? n32 : n73739;
  assign n73741 = pi16 ? n32 : n73740;
  assign n73742 = pi15 ? n73741 : n16352;
  assign n73743 = pi14 ? n27341 : n73742;
  assign n73744 = pi13 ? n73736 : n73743;
  assign n73745 = pi15 ? n73701 : n32;
  assign n73746 = pi14 ? n73697 : n73745;
  assign n73747 = pi20 ? n9667 : n32;
  assign n73748 = pi19 ? n32 : n73747;
  assign n73749 = pi18 ? n32 : n73748;
  assign n73750 = pi17 ? n32 : n73749;
  assign n73751 = pi16 ? n32 : n73750;
  assign n73752 = pi15 ? n15847 : n73751;
  assign n73753 = pi14 ? n73752 : n37574;
  assign n73754 = pi13 ? n73746 : n73753;
  assign n73755 = pi12 ? n73744 : n73754;
  assign n73756 = pi11 ? n73725 : n73755;
  assign n73757 = pi18 ? n32 : n3845;
  assign n73758 = pi17 ? n32 : n73757;
  assign n73759 = pi16 ? n32 : n73758;
  assign n73760 = pi15 ? n73759 : n16319;
  assign n73761 = pi14 ? n73760 : n16378;
  assign n73762 = pi13 ? n73761 : n16322;
  assign n73763 = pi12 ? n73762 : n32;
  assign n73764 = pi11 ? n73763 : n32;
  assign n73765 = pi10 ? n73756 : n73764;
  assign n73766 = pi09 ? n32 : n73765;
  assign n73767 = pi15 ? n73596 : n17278;
  assign n73768 = pi14 ? n73424 : n73767;
  assign n73769 = pi13 ? n73296 : n73768;
  assign n73770 = pi12 ? n32 : n73769;
  assign n73771 = pi19 ? n32 : n13353;
  assign n73772 = pi18 ? n32 : n73771;
  assign n73773 = pi17 ? n32 : n73772;
  assign n73774 = pi16 ? n32 : n73773;
  assign n73775 = pi15 ? n73774 : n16352;
  assign n73776 = pi14 ? n27341 : n73775;
  assign n73777 = pi13 ? n73736 : n73776;
  assign n73778 = pi20 ? n1475 : ~n207;
  assign n73779 = pi19 ? n32 : n73778;
  assign n73780 = pi18 ? n32 : n73779;
  assign n73781 = pi17 ? n32 : n73780;
  assign n73782 = pi16 ? n32 : n73781;
  assign n73783 = pi15 ? n15847 : n73782;
  assign n73784 = pi14 ? n73783 : n73745;
  assign n73785 = pi15 ? n15847 : n16333;
  assign n73786 = pi21 ? n100 : ~n50;
  assign n73787 = pi20 ? n73786 : n32;
  assign n73788 = pi19 ? n32 : n73787;
  assign n73789 = pi18 ? n32 : n73788;
  assign n73790 = pi17 ? n32 : n73789;
  assign n73791 = pi16 ? n32 : n73790;
  assign n73792 = pi15 ? n73791 : n16293;
  assign n73793 = pi14 ? n73785 : n73792;
  assign n73794 = pi13 ? n73784 : n73793;
  assign n73795 = pi12 ? n73777 : n73794;
  assign n73796 = pi11 ? n73770 : n73795;
  assign n73797 = pi14 ? n16457 : n16378;
  assign n73798 = pi13 ? n73797 : n32;
  assign n73799 = pi12 ? n73798 : n32;
  assign n73800 = pi11 ? n73799 : n32;
  assign n73801 = pi10 ? n73796 : n73800;
  assign n73802 = pi09 ? n32 : n73801;
  assign n73803 = pi08 ? n73766 : n73802;
  assign n73804 = pi07 ? n73722 : n73803;
  assign n73805 = pi06 ? n73585 : n73804;
  assign n73806 = pi05 ? n73295 : n73805;
  assign n73807 = pi13 ? n32 : n54461;
  assign n73808 = pi12 ? n32 : n73807;
  assign n73809 = pi11 ? n32 : n73808;
  assign n73810 = pi10 ? n32 : n73809;
  assign n73811 = pi14 ? n32 : n16397;
  assign n73812 = pi19 ? n32 : n65428;
  assign n73813 = pi18 ? n32 : n73812;
  assign n73814 = pi17 ? n32 : n73813;
  assign n73815 = pi16 ? n32 : n73814;
  assign n73816 = pi15 ? n73815 : n16392;
  assign n73817 = pi15 ? n17278 : n68991;
  assign n73818 = pi14 ? n73816 : n73817;
  assign n73819 = pi13 ? n73811 : n73818;
  assign n73820 = pi12 ? n32 : n73819;
  assign n73821 = pi20 ? n518 : n1817;
  assign n73822 = pi19 ? n32 : n73821;
  assign n73823 = pi18 ? n32 : n73822;
  assign n73824 = pi17 ? n32 : n73823;
  assign n73825 = pi16 ? n32 : n73824;
  assign n73826 = pi15 ? n17121 : n73825;
  assign n73827 = pi20 ? n518 : n1445;
  assign n73828 = pi19 ? n32 : n73827;
  assign n73829 = pi18 ? n32 : n73828;
  assign n73830 = pi17 ? n32 : n73829;
  assign n73831 = pi16 ? n32 : n73830;
  assign n73832 = pi20 ? n1817 : ~n1839;
  assign n73833 = pi19 ? n32 : n73832;
  assign n73834 = pi18 ? n32 : n73833;
  assign n73835 = pi17 ? n32 : n73834;
  assign n73836 = pi16 ? n32 : n73835;
  assign n73837 = pi15 ? n73831 : n73836;
  assign n73838 = pi14 ? n73826 : n73837;
  assign n73839 = pi15 ? n25904 : n67879;
  assign n73840 = pi20 ? n1076 : ~n749;
  assign n73841 = pi19 ? n32 : n73840;
  assign n73842 = pi18 ? n32 : n73841;
  assign n73843 = pi17 ? n32 : n73842;
  assign n73844 = pi16 ? n32 : n73843;
  assign n73845 = pi15 ? n67879 : n73844;
  assign n73846 = pi14 ? n73839 : n73845;
  assign n73847 = pi13 ? n73838 : n73846;
  assign n73848 = pi14 ? n16447 : n27557;
  assign n73849 = pi21 ? n32 : ~n50;
  assign n73850 = pi20 ? n73849 : n32;
  assign n73851 = pi19 ? n32 : n73850;
  assign n73852 = pi18 ? n32 : n73851;
  assign n73853 = pi17 ? n32 : n73852;
  assign n73854 = pi16 ? n32 : n73853;
  assign n73855 = pi15 ? n73854 : n16452;
  assign n73856 = pi14 ? n16333 : n73855;
  assign n73857 = pi13 ? n73848 : n73856;
  assign n73858 = pi12 ? n73847 : n73857;
  assign n73859 = pi11 ? n73820 : n73858;
  assign n73860 = pi10 ? n73859 : n16461;
  assign n73861 = pi09 ? n73810 : n73860;
  assign n73862 = pi14 ? n16393 : n24496;
  assign n73863 = pi13 ? n32 : n73862;
  assign n73864 = pi12 ? n32 : n73863;
  assign n73865 = pi11 ? n32 : n73864;
  assign n73866 = pi10 ? n32 : n73865;
  assign n73867 = pi20 ? n8630 : ~n321;
  assign n73868 = pi19 ? n32 : n73867;
  assign n73869 = pi18 ? n32 : n73868;
  assign n73870 = pi17 ? n32 : n73869;
  assign n73871 = pi16 ? n32 : n73870;
  assign n73872 = pi15 ? n16397 : n73871;
  assign n73873 = pi14 ? n32 : n73872;
  assign n73874 = pi13 ? n73873 : n73818;
  assign n73875 = pi12 ? n32 : n73874;
  assign n73876 = pi20 ? n382 : ~n1839;
  assign n73877 = pi19 ? n32 : n73876;
  assign n73878 = pi18 ? n32 : n73877;
  assign n73879 = pi17 ? n32 : n73878;
  assign n73880 = pi16 ? n32 : n73879;
  assign n73881 = pi15 ? n73831 : n73880;
  assign n73882 = pi14 ? n73826 : n73881;
  assign n73883 = pi15 ? n25904 : n16582;
  assign n73884 = pi15 ? n16582 : n16804;
  assign n73885 = pi14 ? n73883 : n73884;
  assign n73886 = pi13 ? n73882 : n73885;
  assign n73887 = pi14 ? n16413 : n25633;
  assign n73888 = pi15 ? n16333 : n27753;
  assign n73889 = pi15 ? n73854 : n16606;
  assign n73890 = pi14 ? n73888 : n73889;
  assign n73891 = pi13 ? n73887 : n73890;
  assign n73892 = pi12 ? n73886 : n73891;
  assign n73893 = pi11 ? n73875 : n73892;
  assign n73894 = pi10 ? n73893 : n32;
  assign n73895 = pi09 ? n73866 : n73894;
  assign n73896 = pi08 ? n73861 : n73895;
  assign n73897 = pi15 ? n15987 : n16397;
  assign n73898 = pi14 ? n24563 : n73897;
  assign n73899 = pi14 ? n25498 : n73817;
  assign n73900 = pi13 ? n73898 : n73899;
  assign n73901 = pi12 ? n32 : n73900;
  assign n73902 = pi15 ? n16606 : n73825;
  assign n73903 = pi20 ? n8630 : ~n518;
  assign n73904 = pi19 ? n32 : n73903;
  assign n73905 = pi18 ? n32 : n73904;
  assign n73906 = pi17 ? n32 : n73905;
  assign n73907 = pi16 ? n32 : n73906;
  assign n73908 = pi20 ? n382 : n16570;
  assign n73909 = pi19 ? n32 : n73908;
  assign n73910 = pi18 ? n32 : n73909;
  assign n73911 = pi17 ? n32 : n73910;
  assign n73912 = pi16 ? n32 : n73911;
  assign n73913 = pi15 ? n73907 : n73912;
  assign n73914 = pi14 ? n73902 : n73913;
  assign n73915 = pi20 ? n8630 : ~n1475;
  assign n73916 = pi19 ? n32 : n73915;
  assign n73917 = pi18 ? n32 : n73916;
  assign n73918 = pi17 ? n32 : n73917;
  assign n73919 = pi16 ? n32 : n73918;
  assign n73920 = pi15 ? n16606 : n73919;
  assign n73921 = pi15 ? n73919 : n16587;
  assign n73922 = pi14 ? n73920 : n73921;
  assign n73923 = pi13 ? n73914 : n73922;
  assign n73924 = pi15 ? n16595 : n16804;
  assign n73925 = pi15 ? n16832 : n16546;
  assign n73926 = pi14 ? n73924 : n73925;
  assign n73927 = pi14 ? n27789 : n16607;
  assign n73928 = pi13 ? n73926 : n73927;
  assign n73929 = pi12 ? n73923 : n73928;
  assign n73930 = pi11 ? n73901 : n73929;
  assign n73931 = pi10 ? n73930 : n32;
  assign n73932 = pi09 ? n73810 : n73931;
  assign n73933 = pi15 ? n17193 : n70243;
  assign n73934 = pi14 ? n16393 : n73933;
  assign n73935 = pi13 ? n73898 : n73934;
  assign n73936 = pi12 ? n32 : n73935;
  assign n73937 = pi15 ? n53963 : n27720;
  assign n73938 = pi14 ? n73902 : n73937;
  assign n73939 = pi15 ? n16606 : n16824;
  assign n73940 = pi15 ? n16824 : n16587;
  assign n73941 = pi14 ? n73939 : n73940;
  assign n73942 = pi13 ? n73938 : n73941;
  assign n73943 = pi14 ? n27789 : n16656;
  assign n73944 = pi13 ? n73926 : n73943;
  assign n73945 = pi12 ? n73942 : n73944;
  assign n73946 = pi11 ? n73936 : n73945;
  assign n73947 = pi10 ? n73946 : n32;
  assign n73948 = pi09 ? n73810 : n73947;
  assign n73949 = pi08 ? n73932 : n73948;
  assign n73950 = pi07 ? n73896 : n73949;
  assign n73951 = pi13 ? n32 : n37913;
  assign n73952 = pi15 ? n17193 : n26515;
  assign n73953 = pi14 ? n16393 : n73952;
  assign n73954 = pi13 ? n17077 : n73953;
  assign n73955 = pi12 ? n73951 : n73954;
  assign n73956 = pi20 ? n3523 : n1445;
  assign n73957 = pi19 ? n32 : n73956;
  assign n73958 = pi18 ? n32 : n73957;
  assign n73959 = pi17 ? n32 : n73958;
  assign n73960 = pi16 ? n32 : n73959;
  assign n73961 = pi15 ? n16606 : n73960;
  assign n73962 = pi15 ? n53963 : n16392;
  assign n73963 = pi14 ? n73961 : n73962;
  assign n73964 = pi20 ? n3523 : ~n1475;
  assign n73965 = pi19 ? n32 : n73964;
  assign n73966 = pi18 ? n32 : n73965;
  assign n73967 = pi17 ? n32 : n73966;
  assign n73968 = pi16 ? n32 : n73967;
  assign n73969 = pi15 ? n73968 : n16824;
  assign n73970 = pi15 ? n16467 : n16711;
  assign n73971 = pi14 ? n73969 : n73970;
  assign n73972 = pi13 ? n73963 : n73971;
  assign n73973 = pi15 ? n68001 : n32;
  assign n73974 = pi20 ? n13792 : ~n141;
  assign n73975 = pi19 ? n32 : n73974;
  assign n73976 = pi18 ? n32 : n73975;
  assign n73977 = pi17 ? n32 : n73976;
  assign n73978 = pi16 ? n32 : n73977;
  assign n73979 = pi15 ? n73978 : n16965;
  assign n73980 = pi14 ? n73973 : n73979;
  assign n73981 = pi15 ? n32 : n16655;
  assign n73982 = pi14 ? n73981 : n32;
  assign n73983 = pi13 ? n73980 : n73982;
  assign n73984 = pi12 ? n73972 : n73983;
  assign n73985 = pi11 ? n73955 : n73984;
  assign n73986 = pi10 ? n73985 : n32;
  assign n73987 = pi09 ? n32 : n73986;
  assign n73988 = pi14 ? n24495 : n16850;
  assign n73989 = pi20 ? n151 : n726;
  assign n73990 = pi19 ? n32 : n73989;
  assign n73991 = pi18 ? n32 : n73990;
  assign n73992 = pi17 ? n32 : n73991;
  assign n73993 = pi16 ? n32 : n73992;
  assign n73994 = pi15 ? n17193 : n73993;
  assign n73995 = pi14 ? n16393 : n73994;
  assign n73996 = pi13 ? n73988 : n73995;
  assign n73997 = pi12 ? n73951 : n73996;
  assign n73998 = pi15 ? n55871 : n17286;
  assign n73999 = pi15 ? n16884 : n16467;
  assign n74000 = pi14 ? n73998 : n73999;
  assign n74001 = pi14 ? n52055 : n73970;
  assign n74002 = pi13 ? n74000 : n74001;
  assign n74003 = pi15 ? n68001 : n24495;
  assign n74004 = pi14 ? n74003 : n25633;
  assign n74005 = pi13 ? n74004 : n16787;
  assign n74006 = pi12 ? n74002 : n74005;
  assign n74007 = pi11 ? n73997 : n74006;
  assign n74008 = pi10 ? n74007 : n32;
  assign n74009 = pi09 ? n32 : n74008;
  assign n74010 = pi08 ? n73987 : n74009;
  assign n74011 = pi20 ? n13792 : n726;
  assign n74012 = pi19 ? n32 : n74011;
  assign n74013 = pi18 ? n32 : n74012;
  assign n74014 = pi17 ? n32 : n74013;
  assign n74015 = pi16 ? n32 : n74014;
  assign n74016 = pi15 ? n17278 : n74015;
  assign n74017 = pi14 ? n26161 : n74016;
  assign n74018 = pi13 ? n17077 : n74017;
  assign n74019 = pi12 ? n73807 : n74018;
  assign n74020 = pi15 ? n16392 : n68001;
  assign n74021 = pi14 ? n52055 : n74020;
  assign n74022 = pi13 ? n74000 : n74021;
  assign n74023 = pi15 ? n17121 : n17039;
  assign n74024 = pi14 ? n74023 : n16838;
  assign n74025 = pi13 ? n74024 : n16841;
  assign n74026 = pi12 ? n74022 : n74025;
  assign n74027 = pi11 ? n74019 : n74026;
  assign n74028 = pi10 ? n74027 : n32;
  assign n74029 = pi09 ? n17493 : n74028;
  assign n74030 = pi20 ? n428 : n623;
  assign n74031 = pi19 ? n32 : n74030;
  assign n74032 = pi18 ? n32 : n74031;
  assign n74033 = pi17 ? n32 : n74032;
  assign n74034 = pi16 ? n32 : n74033;
  assign n74035 = pi15 ? n17278 : n74034;
  assign n74036 = pi14 ? n26161 : n74035;
  assign n74037 = pi13 ? n17077 : n74036;
  assign n74038 = pi12 ? n73807 : n74037;
  assign n74039 = pi15 ? n16890 : n16392;
  assign n74040 = pi14 ? n39087 : n74039;
  assign n74041 = pi14 ? n27616 : n74020;
  assign n74042 = pi13 ? n74040 : n74041;
  assign n74043 = pi15 ? n17002 : n32;
  assign n74044 = pi14 ? n37568 : n74043;
  assign n74045 = pi13 ? n74044 : n32;
  assign n74046 = pi12 ? n74042 : n74045;
  assign n74047 = pi11 ? n74038 : n74046;
  assign n74048 = pi10 ? n74047 : n32;
  assign n74049 = pi09 ? n17493 : n74048;
  assign n74050 = pi08 ? n74029 : n74049;
  assign n74051 = pi07 ? n74010 : n74050;
  assign n74052 = pi06 ? n73950 : n74051;
  assign n74053 = pi15 ? n16850 : n17039;
  assign n74054 = pi14 ? n32 : n74053;
  assign n74055 = pi20 ? n13387 : n220;
  assign n74056 = pi19 ? n32 : n74055;
  assign n74057 = pi18 ? n32 : n74056;
  assign n74058 = pi17 ? n32 : n74057;
  assign n74059 = pi16 ? n32 : n74058;
  assign n74060 = pi15 ? n17036 : n74059;
  assign n74061 = pi20 ? n12019 : ~n2140;
  assign n74062 = pi19 ? n32 : n74061;
  assign n74063 = pi18 ? n32 : n74062;
  assign n74064 = pi17 ? n32 : n74063;
  assign n74065 = pi16 ? n32 : n74064;
  assign n74066 = pi15 ? n74065 : n17039;
  assign n74067 = pi14 ? n74060 : n74066;
  assign n74068 = pi13 ? n74054 : n74067;
  assign n74069 = pi12 ? n32 : n74068;
  assign n74070 = pi20 ? n67 : ~n14844;
  assign n74071 = pi19 ? n32 : n74070;
  assign n74072 = pi18 ? n32 : n74071;
  assign n74073 = pi17 ? n32 : n74072;
  assign n74074 = pi16 ? n32 : n74073;
  assign n74075 = pi20 ? n67 : ~n518;
  assign n74076 = pi19 ? n32 : n74075;
  assign n74077 = pi18 ? n32 : n74076;
  assign n74078 = pi17 ? n32 : n74077;
  assign n74079 = pi16 ? n32 : n74078;
  assign n74080 = pi15 ? n74074 : n74079;
  assign n74081 = pi14 ? n74080 : n25133;
  assign n74082 = pi20 ? n67 : ~n1475;
  assign n74083 = pi19 ? n32 : n74082;
  assign n74084 = pi18 ? n32 : n74083;
  assign n74085 = pi17 ? n32 : n74084;
  assign n74086 = pi16 ? n32 : n74085;
  assign n74087 = pi15 ? n74086 : n16862;
  assign n74088 = pi20 ? n67 : ~n207;
  assign n74089 = pi19 ? n32 : n74088;
  assign n74090 = pi18 ? n32 : n74089;
  assign n74091 = pi17 ? n32 : n74090;
  assign n74092 = pi16 ? n32 : n74091;
  assign n74093 = pi15 ? n17061 : n74092;
  assign n74094 = pi14 ? n74087 : n74093;
  assign n74095 = pi13 ? n74081 : n74094;
  assign n74096 = pi15 ? n36851 : n17036;
  assign n74097 = pi14 ? n74096 : n16974;
  assign n74098 = pi13 ? n74097 : n32;
  assign n74099 = pi12 ? n74095 : n74098;
  assign n74100 = pi11 ? n74069 : n74099;
  assign n74101 = pi10 ? n74100 : n32;
  assign n74102 = pi09 ? n17493 : n74101;
  assign n74103 = pi20 ? n16997 : n220;
  assign n74104 = pi19 ? n32 : n74103;
  assign n74105 = pi18 ? n32 : n74104;
  assign n74106 = pi17 ? n32 : n74105;
  assign n74107 = pi16 ? n32 : n74106;
  assign n74108 = pi15 ? n17036 : n74107;
  assign n74109 = pi20 ? n11403 : ~n2140;
  assign n74110 = pi19 ? n32 : n74109;
  assign n74111 = pi18 ? n32 : n74110;
  assign n74112 = pi17 ? n32 : n74111;
  assign n74113 = pi16 ? n32 : n74112;
  assign n74114 = pi15 ? n74113 : n17039;
  assign n74115 = pi14 ? n74108 : n74114;
  assign n74116 = pi13 ? n74054 : n74115;
  assign n74117 = pi12 ? n32 : n74116;
  assign n74118 = pi15 ? n17325 : n17205;
  assign n74119 = pi14 ? n74118 : n40808;
  assign n74120 = pi15 ? n17216 : n16862;
  assign n74121 = pi15 ? n16862 : n16984;
  assign n74122 = pi14 ? n74120 : n74121;
  assign n74123 = pi13 ? n74119 : n74122;
  assign n74124 = pi12 ? n74123 : n32;
  assign n74125 = pi11 ? n74117 : n74124;
  assign n74126 = pi10 ? n74125 : n32;
  assign n74127 = pi09 ? n17493 : n74126;
  assign n74128 = pi08 ? n74102 : n74127;
  assign n74129 = pi13 ? n32 : n38860;
  assign n74130 = pi20 ? n2077 : n9000;
  assign n74131 = pi19 ? n32 : n74130;
  assign n74132 = pi18 ? n32 : n74131;
  assign n74133 = pi17 ? n32 : n74132;
  assign n74134 = pi16 ? n32 : n74133;
  assign n74135 = pi15 ? n17036 : n74134;
  assign n74136 = pi20 ? n101 : ~n2140;
  assign n74137 = pi19 ? n32 : n74136;
  assign n74138 = pi18 ? n32 : n74137;
  assign n74139 = pi17 ? n32 : n74138;
  assign n74140 = pi16 ? n32 : n74139;
  assign n74141 = pi15 ? n74140 : n32;
  assign n74142 = pi14 ? n74135 : n74141;
  assign n74143 = pi13 ? n74054 : n74142;
  assign n74144 = pi12 ? n74129 : n74143;
  assign n74145 = pi20 ? n428 : n1445;
  assign n74146 = pi19 ? n32 : n74145;
  assign n74147 = pi18 ? n32 : n74146;
  assign n74148 = pi17 ? n32 : n74147;
  assign n74149 = pi16 ? n32 : n74148;
  assign n74150 = pi15 ? n17205 : n74149;
  assign n74151 = pi15 ? n17188 : n74086;
  assign n74152 = pi14 ? n74150 : n74151;
  assign n74153 = pi15 ? n17056 : n17061;
  assign n74154 = pi15 ? n17121 : n17066;
  assign n74155 = pi14 ? n74153 : n74154;
  assign n74156 = pi13 ? n74152 : n74155;
  assign n74157 = pi12 ? n74156 : n17072;
  assign n74158 = pi11 ? n74144 : n74157;
  assign n74159 = pi10 ? n74158 : n32;
  assign n74160 = pi09 ? n17493 : n74159;
  assign n74161 = pi15 ? n16919 : n32;
  assign n74162 = pi14 ? n32 : n74161;
  assign n74163 = pi15 ? n32 : n74140;
  assign n74164 = pi14 ? n74163 : n74141;
  assign n74165 = pi13 ? n74162 : n74164;
  assign n74166 = pi12 ? n32 : n74165;
  assign n74167 = pi15 ? n17188 : n17216;
  assign n74168 = pi14 ? n74150 : n74167;
  assign n74169 = pi14 ? n74153 : n27880;
  assign n74170 = pi13 ? n74168 : n74169;
  assign n74171 = pi12 ? n74170 : n17102;
  assign n74172 = pi11 ? n74166 : n74171;
  assign n74173 = pi10 ? n74172 : n32;
  assign n74174 = pi09 ? n17493 : n74173;
  assign n74175 = pi08 ? n74160 : n74174;
  assign n74176 = pi07 ? n74128 : n74175;
  assign n74177 = pi15 ? n17128 : n32;
  assign n74178 = pi14 ? n32 : n74177;
  assign n74179 = pi15 ? n17193 : n17348;
  assign n74180 = pi14 ? n72676 : n74179;
  assign n74181 = pi13 ? n74178 : n74180;
  assign n74182 = pi12 ? n55942 : n74181;
  assign n74183 = pi15 ? n17251 : n17205;
  assign n74184 = pi14 ? n74183 : n17056;
  assign n74185 = pi15 ? n17228 : n17128;
  assign n74186 = pi14 ? n74185 : n17230;
  assign n74187 = pi13 ? n74184 : n74186;
  assign n74188 = pi12 ? n74187 : n32;
  assign n74189 = pi11 ? n74182 : n74188;
  assign n74190 = pi10 ? n74189 : n32;
  assign n74191 = pi09 ? n17493 : n74190;
  assign n74192 = pi14 ? n40847 : n17178;
  assign n74193 = pi15 ? n17278 : n17325;
  assign n74194 = pi14 ? n72676 : n74193;
  assign n74195 = pi13 ? n74192 : n74194;
  assign n74196 = pi12 ? n55942 : n74195;
  assign n74197 = pi14 ? n74183 : n17222;
  assign n74198 = pi13 ? n74197 : n17231;
  assign n74199 = pi12 ? n74198 : n32;
  assign n74200 = pi11 ? n74196 : n74199;
  assign n74201 = pi10 ? n74200 : n32;
  assign n74202 = pi09 ? n17493 : n74201;
  assign n74203 = pi08 ? n74191 : n74202;
  assign n74204 = pi14 ? n17271 : n32;
  assign n74205 = pi15 ? n17188 : n17193;
  assign n74206 = pi15 ? n17278 : n17152;
  assign n74207 = pi14 ? n74205 : n74206;
  assign n74208 = pi13 ? n74204 : n74207;
  assign n74209 = pi12 ? n32 : n74208;
  assign n74210 = pi15 ? n17331 : n17221;
  assign n74211 = pi14 ? n74183 : n74210;
  assign n74212 = pi13 ? n74211 : n17263;
  assign n74213 = pi12 ? n74212 : n32;
  assign n74214 = pi11 ? n74209 : n74213;
  assign n74215 = pi10 ? n74214 : n32;
  assign n74216 = pi09 ? n17493 : n74215;
  assign n74217 = pi14 ? n72676 : n17494;
  assign n74218 = pi13 ? n74204 : n74217;
  assign n74219 = pi12 ? n32 : n74218;
  assign n74220 = pi15 ? n17286 : n17363;
  assign n74221 = pi14 ? n74220 : n27909;
  assign n74222 = pi13 ? n74221 : n17301;
  assign n74223 = pi12 ? n74222 : n32;
  assign n74224 = pi11 ? n74219 : n74223;
  assign n74225 = pi10 ? n74224 : n32;
  assign n74226 = pi09 ? n17493 : n74225;
  assign n74227 = pi08 ? n74216 : n74226;
  assign n74228 = pi07 ? n74203 : n74227;
  assign n74229 = pi06 ? n74176 : n74228;
  assign n74230 = pi05 ? n74052 : n74229;
  assign n74231 = pi04 ? n73806 : n74230;
  assign n74232 = pi03 ? n72448 : n74231;
  assign n74233 = pi15 ? n17216 : n17261;
  assign n74234 = pi14 ? n27908 : n74233;
  assign n74235 = pi13 ? n74234 : n17301;
  assign n74236 = pi12 ? n74235 : n32;
  assign n74237 = pi11 ? n27970 : n74236;
  assign n74238 = pi10 ? n74237 : n32;
  assign n74239 = pi09 ? n17493 : n74238;
  assign n74240 = pi15 ? n17514 : n17205;
  assign n74241 = pi14 ? n17443 : n74240;
  assign n74242 = pi13 ? n32 : n74241;
  assign n74243 = pi12 ? n32 : n74242;
  assign n74244 = pi15 ? n17348 : n17331;
  assign n74245 = pi20 ? n32 : ~n15799;
  assign n74246 = pi19 ? n32 : n74245;
  assign n74247 = pi18 ? n32 : n74246;
  assign n74248 = pi17 ? n32 : n74247;
  assign n74249 = pi16 ? n32 : n74248;
  assign n74250 = pi15 ? n74249 : n17121;
  assign n74251 = pi14 ? n74244 : n74250;
  assign n74252 = pi13 ? n74251 : n27935;
  assign n74253 = pi12 ? n74252 : n32;
  assign n74254 = pi11 ? n74243 : n74253;
  assign n74255 = pi10 ? n74254 : n32;
  assign n74256 = pi09 ? n17493 : n74255;
  assign n74257 = pi07 ? n74239 : n74256;
  assign n74258 = pi14 ? n27770 : n74240;
  assign n74259 = pi13 ? n32 : n74258;
  assign n74260 = pi12 ? n32 : n74259;
  assign n74261 = pi11 ? n74260 : n74253;
  assign n74262 = pi10 ? n74261 : n32;
  assign n74263 = pi09 ? n17493 : n74262;
  assign n74264 = pi13 ? n74251 : n17413;
  assign n74265 = pi12 ? n74264 : n32;
  assign n74266 = pi11 ? n74260 : n74265;
  assign n74267 = pi10 ? n74266 : n32;
  assign n74268 = pi09 ? n17493 : n74267;
  assign n74269 = pi08 ? n74263 : n74268;
  assign n74270 = pi09 ? n17493 : n27945;
  assign n74271 = pi07 ? n74269 : n74270;
  assign n74272 = pi06 ? n74257 : n74271;
  assign n74273 = pi09 ? n17493 : n27958;
  assign n74274 = pi14 ? n27770 : n27928;
  assign n74275 = pi13 ? n32 : n74274;
  assign n74276 = pi12 ? n32 : n74275;
  assign n74277 = pi11 ? n74276 : n17473;
  assign n74278 = pi10 ? n74277 : n32;
  assign n74279 = pi09 ? n17493 : n74278;
  assign n74280 = pi11 ? n74276 : n17480;
  assign n74281 = pi10 ? n74280 : n32;
  assign n74282 = pi09 ? n17493 : n74281;
  assign n74283 = pi08 ? n74279 : n74282;
  assign n74284 = pi07 ? n74273 : n74283;
  assign n74285 = pi09 ? n17493 : n27972;
  assign n74286 = pi09 ? n17493 : n27975;
  assign n74287 = pi08 ? n74285 : n74286;
  assign n74288 = pi09 ? n17493 : n27983;
  assign n74289 = pi07 ? n74287 : n74288;
  assign n74290 = pi06 ? n74284 : n74289;
  assign n74291 = pi05 ? n74272 : n74290;
  assign n74292 = pi04 ? n74291 : n27998;
  assign n74293 = pi06 ? n32 : n55997;
  assign n74294 = pi05 ? n74293 : n17614;
  assign n74295 = pi16 ? n32 : n42505;
  assign n74296 = pi15 ? n32 : n74295;
  assign n74297 = pi14 ? n74296 : n32;
  assign n74298 = pi13 ? n32 : n74297;
  assign n74299 = pi12 ? n32 : n74298;
  assign n74300 = pi11 ? n32 : n74299;
  assign n74301 = pi10 ? n32 : n74300;
  assign n74302 = pi09 ? n74301 : n32;
  assign n74303 = pi07 ? n74302 : n32;
  assign n74304 = pi06 ? n74303 : n32;
  assign n74305 = pi05 ? n17614 : n74304;
  assign n74306 = pi04 ? n74294 : n74305;
  assign n74307 = pi03 ? n74292 : n74306;
  assign n74308 = pi02 ? n74232 : n74307;
  assign n74309 = pi06 ? n32 : n17586;
  assign n74310 = pi05 ? n32 : n74309;
  assign n74311 = pi18 ? n32 : n17927;
  assign n74312 = pi17 ? n32 : n74311;
  assign n74313 = pi16 ? n32 : n74312;
  assign n74314 = pi15 ? n32 : n74313;
  assign n74315 = pi14 ? n74314 : n32;
  assign n74316 = pi13 ? n32 : n74315;
  assign n74317 = pi12 ? n32 : n74316;
  assign n74318 = pi11 ? n32 : n74317;
  assign n74319 = pi10 ? n32 : n74318;
  assign n74320 = pi09 ? n74319 : n32;
  assign n74321 = pi07 ? n74320 : n17614;
  assign n74322 = pi06 ? n74321 : n17614;
  assign n74323 = pi05 ? n17568 : n74322;
  assign n74324 = pi04 ? n74310 : n74323;
  assign n74325 = pi06 ? n32 : n28005;
  assign n74326 = pi05 ? n74325 : n32;
  assign n74327 = pi04 ? n56006 : n74326;
  assign n74328 = pi03 ? n74324 : n74327;
  assign n74329 = pi02 ? n74328 : n32;
  assign n74330 = pi01 ? n74308 : n74329;
  assign n74331 = pi00 ? n67979 : n74330;
  assign n74332 = pi16 ? n1815 : ~n2144;
  assign n74333 = pi16 ? n1944 : ~n2144;
  assign n74334 = pi15 ? n74332 : n74333;
  assign n74335 = pi16 ? n3356 : ~n2144;
  assign n74336 = pi15 ? n74335 : n56012;
  assign n74337 = pi14 ? n74334 : n74336;
  assign n74338 = pi13 ? n32 : n74337;
  assign n74339 = pi16 ? n1581 : ~n2144;
  assign n74340 = pi15 ? n56014 : n74339;
  assign n74341 = pi14 ? n74340 : n56117;
  assign n74342 = pi14 ? n56019 : n43529;
  assign n74343 = pi13 ? n74341 : n74342;
  assign n74344 = pi12 ? n74338 : n74343;
  assign n74345 = pi14 ? n43529 : n57501;
  assign n74346 = pi15 ? n57501 : n43529;
  assign n74347 = pi14 ? n74346 : n43529;
  assign n74348 = pi13 ? n74345 : n74347;
  assign n74349 = pi15 ? n43529 : n43577;
  assign n74350 = pi14 ? n74349 : n43577;
  assign n74351 = pi15 ? n43577 : n57501;
  assign n74352 = pi14 ? n74351 : n57501;
  assign n74353 = pi13 ? n74350 : n74352;
  assign n74354 = pi12 ? n74348 : n74353;
  assign n74355 = pi11 ? n74344 : n74354;
  assign n74356 = pi14 ? n74346 : n57501;
  assign n74357 = pi13 ? n57501 : n74356;
  assign n74358 = pi14 ? n57501 : n56183;
  assign n74359 = pi13 ? n57501 : n74358;
  assign n74360 = pi12 ? n74357 : n74359;
  assign n74361 = pi16 ? n1233 : ~n1843;
  assign n74362 = pi14 ? n74361 : n29519;
  assign n74363 = pi13 ? n42585 : n74362;
  assign n74364 = pi12 ? n56183 : n74363;
  assign n74365 = pi11 ? n74360 : n74364;
  assign n74366 = pi10 ? n74355 : n74365;
  assign n74367 = pi09 ? n32 : n74366;
  assign n74368 = pi16 ? n2137 : ~n1834;
  assign n74369 = pi15 ? n32 : n74368;
  assign n74370 = pi14 ? n32 : n74369;
  assign n74371 = pi16 ? n1944 : ~n1834;
  assign n74372 = pi16 ? n3356 : ~n1834;
  assign n74373 = pi15 ? n74371 : n74372;
  assign n74374 = pi16 ? n1683 : ~n1834;
  assign n74375 = pi15 ? n74374 : n56014;
  assign n74376 = pi14 ? n74373 : n74375;
  assign n74377 = pi13 ? n74370 : n74376;
  assign n74378 = pi14 ? n56015 : n56019;
  assign n74379 = pi15 ? n56019 : n43577;
  assign n74380 = pi14 ? n74379 : n43577;
  assign n74381 = pi13 ? n74378 : n74380;
  assign n74382 = pi12 ? n74377 : n74381;
  assign n74383 = pi14 ? n58044 : n43529;
  assign n74384 = pi13 ? n43577 : n74383;
  assign n74385 = pi12 ? n43577 : n74384;
  assign n74386 = pi11 ? n74382 : n74385;
  assign n74387 = pi14 ? n74349 : n43529;
  assign n74388 = pi13 ? n43529 : n74387;
  assign n74389 = pi13 ? n43529 : n74345;
  assign n74390 = pi12 ? n74388 : n74389;
  assign n74391 = pi15 ? n30025 : n56183;
  assign n74392 = pi14 ? n57501 : n74391;
  assign n74393 = pi13 ? n74392 : n56183;
  assign n74394 = pi12 ? n74393 : n74363;
  assign n74395 = pi11 ? n74390 : n74394;
  assign n74396 = pi10 ? n74386 : n74395;
  assign n74397 = pi09 ? n32 : n74396;
  assign n74398 = pi08 ? n74367 : n74397;
  assign n74399 = pi07 ? n32 : n74398;
  assign n74400 = pi06 ? n32 : n74399;
  assign n74401 = pi16 ? n2137 : ~n1577;
  assign n74402 = pi15 ? n32 : n74401;
  assign n74403 = pi14 ? n32 : n74402;
  assign n74404 = pi16 ? n1944 : ~n1577;
  assign n74405 = pi16 ? n3356 : ~n1577;
  assign n74406 = pi15 ? n74404 : n74405;
  assign n74407 = pi16 ? n1683 : ~n1577;
  assign n74408 = pi15 ? n74407 : n56212;
  assign n74409 = pi14 ? n74406 : n74408;
  assign n74410 = pi13 ? n74403 : n74409;
  assign n74411 = pi15 ? n56214 : n56324;
  assign n74412 = pi14 ? n74411 : n56324;
  assign n74413 = pi13 ? n74412 : n19100;
  assign n74414 = pi12 ? n74410 : n74413;
  assign n74415 = pi14 ? n19100 : n58044;
  assign n74416 = pi13 ? n74415 : n19100;
  assign n74417 = pi14 ? n19100 : n43577;
  assign n74418 = pi13 ? n56330 : n74417;
  assign n74419 = pi12 ? n74416 : n74418;
  assign n74420 = pi11 ? n74414 : n74419;
  assign n74421 = pi14 ? n43577 : n43529;
  assign n74422 = pi13 ? n43577 : n74421;
  assign n74423 = pi12 ? n19100 : n74422;
  assign n74424 = pi15 ? n57501 : n30025;
  assign n74425 = pi14 ? n43529 : n74424;
  assign n74426 = pi13 ? n74425 : n30025;
  assign n74427 = pi14 ? n42585 : n74361;
  assign n74428 = pi13 ? n56183 : n74427;
  assign n74429 = pi12 ? n74426 : n74428;
  assign n74430 = pi11 ? n74423 : n74429;
  assign n74431 = pi10 ? n74420 : n74430;
  assign n74432 = pi09 ? n32 : n74431;
  assign n74433 = pi16 ? n1944 : ~n1683;
  assign n74434 = pi16 ? n2326 : ~n1683;
  assign n74435 = pi15 ? n74433 : n74434;
  assign n74436 = pi14 ? n32 : n74435;
  assign n74437 = pi16 ? n3356 : ~n1683;
  assign n74438 = pi16 ? n1683 : ~n1683;
  assign n74439 = pi15 ? n74437 : n74438;
  assign n74440 = pi15 ? n56212 : n56214;
  assign n74441 = pi14 ? n74439 : n74440;
  assign n74442 = pi13 ? n74436 : n74441;
  assign n74443 = pi15 ? n56324 : n19100;
  assign n74444 = pi14 ? n56324 : n74443;
  assign n74445 = pi13 ? n74444 : n56330;
  assign n74446 = pi12 ? n74442 : n74445;
  assign n74447 = pi14 ? n56330 : n43933;
  assign n74448 = pi14 ? n43933 : n19100;
  assign n74449 = pi13 ? n43933 : n74448;
  assign n74450 = pi12 ? n74447 : n74449;
  assign n74451 = pi11 ? n74446 : n74450;
  assign n74452 = pi13 ? n19100 : n74417;
  assign n74453 = pi12 ? n56330 : n74452;
  assign n74454 = pi15 ? n43577 : n43529;
  assign n74455 = pi14 ? n74454 : n74424;
  assign n74456 = pi13 ? n74455 : n30025;
  assign n74457 = pi12 ? n74456 : n74428;
  assign n74458 = pi11 ? n74453 : n74457;
  assign n74459 = pi10 ? n74451 : n74458;
  assign n74460 = pi09 ? n32 : n74459;
  assign n74461 = pi08 ? n74432 : n74460;
  assign n74462 = pi16 ? n1944 : ~n1678;
  assign n74463 = pi16 ? n2326 : ~n1678;
  assign n74464 = pi15 ? n74462 : n74463;
  assign n74465 = pi14 ? n32 : n74464;
  assign n74466 = pi16 ? n3356 : ~n1678;
  assign n74467 = pi16 ? n1683 : ~n1678;
  assign n74468 = pi15 ? n74466 : n74467;
  assign n74469 = pi16 ? n1834 : ~n3356;
  assign n74470 = pi15 ? n74469 : n56460;
  assign n74471 = pi14 ? n74468 : n74470;
  assign n74472 = pi13 ? n74465 : n74471;
  assign n74473 = pi14 ? n56462 : n43933;
  assign n74474 = pi13 ? n74473 : n43933;
  assign n74475 = pi12 ? n74472 : n74474;
  assign n74476 = pi15 ? n44289 : n43933;
  assign n74477 = pi14 ? n43933 : n74476;
  assign n74478 = pi14 ? n43933 : n44289;
  assign n74479 = pi13 ? n74477 : n74478;
  assign n74480 = pi15 ? n43787 : n44289;
  assign n74481 = pi14 ? n43787 : n74480;
  assign n74482 = pi14 ? n44289 : n43933;
  assign n74483 = pi13 ? n74481 : n74482;
  assign n74484 = pi12 ? n74479 : n74483;
  assign n74485 = pi11 ? n74475 : n74484;
  assign n74486 = pi15 ? n43933 : n56330;
  assign n74487 = pi14 ? n43933 : n74486;
  assign n74488 = pi13 ? n74487 : n56330;
  assign n74489 = pi15 ? n19100 : n56330;
  assign n74490 = pi14 ? n74489 : n19100;
  assign n74491 = pi13 ? n74490 : n74417;
  assign n74492 = pi12 ? n74488 : n74491;
  assign n74493 = pi15 ? n43529 : n57501;
  assign n74494 = pi14 ? n43577 : n74493;
  assign n74495 = pi13 ? n74494 : n57501;
  assign n74496 = pi15 ? n42585 : n74361;
  assign n74497 = pi14 ? n74391 : n74496;
  assign n74498 = pi13 ? n30025 : n74497;
  assign n74499 = pi12 ? n74495 : n74498;
  assign n74500 = pi11 ? n74492 : n74499;
  assign n74501 = pi10 ? n74485 : n74500;
  assign n74502 = pi09 ? n32 : n74501;
  assign n74503 = pi16 ? n2326 : ~n3356;
  assign n74504 = pi15 ? n32 : n74503;
  assign n74505 = pi16 ? n3352 : ~n3356;
  assign n74506 = pi16 ? n3356 : ~n3356;
  assign n74507 = pi15 ? n74505 : n74506;
  assign n74508 = pi14 ? n74504 : n74507;
  assign n74509 = pi16 ? n1683 : ~n3356;
  assign n74510 = pi15 ? n74509 : n74469;
  assign n74511 = pi15 ? n56460 : n56594;
  assign n74512 = pi14 ? n74510 : n74511;
  assign n74513 = pi13 ? n74508 : n74512;
  assign n74514 = pi15 ? n56462 : n44289;
  assign n74515 = pi14 ? n74514 : n44289;
  assign n74516 = pi15 ? n44289 : n43787;
  assign n74517 = pi14 ? n44289 : n74516;
  assign n74518 = pi13 ? n74515 : n74517;
  assign n74519 = pi12 ? n74513 : n74518;
  assign n74520 = pi14 ? n74516 : n43787;
  assign n74521 = pi13 ? n74520 : n43787;
  assign n74522 = pi15 ? n19778 : n43787;
  assign n74523 = pi14 ? n19778 : n74522;
  assign n74524 = pi14 ? n43787 : n44289;
  assign n74525 = pi13 ? n74523 : n74524;
  assign n74526 = pi12 ? n74521 : n74525;
  assign n74527 = pi11 ? n74519 : n74526;
  assign n74528 = pi14 ? n44289 : n74476;
  assign n74529 = pi13 ? n74528 : n43933;
  assign n74530 = pi14 ? n56330 : n19100;
  assign n74531 = pi13 ? n56330 : n74530;
  assign n74532 = pi12 ? n74529 : n74531;
  assign n74533 = pi14 ? n58044 : n74493;
  assign n74534 = pi13 ? n74533 : n57501;
  assign n74535 = pi14 ? n74391 : n42585;
  assign n74536 = pi13 ? n30025 : n74535;
  assign n74537 = pi12 ? n74534 : n74536;
  assign n74538 = pi11 ? n74532 : n74537;
  assign n74539 = pi10 ? n74527 : n74538;
  assign n74540 = pi09 ? n32 : n74539;
  assign n74541 = pi08 ? n74502 : n74540;
  assign n74542 = pi07 ? n74461 : n74541;
  assign n74543 = pi16 ? n2326 : ~n3352;
  assign n74544 = pi15 ? n32 : n74543;
  assign n74545 = pi16 ? n3352 : ~n3352;
  assign n74546 = pi16 ? n3356 : ~n3352;
  assign n74547 = pi15 ? n74545 : n74546;
  assign n74548 = pi14 ? n74544 : n74547;
  assign n74549 = pi16 ? n1683 : ~n3352;
  assign n74550 = pi16 ? n1834 : ~n2326;
  assign n74551 = pi15 ? n74549 : n74550;
  assign n74552 = pi16 ? n1581 : ~n2326;
  assign n74553 = pi15 ? n74552 : n56717;
  assign n74554 = pi14 ? n74551 : n74553;
  assign n74555 = pi13 ? n74548 : n74554;
  assign n74556 = pi15 ? n43787 : n19778;
  assign n74557 = pi14 ? n74556 : n19778;
  assign n74558 = pi14 ? n19778 : n43787;
  assign n74559 = pi13 ? n74557 : n74558;
  assign n74560 = pi12 ? n74555 : n74559;
  assign n74561 = pi13 ? n74557 : n19778;
  assign n74562 = pi13 ? n19778 : n74558;
  assign n74563 = pi12 ? n74561 : n74562;
  assign n74564 = pi11 ? n74560 : n74563;
  assign n74565 = pi14 ? n74480 : n74476;
  assign n74566 = pi15 ? n43933 : n44289;
  assign n74567 = pi14 ? n74566 : n43933;
  assign n74568 = pi13 ? n74565 : n74567;
  assign n74569 = pi15 ? n56330 : n43933;
  assign n74570 = pi14 ? n74569 : n56330;
  assign n74571 = pi13 ? n74570 : n74530;
  assign n74572 = pi12 ? n74568 : n74571;
  assign n74573 = pi14 ? n19100 : n43529;
  assign n74574 = pi13 ? n74573 : n43529;
  assign n74575 = pi15 ? n57501 : n56183;
  assign n74576 = pi14 ? n74575 : n42585;
  assign n74577 = pi13 ? n57501 : n74576;
  assign n74578 = pi12 ? n74574 : n74577;
  assign n74579 = pi11 ? n74572 : n74578;
  assign n74580 = pi10 ? n74564 : n74579;
  assign n74581 = pi09 ? n32 : n74580;
  assign n74582 = pi16 ? n3352 : ~n2326;
  assign n74583 = pi16 ? n3356 : ~n2326;
  assign n74584 = pi15 ? n74582 : n74583;
  assign n74585 = pi16 ? n1678 : ~n2326;
  assign n74586 = pi15 ? n74585 : n35161;
  assign n74587 = pi14 ? n74584 : n74586;
  assign n74588 = pi15 ? n74550 : n74552;
  assign n74589 = pi15 ? n56717 : n32185;
  assign n74590 = pi14 ? n74588 : n74589;
  assign n74591 = pi13 ? n74587 : n74590;
  assign n74592 = pi15 ? n19778 : n32185;
  assign n74593 = pi14 ? n74592 : n32185;
  assign n74594 = pi15 ? n44537 : n32185;
  assign n74595 = pi14 ? n32185 : n74594;
  assign n74596 = pi13 ? n74593 : n74595;
  assign n74597 = pi12 ? n74591 : n74596;
  assign n74598 = pi15 ? n32185 : n19778;
  assign n74599 = pi14 ? n44537 : n74598;
  assign n74600 = pi14 ? n19778 : n74592;
  assign n74601 = pi13 ? n74599 : n74600;
  assign n74602 = pi14 ? n32185 : n19778;
  assign n74603 = pi13 ? n74602 : n74558;
  assign n74604 = pi12 ? n74601 : n74603;
  assign n74605 = pi11 ? n74597 : n74604;
  assign n74606 = pi13 ? n74481 : n44289;
  assign n74607 = pi14 ? n43933 : n56330;
  assign n74608 = pi13 ? n43933 : n74607;
  assign n74609 = pi12 ? n74606 : n74608;
  assign n74610 = pi15 ? n56183 : n42585;
  assign n74611 = pi14 ? n74575 : n74610;
  assign n74612 = pi13 ? n57501 : n74611;
  assign n74613 = pi12 ? n74574 : n74612;
  assign n74614 = pi11 ? n74609 : n74613;
  assign n74615 = pi10 ? n74605 : n74614;
  assign n74616 = pi09 ? n32 : n74615;
  assign n74617 = pi08 ? n74581 : n74616;
  assign n74618 = pi16 ? n3352 : ~n1944;
  assign n74619 = pi16 ? n3356 : ~n1944;
  assign n74620 = pi15 ? n74618 : n74619;
  assign n74621 = pi16 ? n1678 : ~n1944;
  assign n74622 = pi16 ? n1683 : ~n1944;
  assign n74623 = pi15 ? n74621 : n74622;
  assign n74624 = pi14 ? n74620 : n74623;
  assign n74625 = pi16 ? n1834 : ~n2137;
  assign n74626 = pi16 ? n1581 : ~n2137;
  assign n74627 = pi15 ? n74625 : n74626;
  assign n74628 = pi16 ? n1594 : ~n1815;
  assign n74629 = pi15 ? n74628 : n44537;
  assign n74630 = pi14 ? n74627 : n74629;
  assign n74631 = pi13 ? n74624 : n74630;
  assign n74632 = pi15 ? n29601 : n44537;
  assign n74633 = pi14 ? n44537 : n74632;
  assign n74634 = pi13 ? n44537 : n74633;
  assign n74635 = pi12 ? n74631 : n74634;
  assign n74636 = pi14 ? n74632 : n74594;
  assign n74637 = pi13 ? n74636 : n32185;
  assign n74638 = pi13 ? n32185 : n74602;
  assign n74639 = pi12 ? n74637 : n74638;
  assign n74640 = pi11 ? n74635 : n74639;
  assign n74641 = pi14 ? n74522 : n74480;
  assign n74642 = pi13 ? n74641 : n44289;
  assign n74643 = pi12 ? n74642 : n74608;
  assign n74644 = pi14 ? n56330 : n43577;
  assign n74645 = pi13 ? n74644 : n43577;
  assign n74646 = pi14 ? n43786 : n56183;
  assign n74647 = pi13 ? n43529 : n74646;
  assign n74648 = pi12 ? n74645 : n74647;
  assign n74649 = pi11 ? n74643 : n74648;
  assign n74650 = pi10 ? n74640 : n74649;
  assign n74651 = pi09 ? n32 : n74650;
  assign n74652 = pi16 ? n3356 : ~n1808;
  assign n74653 = pi15 ? n32 : n74652;
  assign n74654 = pi14 ? n32 : n74653;
  assign n74655 = pi13 ? n32 : n74654;
  assign n74656 = pi12 ? n32 : n74655;
  assign n74657 = pi11 ? n32 : n74656;
  assign n74658 = pi10 ? n32 : n74657;
  assign n74659 = pi16 ? n1678 : ~n2137;
  assign n74660 = pi16 ? n1683 : ~n1815;
  assign n74661 = pi15 ? n74659 : n74660;
  assign n74662 = pi16 ? n1577 : ~n2137;
  assign n74663 = pi16 ? n1834 : ~n1815;
  assign n74664 = pi15 ? n74662 : n74663;
  assign n74665 = pi14 ? n74661 : n74664;
  assign n74666 = pi15 ? n74626 : n74628;
  assign n74667 = pi14 ? n74666 : n29601;
  assign n74668 = pi13 ? n74665 : n74667;
  assign n74669 = pi12 ? n74668 : n29601;
  assign n74670 = pi15 ? n32185 : n44537;
  assign n74671 = pi14 ? n32185 : n74670;
  assign n74672 = pi13 ? n74636 : n74671;
  assign n74673 = pi14 ? n44537 : n32185;
  assign n74674 = pi13 ? n74673 : n74602;
  assign n74675 = pi12 ? n74672 : n74674;
  assign n74676 = pi11 ? n74669 : n74675;
  assign n74677 = pi13 ? n74558 : n43787;
  assign n74678 = pi14 ? n74476 : n74486;
  assign n74679 = pi13 ? n44289 : n74678;
  assign n74680 = pi12 ? n74677 : n74679;
  assign n74681 = pi15 ? n56330 : n19100;
  assign n74682 = pi14 ? n74681 : n43577;
  assign n74683 = pi14 ? n43577 : n74454;
  assign n74684 = pi13 ? n74682 : n74683;
  assign n74685 = pi14 ? n74424 : n74391;
  assign n74686 = pi13 ? n43529 : n74685;
  assign n74687 = pi12 ? n74684 : n74686;
  assign n74688 = pi11 ? n74680 : n74687;
  assign n74689 = pi10 ? n74676 : n74688;
  assign n74690 = pi09 ? n74658 : n74689;
  assign n74691 = pi08 ? n74651 : n74690;
  assign n74692 = pi07 ? n74617 : n74691;
  assign n74693 = pi06 ? n74542 : n74692;
  assign n74694 = pi05 ? n74400 : n74693;
  assign n74695 = pi04 ? n32 : n74694;
  assign n74696 = pi16 ? n3356 : ~n3338;
  assign n74697 = pi15 ? n32 : n74696;
  assign n74698 = pi14 ? n32 : n74697;
  assign n74699 = pi13 ? n32 : n74698;
  assign n74700 = pi12 ? n32 : n74699;
  assign n74701 = pi11 ? n32 : n74700;
  assign n74702 = pi10 ? n32 : n74701;
  assign n74703 = pi16 ? n1678 : ~n1815;
  assign n74704 = pi15 ? n74703 : n31687;
  assign n74705 = pi16 ? n1577 : ~n1815;
  assign n74706 = pi16 ? n1834 : ~n1808;
  assign n74707 = pi15 ? n74705 : n74706;
  assign n74708 = pi14 ? n74704 : n74707;
  assign n74709 = pi16 ? n1581 : ~n1808;
  assign n74710 = pi16 ? n1594 : ~n1808;
  assign n74711 = pi15 ? n74709 : n74710;
  assign n74712 = pi14 ? n74711 : n29601;
  assign n74713 = pi13 ? n74708 : n74712;
  assign n74714 = pi13 ? n29601 : n57387;
  assign n74715 = pi12 ? n74713 : n74714;
  assign n74716 = pi15 ? n32806 : n29601;
  assign n74717 = pi14 ? n74716 : n74632;
  assign n74718 = pi13 ? n74717 : n44537;
  assign n74719 = pi13 ? n44537 : n74673;
  assign n74720 = pi12 ? n74718 : n74719;
  assign n74721 = pi11 ? n74715 : n74720;
  assign n74722 = pi14 ? n74476 : n43933;
  assign n74723 = pi13 ? n44289 : n74722;
  assign n74724 = pi12 ? n74677 : n74723;
  assign n74725 = pi14 ? n74486 : n19100;
  assign n74726 = pi13 ? n74725 : n74415;
  assign n74727 = pi14 ? n43786 : n30025;
  assign n74728 = pi13 ? n74683 : n74727;
  assign n74729 = pi12 ? n74726 : n74728;
  assign n74730 = pi11 ? n74724 : n74729;
  assign n74731 = pi10 ? n74721 : n74730;
  assign n74732 = pi09 ? n74702 : n74731;
  assign n74733 = pi16 ? n1678 : ~n3338;
  assign n74734 = pi16 ? n1683 : ~n3338;
  assign n74735 = pi15 ? n74733 : n74734;
  assign n74736 = pi14 ? n32 : n74735;
  assign n74737 = pi13 ? n32 : n74736;
  assign n74738 = pi12 ? n32 : n74737;
  assign n74739 = pi11 ? n32 : n74738;
  assign n74740 = pi10 ? n32 : n74739;
  assign n74741 = pi16 ? n1577 : ~n3338;
  assign n74742 = pi16 ? n1834 : ~n3338;
  assign n74743 = pi15 ? n74741 : n74742;
  assign n74744 = pi16 ? n2144 : ~n1808;
  assign n74745 = pi15 ? n74744 : n74709;
  assign n74746 = pi14 ? n74743 : n74745;
  assign n74747 = pi15 ? n74710 : n32806;
  assign n74748 = pi14 ? n74747 : n32806;
  assign n74749 = pi13 ? n74746 : n74748;
  assign n74750 = pi12 ? n74749 : n32806;
  assign n74751 = pi11 ? n74750 : n74720;
  assign n74752 = pi13 ? n74602 : n19778;
  assign n74753 = pi13 ? n43787 : n74565;
  assign n74754 = pi12 ? n74752 : n74753;
  assign n74755 = pi14 ? n74493 : n30025;
  assign n74756 = pi13 ? n74683 : n74755;
  assign n74757 = pi12 ? n74726 : n74756;
  assign n74758 = pi11 ? n74754 : n74757;
  assign n74759 = pi10 ? n74751 : n74758;
  assign n74760 = pi09 ? n74740 : n74759;
  assign n74761 = pi08 ? n74732 : n74760;
  assign n74762 = pi16 ? n1678 : ~n2540;
  assign n74763 = pi15 ? n74762 : n31857;
  assign n74764 = pi14 ? n32 : n74763;
  assign n74765 = pi13 ? n32 : n74764;
  assign n74766 = pi12 ? n32 : n74765;
  assign n74767 = pi11 ? n32 : n74766;
  assign n74768 = pi10 ? n32 : n74767;
  assign n74769 = pi16 ? n1577 : ~n2540;
  assign n74770 = pi16 ? n1834 : ~n2540;
  assign n74771 = pi15 ? n74769 : n74770;
  assign n74772 = pi16 ? n2144 : ~n3338;
  assign n74773 = pi16 ? n1581 : ~n3338;
  assign n74774 = pi15 ? n74772 : n74773;
  assign n74775 = pi14 ? n74771 : n74774;
  assign n74776 = pi16 ? n1594 : ~n3338;
  assign n74777 = pi15 ? n74776 : n32806;
  assign n74778 = pi14 ? n74777 : n32806;
  assign n74779 = pi13 ? n74775 : n74778;
  assign n74780 = pi15 ? n32806 : n57596;
  assign n74781 = pi14 ? n32806 : n74780;
  assign n74782 = pi13 ? n32806 : n74781;
  assign n74783 = pi12 ? n74779 : n74782;
  assign n74784 = pi15 ? n57596 : n32806;
  assign n74785 = pi14 ? n74784 : n74716;
  assign n74786 = pi13 ? n74785 : n29601;
  assign n74787 = pi13 ? n29601 : n57151;
  assign n74788 = pi12 ? n74786 : n74787;
  assign n74789 = pi11 ? n74783 : n74788;
  assign n74790 = pi14 ? n74480 : n44289;
  assign n74791 = pi13 ? n43787 : n74790;
  assign n74792 = pi12 ? n74752 : n74791;
  assign n74793 = pi14 ? n74476 : n56330;
  assign n74794 = pi14 ? n56330 : n74681;
  assign n74795 = pi13 ? n74793 : n74794;
  assign n74796 = pi14 ? n74493 : n57501;
  assign n74797 = pi13 ? n74415 : n74796;
  assign n74798 = pi12 ? n74795 : n74797;
  assign n74799 = pi11 ? n74792 : n74798;
  assign n74800 = pi10 ? n74789 : n74799;
  assign n74801 = pi09 ? n74768 : n74800;
  assign n74802 = pi15 ? n32 : n31857;
  assign n74803 = pi14 ? n74802 : n74771;
  assign n74804 = pi13 ? n32 : n74803;
  assign n74805 = pi12 ? n32 : n74804;
  assign n74806 = pi11 ? n32 : n74805;
  assign n74807 = pi10 ? n32 : n74806;
  assign n74808 = pi16 ? n2144 : ~n2540;
  assign n74809 = pi16 ? n1581 : ~n2540;
  assign n74810 = pi15 ? n74808 : n74809;
  assign n74811 = pi16 ? n1323 : ~n3338;
  assign n74812 = pi15 ? n74811 : n74776;
  assign n74813 = pi14 ? n74810 : n74812;
  assign n74814 = pi14 ? n74780 : n57596;
  assign n74815 = pi13 ? n74813 : n74814;
  assign n74816 = pi12 ? n74815 : n57596;
  assign n74817 = pi11 ? n74816 : n74788;
  assign n74818 = pi13 ? n74673 : n32185;
  assign n74819 = pi13 ? n19778 : n74481;
  assign n74820 = pi12 ? n74818 : n74819;
  assign n74821 = pi14 ? n74454 : n57501;
  assign n74822 = pi13 ? n19100 : n74821;
  assign n74823 = pi12 ? n74795 : n74822;
  assign n74824 = pi11 ? n74820 : n74823;
  assign n74825 = pi10 ? n74817 : n74824;
  assign n74826 = pi09 ? n74807 : n74825;
  assign n74827 = pi08 ? n74801 : n74826;
  assign n74828 = pi07 ? n74761 : n74827;
  assign n74829 = pi16 ? n1683 : ~n2320;
  assign n74830 = pi15 ? n32 : n74829;
  assign n74831 = pi16 ? n1577 : ~n2320;
  assign n74832 = pi16 ? n1834 : ~n2320;
  assign n74833 = pi15 ? n74831 : n74832;
  assign n74834 = pi14 ? n74830 : n74833;
  assign n74835 = pi13 ? n32 : n74834;
  assign n74836 = pi12 ? n32 : n74835;
  assign n74837 = pi11 ? n32 : n74836;
  assign n74838 = pi10 ? n32 : n74837;
  assign n74839 = pi16 ? n2144 : ~n2320;
  assign n74840 = pi16 ? n1581 : ~n2320;
  assign n74841 = pi15 ? n74839 : n74840;
  assign n74842 = pi16 ? n1323 : ~n2540;
  assign n74843 = pi16 ? n1594 : ~n2540;
  assign n74844 = pi15 ? n74842 : n74843;
  assign n74845 = pi14 ? n74841 : n74844;
  assign n74846 = pi13 ? n74845 : n57596;
  assign n74847 = pi14 ? n57596 : n57755;
  assign n74848 = pi13 ? n57596 : n74847;
  assign n74849 = pi12 ? n74846 : n74848;
  assign n74850 = pi15 ? n57695 : n57596;
  assign n74851 = pi14 ? n74850 : n74784;
  assign n74852 = pi13 ? n74851 : n32806;
  assign n74853 = pi14 ? n32806 : n29601;
  assign n74854 = pi13 ? n32806 : n74853;
  assign n74855 = pi12 ? n74852 : n74854;
  assign n74856 = pi11 ? n74849 : n74855;
  assign n74857 = pi13 ? n19778 : n43787;
  assign n74858 = pi12 ? n74818 : n74857;
  assign n74859 = pi14 ? n74480 : n43933;
  assign n74860 = pi13 ? n74859 : n74487;
  assign n74861 = pi14 ? n74454 : n43529;
  assign n74862 = pi13 ? n74794 : n74861;
  assign n74863 = pi12 ? n74860 : n74862;
  assign n74864 = pi11 ? n74858 : n74863;
  assign n74865 = pi10 ? n74856 : n74864;
  assign n74866 = pi09 ? n74838 : n74865;
  assign n74867 = pi15 ? n32 : n74831;
  assign n74868 = pi15 ? n74832 : n74839;
  assign n74869 = pi14 ? n74867 : n74868;
  assign n74870 = pi13 ? n32 : n74869;
  assign n74871 = pi12 ? n32 : n74870;
  assign n74872 = pi11 ? n32 : n74871;
  assign n74873 = pi10 ? n32 : n74872;
  assign n74874 = pi16 ? n1323 : ~n2320;
  assign n74875 = pi15 ? n74840 : n74874;
  assign n74876 = pi16 ? n1843 : ~n2540;
  assign n74877 = pi15 ? n74843 : n74876;
  assign n74878 = pi14 ? n74875 : n74877;
  assign n74879 = pi13 ? n74878 : n57755;
  assign n74880 = pi12 ? n74879 : n57695;
  assign n74881 = pi11 ? n74880 : n74855;
  assign n74882 = pi13 ? n57151 : n44537;
  assign n74883 = pi13 ? n32185 : n74523;
  assign n74884 = pi12 ? n74882 : n74883;
  assign n74885 = pi13 ? n74794 : n74383;
  assign n74886 = pi12 ? n74860 : n74885;
  assign n74887 = pi11 ? n74884 : n74886;
  assign n74888 = pi10 ? n74881 : n74887;
  assign n74889 = pi09 ? n74873 : n74888;
  assign n74890 = pi08 ? n74866 : n74889;
  assign n74891 = pi16 ? n1577 : ~n1934;
  assign n74892 = pi15 ? n32 : n74891;
  assign n74893 = pi16 ? n1834 : ~n1934;
  assign n74894 = pi16 ? n2144 : ~n1934;
  assign n74895 = pi15 ? n74893 : n74894;
  assign n74896 = pi14 ? n74892 : n74895;
  assign n74897 = pi13 ? n32 : n74896;
  assign n74898 = pi12 ? n32 : n74897;
  assign n74899 = pi11 ? n32 : n74898;
  assign n74900 = pi10 ? n32 : n74899;
  assign n74901 = pi16 ? n1581 : ~n1934;
  assign n74902 = pi16 ? n1323 : ~n1934;
  assign n74903 = pi15 ? n74901 : n74902;
  assign n74904 = pi16 ? n1594 : ~n2320;
  assign n74905 = pi16 ? n1843 : ~n2320;
  assign n74906 = pi15 ? n74904 : n74905;
  assign n74907 = pi14 ? n74903 : n74906;
  assign n74908 = pi13 ? n74907 : n57695;
  assign n74909 = pi14 ? n57695 : n45572;
  assign n74910 = pi13 ? n57695 : n74909;
  assign n74911 = pi12 ? n74908 : n74910;
  assign n74912 = pi14 ? n58990 : n74850;
  assign n74913 = pi13 ? n74912 : n57596;
  assign n74914 = pi14 ? n57596 : n32806;
  assign n74915 = pi13 ? n57596 : n74914;
  assign n74916 = pi12 ? n74913 : n74915;
  assign n74917 = pi11 ? n74911 : n74916;
  assign n74918 = pi14 ? n74598 : n19778;
  assign n74919 = pi13 ? n32185 : n74918;
  assign n74920 = pi12 ? n74882 : n74919;
  assign n74921 = pi14 ? n74522 : n44289;
  assign n74922 = pi13 ? n74921 : n74528;
  assign n74923 = pi14 ? n58044 : n74454;
  assign n74924 = pi13 ? n74487 : n74923;
  assign n74925 = pi12 ? n74922 : n74924;
  assign n74926 = pi11 ? n74920 : n74925;
  assign n74927 = pi10 ? n74917 : n74926;
  assign n74928 = pi09 ? n74900 : n74927;
  assign n74929 = pi15 ? n32 : n74893;
  assign n74930 = pi15 ? n74894 : n74901;
  assign n74931 = pi14 ? n74929 : n74930;
  assign n74932 = pi13 ? n32 : n74931;
  assign n74933 = pi12 ? n32 : n74932;
  assign n74934 = pi11 ? n32 : n74933;
  assign n74935 = pi10 ? n32 : n74934;
  assign n74936 = pi16 ? n1594 : ~n1934;
  assign n74937 = pi15 ? n74902 : n74936;
  assign n74938 = pi16 ? n1471 : ~n2320;
  assign n74939 = pi15 ? n74905 : n74938;
  assign n74940 = pi14 ? n74937 : n74939;
  assign n74941 = pi15 ? n57695 : n45572;
  assign n74942 = pi13 ? n74940 : n74941;
  assign n74943 = pi12 ? n74942 : n45572;
  assign n74944 = pi14 ? n74784 : n74780;
  assign n74945 = pi13 ? n57596 : n74944;
  assign n74946 = pi12 ? n74913 : n74945;
  assign n74947 = pi11 ? n74943 : n74946;
  assign n74948 = pi13 ? n74853 : n29601;
  assign n74949 = pi14 ? n32185 : n74598;
  assign n74950 = pi13 ? n44537 : n74949;
  assign n74951 = pi12 ? n74948 : n74950;
  assign n74952 = pi15 ? n56330 : n43577;
  assign n74953 = pi14 ? n74952 : n74454;
  assign n74954 = pi13 ? n74487 : n74953;
  assign n74955 = pi12 ? n74922 : n74954;
  assign n74956 = pi11 ? n74951 : n74955;
  assign n74957 = pi10 ? n74947 : n74956;
  assign n74958 = pi09 ? n74935 : n74957;
  assign n74959 = pi08 ? n74928 : n74958;
  assign n74960 = pi07 ? n74890 : n74959;
  assign n74961 = pi06 ? n74828 : n74960;
  assign n74962 = pi16 ? n1834 : ~n2306;
  assign n74963 = pi15 ? n32 : n74962;
  assign n74964 = pi16 ? n2144 : ~n2306;
  assign n74965 = pi16 ? n1581 : ~n2306;
  assign n74966 = pi15 ? n74964 : n74965;
  assign n74967 = pi14 ? n74963 : n74966;
  assign n74968 = pi13 ? n32 : n74967;
  assign n74969 = pi12 ? n32 : n74968;
  assign n74970 = pi11 ? n32 : n74969;
  assign n74971 = pi10 ? n32 : n74970;
  assign n74972 = pi16 ? n1323 : ~n2306;
  assign n74973 = pi16 ? n1594 : ~n2306;
  assign n74974 = pi15 ? n74972 : n74973;
  assign n74975 = pi16 ? n1843 : ~n1934;
  assign n74976 = pi16 ? n1471 : ~n1934;
  assign n74977 = pi15 ? n74975 : n74976;
  assign n74978 = pi14 ? n74974 : n74977;
  assign n74979 = pi13 ? n74978 : n45572;
  assign n74980 = pi14 ? n45572 : n58074;
  assign n74981 = pi13 ? n45572 : n74980;
  assign n74982 = pi12 ? n74979 : n74981;
  assign n74983 = pi15 ? n58074 : n45572;
  assign n74984 = pi14 ? n74983 : n58990;
  assign n74985 = pi13 ? n74984 : n57695;
  assign n74986 = pi14 ? n74850 : n57596;
  assign n74987 = pi13 ? n57695 : n74986;
  assign n74988 = pi12 ? n74985 : n74987;
  assign n74989 = pi11 ? n74982 : n74988;
  assign n74990 = pi14 ? n74594 : n32185;
  assign n74991 = pi13 ? n44537 : n74990;
  assign n74992 = pi12 ? n74948 : n74991;
  assign n74993 = pi13 ? n74558 : n74481;
  assign n74994 = pi14 ? n44289 : n74486;
  assign n74995 = pi14 ? n74681 : n58044;
  assign n74996 = pi13 ? n74994 : n74995;
  assign n74997 = pi12 ? n74993 : n74996;
  assign n74998 = pi11 ? n74992 : n74997;
  assign n74999 = pi10 ? n74989 : n74998;
  assign n75000 = pi09 ? n74971 : n74999;
  assign n75001 = pi15 ? n32 : n74964;
  assign n75002 = pi15 ? n74965 : n74972;
  assign n75003 = pi14 ? n75001 : n75002;
  assign n75004 = pi13 ? n32 : n75003;
  assign n75005 = pi12 ? n32 : n75004;
  assign n75006 = pi11 ? n32 : n75005;
  assign n75007 = pi10 ? n32 : n75006;
  assign n75008 = pi16 ? n1843 : ~n2306;
  assign n75009 = pi15 ? n74973 : n75008;
  assign n75010 = pi16 ? n1479 : ~n1934;
  assign n75011 = pi15 ? n74976 : n75010;
  assign n75012 = pi14 ? n75009 : n75011;
  assign n75013 = pi15 ? n45572 : n58074;
  assign n75014 = pi14 ? n45572 : n75013;
  assign n75015 = pi13 ? n75012 : n75014;
  assign n75016 = pi12 ? n75015 : n58074;
  assign n75017 = pi14 ? n57695 : n74941;
  assign n75018 = pi14 ? n57695 : n57755;
  assign n75019 = pi13 ? n75017 : n75018;
  assign n75020 = pi12 ? n74985 : n75019;
  assign n75021 = pi11 ? n75016 : n75020;
  assign n75022 = pi13 ? n74914 : n32806;
  assign n75023 = pi13 ? n29601 : n74673;
  assign n75024 = pi12 ? n75022 : n75023;
  assign n75025 = pi15 ? n43933 : n19100;
  assign n75026 = pi14 ? n75025 : n58044;
  assign n75027 = pi13 ? n74482 : n75026;
  assign n75028 = pi12 ? n74993 : n75027;
  assign n75029 = pi11 ? n75024 : n75028;
  assign n75030 = pi10 ? n75021 : n75029;
  assign n75031 = pi09 ? n75007 : n75030;
  assign n75032 = pi08 ? n75000 : n75031;
  assign n75033 = pi16 ? n2144 : ~n2530;
  assign n75034 = pi15 ? n32 : n75033;
  assign n75035 = pi16 ? n1323 : ~n2530;
  assign n75036 = pi15 ? n30386 : n75035;
  assign n75037 = pi14 ? n75034 : n75036;
  assign n75038 = pi13 ? n32 : n75037;
  assign n75039 = pi12 ? n32 : n75038;
  assign n75040 = pi11 ? n32 : n75039;
  assign n75041 = pi10 ? n32 : n75040;
  assign n75042 = pi16 ? n1594 : ~n2530;
  assign n75043 = pi16 ? n1843 : ~n2530;
  assign n75044 = pi15 ? n75042 : n75043;
  assign n75045 = pi16 ? n1471 : ~n2306;
  assign n75046 = pi16 ? n1479 : ~n2306;
  assign n75047 = pi15 ? n75045 : n75046;
  assign n75048 = pi14 ? n75044 : n75047;
  assign n75049 = pi13 ? n75048 : n58074;
  assign n75050 = pi14 ? n58074 : n46354;
  assign n75051 = pi13 ? n58074 : n75050;
  assign n75052 = pi12 ? n75049 : n75051;
  assign n75053 = pi14 ? n46354 : n74983;
  assign n75054 = pi13 ? n75053 : n45572;
  assign n75055 = pi14 ? n58990 : n57695;
  assign n75056 = pi13 ? n45572 : n75055;
  assign n75057 = pi12 ? n75054 : n75056;
  assign n75058 = pi11 ? n75052 : n75057;
  assign n75059 = pi13 ? n29601 : n44537;
  assign n75060 = pi12 ? n75022 : n75059;
  assign n75061 = pi13 ? n74602 : n74523;
  assign n75062 = pi13 ? n74859 : n74725;
  assign n75063 = pi12 ? n75061 : n75062;
  assign n75064 = pi11 ? n75060 : n75063;
  assign n75065 = pi10 ? n75058 : n75064;
  assign n75066 = pi09 ? n75041 : n75065;
  assign n75067 = pi15 ? n32 : n30386;
  assign n75068 = pi15 ? n75035 : n75042;
  assign n75069 = pi14 ? n75067 : n75068;
  assign n75070 = pi13 ? n32 : n75069;
  assign n75071 = pi12 ? n32 : n75070;
  assign n75072 = pi11 ? n32 : n75071;
  assign n75073 = pi10 ? n32 : n75072;
  assign n75074 = pi16 ? n1471 : ~n2530;
  assign n75075 = pi15 ? n75043 : n75074;
  assign n75076 = pi16 ? n1705 : ~n2306;
  assign n75077 = pi15 ? n75046 : n75076;
  assign n75078 = pi14 ? n75075 : n75077;
  assign n75079 = pi13 ? n75078 : n75050;
  assign n75080 = pi12 ? n75079 : n46354;
  assign n75081 = pi15 ? n46354 : n58074;
  assign n75082 = pi14 ? n75081 : n74983;
  assign n75083 = pi13 ? n75082 : n45572;
  assign n75084 = pi14 ? n45572 : n74941;
  assign n75085 = pi13 ? n75014 : n75084;
  assign n75086 = pi12 ? n75083 : n75085;
  assign n75087 = pi11 ? n75080 : n75086;
  assign n75088 = pi14 ? n57695 : n57596;
  assign n75089 = pi13 ? n75088 : n57596;
  assign n75090 = pi13 ? n32806 : n57151;
  assign n75091 = pi12 ? n75089 : n75090;
  assign n75092 = pi13 ? n74524 : n74725;
  assign n75093 = pi12 ? n75061 : n75092;
  assign n75094 = pi11 ? n75091 : n75093;
  assign n75095 = pi10 ? n75087 : n75094;
  assign n75096 = pi09 ? n75073 : n75095;
  assign n75097 = pi08 ? n75066 : n75096;
  assign n75098 = pi07 ? n75032 : n75097;
  assign n75099 = pi15 ? n32 : n30490;
  assign n75100 = pi16 ? n1323 : ~n2300;
  assign n75101 = pi15 ? n75100 : n30565;
  assign n75102 = pi14 ? n75099 : n75101;
  assign n75103 = pi13 ? n32 : n75102;
  assign n75104 = pi12 ? n32 : n75103;
  assign n75105 = pi11 ? n32 : n75104;
  assign n75106 = pi10 ? n32 : n75105;
  assign n75107 = pi16 ? n1843 : ~n2300;
  assign n75108 = pi16 ? n1471 : ~n2300;
  assign n75109 = pi15 ? n75107 : n75108;
  assign n75110 = pi16 ? n1479 : ~n2530;
  assign n75111 = pi15 ? n75110 : n58318;
  assign n75112 = pi14 ? n75109 : n75111;
  assign n75113 = pi13 ? n75112 : n46354;
  assign n75114 = pi14 ? n46354 : n58400;
  assign n75115 = pi13 ? n46354 : n75114;
  assign n75116 = pi12 ? n75113 : n75115;
  assign n75117 = pi15 ? n58400 : n46354;
  assign n75118 = pi14 ? n75117 : n75081;
  assign n75119 = pi13 ? n75118 : n58074;
  assign n75120 = pi13 ? n58074 : n74984;
  assign n75121 = pi12 ? n75119 : n75120;
  assign n75122 = pi11 ? n75116 : n75121;
  assign n75123 = pi13 ? n74986 : n57596;
  assign n75124 = pi14 ? n32806 : n74716;
  assign n75125 = pi14 ? n29601 : n74632;
  assign n75126 = pi13 ? n75124 : n75125;
  assign n75127 = pi12 ? n75123 : n75126;
  assign n75128 = pi14 ? n74486 : n56330;
  assign n75129 = pi13 ? n74921 : n75128;
  assign n75130 = pi12 ? n74674 : n75129;
  assign n75131 = pi11 ? n75127 : n75130;
  assign n75132 = pi10 ? n75122 : n75131;
  assign n75133 = pi09 ? n75106 : n75132;
  assign n75134 = pi15 ? n32 : n75100;
  assign n75135 = pi15 ? n30565 : n75107;
  assign n75136 = pi14 ? n75134 : n75135;
  assign n75137 = pi13 ? n32 : n75136;
  assign n75138 = pi12 ? n32 : n75137;
  assign n75139 = pi11 ? n32 : n75138;
  assign n75140 = pi10 ? n32 : n75139;
  assign n75141 = pi16 ? n1479 : ~n2300;
  assign n75142 = pi15 ? n75108 : n75141;
  assign n75143 = pi16 ? n1972 : ~n2530;
  assign n75144 = pi15 ? n58318 : n75143;
  assign n75145 = pi14 ? n75142 : n75144;
  assign n75146 = pi13 ? n75145 : n75114;
  assign n75147 = pi12 ? n75146 : n58400;
  assign n75148 = pi14 ? n74983 : n45572;
  assign n75149 = pi13 ? n58074 : n75148;
  assign n75150 = pi12 ? n75119 : n75149;
  assign n75151 = pi11 ? n75147 : n75150;
  assign n75152 = pi13 ? n75055 : n57695;
  assign n75153 = pi14 ? n57596 : n74784;
  assign n75154 = pi13 ? n75153 : n74717;
  assign n75155 = pi12 ? n75152 : n75154;
  assign n75156 = pi13 ? n74641 : n74722;
  assign n75157 = pi12 ? n74674 : n75156;
  assign n75158 = pi11 ? n75155 : n75157;
  assign n75159 = pi10 ? n75151 : n75158;
  assign n75160 = pi09 ? n75140 : n75159;
  assign n75161 = pi08 ? n75133 : n75160;
  assign n75162 = pi16 ? n1323 : ~n3625;
  assign n75163 = pi15 ? n32 : n75162;
  assign n75164 = pi16 ? n1843 : ~n3625;
  assign n75165 = pi15 ? n30679 : n75164;
  assign n75166 = pi14 ? n75163 : n75165;
  assign n75167 = pi13 ? n32 : n75166;
  assign n75168 = pi12 ? n32 : n75167;
  assign n75169 = pi11 ? n32 : n75168;
  assign n75170 = pi10 ? n32 : n75169;
  assign n75171 = pi16 ? n1471 : ~n3625;
  assign n75172 = pi16 ? n1479 : ~n3625;
  assign n75173 = pi15 ? n75171 : n75172;
  assign n75174 = pi16 ? n1972 : ~n2300;
  assign n75175 = pi15 ? n58576 : n75174;
  assign n75176 = pi14 ? n75173 : n75175;
  assign n75177 = pi13 ? n75176 : n58400;
  assign n75178 = pi14 ? n58400 : n35359;
  assign n75179 = pi13 ? n58400 : n75178;
  assign n75180 = pi12 ? n75177 : n75179;
  assign n75181 = pi15 ? n35359 : n58400;
  assign n75182 = pi14 ? n75181 : n75117;
  assign n75183 = pi13 ? n75182 : n46354;
  assign n75184 = pi13 ? n46354 : n75082;
  assign n75185 = pi12 ? n75183 : n75184;
  assign n75186 = pi11 ? n75180 : n75185;
  assign n75187 = pi13 ? n75153 : n74853;
  assign n75188 = pi12 ? n75152 : n75187;
  assign n75189 = pi13 ? n57151 : n74673;
  assign n75190 = pi13 ? n74558 : n74790;
  assign n75191 = pi12 ? n75189 : n75190;
  assign n75192 = pi11 ? n75188 : n75191;
  assign n75193 = pi10 ? n75186 : n75192;
  assign n75194 = pi09 ? n75170 : n75193;
  assign n75195 = pi15 ? n32 : n30679;
  assign n75196 = pi15 ? n75164 : n75171;
  assign n75197 = pi14 ? n75195 : n75196;
  assign n75198 = pi13 ? n32 : n75197;
  assign n75199 = pi12 ? n32 : n75198;
  assign n75200 = pi11 ? n32 : n75199;
  assign n75201 = pi10 ? n32 : n75200;
  assign n75202 = pi15 ? n75172 : n58576;
  assign n75203 = pi16 ? n1972 : ~n3625;
  assign n75204 = pi15 ? n75203 : n58396;
  assign n75205 = pi14 ? n75202 : n75204;
  assign n75206 = pi13 ? n75205 : n75178;
  assign n75207 = pi12 ? n75206 : n35359;
  assign n75208 = pi14 ? n75081 : n58074;
  assign n75209 = pi13 ? n46354 : n75208;
  assign n75210 = pi12 ? n75183 : n75209;
  assign n75211 = pi11 ? n75207 : n75210;
  assign n75212 = pi13 ? n75148 : n45572;
  assign n75213 = pi14 ? n57695 : n74850;
  assign n75214 = pi14 ? n74784 : n32806;
  assign n75215 = pi13 ? n75213 : n75214;
  assign n75216 = pi12 ? n75212 : n75215;
  assign n75217 = pi13 ? n74853 : n57151;
  assign n75218 = pi14 ? n74598 : n74522;
  assign n75219 = pi13 ? n75218 : n74790;
  assign n75220 = pi12 ? n75217 : n75219;
  assign n75221 = pi11 ? n75216 : n75220;
  assign n75222 = pi10 ? n75211 : n75221;
  assign n75223 = pi09 ? n75201 : n75222;
  assign n75224 = pi08 ? n75194 : n75223;
  assign n75225 = pi07 ? n75161 : n75224;
  assign n75226 = pi06 ? n75098 : n75225;
  assign n75227 = pi05 ? n74961 : n75226;
  assign n75228 = pi16 ? n1594 : ~n3788;
  assign n75229 = pi15 ? n32 : n75228;
  assign n75230 = pi16 ? n1843 : ~n3788;
  assign n75231 = pi16 ? n1471 : ~n3788;
  assign n75232 = pi15 ? n75230 : n75231;
  assign n75233 = pi14 ? n75229 : n75232;
  assign n75234 = pi13 ? n32 : n75233;
  assign n75235 = pi12 ? n32 : n75234;
  assign n75236 = pi11 ? n32 : n75235;
  assign n75237 = pi10 ? n32 : n75236;
  assign n75238 = pi16 ? n1479 : ~n3788;
  assign n75239 = pi16 ? n1705 : ~n3788;
  assign n75240 = pi15 ? n75238 : n75239;
  assign n75241 = pi16 ? n1972 : ~n3788;
  assign n75242 = pi15 ? n75241 : n47261;
  assign n75243 = pi14 ? n75240 : n75242;
  assign n75244 = pi13 ? n75243 : n35359;
  assign n75245 = pi14 ? n35359 : n58837;
  assign n75246 = pi13 ? n35359 : n75245;
  assign n75247 = pi12 ? n75244 : n75246;
  assign n75248 = pi15 ? n58837 : n35359;
  assign n75249 = pi14 ? n75248 : n75181;
  assign n75250 = pi13 ? n75249 : n58400;
  assign n75251 = pi13 ? n58400 : n75118;
  assign n75252 = pi12 ? n75250 : n75251;
  assign n75253 = pi11 ? n75247 : n75252;
  assign n75254 = pi13 ? n75213 : n57596;
  assign n75255 = pi12 ? n75212 : n75254;
  assign n75256 = pi14 ? n32806 : n74632;
  assign n75257 = pi13 ? n74914 : n75256;
  assign n75258 = pi14 ? n74594 : n74598;
  assign n75259 = pi14 ? n74522 : n43787;
  assign n75260 = pi13 ? n75258 : n75259;
  assign n75261 = pi12 ? n75257 : n75260;
  assign n75262 = pi11 ? n75255 : n75261;
  assign n75263 = pi10 ? n75253 : n75262;
  assign n75264 = pi09 ? n75237 : n75263;
  assign n75265 = pi15 ? n32 : n75230;
  assign n75266 = pi15 ? n75231 : n75238;
  assign n75267 = pi14 ? n75265 : n75266;
  assign n75268 = pi13 ? n32 : n75267;
  assign n75269 = pi12 ? n32 : n75268;
  assign n75270 = pi11 ? n32 : n75269;
  assign n75271 = pi10 ? n32 : n75270;
  assign n75272 = pi15 ? n75239 : n75241;
  assign n75273 = pi16 ? n1214 : ~n3788;
  assign n75274 = pi16 ? n931 : ~n3625;
  assign n75275 = pi15 ? n75273 : n75274;
  assign n75276 = pi14 ? n75272 : n75275;
  assign n75277 = pi13 ? n75276 : n75245;
  assign n75278 = pi12 ? n75277 : n58837;
  assign n75279 = pi14 ? n58400 : n75181;
  assign n75280 = pi13 ? n75279 : n75117;
  assign n75281 = pi12 ? n75250 : n75280;
  assign n75282 = pi11 ? n75278 : n75281;
  assign n75283 = pi14 ? n45572 : n58990;
  assign n75284 = pi13 ? n75283 : n74986;
  assign n75285 = pi12 ? n58074 : n75284;
  assign n75286 = pi13 ? n74914 : n74853;
  assign n75287 = pi15 ? n29601 : n32185;
  assign n75288 = pi14 ? n75287 : n32185;
  assign n75289 = pi15 ? n32185 : n43787;
  assign n75290 = pi14 ? n75289 : n43787;
  assign n75291 = pi13 ? n75288 : n75290;
  assign n75292 = pi12 ? n75286 : n75291;
  assign n75293 = pi11 ? n75285 : n75292;
  assign n75294 = pi10 ? n75282 : n75293;
  assign n75295 = pi09 ? n75271 : n75294;
  assign n75296 = pi08 ? n75264 : n75295;
  assign n75297 = pi16 ? n1843 : ~n2654;
  assign n75298 = pi15 ? n32 : n75297;
  assign n75299 = pi16 ? n1479 : ~n2654;
  assign n75300 = pi15 ? n59131 : n75299;
  assign n75301 = pi14 ? n75298 : n75300;
  assign n75302 = pi13 ? n32 : n75301;
  assign n75303 = pi12 ? n32 : n75302;
  assign n75304 = pi11 ? n32 : n75303;
  assign n75305 = pi10 ? n32 : n75304;
  assign n75306 = pi16 ? n1705 : ~n2654;
  assign n75307 = pi16 ? n1972 : ~n2654;
  assign n75308 = pi15 ? n75306 : n75307;
  assign n75309 = pi16 ? n931 : ~n3788;
  assign n75310 = pi15 ? n47264 : n75309;
  assign n75311 = pi14 ? n75308 : n75310;
  assign n75312 = pi13 ? n75311 : n58837;
  assign n75313 = pi14 ? n58837 : n46655;
  assign n75314 = pi13 ? n58837 : n75313;
  assign n75315 = pi12 ? n75312 : n75314;
  assign n75316 = pi15 ? n46655 : n58837;
  assign n75317 = pi14 ? n75316 : n75248;
  assign n75318 = pi13 ? n75317 : n35359;
  assign n75319 = pi13 ? n35359 : n75182;
  assign n75320 = pi12 ? n75318 : n75319;
  assign n75321 = pi11 ? n75315 : n75320;
  assign n75322 = pi14 ? n58074 : n74983;
  assign n75323 = pi13 ? n75322 : n75055;
  assign n75324 = pi12 ? n46354 : n75323;
  assign n75325 = pi14 ? n57596 : n74716;
  assign n75326 = pi13 ? n75088 : n75325;
  assign n75327 = pi14 ? n74632 : n32185;
  assign n75328 = pi13 ? n75327 : n74918;
  assign n75329 = pi12 ? n75326 : n75328;
  assign n75330 = pi11 ? n75324 : n75329;
  assign n75331 = pi10 ? n75321 : n75330;
  assign n75332 = pi09 ? n75305 : n75331;
  assign n75333 = pi15 ? n32 : n59131;
  assign n75334 = pi15 ? n75299 : n75306;
  assign n75335 = pi14 ? n75333 : n75334;
  assign n75336 = pi13 ? n32 : n75335;
  assign n75337 = pi12 ? n32 : n75336;
  assign n75338 = pi11 ? n32 : n75337;
  assign n75339 = pi10 ? n32 : n75338;
  assign n75340 = pi15 ? n75307 : n47264;
  assign n75341 = pi16 ? n931 : ~n2654;
  assign n75342 = pi15 ? n75341 : n46774;
  assign n75343 = pi14 ? n75340 : n75342;
  assign n75344 = pi13 ? n75343 : n75313;
  assign n75345 = pi12 ? n75344 : n46655;
  assign n75346 = pi14 ? n35359 : n75248;
  assign n75347 = pi13 ? n75346 : n75181;
  assign n75348 = pi12 ? n75318 : n75347;
  assign n75349 = pi11 ? n75345 : n75348;
  assign n75350 = pi15 ? n46354 : n45572;
  assign n75351 = pi14 ? n46354 : n75350;
  assign n75352 = pi13 ? n75351 : n75283;
  assign n75353 = pi12 ? n58400 : n75352;
  assign n75354 = pi13 ? n75088 : n74914;
  assign n75355 = pi14 ? n74632 : n44537;
  assign n75356 = pi13 ? n75355 : n74918;
  assign n75357 = pi12 ? n75354 : n75356;
  assign n75358 = pi11 ? n75353 : n75357;
  assign n75359 = pi10 ? n75349 : n75358;
  assign n75360 = pi09 ? n75339 : n75359;
  assign n75361 = pi08 ? n75332 : n75360;
  assign n75362 = pi07 ? n75296 : n75361;
  assign n75363 = pi15 ? n32 : n59230;
  assign n75364 = pi16 ? n1479 : ~n2426;
  assign n75365 = pi16 ? n1705 : ~n2426;
  assign n75366 = pi15 ? n75364 : n75365;
  assign n75367 = pi14 ? n75363 : n75366;
  assign n75368 = pi13 ? n32 : n75367;
  assign n75369 = pi12 ? n32 : n75368;
  assign n75370 = pi11 ? n32 : n75369;
  assign n75371 = pi10 ? n32 : n75370;
  assign n75372 = pi16 ? n1972 : ~n2426;
  assign n75373 = pi15 ? n75372 : n47341;
  assign n75374 = pi16 ? n931 : ~n2426;
  assign n75375 = pi15 ? n75374 : n46441;
  assign n75376 = pi14 ? n75373 : n75375;
  assign n75377 = pi13 ? n75376 : n46655;
  assign n75378 = pi15 ? n46655 : n60033;
  assign n75379 = pi14 ? n75378 : n60033;
  assign n75380 = pi13 ? n46655 : n75379;
  assign n75381 = pi12 ? n75377 : n75380;
  assign n75382 = pi14 ? n60034 : n58837;
  assign n75383 = pi13 ? n75382 : n58837;
  assign n75384 = pi13 ? n58837 : n75249;
  assign n75385 = pi12 ? n75383 : n75384;
  assign n75386 = pi11 ? n75381 : n75385;
  assign n75387 = pi14 ? n46354 : n75081;
  assign n75388 = pi13 ? n75387 : n45572;
  assign n75389 = pi12 ? n58400 : n75388;
  assign n75390 = pi14 ? n45572 : n57695;
  assign n75391 = pi14 ? n57695 : n32806;
  assign n75392 = pi13 ? n75390 : n75391;
  assign n75393 = pi15 ? n32806 : n44537;
  assign n75394 = pi14 ? n75393 : n44537;
  assign n75395 = pi13 ? n75394 : n74990;
  assign n75396 = pi12 ? n75392 : n75395;
  assign n75397 = pi11 ? n75389 : n75396;
  assign n75398 = pi10 ? n75386 : n75397;
  assign n75399 = pi09 ? n75371 : n75398;
  assign n75400 = pi14 ? n46655 : n60033;
  assign n75401 = pi13 ? n75376 : n75400;
  assign n75402 = pi12 ? n75401 : n60033;
  assign n75403 = pi14 ? n60034 : n46655;
  assign n75404 = pi13 ? n75403 : n46655;
  assign n75405 = pi13 ? n46655 : n75317;
  assign n75406 = pi12 ? n75404 : n75405;
  assign n75407 = pi11 ? n75402 : n75406;
  assign n75408 = pi14 ? n58400 : n75081;
  assign n75409 = pi14 ? n58074 : n45572;
  assign n75410 = pi13 ? n75408 : n75409;
  assign n75411 = pi12 ? n35359 : n75410;
  assign n75412 = pi13 ? n75390 : n75088;
  assign n75413 = pi14 ? n74716 : n29601;
  assign n75414 = pi13 ? n75413 : n74990;
  assign n75415 = pi12 ? n75412 : n75414;
  assign n75416 = pi11 ? n75411 : n75415;
  assign n75417 = pi10 ? n75407 : n75416;
  assign n75418 = pi09 ? n75371 : n75417;
  assign n75419 = pi08 ? n75399 : n75418;
  assign n75420 = pi16 ? n1479 : ~n2120;
  assign n75421 = pi15 ? n32 : n75420;
  assign n75422 = pi16 ? n1705 : ~n2120;
  assign n75423 = pi15 ? n75420 : n75422;
  assign n75424 = pi14 ? n75421 : n75423;
  assign n75425 = pi13 ? n32 : n75424;
  assign n75426 = pi12 ? n32 : n75425;
  assign n75427 = pi11 ? n32 : n75426;
  assign n75428 = pi10 ? n32 : n75427;
  assign n75429 = pi15 ? n37160 : n47471;
  assign n75430 = pi16 ? n931 : ~n2120;
  assign n75431 = pi15 ? n75430 : n46991;
  assign n75432 = pi14 ? n75429 : n75431;
  assign n75433 = pi13 ? n75432 : n60033;
  assign n75434 = pi15 ? n60033 : n36601;
  assign n75435 = pi14 ? n75434 : n36601;
  assign n75436 = pi13 ? n60033 : n75435;
  assign n75437 = pi12 ? n75433 : n75436;
  assign n75438 = pi15 ? n36601 : n60033;
  assign n75439 = pi14 ? n75438 : n60033;
  assign n75440 = pi13 ? n75439 : n60033;
  assign n75441 = pi15 ? n60033 : n58837;
  assign n75442 = pi14 ? n75441 : n58837;
  assign n75443 = pi13 ? n60033 : n75442;
  assign n75444 = pi12 ? n75440 : n75443;
  assign n75445 = pi11 ? n75437 : n75444;
  assign n75446 = pi14 ? n75248 : n35359;
  assign n75447 = pi13 ? n75446 : n35359;
  assign n75448 = pi15 ? n58400 : n58074;
  assign n75449 = pi14 ? n58400 : n75448;
  assign n75450 = pi13 ? n75449 : n58074;
  assign n75451 = pi12 ? n75447 : n75450;
  assign n75452 = pi14 ? n58990 : n57596;
  assign n75453 = pi13 ? n75409 : n75452;
  assign n75454 = pi13 ? n75413 : n75355;
  assign n75455 = pi12 ? n75453 : n75454;
  assign n75456 = pi11 ? n75451 : n75455;
  assign n75457 = pi10 ? n75445 : n75456;
  assign n75458 = pi09 ? n75428 : n75457;
  assign n75459 = pi14 ? n60033 : n36601;
  assign n75460 = pi13 ? n75432 : n75459;
  assign n75461 = pi15 ? n36601 : n59560;
  assign n75462 = pi15 ? n59560 : n36601;
  assign n75463 = pi14 ? n75461 : n75462;
  assign n75464 = pi13 ? n36601 : n75463;
  assign n75465 = pi12 ? n75460 : n75464;
  assign n75466 = pi13 ? n60033 : n75382;
  assign n75467 = pi12 ? n75440 : n75466;
  assign n75468 = pi11 ? n75465 : n75467;
  assign n75469 = pi14 ? n35359 : n75117;
  assign n75470 = pi14 ? n46354 : n58074;
  assign n75471 = pi13 ? n75469 : n75470;
  assign n75472 = pi12 ? n58837 : n75471;
  assign n75473 = pi14 ? n45572 : n74850;
  assign n75474 = pi13 ? n75409 : n75473;
  assign n75475 = pi13 ? n74853 : n75355;
  assign n75476 = pi12 ? n75474 : n75475;
  assign n75477 = pi11 ? n75472 : n75476;
  assign n75478 = pi10 ? n75468 : n75477;
  assign n75479 = pi09 ? n75428 : n75478;
  assign n75480 = pi08 ? n75458 : n75479;
  assign n75481 = pi07 ? n75419 : n75480;
  assign n75482 = pi06 ? n75362 : n75481;
  assign n75483 = pi16 ? n1479 : ~n2415;
  assign n75484 = pi15 ? n32 : n75483;
  assign n75485 = pi16 ? n1705 : ~n2415;
  assign n75486 = pi14 ? n75484 : n75485;
  assign n75487 = pi13 ? n32 : n75486;
  assign n75488 = pi12 ? n32 : n75487;
  assign n75489 = pi11 ? n32 : n75488;
  assign n75490 = pi10 ? n32 : n75489;
  assign n75491 = pi16 ? n1972 : ~n2415;
  assign n75492 = pi15 ? n75491 : n61887;
  assign n75493 = pi16 ? n931 : ~n2415;
  assign n75494 = pi15 ? n75493 : n47256;
  assign n75495 = pi14 ? n75492 : n75494;
  assign n75496 = pi14 ? n36601 : n59560;
  assign n75497 = pi13 ? n75495 : n75496;
  assign n75498 = pi15 ? n59560 : n34044;
  assign n75499 = pi14 ? n75498 : n59560;
  assign n75500 = pi13 ? n59560 : n75499;
  assign n75501 = pi12 ? n75497 : n75500;
  assign n75502 = pi14 ? n75462 : n36601;
  assign n75503 = pi13 ? n75502 : n36601;
  assign n75504 = pi13 ? n36601 : n75403;
  assign n75505 = pi12 ? n75503 : n75504;
  assign n75506 = pi11 ? n75501 : n75505;
  assign n75507 = pi15 ? n35359 : n46354;
  assign n75508 = pi14 ? n35359 : n75507;
  assign n75509 = pi13 ? n75508 : n46354;
  assign n75510 = pi12 ? n58837 : n75509;
  assign n75511 = pi14 ? n74983 : n57695;
  assign n75512 = pi13 ? n75470 : n75511;
  assign n75513 = pi13 ? n75214 : n75413;
  assign n75514 = pi12 ? n75512 : n75513;
  assign n75515 = pi11 ? n75510 : n75514;
  assign n75516 = pi10 ? n75506 : n75515;
  assign n75517 = pi09 ? n75490 : n75516;
  assign n75518 = pi16 ? n1705 : ~n2409;
  assign n75519 = pi15 ? n75518 : n75485;
  assign n75520 = pi14 ? n75484 : n75519;
  assign n75521 = pi13 ? n32 : n75520;
  assign n75522 = pi12 ? n32 : n75521;
  assign n75523 = pi11 ? n32 : n75522;
  assign n75524 = pi10 ? n32 : n75523;
  assign n75525 = pi16 ? n1972 : ~n2409;
  assign n75526 = pi15 ? n75525 : n61887;
  assign n75527 = pi14 ? n75526 : n75494;
  assign n75528 = pi14 ? n75498 : n34044;
  assign n75529 = pi13 ? n75527 : n75528;
  assign n75530 = pi14 ? n34044 : n61073;
  assign n75531 = pi13 ? n34044 : n75530;
  assign n75532 = pi12 ? n75529 : n75531;
  assign n75533 = pi14 ? n59560 : n75462;
  assign n75534 = pi13 ? n75533 : n36601;
  assign n75535 = pi14 ? n47101 : n46655;
  assign n75536 = pi13 ? n36601 : n75535;
  assign n75537 = pi12 ? n75534 : n75536;
  assign n75538 = pi11 ? n75532 : n75537;
  assign n75539 = pi14 ? n75248 : n58400;
  assign n75540 = pi13 ? n75539 : n46354;
  assign n75541 = pi12 ? n46655 : n75540;
  assign n75542 = pi13 ? n75214 : n74717;
  assign n75543 = pi12 ? n75512 : n75542;
  assign n75544 = pi11 ? n75541 : n75543;
  assign n75545 = pi10 ? n75538 : n75544;
  assign n75546 = pi09 ? n75524 : n75545;
  assign n75547 = pi08 ? n75517 : n75546;
  assign n75548 = pi16 ? n1479 : ~n2409;
  assign n75549 = pi15 ? n32 : n75548;
  assign n75550 = pi16 ? n1705 : ~n2293;
  assign n75551 = pi15 ? n75550 : n75525;
  assign n75552 = pi14 ? n75549 : n75551;
  assign n75553 = pi13 ? n32 : n75552;
  assign n75554 = pi12 ? n32 : n75553;
  assign n75555 = pi11 ? n32 : n75554;
  assign n75556 = pi10 ? n32 : n75555;
  assign n75557 = pi16 ? n1972 : ~n2293;
  assign n75558 = pi15 ? n75557 : n59715;
  assign n75559 = pi16 ? n931 : ~n2409;
  assign n75560 = pi15 ? n75559 : n60402;
  assign n75561 = pi14 ? n75558 : n75560;
  assign n75562 = pi13 ? n75561 : n34044;
  assign n75563 = pi15 ? n34044 : n59901;
  assign n75564 = pi15 ? n59901 : n34044;
  assign n75565 = pi14 ? n75563 : n75564;
  assign n75566 = pi13 ? n34044 : n75565;
  assign n75567 = pi12 ? n75562 : n75566;
  assign n75568 = pi13 ? n59560 : n75439;
  assign n75569 = pi12 ? n59560 : n75568;
  assign n75570 = pi11 ? n75567 : n75569;
  assign n75571 = pi14 ? n58837 : n75181;
  assign n75572 = pi13 ? n75571 : n58400;
  assign n75573 = pi12 ? n46655 : n75572;
  assign n75574 = pi14 ? n58400 : n46354;
  assign n75575 = pi14 ? n58074 : n58990;
  assign n75576 = pi13 ? n75574 : n75575;
  assign n75577 = pi13 ? n57596 : n74785;
  assign n75578 = pi12 ? n75576 : n75577;
  assign n75579 = pi11 ? n75573 : n75578;
  assign n75580 = pi10 ? n75570 : n75579;
  assign n75581 = pi09 ? n75556 : n75580;
  assign n75582 = pi16 ? n1479 : ~n2293;
  assign n75583 = pi15 ? n32 : n75582;
  assign n75584 = pi15 ? n75550 : n75557;
  assign n75585 = pi14 ? n75583 : n75584;
  assign n75586 = pi13 ? n32 : n75585;
  assign n75587 = pi12 ? n32 : n75586;
  assign n75588 = pi11 ? n32 : n75587;
  assign n75589 = pi10 ? n32 : n75588;
  assign n75590 = pi15 ? n75559 : n34146;
  assign n75591 = pi14 ? n75558 : n75590;
  assign n75592 = pi14 ? n75563 : n59901;
  assign n75593 = pi13 ? n75591 : n75592;
  assign n75594 = pi14 ? n59901 : n75564;
  assign n75595 = pi13 ? n59901 : n75594;
  assign n75596 = pi12 ? n75593 : n75595;
  assign n75597 = pi13 ? n75530 : n59560;
  assign n75598 = pi15 ? n59560 : n60033;
  assign n75599 = pi14 ? n75598 : n60033;
  assign n75600 = pi13 ? n59560 : n75599;
  assign n75601 = pi12 ? n75597 : n75600;
  assign n75602 = pi11 ? n75596 : n75601;
  assign n75603 = pi14 ? n75316 : n35359;
  assign n75604 = pi13 ? n75603 : n58400;
  assign n75605 = pi12 ? n60033 : n75604;
  assign n75606 = pi14 ? n75081 : n58990;
  assign n75607 = pi13 ? n75574 : n75606;
  assign n75608 = pi13 ? n74986 : n74785;
  assign n75609 = pi12 ? n75607 : n75608;
  assign n75610 = pi11 ? n75605 : n75609;
  assign n75611 = pi10 ? n75602 : n75610;
  assign n75612 = pi09 ? n75589 : n75611;
  assign n75613 = pi08 ? n75581 : n75612;
  assign n75614 = pi07 ? n75547 : n75613;
  assign n75615 = pi16 ? n1705 : ~n3769;
  assign n75616 = pi15 ? n32 : n75615;
  assign n75617 = pi16 ? n1972 : ~n3769;
  assign n75618 = pi15 ? n75615 : n75617;
  assign n75619 = pi14 ? n75616 : n75618;
  assign n75620 = pi13 ? n32 : n75619;
  assign n75621 = pi12 ? n32 : n75620;
  assign n75622 = pi11 ? n32 : n75621;
  assign n75623 = pi10 ? n32 : n75622;
  assign n75624 = pi15 ? n48747 : n59799;
  assign n75625 = pi16 ? n931 : ~n2293;
  assign n75626 = pi15 ? n75625 : n60814;
  assign n75627 = pi14 ? n75624 : n75626;
  assign n75628 = pi13 ? n75627 : n59901;
  assign n75629 = pi15 ? n59901 : n60190;
  assign n75630 = pi14 ? n75629 : n61070;
  assign n75631 = pi13 ? n59901 : n75630;
  assign n75632 = pi12 ? n75628 : n75631;
  assign n75633 = pi14 ? n75462 : n75438;
  assign n75634 = pi13 ? n34044 : n75633;
  assign n75635 = pi12 ? n34044 : n75634;
  assign n75636 = pi11 ? n75632 : n75635;
  assign n75637 = pi14 ? n46655 : n75248;
  assign n75638 = pi13 ? n75637 : n35359;
  assign n75639 = pi12 ? n60033 : n75638;
  assign n75640 = pi13 ? n75469 : n75053;
  assign n75641 = pi13 ? n57695 : n74851;
  assign n75642 = pi12 ? n75640 : n75641;
  assign n75643 = pi11 ? n75639 : n75642;
  assign n75644 = pi10 ? n75636 : n75643;
  assign n75645 = pi09 ? n75623 : n75644;
  assign n75646 = pi14 ? n48747 : n75626;
  assign n75647 = pi14 ? n75629 : n60190;
  assign n75648 = pi13 ? n75646 : n75647;
  assign n75649 = pi14 ? n60190 : n61070;
  assign n75650 = pi13 ? n60190 : n75649;
  assign n75651 = pi12 ? n75648 : n75650;
  assign n75652 = pi13 ? n75594 : n34044;
  assign n75653 = pi15 ? n34044 : n36601;
  assign n75654 = pi14 ? n75653 : n36601;
  assign n75655 = pi13 ? n34044 : n75654;
  assign n75656 = pi12 ? n75652 : n75655;
  assign n75657 = pi11 ? n75651 : n75656;
  assign n75658 = pi13 ? n75382 : n35359;
  assign n75659 = pi12 ? n36601 : n75658;
  assign n75660 = pi14 ? n35359 : n58400;
  assign n75661 = pi14 ? n75117 : n74983;
  assign n75662 = pi13 ? n75660 : n75661;
  assign n75663 = pi13 ? n75055 : n74851;
  assign n75664 = pi12 ? n75662 : n75663;
  assign n75665 = pi11 ? n75659 : n75664;
  assign n75666 = pi10 ? n75657 : n75665;
  assign n75667 = pi09 ? n75623 : n75666;
  assign n75668 = pi08 ? n75645 : n75667;
  assign n75669 = pi16 ? n1705 : ~n2756;
  assign n75670 = pi15 ? n32 : n75669;
  assign n75671 = pi16 ? n1972 : ~n2756;
  assign n75672 = pi14 ? n75670 : n75671;
  assign n75673 = pi13 ? n32 : n75672;
  assign n75674 = pi12 ? n32 : n75673;
  assign n75675 = pi11 ? n32 : n75674;
  assign n75676 = pi10 ? n32 : n75675;
  assign n75677 = pi16 ? n931 : ~n2756;
  assign n75678 = pi15 ? n45903 : n75677;
  assign n75679 = pi16 ? n931 : ~n3769;
  assign n75680 = pi15 ? n75679 : n47710;
  assign n75681 = pi14 ? n75678 : n75680;
  assign n75682 = pi13 ? n75681 : n60190;
  assign n75683 = pi15 ? n60190 : n61238;
  assign n75684 = pi14 ? n75683 : n61239;
  assign n75685 = pi13 ? n60190 : n75684;
  assign n75686 = pi12 ? n75682 : n75685;
  assign n75687 = pi14 ? n61073 : n75462;
  assign n75688 = pi13 ? n59901 : n75687;
  assign n75689 = pi12 ? n59901 : n75688;
  assign n75690 = pi11 ? n75686 : n75689;
  assign n75691 = pi14 ? n60033 : n58837;
  assign n75692 = pi13 ? n75691 : n58837;
  assign n75693 = pi12 ? n36601 : n75692;
  assign n75694 = pi14 ? n58837 : n58400;
  assign n75695 = pi14 ? n75117 : n75350;
  assign n75696 = pi13 ? n75694 : n75695;
  assign n75697 = pi15 ? n57695 : n32806;
  assign n75698 = pi14 ? n58990 : n75697;
  assign n75699 = pi13 ? n45572 : n75698;
  assign n75700 = pi12 ? n75696 : n75699;
  assign n75701 = pi11 ? n75693 : n75700;
  assign n75702 = pi10 ? n75690 : n75701;
  assign n75703 = pi09 ? n75676 : n75702;
  assign n75704 = pi15 ? n32 : n75671;
  assign n75705 = pi14 ? n75704 : n75671;
  assign n75706 = pi13 ? n32 : n75705;
  assign n75707 = pi12 ? n32 : n75706;
  assign n75708 = pi11 ? n32 : n75707;
  assign n75709 = pi10 ? n32 : n75708;
  assign n75710 = pi14 ? n75678 : n47710;
  assign n75711 = pi14 ? n75683 : n61238;
  assign n75712 = pi13 ? n75710 : n75711;
  assign n75713 = pi13 ? n61238 : n61240;
  assign n75714 = pi12 ? n75712 : n75713;
  assign n75715 = pi14 ? n60190 : n59901;
  assign n75716 = pi13 ? n75715 : n59901;
  assign n75717 = pi15 ? n59901 : n59560;
  assign n75718 = pi14 ? n75717 : n59560;
  assign n75719 = pi13 ? n59901 : n75718;
  assign n75720 = pi12 ? n75716 : n75719;
  assign n75721 = pi11 ? n75714 : n75720;
  assign n75722 = pi14 ? n60033 : n46655;
  assign n75723 = pi13 ? n75722 : n58837;
  assign n75724 = pi12 ? n59560 : n75723;
  assign n75725 = pi14 ? n58837 : n35359;
  assign n75726 = pi14 ? n75507 : n75081;
  assign n75727 = pi13 ? n75725 : n75726;
  assign n75728 = pi13 ? n75148 : n74912;
  assign n75729 = pi12 ? n75727 : n75728;
  assign n75730 = pi11 ? n75724 : n75729;
  assign n75731 = pi10 ? n75721 : n75730;
  assign n75732 = pi09 ? n75709 : n75731;
  assign n75733 = pi08 ? n75703 : n75732;
  assign n75734 = pi07 ? n75668 : n75733;
  assign n75735 = pi06 ? n75614 : n75734;
  assign n75736 = pi05 ? n75482 : n75735;
  assign n75737 = pi04 ? n75227 : n75736;
  assign n75738 = pi03 ? n74695 : n75737;
  assign n75739 = pi16 ? n1972 : ~n2518;
  assign n75740 = pi15 ? n32 : n75739;
  assign n75741 = pi15 ? n75739 : n46036;
  assign n75742 = pi14 ? n75740 : n75741;
  assign n75743 = pi13 ? n32 : n75742;
  assign n75744 = pi12 ? n32 : n75743;
  assign n75745 = pi11 ? n32 : n75744;
  assign n75746 = pi10 ? n32 : n75745;
  assign n75747 = pi16 ? n931 : ~n2518;
  assign n75748 = pi15 ? n46036 : n75747;
  assign n75749 = pi15 ? n60189 : n61238;
  assign n75750 = pi14 ? n75748 : n75749;
  assign n75751 = pi13 ? n75750 : n61238;
  assign n75752 = pi14 ? n61506 : n61238;
  assign n75753 = pi13 ? n61238 : n75752;
  assign n75754 = pi12 ? n75751 : n75753;
  assign n75755 = pi14 ? n75564 : n61073;
  assign n75756 = pi13 ? n60190 : n75755;
  assign n75757 = pi12 ? n60190 : n75756;
  assign n75758 = pi11 ? n75754 : n75757;
  assign n75759 = pi14 ? n36601 : n46655;
  assign n75760 = pi13 ? n75759 : n46655;
  assign n75761 = pi12 ? n59560 : n75760;
  assign n75762 = pi14 ? n46655 : n35359;
  assign n75763 = pi13 ? n75762 : n75726;
  assign n75764 = pi14 ? n74983 : n74850;
  assign n75765 = pi13 ? n58074 : n75764;
  assign n75766 = pi12 ? n75763 : n75765;
  assign n75767 = pi11 ? n75761 : n75766;
  assign n75768 = pi10 ? n75758 : n75767;
  assign n75769 = pi09 ? n75746 : n75768;
  assign n75770 = pi14 ? n75740 : n46036;
  assign n75771 = pi13 ? n32 : n75770;
  assign n75772 = pi12 ? n32 : n75771;
  assign n75773 = pi11 ? n32 : n75772;
  assign n75774 = pi10 ? n32 : n75773;
  assign n75775 = pi15 ? n61238 : n61506;
  assign n75776 = pi14 ? n75775 : n61506;
  assign n75777 = pi13 ? n75750 : n75776;
  assign n75778 = pi15 ? n61506 : n61238;
  assign n75779 = pi14 ? n61506 : n75778;
  assign n75780 = pi13 ? n61506 : n75779;
  assign n75781 = pi12 ? n75777 : n75780;
  assign n75782 = pi14 ? n61238 : n60190;
  assign n75783 = pi13 ? n75782 : n60190;
  assign n75784 = pi15 ? n60190 : n34044;
  assign n75785 = pi14 ? n75784 : n34044;
  assign n75786 = pi13 ? n60190 : n75785;
  assign n75787 = pi12 ? n75783 : n75786;
  assign n75788 = pi11 ? n75781 : n75787;
  assign n75789 = pi14 ? n36601 : n60033;
  assign n75790 = pi13 ? n75789 : n46655;
  assign n75791 = pi12 ? n34044 : n75790;
  assign n75792 = pi14 ? n46655 : n58837;
  assign n75793 = pi15 ? n58837 : n58400;
  assign n75794 = pi14 ? n75793 : n75117;
  assign n75795 = pi13 ? n75792 : n75794;
  assign n75796 = pi12 ? n75795 : n75120;
  assign n75797 = pi11 ? n75791 : n75796;
  assign n75798 = pi10 ? n75788 : n75797;
  assign n75799 = pi09 ? n75774 : n75798;
  assign n75800 = pi08 ? n75769 : n75799;
  assign n75801 = pi16 ? n1972 : ~n2749;
  assign n75802 = pi15 ? n32 : n75801;
  assign n75803 = pi16 ? n1214 : ~n2749;
  assign n75804 = pi14 ? n75802 : n75803;
  assign n75805 = pi13 ? n32 : n75804;
  assign n75806 = pi12 ? n32 : n75805;
  assign n75807 = pi11 ? n32 : n75806;
  assign n75808 = pi10 ? n32 : n75807;
  assign n75809 = pi16 ? n931 : ~n2749;
  assign n75810 = pi15 ? n61329 : n61506;
  assign n75811 = pi14 ? n75809 : n75810;
  assign n75812 = pi13 ? n75811 : n61506;
  assign n75813 = pi13 ? n61506 : n61508;
  assign n75814 = pi12 ? n75812 : n75813;
  assign n75815 = pi14 ? n61070 : n75564;
  assign n75816 = pi13 ? n61240 : n75815;
  assign n75817 = pi12 ? n61238 : n75816;
  assign n75818 = pi11 ? n75814 : n75817;
  assign n75819 = pi13 ? n75789 : n60033;
  assign n75820 = pi12 ? n34044 : n75819;
  assign n75821 = pi13 ? n75382 : n75794;
  assign n75822 = pi14 ? n75350 : n58990;
  assign n75823 = pi13 ? n46354 : n75822;
  assign n75824 = pi12 ? n75821 : n75823;
  assign n75825 = pi11 ? n75820 : n75824;
  assign n75826 = pi10 ? n75818 : n75825;
  assign n75827 = pi09 ? n75808 : n75826;
  assign n75828 = pi15 ? n32 : n75803;
  assign n75829 = pi15 ? n75803 : n75809;
  assign n75830 = pi14 ? n75828 : n75829;
  assign n75831 = pi13 ? n32 : n75830;
  assign n75832 = pi12 ? n32 : n75831;
  assign n75833 = pi11 ? n32 : n75832;
  assign n75834 = pi10 ? n32 : n75833;
  assign n75835 = pi15 ? n75809 : n61629;
  assign n75836 = pi14 ? n75835 : n75810;
  assign n75837 = pi15 ? n61506 : n61505;
  assign n75838 = pi14 ? n75837 : n61505;
  assign n75839 = pi13 ? n75836 : n75838;
  assign n75840 = pi14 ? n61505 : n61507;
  assign n75841 = pi13 ? n61505 : n75840;
  assign n75842 = pi12 ? n75839 : n75841;
  assign n75843 = pi13 ? n75752 : n61238;
  assign n75844 = pi15 ? n61238 : n59901;
  assign n75845 = pi14 ? n75844 : n59901;
  assign n75846 = pi13 ? n61238 : n75845;
  assign n75847 = pi12 ? n75843 : n75846;
  assign n75848 = pi11 ? n75842 : n75847;
  assign n75849 = pi14 ? n59560 : n75438;
  assign n75850 = pi13 ? n75849 : n60033;
  assign n75851 = pi12 ? n59901 : n75850;
  assign n75852 = pi14 ? n75248 : n75117;
  assign n75853 = pi13 ? n75722 : n75852;
  assign n75854 = pi12 ? n75853 : n75184;
  assign n75855 = pi11 ? n75851 : n75854;
  assign n75856 = pi10 ? n75848 : n75855;
  assign n75857 = pi09 ? n75834 : n75856;
  assign n75858 = pi08 ? n75827 : n75857;
  assign n75859 = pi07 ? n75800 : n75858;
  assign n75860 = pi16 ? n1214 : ~n2513;
  assign n75861 = pi15 ? n32 : n75860;
  assign n75862 = pi16 ? n931 : ~n2513;
  assign n75863 = pi15 ? n75860 : n75862;
  assign n75864 = pi14 ? n75861 : n75863;
  assign n75865 = pi13 ? n32 : n75864;
  assign n75866 = pi12 ? n32 : n75865;
  assign n75867 = pi11 ? n32 : n75866;
  assign n75868 = pi10 ? n32 : n75867;
  assign n75869 = pi15 ? n75862 : n61868;
  assign n75870 = pi15 ? n61629 : n61505;
  assign n75871 = pi14 ? n75869 : n75870;
  assign n75872 = pi13 ? n75871 : n61505;
  assign n75873 = pi13 ? n61505 : n61712;
  assign n75874 = pi12 ? n75872 : n75873;
  assign n75875 = pi14 ? n61239 : n61070;
  assign n75876 = pi13 ? n61506 : n75875;
  assign n75877 = pi12 ? n61506 : n75876;
  assign n75878 = pi11 ? n75874 : n75877;
  assign n75879 = pi14 ? n59560 : n36601;
  assign n75880 = pi13 ? n75879 : n36601;
  assign n75881 = pi12 ? n59901 : n75880;
  assign n75882 = pi13 ? n75722 : n75539;
  assign n75883 = pi14 ? n75448 : n74983;
  assign n75884 = pi13 ? n58400 : n75883;
  assign n75885 = pi12 ? n75882 : n75884;
  assign n75886 = pi11 ? n75881 : n75885;
  assign n75887 = pi10 ? n75878 : n75886;
  assign n75888 = pi09 ? n75868 : n75887;
  assign n75889 = pi15 ? n61505 : n61710;
  assign n75890 = pi14 ? n75889 : n61710;
  assign n75891 = pi13 ? n75871 : n75890;
  assign n75892 = pi14 ? n61710 : n61505;
  assign n75893 = pi13 ? n61710 : n75892;
  assign n75894 = pi12 ? n75891 : n75893;
  assign n75895 = pi14 ? n61505 : n61506;
  assign n75896 = pi13 ? n75895 : n61506;
  assign n75897 = pi14 ? n61239 : n60190;
  assign n75898 = pi13 ? n75779 : n75897;
  assign n75899 = pi12 ? n75896 : n75898;
  assign n75900 = pi11 ? n75894 : n75899;
  assign n75901 = pi14 ? n61073 : n36601;
  assign n75902 = pi13 ? n75901 : n36601;
  assign n75903 = pi12 ? n75650 : n75902;
  assign n75904 = pi14 ? n75316 : n75181;
  assign n75905 = pi13 ? n75789 : n75904;
  assign n75906 = pi12 ? n75905 : n75251;
  assign n75907 = pi11 ? n75903 : n75906;
  assign n75908 = pi10 ? n75900 : n75907;
  assign n75909 = pi09 ? n75868 : n75908;
  assign n75910 = pi08 ? n75888 : n75909;
  assign n75911 = pi15 ? n32 : n62102;
  assign n75912 = pi16 ? n931 : ~n2629;
  assign n75913 = pi15 ? n62102 : n75912;
  assign n75914 = pi14 ? n75911 : n75913;
  assign n75915 = pi13 ? n32 : n75914;
  assign n75916 = pi12 ? n32 : n75915;
  assign n75917 = pi11 ? n32 : n75916;
  assign n75918 = pi10 ? n32 : n75917;
  assign n75919 = pi15 ? n75912 : n62213;
  assign n75920 = pi15 ? n61868 : n61710;
  assign n75921 = pi14 ? n75919 : n75920;
  assign n75922 = pi13 ? n75921 : n61710;
  assign n75923 = pi12 ? n75922 : n61710;
  assign n75924 = pi14 ? n75778 : n60190;
  assign n75925 = pi13 ? n75840 : n75924;
  assign n75926 = pi12 ? n61505 : n75925;
  assign n75927 = pi11 ? n75923 : n75926;
  assign n75928 = pi14 ? n61073 : n59560;
  assign n75929 = pi13 ? n75928 : n59560;
  assign n75930 = pi12 ? n75650 : n75929;
  assign n75931 = pi14 ? n36601 : n60034;
  assign n75932 = pi13 ? n75931 : n75446;
  assign n75933 = pi14 ? n35359 : n75181;
  assign n75934 = pi13 ? n75933 : n75661;
  assign n75935 = pi12 ? n75932 : n75934;
  assign n75936 = pi11 ? n75930 : n75935;
  assign n75937 = pi10 ? n75927 : n75936;
  assign n75938 = pi09 ? n75918 : n75937;
  assign n75939 = pi13 ? n75921 : n62214;
  assign n75940 = pi15 ? n62214 : n61710;
  assign n75941 = pi14 ? n62214 : n75940;
  assign n75942 = pi13 ? n62214 : n75941;
  assign n75943 = pi12 ? n75939 : n75942;
  assign n75944 = pi13 ? n75892 : n61505;
  assign n75945 = pi14 ? n75778 : n61238;
  assign n75946 = pi13 ? n75840 : n75945;
  assign n75947 = pi12 ? n75944 : n75946;
  assign n75948 = pi11 ? n75943 : n75947;
  assign n75949 = pi14 ? n75564 : n59560;
  assign n75950 = pi13 ? n75949 : n59560;
  assign n75951 = pi12 ? n75713 : n75950;
  assign n75952 = pi13 ? n75849 : n75603;
  assign n75953 = pi13 ? n35359 : n75726;
  assign n75954 = pi12 ? n75952 : n75953;
  assign n75955 = pi11 ? n75951 : n75954;
  assign n75956 = pi10 ? n75948 : n75955;
  assign n75957 = pi09 ? n75918 : n75956;
  assign n75958 = pi08 ? n75938 : n75957;
  assign n75959 = pi07 ? n75910 : n75958;
  assign n75960 = pi06 ? n75859 : n75959;
  assign n75961 = pi15 ? n32 : n62210;
  assign n75962 = pi16 ? n931 : ~n3946;
  assign n75963 = pi15 ? n62210 : n75962;
  assign n75964 = pi14 ? n75961 : n75963;
  assign n75965 = pi13 ? n32 : n75964;
  assign n75966 = pi12 ? n32 : n75965;
  assign n75967 = pi11 ? n32 : n75966;
  assign n75968 = pi10 ? n32 : n75967;
  assign n75969 = pi15 ? n75962 : n62813;
  assign n75970 = pi14 ? n75969 : n62215;
  assign n75971 = pi13 ? n75970 : n62214;
  assign n75972 = pi12 ? n75971 : n75942;
  assign n75973 = pi14 ? n61507 : n61238;
  assign n75974 = pi13 ? n61985 : n75973;
  assign n75975 = pi12 ? n61710 : n75974;
  assign n75976 = pi11 ? n75972 : n75975;
  assign n75977 = pi14 ? n75564 : n34044;
  assign n75978 = pi13 ? n75977 : n75530;
  assign n75979 = pi12 ? n75713 : n75978;
  assign n75980 = pi14 ? n75316 : n58837;
  assign n75981 = pi13 ? n75849 : n75980;
  assign n75982 = pi12 ? n75981 : n75727;
  assign n75983 = pi11 ? n75979 : n75982;
  assign n75984 = pi10 ? n75976 : n75983;
  assign n75985 = pi09 ? n75968 : n75984;
  assign n75986 = pi15 ? n62813 : n62214;
  assign n75987 = pi14 ? n75969 : n75986;
  assign n75988 = pi16 ? n1233 : ~n3946;
  assign n75989 = pi13 ? n75987 : n75988;
  assign n75990 = pi15 ? n75988 : n62214;
  assign n75991 = pi14 ? n75988 : n75990;
  assign n75992 = pi13 ? n75988 : n75991;
  assign n75993 = pi12 ? n75989 : n75992;
  assign n75994 = pi14 ? n62214 : n61710;
  assign n75995 = pi13 ? n75994 : n61710;
  assign n75996 = pi13 ? n61985 : n61508;
  assign n75997 = pi12 ? n75995 : n75996;
  assign n75998 = pi11 ? n75993 : n75997;
  assign n75999 = pi14 ? n61070 : n34044;
  assign n76000 = pi13 ? n75999 : n34044;
  assign n76001 = pi12 ? n75780 : n76000;
  assign n76002 = pi13 ? n75901 : n75382;
  assign n76003 = pi14 ? n75793 : n75081;
  assign n76004 = pi13 ? n58837 : n76003;
  assign n76005 = pi12 ? n76002 : n76004;
  assign n76006 = pi11 ? n76001 : n76005;
  assign n76007 = pi10 ? n75998 : n76006;
  assign n76008 = pi09 ? n75968 : n76007;
  assign n76009 = pi08 ? n75985 : n76008;
  assign n76010 = pi15 ? n32 : n62671;
  assign n76011 = pi16 ? n931 : ~n4100;
  assign n76012 = pi15 ? n62671 : n76011;
  assign n76013 = pi14 ? n76010 : n76012;
  assign n76014 = pi13 ? n32 : n76013;
  assign n76015 = pi12 ? n32 : n76014;
  assign n76016 = pi11 ? n32 : n76015;
  assign n76017 = pi10 ? n32 : n76016;
  assign n76018 = pi16 ? n1135 : ~n4100;
  assign n76019 = pi15 ? n76011 : n76018;
  assign n76020 = pi15 ? n76018 : n75988;
  assign n76021 = pi14 ? n76019 : n76020;
  assign n76022 = pi13 ? n76021 : n75988;
  assign n76023 = pi12 ? n76022 : n75992;
  assign n76024 = pi14 ? n61711 : n61506;
  assign n76025 = pi13 ? n75941 : n76024;
  assign n76026 = pi12 ? n62214 : n76025;
  assign n76027 = pi11 ? n76023 : n76026;
  assign n76028 = pi14 ? n61070 : n59901;
  assign n76029 = pi14 ? n59901 : n34044;
  assign n76030 = pi13 ? n76028 : n76029;
  assign n76031 = pi12 ? n75780 : n76030;
  assign n76032 = pi13 ? n75901 : n75403;
  assign n76033 = pi13 ? n75792 : n76003;
  assign n76034 = pi12 ? n76032 : n76033;
  assign n76035 = pi11 ? n76031 : n76034;
  assign n76036 = pi10 ? n76027 : n76035;
  assign n76037 = pi09 ? n76017 : n76036;
  assign n76038 = pi16 ? n1233 : ~n4100;
  assign n76039 = pi15 ? n76038 : n75988;
  assign n76040 = pi14 ? n76039 : n76038;
  assign n76041 = pi13 ? n76021 : n76040;
  assign n76042 = pi14 ? n76038 : n76039;
  assign n76043 = pi13 ? n76038 : n76042;
  assign n76044 = pi12 ? n76041 : n76043;
  assign n76045 = pi14 ? n75988 : n62214;
  assign n76046 = pi13 ? n76045 : n62214;
  assign n76047 = pi13 ? n75941 : n61712;
  assign n76048 = pi12 ? n76046 : n76047;
  assign n76049 = pi11 ? n76044 : n76048;
  assign n76050 = pi13 ? n61505 : n61508;
  assign n76051 = pi14 ? n61239 : n59901;
  assign n76052 = pi13 ? n76051 : n59901;
  assign n76053 = pi12 ? n76050 : n76052;
  assign n76054 = pi14 ? n75564 : n75462;
  assign n76055 = pi14 ? n75438 : n46655;
  assign n76056 = pi13 ? n76054 : n76055;
  assign n76057 = pi13 ? n46655 : n75852;
  assign n76058 = pi12 ? n76056 : n76057;
  assign n76059 = pi11 ? n76053 : n76058;
  assign n76060 = pi10 ? n76049 : n76059;
  assign n76061 = pi09 ? n76017 : n76060;
  assign n76062 = pi08 ? n76037 : n76061;
  assign n76063 = pi07 ? n76009 : n76062;
  assign n76064 = pi16 ? n1214 : ~n2860;
  assign n76065 = pi15 ? n32 : n76064;
  assign n76066 = pi16 ? n931 : ~n2860;
  assign n76067 = pi15 ? n76064 : n76066;
  assign n76068 = pi14 ? n76065 : n76067;
  assign n76069 = pi13 ? n32 : n76068;
  assign n76070 = pi12 ? n32 : n76069;
  assign n76071 = pi11 ? n32 : n76070;
  assign n76072 = pi10 ? n32 : n76071;
  assign n76073 = pi15 ? n76066 : n62922;
  assign n76074 = pi15 ? n62922 : n76038;
  assign n76075 = pi14 ? n76073 : n76074;
  assign n76076 = pi13 ? n76075 : n76038;
  assign n76077 = pi12 ? n76076 : n76043;
  assign n76078 = pi14 ? n75940 : n61505;
  assign n76079 = pi13 ? n75991 : n76078;
  assign n76080 = pi12 ? n75988 : n76079;
  assign n76081 = pi11 ? n76077 : n76080;
  assign n76082 = pi13 ? n75897 : n75715;
  assign n76083 = pi12 ? n76050 : n76082;
  assign n76084 = pi13 ? n76054 : n75439;
  assign n76085 = pi13 ? n75403 : n75852;
  assign n76086 = pi12 ? n76084 : n76085;
  assign n76087 = pi11 ? n76083 : n76086;
  assign n76088 = pi10 ? n76081 : n76087;
  assign n76089 = pi09 ? n76072 : n76088;
  assign n76090 = pi16 ? n1233 : ~n2860;
  assign n76091 = pi15 ? n76090 : n76038;
  assign n76092 = pi14 ? n76091 : n76090;
  assign n76093 = pi13 ? n76075 : n76092;
  assign n76094 = pi14 ? n76090 : n76091;
  assign n76095 = pi13 ? n76090 : n76094;
  assign n76096 = pi12 ? n76093 : n76095;
  assign n76097 = pi14 ? n76038 : n75988;
  assign n76098 = pi13 ? n76097 : n75988;
  assign n76099 = pi14 ? n75940 : n61710;
  assign n76100 = pi13 ? n75991 : n76099;
  assign n76101 = pi12 ? n76098 : n76100;
  assign n76102 = pi11 ? n76096 : n76101;
  assign n76103 = pi13 ? n61710 : n61712;
  assign n76104 = pi13 ? n75924 : n60190;
  assign n76105 = pi12 ? n76103 : n76104;
  assign n76106 = pi14 ? n59901 : n61073;
  assign n76107 = pi13 ? n76106 : n75599;
  assign n76108 = pi14 ? n60033 : n60034;
  assign n76109 = pi13 ? n76108 : n75904;
  assign n76110 = pi12 ? n76107 : n76109;
  assign n76111 = pi11 ? n76105 : n76110;
  assign n76112 = pi10 ? n76102 : n76111;
  assign n76113 = pi09 ? n76072 : n76112;
  assign n76114 = pi08 ? n76089 : n76113;
  assign n76115 = pi15 ? n32 : n63127;
  assign n76116 = pi16 ? n931 : ~n2624;
  assign n76117 = pi15 ? n63127 : n76116;
  assign n76118 = pi14 ? n76115 : n76117;
  assign n76119 = pi13 ? n32 : n76118;
  assign n76120 = pi12 ? n32 : n76119;
  assign n76121 = pi11 ? n32 : n76120;
  assign n76122 = pi10 ? n32 : n76121;
  assign n76123 = pi16 ? n1135 : ~n2624;
  assign n76124 = pi15 ? n76116 : n76123;
  assign n76125 = pi15 ? n76123 : n76090;
  assign n76126 = pi14 ? n76124 : n76125;
  assign n76127 = pi13 ? n76126 : n76090;
  assign n76128 = pi12 ? n76127 : n76095;
  assign n76129 = pi14 ? n76039 : n75988;
  assign n76130 = pi14 ? n75990 : n61710;
  assign n76131 = pi13 ? n76129 : n76130;
  assign n76132 = pi12 ? n76038 : n76131;
  assign n76133 = pi11 ? n76128 : n76132;
  assign n76134 = pi14 ? n61711 : n61507;
  assign n76135 = pi13 ? n61710 : n76134;
  assign n76136 = pi13 ? n75945 : n75897;
  assign n76137 = pi12 ? n76135 : n76136;
  assign n76138 = pi13 ? n76106 : n75502;
  assign n76139 = pi12 ? n76138 : n76109;
  assign n76140 = pi11 ? n76137 : n76139;
  assign n76141 = pi10 ? n76133 : n76140;
  assign n76142 = pi09 ? n76122 : n76141;
  assign n76143 = pi16 ? n1233 : ~n2624;
  assign n76144 = pi14 ? n76090 : n76143;
  assign n76145 = pi13 ? n76126 : n76144;
  assign n76146 = pi15 ? n76143 : n76090;
  assign n76147 = pi14 ? n76143 : n76146;
  assign n76148 = pi13 ? n76143 : n76147;
  assign n76149 = pi12 ? n76145 : n76148;
  assign n76150 = pi14 ? n76090 : n76038;
  assign n76151 = pi13 ? n76150 : n76038;
  assign n76152 = pi14 ? n75990 : n62214;
  assign n76153 = pi13 ? n76129 : n76152;
  assign n76154 = pi12 ? n76151 : n76153;
  assign n76155 = pi11 ? n76149 : n76154;
  assign n76156 = pi13 ? n62214 : n61985;
  assign n76157 = pi15 ? n61505 : n61238;
  assign n76158 = pi14 ? n76157 : n61238;
  assign n76159 = pi13 ? n76158 : n61240;
  assign n76160 = pi12 ? n76156 : n76159;
  assign n76161 = pi14 ? n60190 : n75564;
  assign n76162 = pi13 ? n76161 : n75502;
  assign n76163 = pi14 ? n36601 : n75438;
  assign n76164 = pi14 ? n60034 : n75181;
  assign n76165 = pi13 ? n76163 : n76164;
  assign n76166 = pi12 ? n76162 : n76165;
  assign n76167 = pi11 ? n76160 : n76166;
  assign n76168 = pi10 ? n76155 : n76167;
  assign n76169 = pi09 ? n76122 : n76168;
  assign n76170 = pi08 ? n76142 : n76169;
  assign n76171 = pi07 ? n76114 : n76170;
  assign n76172 = pi06 ? n76063 : n76171;
  assign n76173 = pi05 ? n75960 : n76172;
  assign n76174 = pi16 ? n1214 : ~n2856;
  assign n76175 = pi15 ? n32 : n76174;
  assign n76176 = pi16 ? n931 : ~n2856;
  assign n76177 = pi15 ? n76174 : n76176;
  assign n76178 = pi14 ? n76175 : n76177;
  assign n76179 = pi13 ? n32 : n76178;
  assign n76180 = pi12 ? n32 : n76179;
  assign n76181 = pi11 ? n32 : n76180;
  assign n76182 = pi10 ? n32 : n76181;
  assign n76183 = pi16 ? n1135 : ~n2856;
  assign n76184 = pi15 ? n76176 : n76183;
  assign n76185 = pi15 ? n76183 : n76143;
  assign n76186 = pi14 ? n76184 : n76185;
  assign n76187 = pi13 ? n76186 : n76143;
  assign n76188 = pi12 ? n76187 : n76148;
  assign n76189 = pi14 ? n76091 : n76038;
  assign n76190 = pi14 ? n76039 : n62214;
  assign n76191 = pi13 ? n76189 : n76190;
  assign n76192 = pi12 ? n76090 : n76191;
  assign n76193 = pi11 ? n76188 : n76192;
  assign n76194 = pi13 ? n61508 : n61240;
  assign n76195 = pi12 ? n76156 : n76194;
  assign n76196 = pi13 ? n76161 : n75533;
  assign n76197 = pi12 ? n76196 : n76165;
  assign n76198 = pi11 ? n76195 : n76197;
  assign n76199 = pi10 ? n76193 : n76198;
  assign n76200 = pi09 ? n76182 : n76199;
  assign n76201 = pi14 ? n76175 : n76176;
  assign n76202 = pi13 ? n32 : n76201;
  assign n76203 = pi12 ? n32 : n76202;
  assign n76204 = pi11 ? n32 : n76203;
  assign n76205 = pi10 ? n32 : n76204;
  assign n76206 = pi16 ? n1233 : ~n2856;
  assign n76207 = pi14 ? n76143 : n76206;
  assign n76208 = pi13 ? n76186 : n76207;
  assign n76209 = pi15 ? n76206 : n76143;
  assign n76210 = pi14 ? n76209 : n76143;
  assign n76211 = pi13 ? n76206 : n76210;
  assign n76212 = pi12 ? n76208 : n76211;
  assign n76213 = pi14 ? n76143 : n76090;
  assign n76214 = pi13 ? n76213 : n76090;
  assign n76215 = pi13 ? n76189 : n76129;
  assign n76216 = pi12 ? n76214 : n76215;
  assign n76217 = pi11 ? n76212 : n76216;
  assign n76218 = pi13 ? n75988 : n75941;
  assign n76219 = pi15 ? n61710 : n61506;
  assign n76220 = pi14 ? n76219 : n61506;
  assign n76221 = pi13 ? n76220 : n75779;
  assign n76222 = pi12 ? n76218 : n76221;
  assign n76223 = pi14 ? n61238 : n61070;
  assign n76224 = pi13 ? n76223 : n75928;
  assign n76225 = pi14 ? n75438 : n75248;
  assign n76226 = pi13 ? n75879 : n76225;
  assign n76227 = pi12 ? n76224 : n76226;
  assign n76228 = pi11 ? n76222 : n76227;
  assign n76229 = pi10 ? n76217 : n76228;
  assign n76230 = pi09 ? n76205 : n76229;
  assign n76231 = pi08 ? n76200 : n76230;
  assign n76232 = pi16 ? n931 : ~n2617;
  assign n76233 = pi15 ? n32 : n76232;
  assign n76234 = pi14 ? n76233 : n76232;
  assign n76235 = pi13 ? n32 : n76234;
  assign n76236 = pi12 ? n32 : n76235;
  assign n76237 = pi11 ? n32 : n76236;
  assign n76238 = pi10 ? n32 : n76237;
  assign n76239 = pi16 ? n1135 : ~n2617;
  assign n76240 = pi15 ? n76239 : n76206;
  assign n76241 = pi14 ? n76239 : n76240;
  assign n76242 = pi13 ? n76241 : n76206;
  assign n76243 = pi15 ? n76143 : n76206;
  assign n76244 = pi14 ? n76209 : n76243;
  assign n76245 = pi13 ? n76206 : n76244;
  assign n76246 = pi12 ? n76242 : n76245;
  assign n76247 = pi15 ? n76090 : n75988;
  assign n76248 = pi14 ? n76247 : n75988;
  assign n76249 = pi13 ? n76090 : n76248;
  assign n76250 = pi12 ? n76143 : n76249;
  assign n76251 = pi11 ? n76246 : n76250;
  assign n76252 = pi13 ? n75991 : n75941;
  assign n76253 = pi13 ? n75840 : n75779;
  assign n76254 = pi12 ? n76252 : n76253;
  assign n76255 = pi14 ? n61238 : n75564;
  assign n76256 = pi14 ? n34044 : n59560;
  assign n76257 = pi13 ? n76255 : n76256;
  assign n76258 = pi13 ? n75502 : n76225;
  assign n76259 = pi12 ? n76257 : n76258;
  assign n76260 = pi11 ? n76254 : n76259;
  assign n76261 = pi10 ? n76251 : n76260;
  assign n76262 = pi09 ? n76238 : n76261;
  assign n76263 = pi16 ? n1233 : ~n2617;
  assign n76264 = pi15 ? n76206 : n76263;
  assign n76265 = pi14 ? n76264 : n76263;
  assign n76266 = pi13 ? n76241 : n76265;
  assign n76267 = pi15 ? n76263 : n76206;
  assign n76268 = pi14 ? n76267 : n76206;
  assign n76269 = pi13 ? n76263 : n76268;
  assign n76270 = pi12 ? n76266 : n76269;
  assign n76271 = pi14 ? n76206 : n76143;
  assign n76272 = pi13 ? n76271 : n76143;
  assign n76273 = pi13 ? n76090 : n76189;
  assign n76274 = pi12 ? n76272 : n76273;
  assign n76275 = pi11 ? n76270 : n76274;
  assign n76276 = pi13 ? n76042 : n75991;
  assign n76277 = pi13 ? n61712 : n75895;
  assign n76278 = pi12 ? n76276 : n76277;
  assign n76279 = pi14 ? n61506 : n61070;
  assign n76280 = pi13 ? n76279 : n34044;
  assign n76281 = pi14 ? n75598 : n75248;
  assign n76282 = pi13 ? n59560 : n76281;
  assign n76283 = pi12 ? n76280 : n76282;
  assign n76284 = pi11 ? n76278 : n76283;
  assign n76285 = pi10 ? n76275 : n76284;
  assign n76286 = pi09 ? n76238 : n76285;
  assign n76287 = pi08 ? n76262 : n76286;
  assign n76288 = pi07 ? n76231 : n76287;
  assign n76289 = pi16 ? n931 : ~n2745;
  assign n76290 = pi15 ? n32 : n76289;
  assign n76291 = pi14 ? n76290 : n76289;
  assign n76292 = pi13 ? n32 : n76291;
  assign n76293 = pi12 ? n32 : n76292;
  assign n76294 = pi11 ? n32 : n76293;
  assign n76295 = pi10 ? n32 : n76294;
  assign n76296 = pi16 ? n1135 : ~n2745;
  assign n76297 = pi15 ? n76296 : n76263;
  assign n76298 = pi14 ? n76296 : n76297;
  assign n76299 = pi13 ? n76298 : n76263;
  assign n76300 = pi14 ? n76267 : n76264;
  assign n76301 = pi13 ? n76263 : n76300;
  assign n76302 = pi12 ? n76299 : n76301;
  assign n76303 = pi15 ? n76143 : n76038;
  assign n76304 = pi14 ? n76303 : n76038;
  assign n76305 = pi13 ? n76143 : n76304;
  assign n76306 = pi12 ? n76206 : n76305;
  assign n76307 = pi11 ? n76302 : n76306;
  assign n76308 = pi13 ? n61985 : n75895;
  assign n76309 = pi12 ? n76276 : n76308;
  assign n76310 = pi13 ? n76279 : n75977;
  assign n76311 = pi13 ? n75928 : n76281;
  assign n76312 = pi12 ? n76310 : n76311;
  assign n76313 = pi11 ? n76309 : n76312;
  assign n76314 = pi10 ? n76307 : n76313;
  assign n76315 = pi09 ? n76295 : n76314;
  assign n76316 = pi15 ? n76239 : n76263;
  assign n76317 = pi14 ? n76296 : n76316;
  assign n76318 = pi16 ? n1233 : ~n2745;
  assign n76319 = pi15 ? n76263 : n76318;
  assign n76320 = pi14 ? n76319 : n76318;
  assign n76321 = pi13 ? n76317 : n76320;
  assign n76322 = pi15 ? n76318 : n76263;
  assign n76323 = pi14 ? n76322 : n76263;
  assign n76324 = pi13 ? n76318 : n76323;
  assign n76325 = pi12 ? n76321 : n76324;
  assign n76326 = pi14 ? n76263 : n76206;
  assign n76327 = pi13 ? n76326 : n76206;
  assign n76328 = pi14 ? n76146 : n76090;
  assign n76329 = pi13 ? n76143 : n76328;
  assign n76330 = pi12 ? n76327 : n76329;
  assign n76331 = pi11 ? n76325 : n76330;
  assign n76332 = pi13 ? n76094 : n76042;
  assign n76333 = pi13 ? n76099 : n61712;
  assign n76334 = pi12 ? n76332 : n76333;
  assign n76335 = pi14 ? n61505 : n61239;
  assign n76336 = pi13 ? n76335 : n59901;
  assign n76337 = pi14 ? n75653 : n75316;
  assign n76338 = pi13 ? n75977 : n76337;
  assign n76339 = pi12 ? n76336 : n76338;
  assign n76340 = pi11 ? n76334 : n76339;
  assign n76341 = pi10 ? n76331 : n76340;
  assign n76342 = pi09 ? n76295 : n76341;
  assign n76343 = pi08 ? n76315 : n76342;
  assign n76344 = pi16 ? n931 : ~n2732;
  assign n76345 = pi15 ? n32 : n76344;
  assign n76346 = pi14 ? n76345 : n76344;
  assign n76347 = pi13 ? n32 : n76346;
  assign n76348 = pi12 ? n32 : n76347;
  assign n76349 = pi11 ? n32 : n76348;
  assign n76350 = pi10 ? n32 : n76349;
  assign n76351 = pi16 ? n1135 : ~n2732;
  assign n76352 = pi15 ? n76296 : n76318;
  assign n76353 = pi14 ? n76351 : n76352;
  assign n76354 = pi13 ? n76353 : n76318;
  assign n76355 = pi14 ? n76322 : n76319;
  assign n76356 = pi13 ? n76318 : n76355;
  assign n76357 = pi12 ? n76354 : n76356;
  assign n76358 = pi15 ? n76206 : n76090;
  assign n76359 = pi14 ? n76358 : n76090;
  assign n76360 = pi13 ? n76206 : n76359;
  assign n76361 = pi12 ? n76263 : n76360;
  assign n76362 = pi11 ? n76357 : n76361;
  assign n76363 = pi13 ? n75994 : n75892;
  assign n76364 = pi12 ? n76332 : n76363;
  assign n76365 = pi15 ? n61506 : n60190;
  assign n76366 = pi14 ? n61505 : n76365;
  assign n76367 = pi13 ? n76366 : n59901;
  assign n76368 = pi15 ? n59901 : n36601;
  assign n76369 = pi14 ? n76368 : n75441;
  assign n76370 = pi13 ? n59901 : n76369;
  assign n76371 = pi12 ? n76367 : n76370;
  assign n76372 = pi11 ? n76364 : n76371;
  assign n76373 = pi10 ? n76362 : n76372;
  assign n76374 = pi09 ? n76350 : n76373;
  assign n76375 = pi16 ? n1233 : ~n2732;
  assign n76376 = pi15 ? n76318 : n76375;
  assign n76377 = pi14 ? n76376 : n76375;
  assign n76378 = pi13 ? n76353 : n76377;
  assign n76379 = pi15 ? n76375 : n76318;
  assign n76380 = pi14 ? n76379 : n76318;
  assign n76381 = pi13 ? n76375 : n76380;
  assign n76382 = pi12 ? n76378 : n76381;
  assign n76383 = pi14 ? n76318 : n76263;
  assign n76384 = pi13 ? n76383 : n76263;
  assign n76385 = pi12 ? n76384 : n76211;
  assign n76386 = pi11 ? n76382 : n76385;
  assign n76387 = pi13 ? n76213 : n76094;
  assign n76388 = pi13 ? n62214 : n75994;
  assign n76389 = pi12 ? n76387 : n76388;
  assign n76390 = pi14 ? n61710 : n76365;
  assign n76391 = pi13 ? n76390 : n60190;
  assign n76392 = pi14 ? n76368 : n46655;
  assign n76393 = pi13 ? n59901 : n76392;
  assign n76394 = pi12 ? n76391 : n76393;
  assign n76395 = pi11 ? n76389 : n76394;
  assign n76396 = pi10 ? n76386 : n76395;
  assign n76397 = pi09 ? n76350 : n76396;
  assign n76398 = pi08 ? n76374 : n76397;
  assign n76399 = pi07 ? n76343 : n76398;
  assign n76400 = pi06 ? n76288 : n76399;
  assign n76401 = pi16 ? n931 : ~n2725;
  assign n76402 = pi15 ? n32 : n76401;
  assign n76403 = pi14 ? n76402 : n76401;
  assign n76404 = pi13 ? n32 : n76403;
  assign n76405 = pi12 ? n32 : n76404;
  assign n76406 = pi11 ? n32 : n76405;
  assign n76407 = pi10 ? n32 : n76406;
  assign n76408 = pi16 ? n1135 : ~n2725;
  assign n76409 = pi15 ? n76351 : n76375;
  assign n76410 = pi14 ? n76408 : n76409;
  assign n76411 = pi13 ? n76410 : n76375;
  assign n76412 = pi14 ? n76379 : n76376;
  assign n76413 = pi13 ? n76375 : n76412;
  assign n76414 = pi12 ? n76411 : n76413;
  assign n76415 = pi15 ? n76263 : n76143;
  assign n76416 = pi14 ? n76415 : n76143;
  assign n76417 = pi13 ? n76263 : n76416;
  assign n76418 = pi12 ? n76318 : n76417;
  assign n76419 = pi11 ? n76414 : n76418;
  assign n76420 = pi13 ? n76152 : n62214;
  assign n76421 = pi12 ? n76214 : n76420;
  assign n76422 = pi14 ? n62214 : n76157;
  assign n76423 = pi13 ? n76422 : n60190;
  assign n76424 = pi13 ? n60190 : n76392;
  assign n76425 = pi12 ? n76423 : n76424;
  assign n76426 = pi11 ? n76421 : n76425;
  assign n76427 = pi10 ? n76419 : n76426;
  assign n76428 = pi09 ? n76407 : n76427;
  assign n76429 = pi16 ? n1233 : ~n2725;
  assign n76430 = pi15 ? n76375 : n76429;
  assign n76431 = pi14 ? n76430 : n76429;
  assign n76432 = pi13 ? n76410 : n76431;
  assign n76433 = pi15 ? n76429 : n76375;
  assign n76434 = pi14 ? n76433 : n76375;
  assign n76435 = pi13 ? n76429 : n76434;
  assign n76436 = pi12 ? n76432 : n76435;
  assign n76437 = pi14 ? n76375 : n76318;
  assign n76438 = pi13 ? n76437 : n76318;
  assign n76439 = pi12 ? n76438 : n76269;
  assign n76440 = pi11 ? n76436 : n76439;
  assign n76441 = pi14 ? n76206 : n76209;
  assign n76442 = pi13 ? n76441 : n76147;
  assign n76443 = pi13 ? n75988 : n76152;
  assign n76444 = pi12 ? n76442 : n76443;
  assign n76445 = pi13 ? n76422 : n61238;
  assign n76446 = pi14 ? n76368 : n60033;
  assign n76447 = pi13 ? n60190 : n76446;
  assign n76448 = pi12 ? n76445 : n76447;
  assign n76449 = pi11 ? n76444 : n76448;
  assign n76450 = pi10 ? n76440 : n76449;
  assign n76451 = pi09 ? n76407 : n76450;
  assign n76452 = pi08 ? n76428 : n76451;
  assign n76453 = pi16 ? n931 : ~n4246;
  assign n76454 = pi15 ? n32 : n76453;
  assign n76455 = pi14 ? n76454 : n76453;
  assign n76456 = pi13 ? n32 : n76455;
  assign n76457 = pi12 ? n32 : n76456;
  assign n76458 = pi11 ? n32 : n76457;
  assign n76459 = pi10 ? n32 : n76458;
  assign n76460 = pi16 ? n1135 : ~n4246;
  assign n76461 = pi15 ? n76408 : n76429;
  assign n76462 = pi14 ? n76460 : n76461;
  assign n76463 = pi13 ? n76462 : n76429;
  assign n76464 = pi14 ? n76433 : n76430;
  assign n76465 = pi13 ? n76429 : n76464;
  assign n76466 = pi12 ? n76463 : n76465;
  assign n76467 = pi14 ? n76375 : n76379;
  assign n76468 = pi13 ? n76375 : n76467;
  assign n76469 = pi15 ? n76318 : n76206;
  assign n76470 = pi14 ? n76469 : n76206;
  assign n76471 = pi13 ? n76318 : n76470;
  assign n76472 = pi12 ? n76468 : n76471;
  assign n76473 = pi11 ? n76466 : n76472;
  assign n76474 = pi13 ? n76206 : n76441;
  assign n76475 = pi13 ? n76129 : n75988;
  assign n76476 = pi12 ? n76474 : n76475;
  assign n76477 = pi14 ? n75990 : n76157;
  assign n76478 = pi13 ? n76477 : n61238;
  assign n76479 = pi13 ? n61240 : n76446;
  assign n76480 = pi12 ? n76478 : n76479;
  assign n76481 = pi11 ? n76476 : n76480;
  assign n76482 = pi10 ? n76473 : n76481;
  assign n76483 = pi09 ? n76459 : n76482;
  assign n76484 = pi16 ? n1233 : ~n4246;
  assign n76485 = pi15 ? n76429 : n76484;
  assign n76486 = pi14 ? n76485 : n76484;
  assign n76487 = pi13 ? n76462 : n76486;
  assign n76488 = pi15 ? n76484 : n76429;
  assign n76489 = pi14 ? n76488 : n76429;
  assign n76490 = pi13 ? n76484 : n76489;
  assign n76491 = pi12 ? n76487 : n76490;
  assign n76492 = pi14 ? n76429 : n76375;
  assign n76493 = pi13 ? n76492 : n76467;
  assign n76494 = pi15 ? n76375 : n76263;
  assign n76495 = pi14 ? n76494 : n76263;
  assign n76496 = pi13 ? n76377 : n76495;
  assign n76497 = pi12 ? n76493 : n76496;
  assign n76498 = pi11 ? n76491 : n76497;
  assign n76499 = pi13 ? n76326 : n76441;
  assign n76500 = pi13 ? n76038 : n76129;
  assign n76501 = pi12 ? n76499 : n76500;
  assign n76502 = pi14 ? n75990 : n61507;
  assign n76503 = pi13 ? n76502 : n75779;
  assign n76504 = pi14 ? n76368 : n36601;
  assign n76505 = pi13 ? n61240 : n76504;
  assign n76506 = pi12 ? n76503 : n76505;
  assign n76507 = pi11 ? n76501 : n76506;
  assign n76508 = pi10 ? n76498 : n76507;
  assign n76509 = pi09 ? n76459 : n76508;
  assign n76510 = pi08 ? n76483 : n76509;
  assign n76511 = pi07 ? n76452 : n76510;
  assign n76512 = pi16 ? n1214 : ~n3068;
  assign n76513 = pi15 ? n32 : n76512;
  assign n76514 = pi16 ? n931 : ~n3068;
  assign n76515 = pi14 ? n76513 : n76514;
  assign n76516 = pi13 ? n32 : n76515;
  assign n76517 = pi12 ? n32 : n76516;
  assign n76518 = pi11 ? n32 : n76517;
  assign n76519 = pi10 ? n32 : n76518;
  assign n76520 = pi16 ? n1135 : ~n3068;
  assign n76521 = pi15 ? n76460 : n76484;
  assign n76522 = pi14 ? n76520 : n76521;
  assign n76523 = pi13 ? n76522 : n76484;
  assign n76524 = pi14 ? n76488 : n76485;
  assign n76525 = pi13 ? n76484 : n76524;
  assign n76526 = pi12 ? n76523 : n76525;
  assign n76527 = pi13 ? n76489 : n76429;
  assign n76528 = pi13 ? n76375 : n76495;
  assign n76529 = pi12 ? n76527 : n76528;
  assign n76530 = pi11 ? n76526 : n76529;
  assign n76531 = pi14 ? n76263 : n76209;
  assign n76532 = pi13 ? n76263 : n76531;
  assign n76533 = pi12 ? n76532 : n76038;
  assign n76534 = pi13 ? n76502 : n61506;
  assign n76535 = pi14 ? n61506 : n61239;
  assign n76536 = pi13 ? n76535 : n76504;
  assign n76537 = pi12 ? n76534 : n76536;
  assign n76538 = pi11 ? n76533 : n76537;
  assign n76539 = pi10 ? n76530 : n76538;
  assign n76540 = pi09 ? n76519 : n76539;
  assign n76541 = pi16 ? n1323 : ~n3068;
  assign n76542 = pi15 ? n32 : n76541;
  assign n76543 = pi14 ? n76542 : n76514;
  assign n76544 = pi13 ? n32 : n76543;
  assign n76545 = pi12 ? n32 : n76544;
  assign n76546 = pi11 ? n32 : n76545;
  assign n76547 = pi10 ? n32 : n76546;
  assign n76548 = pi16 ? n1233 : ~n3068;
  assign n76549 = pi15 ? n76484 : n76548;
  assign n76550 = pi14 ? n76549 : n76548;
  assign n76551 = pi13 ? n76522 : n76550;
  assign n76552 = pi15 ? n76548 : n76484;
  assign n76553 = pi14 ? n76552 : n76484;
  assign n76554 = pi13 ? n76548 : n76553;
  assign n76555 = pi12 ? n76551 : n76554;
  assign n76556 = pi14 ? n76484 : n76429;
  assign n76557 = pi13 ? n76556 : n76429;
  assign n76558 = pi15 ? n76429 : n76318;
  assign n76559 = pi14 ? n76558 : n76318;
  assign n76560 = pi13 ? n76429 : n76559;
  assign n76561 = pi12 ? n76557 : n76560;
  assign n76562 = pi11 ? n76555 : n76561;
  assign n76563 = pi13 ? n76383 : n76531;
  assign n76564 = pi13 ? n76090 : n76038;
  assign n76565 = pi12 ? n76563 : n76564;
  assign n76566 = pi14 ? n75990 : n61505;
  assign n76567 = pi13 ? n76566 : n75895;
  assign n76568 = pi13 ? n76535 : n75718;
  assign n76569 = pi12 ? n76567 : n76568;
  assign n76570 = pi11 ? n76565 : n76569;
  assign n76571 = pi10 ? n76562 : n76570;
  assign n76572 = pi09 ? n76547 : n76571;
  assign n76573 = pi08 ? n76540 : n76572;
  assign n76574 = pi16 ? n1323 : ~n2851;
  assign n76575 = pi15 ? n32 : n76574;
  assign n76576 = pi16 ? n1471 : ~n2851;
  assign n76577 = pi16 ? n1479 : ~n2851;
  assign n76578 = pi15 ? n76576 : n76577;
  assign n76579 = pi14 ? n76575 : n76578;
  assign n76580 = pi13 ? n32 : n76579;
  assign n76581 = pi12 ? n32 : n76580;
  assign n76582 = pi11 ? n32 : n76581;
  assign n76583 = pi10 ? n32 : n76582;
  assign n76584 = pi16 ? n931 : ~n2851;
  assign n76585 = pi16 ? n1135 : ~n2851;
  assign n76586 = pi15 ? n76584 : n76585;
  assign n76587 = pi15 ? n76520 : n76548;
  assign n76588 = pi14 ? n76586 : n76587;
  assign n76589 = pi13 ? n76588 : n76548;
  assign n76590 = pi13 ? n76548 : n76550;
  assign n76591 = pi12 ? n76589 : n76590;
  assign n76592 = pi14 ? n76548 : n76484;
  assign n76593 = pi14 ? n76484 : n76488;
  assign n76594 = pi13 ? n76592 : n76593;
  assign n76595 = pi13 ? n76429 : n76380;
  assign n76596 = pi12 ? n76594 : n76595;
  assign n76597 = pi11 ? n76591 : n76596;
  assign n76598 = pi14 ? n76322 : n76206;
  assign n76599 = pi13 ? n76318 : n76598;
  assign n76600 = pi12 ? n76599 : n76090;
  assign n76601 = pi14 ? n76039 : n61505;
  assign n76602 = pi13 ? n76601 : n61505;
  assign n76603 = pi14 ? n61505 : n75778;
  assign n76604 = pi15 ? n60190 : n59560;
  assign n76605 = pi14 ? n76604 : n59560;
  assign n76606 = pi13 ? n76603 : n76605;
  assign n76607 = pi12 ? n76602 : n76606;
  assign n76608 = pi11 ? n76600 : n76607;
  assign n76609 = pi10 ? n76597 : n76608;
  assign n76610 = pi09 ? n76583 : n76609;
  assign n76611 = pi16 ? n1577 : ~n2851;
  assign n76612 = pi15 ? n32 : n76611;
  assign n76613 = pi16 ? n1581 : ~n2851;
  assign n76614 = pi15 ? n76613 : n76574;
  assign n76615 = pi14 ? n76612 : n76614;
  assign n76616 = pi13 ? n32 : n76615;
  assign n76617 = pi12 ? n32 : n76616;
  assign n76618 = pi11 ? n32 : n76617;
  assign n76619 = pi10 ? n32 : n76618;
  assign n76620 = pi16 ? n1594 : ~n2851;
  assign n76621 = pi15 ? n76620 : n76585;
  assign n76622 = pi14 ? n76621 : n76587;
  assign n76623 = pi16 ? n1233 : ~n2851;
  assign n76624 = pi15 ? n76548 : n76623;
  assign n76625 = pi14 ? n76624 : n76623;
  assign n76626 = pi13 ? n76622 : n76625;
  assign n76627 = pi15 ? n76623 : n76548;
  assign n76628 = pi14 ? n76627 : n76548;
  assign n76629 = pi13 ? n76623 : n76628;
  assign n76630 = pi12 ? n76626 : n76629;
  assign n76631 = pi13 ? n76592 : n76484;
  assign n76632 = pi13 ? n76593 : n76434;
  assign n76633 = pi12 ? n76631 : n76632;
  assign n76634 = pi11 ? n76630 : n76633;
  assign n76635 = pi14 ? n76322 : n76209;
  assign n76636 = pi13 ? n76380 : n76635;
  assign n76637 = pi13 ? n76147 : n76094;
  assign n76638 = pi12 ? n76636 : n76637;
  assign n76639 = pi13 ? n76130 : n61712;
  assign n76640 = pi14 ? n61507 : n61239;
  assign n76641 = pi13 ? n76640 : n75949;
  assign n76642 = pi12 ? n76639 : n76641;
  assign n76643 = pi11 ? n76638 : n76642;
  assign n76644 = pi10 ? n76634 : n76643;
  assign n76645 = pi09 ? n76619 : n76644;
  assign n76646 = pi08 ? n76610 : n76645;
  assign n76647 = pi07 ? n76573 : n76646;
  assign n76648 = pi06 ? n76511 : n76647;
  assign n76649 = pi05 ? n76400 : n76648;
  assign n76650 = pi04 ? n76173 : n76649;
  assign n76651 = pi16 ? n1678 : ~n2840;
  assign n76652 = pi15 ? n32 : n76651;
  assign n76653 = pi16 ? n1683 : ~n2840;
  assign n76654 = pi16 ? n1323 : ~n2840;
  assign n76655 = pi15 ? n76653 : n76654;
  assign n76656 = pi14 ? n76652 : n76655;
  assign n76657 = pi13 ? n32 : n76656;
  assign n76658 = pi12 ? n32 : n76657;
  assign n76659 = pi11 ? n32 : n76658;
  assign n76660 = pi10 ? n32 : n76659;
  assign n76661 = pi16 ? n1594 : ~n2840;
  assign n76662 = pi16 ? n1479 : ~n2840;
  assign n76663 = pi15 ? n76661 : n76662;
  assign n76664 = pi16 ? n1705 : ~n2851;
  assign n76665 = pi15 ? n76664 : n76585;
  assign n76666 = pi14 ? n76663 : n76665;
  assign n76667 = pi13 ? n76666 : n76623;
  assign n76668 = pi12 ? n76667 : n76623;
  assign n76669 = pi14 ? n76623 : n76548;
  assign n76670 = pi14 ? n76548 : n76552;
  assign n76671 = pi13 ? n76669 : n76670;
  assign n76672 = pi12 ? n76671 : n76632;
  assign n76673 = pi11 ? n76668 : n76672;
  assign n76674 = pi14 ? n76379 : n76415;
  assign n76675 = pi13 ? n76375 : n76674;
  assign n76676 = pi12 ? n76675 : n76148;
  assign n76677 = pi14 ? n76039 : n61710;
  assign n76678 = pi13 ? n76677 : n61710;
  assign n76679 = pi14 ? n61711 : n75778;
  assign n76680 = pi13 ? n76679 : n75785;
  assign n76681 = pi12 ? n76678 : n76680;
  assign n76682 = pi11 ? n76676 : n76681;
  assign n76683 = pi10 ? n76673 : n76682;
  assign n76684 = pi09 ? n76660 : n76683;
  assign n76685 = pi16 ? n1808 : ~n2840;
  assign n76686 = pi15 ? n32 : n76685;
  assign n76687 = pi16 ? n1815 : ~n2840;
  assign n76688 = pi15 ? n76687 : n76653;
  assign n76689 = pi14 ? n76686 : n76688;
  assign n76690 = pi13 ? n32 : n76689;
  assign n76691 = pi12 ? n32 : n76690;
  assign n76692 = pi11 ? n32 : n76691;
  assign n76693 = pi10 ? n32 : n76692;
  assign n76694 = pi16 ? n1834 : ~n2840;
  assign n76695 = pi15 ? n76694 : n76654;
  assign n76696 = pi16 ? n1843 : ~n2851;
  assign n76697 = pi15 ? n76620 : n76696;
  assign n76698 = pi14 ? n76695 : n76697;
  assign n76699 = pi16 ? n1233 : ~n2840;
  assign n76700 = pi13 ? n76698 : n76699;
  assign n76701 = pi15 ? n76699 : n76623;
  assign n76702 = pi14 ? n76701 : n76623;
  assign n76703 = pi13 ? n76699 : n76702;
  assign n76704 = pi12 ? n76700 : n76703;
  assign n76705 = pi13 ? n76669 : n76548;
  assign n76706 = pi13 ? n76670 : n76429;
  assign n76707 = pi12 ? n76705 : n76706;
  assign n76708 = pi11 ? n76704 : n76707;
  assign n76709 = pi14 ? n76379 : n76267;
  assign n76710 = pi13 ? n76434 : n76709;
  assign n76711 = pi12 ? n76710 : n76442;
  assign n76712 = pi13 ? n76190 : n61710;
  assign n76713 = pi12 ? n76712 : n76680;
  assign n76714 = pi11 ? n76711 : n76713;
  assign n76715 = pi10 ? n76708 : n76714;
  assign n76716 = pi09 ? n76693 : n76715;
  assign n76717 = pi08 ? n76684 : n76716;
  assign n76718 = pi16 ? n1934 : ~n2837;
  assign n76719 = pi15 ? n32 : n76718;
  assign n76720 = pi16 ? n1815 : ~n2837;
  assign n76721 = pi16 ? n1944 : ~n2837;
  assign n76722 = pi15 ? n76720 : n76721;
  assign n76723 = pi14 ? n76719 : n76722;
  assign n76724 = pi13 ? n32 : n76723;
  assign n76725 = pi12 ? n32 : n76724;
  assign n76726 = pi11 ? n32 : n76725;
  assign n76727 = pi10 ? n32 : n76726;
  assign n76728 = pi16 ? n1683 : ~n2837;
  assign n76729 = pi16 ? n1577 : ~n2837;
  assign n76730 = pi15 ? n76728 : n76729;
  assign n76731 = pi16 ? n1594 : ~n2837;
  assign n76732 = pi16 ? n1471 : ~n2840;
  assign n76733 = pi15 ? n76731 : n76732;
  assign n76734 = pi14 ? n76730 : n76733;
  assign n76735 = pi16 ? n1705 : ~n2840;
  assign n76736 = pi16 ? n1972 : ~n2840;
  assign n76737 = pi15 ? n76735 : n76736;
  assign n76738 = pi16 ? n1135 : ~n2840;
  assign n76739 = pi15 ? n76738 : n76699;
  assign n76740 = pi14 ? n76737 : n76739;
  assign n76741 = pi13 ? n76734 : n76740;
  assign n76742 = pi12 ? n76741 : n76699;
  assign n76743 = pi14 ? n76699 : n76623;
  assign n76744 = pi14 ? n76623 : n76627;
  assign n76745 = pi13 ? n76743 : n76744;
  assign n76746 = pi12 ? n76745 : n76706;
  assign n76747 = pi11 ? n76742 : n76746;
  assign n76748 = pi14 ? n76433 : n76469;
  assign n76749 = pi13 ? n76429 : n76748;
  assign n76750 = pi12 ? n76749 : n76474;
  assign n76751 = pi14 ? n76091 : n62214;
  assign n76752 = pi13 ? n76751 : n62214;
  assign n76753 = pi14 ? n61710 : n61507;
  assign n76754 = pi15 ? n61238 : n34044;
  assign n76755 = pi14 ? n76754 : n34044;
  assign n76756 = pi13 ? n76753 : n76755;
  assign n76757 = pi12 ? n76752 : n76756;
  assign n76758 = pi11 ? n76750 : n76757;
  assign n76759 = pi10 ? n76747 : n76758;
  assign n76760 = pi09 ? n76727 : n76759;
  assign n76761 = pi16 ? n2120 : ~n2837;
  assign n76762 = pi15 ? n32 : n76761;
  assign n76763 = pi16 ? n1808 : ~n2837;
  assign n76764 = pi15 ? n76718 : n76763;
  assign n76765 = pi14 ? n76762 : n76764;
  assign n76766 = pi13 ? n32 : n76765;
  assign n76767 = pi12 ? n32 : n76766;
  assign n76768 = pi11 ? n32 : n76767;
  assign n76769 = pi10 ? n32 : n76768;
  assign n76770 = pi16 ? n2137 : ~n2837;
  assign n76771 = pi15 ? n76720 : n76770;
  assign n76772 = pi16 ? n2144 : ~n2840;
  assign n76773 = pi15 ? n76729 : n76772;
  assign n76774 = pi14 ? n76771 : n76773;
  assign n76775 = pi16 ? n1843 : ~n2837;
  assign n76776 = pi15 ? n76731 : n76775;
  assign n76777 = pi16 ? n1233 : ~n2837;
  assign n76778 = pi15 ? n76775 : n76777;
  assign n76779 = pi14 ? n76776 : n76778;
  assign n76780 = pi13 ? n76774 : n76779;
  assign n76781 = pi15 ? n76777 : n76699;
  assign n76782 = pi14 ? n76781 : n76699;
  assign n76783 = pi13 ? n76777 : n76782;
  assign n76784 = pi12 ? n76780 : n76783;
  assign n76785 = pi13 ? n76702 : n76623;
  assign n76786 = pi13 ? n76744 : n76484;
  assign n76787 = pi12 ? n76785 : n76786;
  assign n76788 = pi11 ? n76784 : n76787;
  assign n76789 = pi14 ? n76433 : n76322;
  assign n76790 = pi13 ? n76489 : n76789;
  assign n76791 = pi12 ? n76790 : n76499;
  assign n76792 = pi13 ? n76753 : n75845;
  assign n76793 = pi12 ? n76752 : n76792;
  assign n76794 = pi11 ? n76791 : n76793;
  assign n76795 = pi10 ? n76788 : n76794;
  assign n76796 = pi09 ? n76769 : n76795;
  assign n76797 = pi08 ? n76760 : n76796;
  assign n76798 = pi07 ? n76717 : n76797;
  assign n76799 = pi16 ? n2293 : ~n3061;
  assign n76800 = pi15 ? n32 : n76799;
  assign n76801 = pi16 ? n2300 : ~n3061;
  assign n76802 = pi16 ? n2306 : ~n3061;
  assign n76803 = pi15 ? n76801 : n76802;
  assign n76804 = pi14 ? n76800 : n76803;
  assign n76805 = pi13 ? n32 : n76804;
  assign n76806 = pi12 ? n32 : n76805;
  assign n76807 = pi11 ? n32 : n76806;
  assign n76808 = pi10 ? n32 : n76807;
  assign n76809 = pi16 ? n1934 : ~n3061;
  assign n76810 = pi16 ? n2320 : ~n3061;
  assign n76811 = pi15 ? n76809 : n76810;
  assign n76812 = pi16 ? n2137 : ~n3061;
  assign n76813 = pi16 ? n2326 : ~n2837;
  assign n76814 = pi15 ? n76812 : n76813;
  assign n76815 = pi14 ? n76811 : n76814;
  assign n76816 = pi16 ? n1834 : ~n2837;
  assign n76817 = pi15 ? n76729 : n76816;
  assign n76818 = pi16 ? n1471 : ~n2837;
  assign n76819 = pi15 ? n76775 : n76818;
  assign n76820 = pi14 ? n76817 : n76819;
  assign n76821 = pi13 ? n76815 : n76820;
  assign n76822 = pi16 ? n1705 : ~n2837;
  assign n76823 = pi16 ? n1972 : ~n2837;
  assign n76824 = pi15 ? n76822 : n76823;
  assign n76825 = pi16 ? n1135 : ~n2837;
  assign n76826 = pi15 ? n76825 : n76777;
  assign n76827 = pi14 ? n76824 : n76826;
  assign n76828 = pi13 ? n76827 : n76777;
  assign n76829 = pi12 ? n76821 : n76828;
  assign n76830 = pi14 ? n76699 : n76701;
  assign n76831 = pi13 ? n76782 : n76830;
  assign n76832 = pi12 ? n76831 : n76786;
  assign n76833 = pi11 ? n76829 : n76832;
  assign n76834 = pi15 ? n76484 : n76375;
  assign n76835 = pi14 ? n76834 : n76322;
  assign n76836 = pi13 ? n76484 : n76835;
  assign n76837 = pi12 ? n76836 : n76532;
  assign n76838 = pi14 ? n75940 : n61507;
  assign n76839 = pi13 ? n76838 : n76028;
  assign n76840 = pi12 ? n76752 : n76839;
  assign n76841 = pi11 ? n76837 : n76840;
  assign n76842 = pi10 ? n76833 : n76841;
  assign n76843 = pi09 ? n76808 : n76842;
  assign n76844 = pi16 ? n2409 : ~n3061;
  assign n76845 = pi16 ? n2415 : ~n3061;
  assign n76846 = pi15 ? n76844 : n76845;
  assign n76847 = pi14 ? n76800 : n76846;
  assign n76848 = pi13 ? n32 : n76847;
  assign n76849 = pi12 ? n32 : n76848;
  assign n76850 = pi11 ? n32 : n76849;
  assign n76851 = pi10 ? n32 : n76850;
  assign n76852 = pi16 ? n2120 : ~n3061;
  assign n76853 = pi16 ? n2426 : ~n3061;
  assign n76854 = pi15 ? n76852 : n76853;
  assign n76855 = pi15 ? n76810 : n76720;
  assign n76856 = pi14 ? n76854 : n76855;
  assign n76857 = pi16 ? n1944 : ~n3061;
  assign n76858 = pi15 ? n76812 : n76857;
  assign n76859 = pi16 ? n1834 : ~n3061;
  assign n76860 = pi16 ? n2144 : ~n3061;
  assign n76861 = pi15 ? n76859 : n76860;
  assign n76862 = pi14 ? n76858 : n76861;
  assign n76863 = pi13 ? n76856 : n76862;
  assign n76864 = pi16 ? n1594 : ~n3061;
  assign n76865 = pi16 ? n1843 : ~n3061;
  assign n76866 = pi15 ? n76864 : n76865;
  assign n76867 = pi16 ? n1233 : ~n3061;
  assign n76868 = pi15 ? n76865 : n76867;
  assign n76869 = pi14 ? n76866 : n76868;
  assign n76870 = pi15 ? n76867 : n76777;
  assign n76871 = pi14 ? n76870 : n76777;
  assign n76872 = pi13 ? n76869 : n76871;
  assign n76873 = pi12 ? n76863 : n76872;
  assign n76874 = pi13 ? n76782 : n76699;
  assign n76875 = pi13 ? n76830 : n76548;
  assign n76876 = pi12 ? n76874 : n76875;
  assign n76877 = pi11 ? n76873 : n76876;
  assign n76878 = pi14 ? n76488 : n76379;
  assign n76879 = pi13 ? n76484 : n76878;
  assign n76880 = pi13 ? n76263 : n76326;
  assign n76881 = pi12 ? n76879 : n76880;
  assign n76882 = pi14 ? n76146 : n75988;
  assign n76883 = pi13 ? n76882 : n75988;
  assign n76884 = pi14 ? n62214 : n76219;
  assign n76885 = pi13 ? n76884 : n75897;
  assign n76886 = pi12 ? n76883 : n76885;
  assign n76887 = pi11 ? n76881 : n76886;
  assign n76888 = pi10 ? n76877 : n76887;
  assign n76889 = pi09 ? n76851 : n76888;
  assign n76890 = pi08 ? n76843 : n76889;
  assign n76891 = pi16 ? n2513 : ~n2832;
  assign n76892 = pi15 ? n32 : n76891;
  assign n76893 = pi16 ? n2518 : ~n2832;
  assign n76894 = pi14 ? n76892 : n76893;
  assign n76895 = pi13 ? n32 : n76894;
  assign n76896 = pi12 ? n32 : n76895;
  assign n76897 = pi11 ? n32 : n76896;
  assign n76898 = pi10 ? n32 : n76897;
  assign n76899 = pi16 ? n2293 : ~n2832;
  assign n76900 = pi16 ? n2409 : ~n2832;
  assign n76901 = pi15 ? n76899 : n76900;
  assign n76902 = pi16 ? n2530 : ~n2832;
  assign n76903 = pi15 ? n76902 : n76809;
  assign n76904 = pi14 ? n76901 : n76903;
  assign n76905 = pi16 ? n2540 : ~n3061;
  assign n76906 = pi15 ? n76810 : n76905;
  assign n76907 = pi16 ? n2326 : ~n3061;
  assign n76908 = pi15 ? n76857 : n76907;
  assign n76909 = pi14 ? n76906 : n76908;
  assign n76910 = pi13 ? n76904 : n76909;
  assign n76911 = pi16 ? n1577 : ~n3061;
  assign n76912 = pi15 ? n76911 : n76859;
  assign n76913 = pi16 ? n1471 : ~n3061;
  assign n76914 = pi15 ? n76865 : n76913;
  assign n76915 = pi14 ? n76912 : n76914;
  assign n76916 = pi16 ? n1705 : ~n3061;
  assign n76917 = pi16 ? n1972 : ~n3061;
  assign n76918 = pi15 ? n76916 : n76917;
  assign n76919 = pi16 ? n1135 : ~n3061;
  assign n76920 = pi15 ? n76919 : n76867;
  assign n76921 = pi14 ? n76918 : n76920;
  assign n76922 = pi13 ? n76915 : n76921;
  assign n76923 = pi12 ? n76910 : n76922;
  assign n76924 = pi14 ? n76777 : n76781;
  assign n76925 = pi13 ? n76871 : n76924;
  assign n76926 = pi12 ? n76925 : n76875;
  assign n76927 = pi11 ? n76923 : n76926;
  assign n76928 = pi13 ? n76548 : n76878;
  assign n76929 = pi14 ? n76263 : n76267;
  assign n76930 = pi13 ? n76263 : n76929;
  assign n76931 = pi12 ? n76928 : n76930;
  assign n76932 = pi11 ? n76931 : n76886;
  assign n76933 = pi10 ? n76927 : n76932;
  assign n76934 = pi09 ? n76898 : n76933;
  assign n76935 = pi16 ? n2617 : ~n2832;
  assign n76936 = pi15 ? n32 : n76935;
  assign n76937 = pi16 ? n2624 : ~n2832;
  assign n76938 = pi16 ? n2629 : ~n2832;
  assign n76939 = pi15 ? n76937 : n76938;
  assign n76940 = pi14 ? n76936 : n76939;
  assign n76941 = pi13 ? n32 : n76940;
  assign n76942 = pi12 ? n32 : n76941;
  assign n76943 = pi11 ? n32 : n76942;
  assign n76944 = pi10 ? n32 : n76943;
  assign n76945 = pi15 ? n76891 : n76900;
  assign n76946 = pi16 ? n2415 : ~n2832;
  assign n76947 = pi15 ? n76946 : n76852;
  assign n76948 = pi14 ? n76945 : n76947;
  assign n76949 = pi16 ? n2426 : ~n2832;
  assign n76950 = pi16 ? n2654 : ~n2832;
  assign n76951 = pi15 ? n76949 : n76950;
  assign n76952 = pi16 ? n2540 : ~n2832;
  assign n76953 = pi16 ? n1815 : ~n2832;
  assign n76954 = pi15 ? n76952 : n76953;
  assign n76955 = pi14 ? n76951 : n76954;
  assign n76956 = pi13 ? n76948 : n76955;
  assign n76957 = pi16 ? n2137 : ~n2832;
  assign n76958 = pi16 ? n1944 : ~n2832;
  assign n76959 = pi15 ? n76957 : n76958;
  assign n76960 = pi16 ? n1834 : ~n2832;
  assign n76961 = pi16 ? n2144 : ~n2832;
  assign n76962 = pi15 ? n76960 : n76961;
  assign n76963 = pi14 ? n76959 : n76962;
  assign n76964 = pi16 ? n1594 : ~n2832;
  assign n76965 = pi15 ? n76964 : n76865;
  assign n76966 = pi14 ? n76965 : n76868;
  assign n76967 = pi13 ? n76963 : n76966;
  assign n76968 = pi12 ? n76956 : n76967;
  assign n76969 = pi13 ? n76871 : n76777;
  assign n76970 = pi13 ? n76924 : n76669;
  assign n76971 = pi12 ? n76969 : n76970;
  assign n76972 = pi11 ? n76968 : n76971;
  assign n76973 = pi14 ? n76484 : n76433;
  assign n76974 = pi13 ? n76548 : n76973;
  assign n76975 = pi13 ? n76318 : n76383;
  assign n76976 = pi12 ? n76974 : n76975;
  assign n76977 = pi14 ? n76358 : n76038;
  assign n76978 = pi13 ? n76977 : n76042;
  assign n76979 = pi14 ? n75990 : n61711;
  assign n76980 = pi14 ? n75778 : n61239;
  assign n76981 = pi13 ? n76979 : n76980;
  assign n76982 = pi12 ? n76978 : n76981;
  assign n76983 = pi11 ? n76976 : n76982;
  assign n76984 = pi10 ? n76972 : n76983;
  assign n76985 = pi09 ? n76944 : n76984;
  assign n76986 = pi08 ? n76934 : n76985;
  assign n76987 = pi07 ? n76890 : n76986;
  assign n76988 = pi06 ? n76798 : n76987;
  assign n76989 = pi16 ? n2725 : ~n3183;
  assign n76990 = pi15 ? n32 : n76989;
  assign n76991 = pi16 ? n2732 : ~n3183;
  assign n76992 = pi14 ? n76990 : n76991;
  assign n76993 = pi13 ? n32 : n76992;
  assign n76994 = pi12 ? n32 : n76993;
  assign n76995 = pi11 ? n32 : n76994;
  assign n76996 = pi10 ? n32 : n76995;
  assign n76997 = pi16 ? n2745 : ~n3183;
  assign n76998 = pi16 ? n2749 : ~n3183;
  assign n76999 = pi15 ? n76997 : n76998;
  assign n77000 = pi16 ? n2756 : ~n3183;
  assign n77001 = pi16 ? n2756 : ~n2832;
  assign n77002 = pi15 ? n77000 : n77001;
  assign n77003 = pi14 ? n76999 : n77002;
  assign n77004 = pi15 ? n76900 : n76946;
  assign n77005 = pi16 ? n2306 : ~n2832;
  assign n77006 = pi16 ? n1934 : ~n2832;
  assign n77007 = pi15 ? n77005 : n77006;
  assign n77008 = pi14 ? n77004 : n77007;
  assign n77009 = pi13 ? n77003 : n77008;
  assign n77010 = pi16 ? n2320 : ~n2832;
  assign n77011 = pi15 ? n77010 : n76952;
  assign n77012 = pi16 ? n2326 : ~n2832;
  assign n77013 = pi15 ? n76958 : n77012;
  assign n77014 = pi14 ? n77011 : n77013;
  assign n77015 = pi16 ? n1577 : ~n2832;
  assign n77016 = pi15 ? n77015 : n76960;
  assign n77017 = pi16 ? n1843 : ~n2832;
  assign n77018 = pi16 ? n1471 : ~n2832;
  assign n77019 = pi15 ? n77017 : n77018;
  assign n77020 = pi14 ? n77016 : n77019;
  assign n77021 = pi13 ? n77014 : n77020;
  assign n77022 = pi12 ? n77009 : n77021;
  assign n77023 = pi16 ? n1705 : ~n2832;
  assign n77024 = pi15 ? n77023 : n76916;
  assign n77025 = pi16 ? n931 : ~n3061;
  assign n77026 = pi15 ? n77025 : n76919;
  assign n77027 = pi14 ? n77024 : n77026;
  assign n77028 = pi14 ? n76867 : n76777;
  assign n77029 = pi13 ? n77027 : n77028;
  assign n77030 = pi12 ? n77029 : n76970;
  assign n77031 = pi11 ? n77022 : n77030;
  assign n77032 = pi14 ? n76552 : n76433;
  assign n77033 = pi13 ? n76548 : n77032;
  assign n77034 = pi12 ? n77033 : n76975;
  assign n77035 = pi13 ? n76979 : n75945;
  assign n77036 = pi12 ? n76978 : n77035;
  assign n77037 = pi11 ? n77034 : n77036;
  assign n77038 = pi10 ? n77031 : n77037;
  assign n77039 = pi09 ? n76996 : n77038;
  assign n77040 = pi16 ? n2832 : ~n3183;
  assign n77041 = pi15 ? n32 : n77040;
  assign n77042 = pi16 ? n2837 : ~n3183;
  assign n77043 = pi16 ? n2840 : ~n3183;
  assign n77044 = pi15 ? n77042 : n77043;
  assign n77045 = pi14 ? n77041 : n77044;
  assign n77046 = pi13 ? n32 : n77045;
  assign n77047 = pi12 ? n32 : n77046;
  assign n77048 = pi11 ? n32 : n77047;
  assign n77049 = pi10 ? n32 : n77048;
  assign n77050 = pi16 ? n2851 : ~n3183;
  assign n77051 = pi16 ? n2856 : ~n3183;
  assign n77052 = pi15 ? n77050 : n77051;
  assign n77053 = pi16 ? n2860 : ~n3183;
  assign n77054 = pi15 ? n77053 : n76891;
  assign n77055 = pi14 ? n77052 : n77054;
  assign n77056 = pi16 ? n2415 : ~n3183;
  assign n77057 = pi15 ? n76998 : n77056;
  assign n77058 = pi16 ? n2120 : ~n3183;
  assign n77059 = pi15 ? n77056 : n77058;
  assign n77060 = pi14 ? n77057 : n77059;
  assign n77061 = pi13 ? n77055 : n77060;
  assign n77062 = pi16 ? n2426 : ~n3183;
  assign n77063 = pi16 ? n2654 : ~n3183;
  assign n77064 = pi15 ? n77062 : n77063;
  assign n77065 = pi16 ? n2540 : ~n3183;
  assign n77066 = pi16 ? n1815 : ~n3183;
  assign n77067 = pi15 ? n77065 : n77066;
  assign n77068 = pi14 ? n77064 : n77067;
  assign n77069 = pi16 ? n2137 : ~n3183;
  assign n77070 = pi15 ? n77069 : n76958;
  assign n77071 = pi14 ? n77070 : n76962;
  assign n77072 = pi13 ? n77068 : n77071;
  assign n77073 = pi12 ? n77061 : n77072;
  assign n77074 = pi15 ? n76964 : n76864;
  assign n77075 = pi14 ? n77074 : n76866;
  assign n77076 = pi16 ? n1479 : ~n3061;
  assign n77077 = pi16 ? n1214 : ~n3061;
  assign n77078 = pi15 ? n77077 : n77025;
  assign n77079 = pi14 ? n77076 : n77078;
  assign n77080 = pi13 ? n77075 : n77079;
  assign n77081 = pi13 ? n77028 : n76743;
  assign n77082 = pi12 ? n77080 : n77081;
  assign n77083 = pi11 ? n77073 : n77082;
  assign n77084 = pi14 ? n76548 : n76834;
  assign n77085 = pi13 ? n76623 : n77084;
  assign n77086 = pi14 ? n76379 : n76322;
  assign n77087 = pi13 ? n76375 : n77086;
  assign n77088 = pi12 ? n77085 : n77087;
  assign n77089 = pi14 ? n76209 : n76090;
  assign n77090 = pi13 ? n77089 : n76189;
  assign n77091 = pi13 ? n76130 : n75973;
  assign n77092 = pi12 ? n77090 : n77091;
  assign n77093 = pi11 ? n77088 : n77092;
  assign n77094 = pi10 ? n77083 : n77093;
  assign n77095 = pi09 ? n77049 : n77094;
  assign n77096 = pi08 ? n77039 : n77095;
  assign n77097 = pi16 ? n2953 : ~n2964;
  assign n77098 = pi15 ? n32 : n77097;
  assign n77099 = pi16 ? n2958 : ~n2964;
  assign n77100 = pi16 ? n2964 : ~n2964;
  assign n77101 = pi15 ? n77099 : n77100;
  assign n77102 = pi14 ? n77098 : n77101;
  assign n77103 = pi13 ? n32 : n77102;
  assign n77104 = pi12 ? n32 : n77103;
  assign n77105 = pi11 ? n32 : n77104;
  assign n77106 = pi10 ? n32 : n77105;
  assign n77107 = pi16 ? n2732 : ~n2964;
  assign n77108 = pi15 ? n77100 : n77107;
  assign n77109 = pi16 ? n2745 : ~n2964;
  assign n77110 = pi15 ? n77109 : n76997;
  assign n77111 = pi14 ? n77108 : n77110;
  assign n77112 = pi16 ? n2617 : ~n3183;
  assign n77113 = pi16 ? n2518 : ~n3183;
  assign n77114 = pi15 ? n77112 : n77113;
  assign n77115 = pi14 ? n77114 : n77000;
  assign n77116 = pi13 ? n77111 : n77115;
  assign n77117 = pi16 ? n2409 : ~n3183;
  assign n77118 = pi15 ? n77117 : n77056;
  assign n77119 = pi16 ? n2306 : ~n3183;
  assign n77120 = pi16 ? n1934 : ~n3183;
  assign n77121 = pi15 ? n77119 : n77120;
  assign n77122 = pi14 ? n77118 : n77121;
  assign n77123 = pi16 ? n2320 : ~n3183;
  assign n77124 = pi15 ? n77123 : n77065;
  assign n77125 = pi16 ? n1944 : ~n3183;
  assign n77126 = pi16 ? n2326 : ~n3183;
  assign n77127 = pi15 ? n77125 : n77126;
  assign n77128 = pi14 ? n77124 : n77127;
  assign n77129 = pi13 ? n77122 : n77128;
  assign n77130 = pi12 ? n77116 : n77129;
  assign n77131 = pi16 ? n1577 : ~n3183;
  assign n77132 = pi15 ? n77131 : n77015;
  assign n77133 = pi14 ? n77132 : n77016;
  assign n77134 = pi16 ? n1323 : ~n3061;
  assign n77135 = pi15 ? n77134 : n76864;
  assign n77136 = pi14 ? n77134 : n77135;
  assign n77137 = pi13 ? n77133 : n77136;
  assign n77138 = pi16 ? n1214 : ~n2837;
  assign n77139 = pi15 ? n76917 : n77138;
  assign n77140 = pi14 ? n76913 : n77139;
  assign n77141 = pi16 ? n931 : ~n2840;
  assign n77142 = pi15 ? n76585 : n76623;
  assign n77143 = pi14 ? n77141 : n77142;
  assign n77144 = pi13 ? n77140 : n77143;
  assign n77145 = pi12 ? n77137 : n77144;
  assign n77146 = pi11 ? n77130 : n77145;
  assign n77147 = pi12 ? n77085 : n76381;
  assign n77148 = pi13 ? n77089 : n76150;
  assign n77149 = pi14 ? n61507 : n75778;
  assign n77150 = pi13 ? n76677 : n77149;
  assign n77151 = pi12 ? n77148 : n77150;
  assign n77152 = pi11 ? n77147 : n77151;
  assign n77153 = pi10 ? n77146 : n77152;
  assign n77154 = pi09 ? n77106 : n77153;
  assign n77155 = pi16 ? n3047 : ~n2964;
  assign n77156 = pi15 ? n32 : n77155;
  assign n77157 = pi16 ? n3051 : ~n2964;
  assign n77158 = pi14 ? n77156 : n77157;
  assign n77159 = pi13 ? n32 : n77158;
  assign n77160 = pi12 ? n32 : n77159;
  assign n77161 = pi11 ? n32 : n77160;
  assign n77162 = pi10 ? n32 : n77161;
  assign n77163 = pi16 ? n3061 : ~n2964;
  assign n77164 = pi15 ? n77097 : n77163;
  assign n77165 = pi16 ? n2840 : ~n2964;
  assign n77166 = pi15 ? n77165 : n77050;
  assign n77167 = pi14 ? n77164 : n77166;
  assign n77168 = pi16 ? n3068 : ~n2964;
  assign n77169 = pi16 ? n2624 : ~n2964;
  assign n77170 = pi15 ? n77168 : n77169;
  assign n77171 = pi16 ? n2860 : ~n2964;
  assign n77172 = pi16 ? n2513 : ~n2964;
  assign n77173 = pi15 ? n77171 : n77172;
  assign n77174 = pi14 ? n77170 : n77173;
  assign n77175 = pi13 ? n77167 : n77174;
  assign n77176 = pi16 ? n2749 : ~n2964;
  assign n77177 = pi16 ? n2415 : ~n2964;
  assign n77178 = pi15 ? n77176 : n77177;
  assign n77179 = pi16 ? n2120 : ~n2964;
  assign n77180 = pi15 ? n77177 : n77179;
  assign n77181 = pi14 ? n77178 : n77180;
  assign n77182 = pi13 ? n77181 : n77068;
  assign n77183 = pi12 ? n77175 : n77182;
  assign n77184 = pi15 ? n77069 : n76957;
  assign n77185 = pi14 ? n77184 : n76959;
  assign n77186 = pi16 ? n1683 : ~n3061;
  assign n77187 = pi15 ? n77186 : n76911;
  assign n77188 = pi14 ? n77186 : n77187;
  assign n77189 = pi13 ? n77185 : n77188;
  assign n77190 = pi16 ? n1581 : ~n3061;
  assign n77191 = pi15 ? n77190 : n77134;
  assign n77192 = pi14 ? n77190 : n77191;
  assign n77193 = pi15 ? n76731 : n76661;
  assign n77194 = pi15 ? n76662 : n76735;
  assign n77195 = pi14 ? n77193 : n77194;
  assign n77196 = pi13 ? n77192 : n77195;
  assign n77197 = pi12 ? n77189 : n77196;
  assign n77198 = pi11 ? n77183 : n77197;
  assign n77199 = pi16 ? n1214 : ~n2840;
  assign n77200 = pi15 ? n77199 : n76584;
  assign n77201 = pi14 ? n76736 : n77200;
  assign n77202 = pi15 ? n76585 : n76520;
  assign n77203 = pi14 ? n77202 : n76488;
  assign n77204 = pi13 ? n77201 : n77203;
  assign n77205 = pi14 ? n76429 : n76433;
  assign n77206 = pi14 ? n76375 : n76322;
  assign n77207 = pi13 ? n77205 : n77206;
  assign n77208 = pi12 ? n77204 : n77207;
  assign n77209 = pi13 ? n76271 : n76094;
  assign n77210 = pi14 ? n75990 : n75940;
  assign n77211 = pi13 ? n77210 : n61508;
  assign n77212 = pi12 ? n77209 : n77211;
  assign n77213 = pi11 ? n77208 : n77212;
  assign n77214 = pi10 ? n77198 : n77213;
  assign n77215 = pi09 ? n77162 : n77214;
  assign n77216 = pi08 ? n77154 : n77215;
  assign n77217 = pi07 ? n77096 : n77216;
  assign n77218 = pi16 ? n3156 : ~n2958;
  assign n77219 = pi15 ? n32 : n77218;
  assign n77220 = pi16 ? n3161 : ~n2958;
  assign n77221 = pi16 ? n3165 : ~n2958;
  assign n77222 = pi15 ? n77220 : n77221;
  assign n77223 = pi14 ? n77219 : n77222;
  assign n77224 = pi13 ? n32 : n77223;
  assign n77225 = pi12 ? n32 : n77224;
  assign n77226 = pi11 ? n32 : n77225;
  assign n77227 = pi10 ? n32 : n77226;
  assign n77228 = pi16 ? n2953 : ~n2958;
  assign n77229 = pi16 ? n3176 : ~n2958;
  assign n77230 = pi15 ? n77228 : n77229;
  assign n77231 = pi16 ? n2964 : ~n2958;
  assign n77232 = pi16 ? n3183 : ~n2964;
  assign n77233 = pi15 ? n77231 : n77232;
  assign n77234 = pi14 ? n77230 : n77233;
  assign n77235 = pi15 ? n77232 : n77109;
  assign n77236 = pi14 ? n77235 : n77109;
  assign n77237 = pi13 ? n77234 : n77236;
  assign n77238 = pi16 ? n2617 : ~n2964;
  assign n77239 = pi16 ? n2518 : ~n2964;
  assign n77240 = pi15 ? n77238 : n77239;
  assign n77241 = pi16 ? n2756 : ~n2964;
  assign n77242 = pi14 ? n77240 : n77241;
  assign n77243 = pi16 ? n2409 : ~n2964;
  assign n77244 = pi15 ? n77243 : n77177;
  assign n77245 = pi16 ? n2306 : ~n2964;
  assign n77246 = pi16 ? n1934 : ~n2964;
  assign n77247 = pi15 ? n77245 : n77246;
  assign n77248 = pi14 ? n77244 : n77247;
  assign n77249 = pi13 ? n77242 : n77248;
  assign n77250 = pi12 ? n77237 : n77249;
  assign n77251 = pi16 ? n1808 : ~n3183;
  assign n77252 = pi15 ? n77123 : n77251;
  assign n77253 = pi14 ? n77123 : n77252;
  assign n77254 = pi15 ? n76953 : n76957;
  assign n77255 = pi14 ? n76953 : n77254;
  assign n77256 = pi13 ? n77253 : n77255;
  assign n77257 = pi16 ? n1678 : ~n2832;
  assign n77258 = pi16 ? n1678 : ~n3061;
  assign n77259 = pi15 ? n77258 : n77186;
  assign n77260 = pi14 ? n77257 : n77259;
  assign n77261 = pi15 ? n76816 : n76694;
  assign n77262 = pi15 ? n76694 : n76772;
  assign n77263 = pi14 ? n77261 : n77262;
  assign n77264 = pi13 ? n77260 : n77263;
  assign n77265 = pi12 ? n77256 : n77264;
  assign n77266 = pi11 ? n77250 : n77265;
  assign n77267 = pi16 ? n1581 : ~n2840;
  assign n77268 = pi16 ? n1843 : ~n2840;
  assign n77269 = pi15 ? n77268 : n76576;
  assign n77270 = pi14 ? n77267 : n77269;
  assign n77271 = pi16 ? n1705 : ~n4246;
  assign n77272 = pi16 ? n1705 : ~n2725;
  assign n77273 = pi15 ? n77271 : n77272;
  assign n77274 = pi14 ? n76577 : n77273;
  assign n77275 = pi13 ? n77270 : n77274;
  assign n77276 = pi16 ? n1972 : ~n2725;
  assign n77277 = pi16 ? n1214 : ~n2725;
  assign n77278 = pi14 ? n77276 : n77277;
  assign n77279 = pi13 ? n77278 : n76467;
  assign n77280 = pi12 ? n77275 : n77279;
  assign n77281 = pi14 ? n76146 : n76091;
  assign n77282 = pi13 ? n76271 : n77281;
  assign n77283 = pi15 ? n62214 : n61868;
  assign n77284 = pi14 ? n76039 : n77283;
  assign n77285 = pi15 ? n61868 : n61629;
  assign n77286 = pi15 ? n61329 : n75739;
  assign n77287 = pi14 ? n77285 : n77286;
  assign n77288 = pi13 ? n77284 : n77287;
  assign n77289 = pi12 ? n77282 : n77288;
  assign n77290 = pi11 ? n77280 : n77289;
  assign n77291 = pi10 ? n77266 : n77290;
  assign n77292 = pi09 ? n77227 : n77291;
  assign n77293 = pi16 ? n32 : ~n2958;
  assign n77294 = pi15 ? n32 : n77293;
  assign n77295 = pi16 ? n3283 : ~n2958;
  assign n77296 = pi15 ? n77295 : n77221;
  assign n77297 = pi14 ? n77294 : n77296;
  assign n77298 = pi13 ? n32 : n77297;
  assign n77299 = pi12 ? n32 : n77298;
  assign n77300 = pi11 ? n32 : n77299;
  assign n77301 = pi10 ? n32 : n77300;
  assign n77302 = pi16 ? n3047 : ~n2958;
  assign n77303 = pi16 ? n3293 : ~n2958;
  assign n77304 = pi15 ? n77302 : n77303;
  assign n77305 = pi14 ? n77304 : n77228;
  assign n77306 = pi16 ? n2837 : ~n2958;
  assign n77307 = pi15 ? n77229 : n77306;
  assign n77308 = pi16 ? n2840 : ~n2958;
  assign n77309 = pi16 ? n2851 : ~n2958;
  assign n77310 = pi15 ? n77308 : n77309;
  assign n77311 = pi14 ? n77307 : n77310;
  assign n77312 = pi13 ? n77305 : n77311;
  assign n77313 = pi16 ? n3068 : ~n2958;
  assign n77314 = pi16 ? n2624 : ~n2958;
  assign n77315 = pi15 ? n77313 : n77314;
  assign n77316 = pi16 ? n2860 : ~n2958;
  assign n77317 = pi15 ? n77316 : n77172;
  assign n77318 = pi14 ? n77315 : n77317;
  assign n77319 = pi13 ? n77318 : n77181;
  assign n77320 = pi12 ? n77312 : n77319;
  assign n77321 = pi16 ? n2426 : ~n2964;
  assign n77322 = pi15 ? n77321 : n77062;
  assign n77323 = pi16 ? n2530 : ~n3183;
  assign n77324 = pi15 ? n77323 : n77119;
  assign n77325 = pi14 ? n77322 : n77324;
  assign n77326 = pi16 ? n3338 : ~n2832;
  assign n77327 = pi15 ? n77006 : n77326;
  assign n77328 = pi14 ? n77006 : n77327;
  assign n77329 = pi13 ? n77325 : n77328;
  assign n77330 = pi16 ? n1808 : ~n2832;
  assign n77331 = pi15 ? n77330 : n76953;
  assign n77332 = pi14 ? n77330 : n77331;
  assign n77333 = pi16 ? n3352 : ~n3061;
  assign n77334 = pi16 ? n3352 : ~n2837;
  assign n77335 = pi15 ? n77333 : n77334;
  assign n77336 = pi16 ? n3356 : ~n2837;
  assign n77337 = pi15 ? n77334 : n77336;
  assign n77338 = pi14 ? n77335 : n77337;
  assign n77339 = pi13 ? n77332 : n77338;
  assign n77340 = pi12 ? n77329 : n77339;
  assign n77341 = pi11 ? n77320 : n77340;
  assign n77342 = pi16 ? n1577 : ~n2840;
  assign n77343 = pi15 ? n76653 : n77342;
  assign n77344 = pi14 ? n76728 : n77343;
  assign n77345 = pi16 ? n1834 : ~n2851;
  assign n77346 = pi15 ? n76694 : n77345;
  assign n77347 = pi16 ? n1323 : ~n4246;
  assign n77348 = pi15 ? n76541 : n77347;
  assign n77349 = pi14 ? n77346 : n77348;
  assign n77350 = pi13 ? n77344 : n77349;
  assign n77351 = pi16 ? n1594 : ~n4246;
  assign n77352 = pi16 ? n1843 : ~n4246;
  assign n77353 = pi16 ? n1843 : ~n2725;
  assign n77354 = pi15 ? n77352 : n77353;
  assign n77355 = pi14 ? n77351 : n77354;
  assign n77356 = pi16 ? n1471 : ~n2725;
  assign n77357 = pi16 ? n1479 : ~n2732;
  assign n77358 = pi16 ? n1479 : ~n2745;
  assign n77359 = pi15 ? n77357 : n77358;
  assign n77360 = pi14 ? n77356 : n77359;
  assign n77361 = pi13 ? n77355 : n77360;
  assign n77362 = pi12 ? n77350 : n77361;
  assign n77363 = pi15 ? n76232 : n76239;
  assign n77364 = pi15 ? n76183 : n76123;
  assign n77365 = pi14 ? n77363 : n77364;
  assign n77366 = pi16 ? n1705 : ~n2624;
  assign n77367 = pi16 ? n1705 : ~n2860;
  assign n77368 = pi15 ? n77366 : n77367;
  assign n77369 = pi14 ? n76116 : n77368;
  assign n77370 = pi13 ? n77365 : n77369;
  assign n77371 = pi16 ? n1705 : ~n4100;
  assign n77372 = pi16 ? n1705 : ~n3946;
  assign n77373 = pi15 ? n77371 : n77372;
  assign n77374 = pi16 ? n1972 : ~n3946;
  assign n77375 = pi16 ? n1479 : ~n2629;
  assign n77376 = pi15 ? n77374 : n77375;
  assign n77377 = pi14 ? n77373 : n77376;
  assign n77378 = pi16 ? n1479 : ~n2513;
  assign n77379 = pi16 ? n1594 : ~n2749;
  assign n77380 = pi15 ? n77378 : n77379;
  assign n77381 = pi14 ? n77380 : n77379;
  assign n77382 = pi13 ? n77377 : n77381;
  assign n77383 = pi12 ? n77370 : n77382;
  assign n77384 = pi11 ? n77362 : n77383;
  assign n77385 = pi10 ? n77341 : n77384;
  assign n77386 = pi09 ? n77301 : n77385;
  assign n77387 = pi08 ? n77292 : n77386;
  assign n77388 = pi17 ? n2005 : ~n3175;
  assign n77389 = pi16 ? n32 : n77388;
  assign n77390 = pi15 ? n32 : n77389;
  assign n77391 = pi17 ? n1028 : ~n3175;
  assign n77392 = pi16 ? n32 : n77391;
  assign n77393 = pi16 ? n3283 : ~n3176;
  assign n77394 = pi15 ? n77392 : n77393;
  assign n77395 = pi14 ? n77390 : n77394;
  assign n77396 = pi13 ? n32 : n77395;
  assign n77397 = pi12 ? n32 : n77396;
  assign n77398 = pi11 ? n32 : n77397;
  assign n77399 = pi10 ? n32 : n77398;
  assign n77400 = pi16 ? n3156 : ~n3176;
  assign n77401 = pi16 ? n3438 : ~n3176;
  assign n77402 = pi15 ? n77400 : n77401;
  assign n77403 = pi16 ? n3165 : ~n3176;
  assign n77404 = pi15 ? n77403 : n77302;
  assign n77405 = pi14 ? n77402 : n77404;
  assign n77406 = pi16 ? n2958 : ~n2958;
  assign n77407 = pi15 ? n77229 : n77406;
  assign n77408 = pi16 ? n3183 : ~n2958;
  assign n77409 = pi15 ? n77231 : n77408;
  assign n77410 = pi14 ? n77407 : n77409;
  assign n77411 = pi13 ? n77405 : n77410;
  assign n77412 = pi16 ? n2745 : ~n2958;
  assign n77413 = pi15 ? n77408 : n77412;
  assign n77414 = pi15 ? n77412 : n77109;
  assign n77415 = pi14 ? n77413 : n77414;
  assign n77416 = pi16 ? n2518 : ~n2958;
  assign n77417 = pi15 ? n77238 : n77416;
  assign n77418 = pi16 ? n2756 : ~n2958;
  assign n77419 = pi15 ? n77241 : n77418;
  assign n77420 = pi14 ? n77417 : n77419;
  assign n77421 = pi13 ? n77415 : n77420;
  assign n77422 = pi12 ? n77411 : n77421;
  assign n77423 = pi14 ? n77243 : n77244;
  assign n77424 = pi16 ? n2300 : ~n3183;
  assign n77425 = pi15 ? n77424 : n77323;
  assign n77426 = pi14 ? n77058 : n77425;
  assign n77427 = pi13 ? n77423 : n77426;
  assign n77428 = pi15 ? n77005 : n76952;
  assign n77429 = pi14 ? n77119 : n77428;
  assign n77430 = pi16 ? n2540 : ~n2837;
  assign n77431 = pi15 ? n76905 : n77430;
  assign n77432 = pi16 ? n3338 : ~n2837;
  assign n77433 = pi15 ? n77430 : n77432;
  assign n77434 = pi14 ? n77431 : n77433;
  assign n77435 = pi13 ? n77429 : n77434;
  assign n77436 = pi12 ? n77427 : n77435;
  assign n77437 = pi11 ? n77422 : n77436;
  assign n77438 = pi16 ? n2326 : ~n2840;
  assign n77439 = pi15 ? n76721 : n77438;
  assign n77440 = pi14 ? n76721 : n77439;
  assign n77441 = pi16 ? n3356 : ~n2840;
  assign n77442 = pi16 ? n3356 : ~n3068;
  assign n77443 = pi16 ? n3356 : ~n4246;
  assign n77444 = pi15 ? n77442 : n77443;
  assign n77445 = pi14 ? n77441 : n77444;
  assign n77446 = pi13 ? n77440 : n77445;
  assign n77447 = pi16 ? n1678 : ~n4246;
  assign n77448 = pi16 ? n1834 : ~n4246;
  assign n77449 = pi14 ? n77447 : n77448;
  assign n77450 = pi16 ? n2144 : ~n2725;
  assign n77451 = pi16 ? n1581 : ~n2732;
  assign n77452 = pi14 ? n77450 : n77451;
  assign n77453 = pi13 ? n77449 : n77452;
  assign n77454 = pi12 ? n77446 : n77453;
  assign n77455 = pi16 ? n1323 : ~n2617;
  assign n77456 = pi16 ? n1479 : ~n2617;
  assign n77457 = pi15 ? n77455 : n77456;
  assign n77458 = pi16 ? n1479 : ~n2856;
  assign n77459 = pi14 ? n77457 : n77458;
  assign n77460 = pi16 ? n1323 : ~n2856;
  assign n77461 = pi16 ? n1323 : ~n2624;
  assign n77462 = pi15 ? n77460 : n77461;
  assign n77463 = pi16 ? n1323 : ~n2860;
  assign n77464 = pi15 ? n77461 : n77463;
  assign n77465 = pi14 ? n77462 : n77464;
  assign n77466 = pi13 ? n77459 : n77465;
  assign n77467 = pi16 ? n1323 : ~n4100;
  assign n77468 = pi16 ? n1594 : ~n3946;
  assign n77469 = pi16 ? n1577 : ~n2629;
  assign n77470 = pi15 ? n77468 : n77469;
  assign n77471 = pi14 ? n77467 : n77470;
  assign n77472 = pi16 ? n1577 : ~n2513;
  assign n77473 = pi15 ? n77469 : n77472;
  assign n77474 = pi16 ? n1577 : ~n2749;
  assign n77475 = pi14 ? n77473 : n77474;
  assign n77476 = pi13 ? n77471 : n77475;
  assign n77477 = pi12 ? n77466 : n77476;
  assign n77478 = pi11 ? n77454 : n77477;
  assign n77479 = pi10 ? n77437 : n77478;
  assign n77480 = pi09 ? n77399 : n77479;
  assign n77481 = pi17 ? n3553 : ~n3175;
  assign n77482 = pi16 ? n32 : n77481;
  assign n77483 = pi15 ? n32 : n77482;
  assign n77484 = pi17 ? n3557 : ~n3175;
  assign n77485 = pi16 ? n32 : n77484;
  assign n77486 = pi15 ? n77392 : n77485;
  assign n77487 = pi14 ? n77483 : n77486;
  assign n77488 = pi13 ? n32 : n77487;
  assign n77489 = pi12 ? n32 : n77488;
  assign n77490 = pi11 ? n32 : n77489;
  assign n77491 = pi10 ? n32 : n77490;
  assign n77492 = pi16 ? n32 : ~n3176;
  assign n77493 = pi16 ? n3570 : ~n3176;
  assign n77494 = pi15 ? n77492 : n77493;
  assign n77495 = pi16 ? n3047 : ~n3176;
  assign n77496 = pi15 ? n77400 : n77495;
  assign n77497 = pi14 ? n77494 : n77496;
  assign n77498 = pi16 ? n3588 : ~n3176;
  assign n77499 = pi15 ? n77303 : n77498;
  assign n77500 = pi16 ? n2953 : ~n3176;
  assign n77501 = pi14 ? n77499 : n77500;
  assign n77502 = pi13 ? n77497 : n77501;
  assign n77503 = pi16 ? n3176 : ~n3176;
  assign n77504 = pi16 ? n2837 : ~n3176;
  assign n77505 = pi15 ? n77503 : n77504;
  assign n77506 = pi16 ? n2840 : ~n3176;
  assign n77507 = pi15 ? n77506 : n77309;
  assign n77508 = pi14 ? n77505 : n77507;
  assign n77509 = pi16 ? n2513 : ~n2958;
  assign n77510 = pi15 ? n77316 : n77509;
  assign n77511 = pi14 ? n77315 : n77510;
  assign n77512 = pi13 ? n77508 : n77511;
  assign n77513 = pi12 ? n77502 : n77512;
  assign n77514 = pi16 ? n2749 : ~n2958;
  assign n77515 = pi15 ? n77514 : n77176;
  assign n77516 = pi14 ? n77515 : n77239;
  assign n77517 = pi16 ? n2293 : ~n3183;
  assign n77518 = pi15 ? n77517 : n77117;
  assign n77519 = pi14 ? n77517 : n77518;
  assign n77520 = pi13 ? n77516 : n77519;
  assign n77521 = pi16 ? n3625 : ~n3183;
  assign n77522 = pi15 ? n77521 : n77424;
  assign n77523 = pi14 ? n77056 : n77522;
  assign n77524 = pi15 ? n76801 : n76809;
  assign n77525 = pi14 ? n76801 : n77524;
  assign n77526 = pi13 ? n77523 : n77525;
  assign n77527 = pi12 ? n77520 : n77526;
  assign n77528 = pi11 ? n77513 : n77527;
  assign n77529 = pi16 ? n2320 : ~n2837;
  assign n77530 = pi15 ? n76718 : n77529;
  assign n77531 = pi14 ? n76809 : n77530;
  assign n77532 = pi15 ? n76720 : n76687;
  assign n77533 = pi16 ? n1815 : ~n2851;
  assign n77534 = pi16 ? n1815 : ~n3068;
  assign n77535 = pi15 ? n77533 : n77534;
  assign n77536 = pi14 ? n77532 : n77535;
  assign n77537 = pi13 ? n77531 : n77536;
  assign n77538 = pi16 ? n1944 : ~n3068;
  assign n77539 = pi16 ? n1944 : ~n4246;
  assign n77540 = pi14 ? n77538 : n77539;
  assign n77541 = pi16 ? n2326 : ~n4246;
  assign n77542 = pi15 ? n77447 : n77541;
  assign n77543 = pi16 ? n1678 : ~n2725;
  assign n77544 = pi16 ? n1678 : ~n2732;
  assign n77545 = pi15 ? n77543 : n77544;
  assign n77546 = pi14 ? n77542 : n77545;
  assign n77547 = pi13 ? n77540 : n77546;
  assign n77548 = pi12 ? n77537 : n77547;
  assign n77549 = pi16 ? n1683 : ~n2745;
  assign n77550 = pi16 ? n1577 : ~n2745;
  assign n77551 = pi15 ? n77549 : n77550;
  assign n77552 = pi16 ? n1577 : ~n2856;
  assign n77553 = pi14 ? n77551 : n77552;
  assign n77554 = pi16 ? n1683 : ~n2856;
  assign n77555 = pi16 ? n3352 : ~n2856;
  assign n77556 = pi16 ? n3352 : ~n2624;
  assign n77557 = pi15 ? n77555 : n77556;
  assign n77558 = pi14 ? n77554 : n77557;
  assign n77559 = pi13 ? n77553 : n77558;
  assign n77560 = pi16 ? n3352 : ~n2860;
  assign n77561 = pi16 ? n3352 : ~n4100;
  assign n77562 = pi15 ? n77560 : n77561;
  assign n77563 = pi16 ? n3356 : ~n4100;
  assign n77564 = pi15 ? n77563 : n61951;
  assign n77565 = pi14 ? n77562 : n77564;
  assign n77566 = pi16 ? n2326 : ~n2629;
  assign n77567 = pi16 ? n1815 : ~n2513;
  assign n77568 = pi15 ? n77566 : n77567;
  assign n77569 = pi16 ? n2137 : ~n2513;
  assign n77570 = pi16 ? n2137 : ~n2749;
  assign n77571 = pi15 ? n77569 : n77570;
  assign n77572 = pi14 ? n77568 : n77571;
  assign n77573 = pi13 ? n77565 : n77572;
  assign n77574 = pi12 ? n77559 : n77573;
  assign n77575 = pi11 ? n77548 : n77574;
  assign n77576 = pi10 ? n77528 : n77575;
  assign n77577 = pi09 ? n77491 : n77576;
  assign n77578 = pi08 ? n77480 : n77577;
  assign n77579 = pi07 ? n77387 : n77578;
  assign n77580 = pi06 ? n77217 : n77579;
  assign n77581 = pi05 ? n76988 : n77580;
  assign n77582 = pi17 ? n1219 : ~n2952;
  assign n77583 = pi16 ? n32 : n77582;
  assign n77584 = pi15 ? n32 : n77583;
  assign n77585 = pi17 ? n1726 : ~n2952;
  assign n77586 = pi16 ? n32 : n77585;
  assign n77587 = pi17 ? n3704 : ~n2952;
  assign n77588 = pi16 ? n32 : n77587;
  assign n77589 = pi15 ? n77586 : n77588;
  assign n77590 = pi14 ? n77584 : n77589;
  assign n77591 = pi13 ? n32 : n77590;
  assign n77592 = pi12 ? n32 : n77591;
  assign n77593 = pi11 ? n32 : n77592;
  assign n77594 = pi10 ? n32 : n77593;
  assign n77595 = pi17 ? n2005 : ~n2952;
  assign n77596 = pi16 ? n32 : n77595;
  assign n77597 = pi17 ? n3715 : ~n2952;
  assign n77598 = pi16 ? n32 : n77597;
  assign n77599 = pi15 ? n77596 : n77598;
  assign n77600 = pi17 ? n3719 : ~n3175;
  assign n77601 = pi16 ? n32 : n77600;
  assign n77602 = pi15 ? n77601 : n77400;
  assign n77603 = pi14 ? n77599 : n77602;
  assign n77604 = pi16 ? n3729 : ~n3176;
  assign n77605 = pi15 ? n77401 : n77604;
  assign n77606 = pi15 ? n77403 : n77495;
  assign n77607 = pi14 ? n77605 : n77606;
  assign n77608 = pi13 ? n77603 : n77607;
  assign n77609 = pi16 ? n2958 : ~n3176;
  assign n77610 = pi15 ? n77503 : n77609;
  assign n77611 = pi16 ? n2964 : ~n3176;
  assign n77612 = pi15 ? n77611 : n77408;
  assign n77613 = pi14 ? n77610 : n77612;
  assign n77614 = pi16 ? n2745 : ~n3176;
  assign n77615 = pi15 ? n77408 : n77614;
  assign n77616 = pi15 ? n77412 : n77614;
  assign n77617 = pi14 ? n77615 : n77616;
  assign n77618 = pi13 ? n77613 : n77617;
  assign n77619 = pi12 ? n77608 : n77618;
  assign n77620 = pi16 ? n2617 : ~n2958;
  assign n77621 = pi16 ? n2856 : ~n2958;
  assign n77622 = pi15 ? n77620 : n77621;
  assign n77623 = pi16 ? n2629 : ~n2958;
  assign n77624 = pi15 ? n77314 : n77623;
  assign n77625 = pi14 ? n77622 : n77624;
  assign n77626 = pi14 ? n77172 : n77176;
  assign n77627 = pi13 ? n77625 : n77626;
  assign n77628 = pi16 ? n3769 : ~n2964;
  assign n77629 = pi16 ? n3769 : ~n3183;
  assign n77630 = pi15 ? n77629 : n77517;
  assign n77631 = pi14 ? n77628 : n77630;
  assign n77632 = pi16 ? n2654 : ~n3061;
  assign n77633 = pi16 ? n3788 : ~n3061;
  assign n77634 = pi15 ? n77632 : n77633;
  assign n77635 = pi14 ? n76799 : n77634;
  assign n77636 = pi13 ? n77631 : n77635;
  assign n77637 = pi12 ? n77627 : n77636;
  assign n77638 = pi11 ? n77619 : n77637;
  assign n77639 = pi16 ? n2530 : ~n2837;
  assign n77640 = pi15 ? n77633 : n77639;
  assign n77641 = pi14 ? n77633 : n77640;
  assign n77642 = pi16 ? n2530 : ~n2840;
  assign n77643 = pi15 ? n77639 : n77642;
  assign n77644 = pi16 ? n2530 : ~n2851;
  assign n77645 = pi16 ? n2530 : ~n3068;
  assign n77646 = pi15 ? n77644 : n77645;
  assign n77647 = pi14 ? n77643 : n77646;
  assign n77648 = pi13 ? n77641 : n77647;
  assign n77649 = pi16 ? n2540 : ~n3068;
  assign n77650 = pi16 ? n1808 : ~n4246;
  assign n77651 = pi16 ? n1808 : ~n2732;
  assign n77652 = pi14 ? n77650 : n77651;
  assign n77653 = pi13 ? n77649 : n77652;
  assign n77654 = pi12 ? n77648 : n77653;
  assign n77655 = pi16 ? n2326 : ~n2745;
  assign n77656 = pi16 ? n2326 : ~n2617;
  assign n77657 = pi14 ? n77655 : n77656;
  assign n77658 = pi16 ? n1815 : ~n2617;
  assign n77659 = pi16 ? n1815 : ~n2856;
  assign n77660 = pi15 ? n77658 : n77659;
  assign n77661 = pi15 ? n63211 : n62810;
  assign n77662 = pi14 ? n77660 : n77661;
  assign n77663 = pi13 ? n77657 : n77662;
  assign n77664 = pi16 ? n1815 : ~n4100;
  assign n77665 = pi16 ? n2320 : ~n3946;
  assign n77666 = pi15 ? n77664 : n77665;
  assign n77667 = pi14 ? n62811 : n77666;
  assign n77668 = pi15 ? n77665 : n65897;
  assign n77669 = pi16 ? n2320 : ~n2513;
  assign n77670 = pi16 ? n2320 : ~n2749;
  assign n77671 = pi15 ? n77669 : n77670;
  assign n77672 = pi14 ? n77668 : n77671;
  assign n77673 = pi13 ? n77667 : n77672;
  assign n77674 = pi12 ? n77663 : n77673;
  assign n77675 = pi11 ? n77654 : n77674;
  assign n77676 = pi10 ? n77638 : n77675;
  assign n77677 = pi09 ? n77594 : n77676;
  assign n77678 = pi17 ? n4037 : ~n2952;
  assign n77679 = pi16 ? n32 : n77678;
  assign n77680 = pi15 ? n32 : n77679;
  assign n77681 = pi17 ? n3855 : ~n2952;
  assign n77682 = pi16 ? n32 : n77681;
  assign n77683 = pi17 ? n1227 : ~n2952;
  assign n77684 = pi16 ? n32 : n77683;
  assign n77685 = pi15 ? n77682 : n77684;
  assign n77686 = pi14 ? n77680 : n77685;
  assign n77687 = pi13 ? n32 : n77686;
  assign n77688 = pi12 ? n32 : n77687;
  assign n77689 = pi11 ? n32 : n77688;
  assign n77690 = pi10 ? n32 : n77689;
  assign n77691 = pi17 ? n3553 : ~n2952;
  assign n77692 = pi16 ? n32 : n77691;
  assign n77693 = pi15 ? n77692 : n77586;
  assign n77694 = pi16 ? n32 : ~n2953;
  assign n77695 = pi15 ? n77601 : n77694;
  assign n77696 = pi14 ? n77693 : n77695;
  assign n77697 = pi16 ? n3283 : ~n2953;
  assign n77698 = pi15 ? n77493 : n77697;
  assign n77699 = pi16 ? n3156 : ~n2953;
  assign n77700 = pi16 ? n3047 : ~n2953;
  assign n77701 = pi15 ? n77699 : n77700;
  assign n77702 = pi14 ? n77698 : n77701;
  assign n77703 = pi13 ? n77696 : n77702;
  assign n77704 = pi16 ? n3293 : ~n2953;
  assign n77705 = pi16 ? n3588 : ~n2953;
  assign n77706 = pi15 ? n77704 : n77705;
  assign n77707 = pi16 ? n2953 : ~n2953;
  assign n77708 = pi15 ? n77707 : n77500;
  assign n77709 = pi14 ? n77706 : n77708;
  assign n77710 = pi16 ? n2851 : ~n3176;
  assign n77711 = pi15 ? n77506 : n77710;
  assign n77712 = pi14 ? n77505 : n77711;
  assign n77713 = pi13 ? n77709 : n77712;
  assign n77714 = pi12 ? n77703 : n77713;
  assign n77715 = pi16 ? n3068 : ~n3176;
  assign n77716 = pi16 ? n2732 : ~n2958;
  assign n77717 = pi15 ? n77715 : n77716;
  assign n77718 = pi14 ? n77717 : n77716;
  assign n77719 = pi15 ? n77109 : n77238;
  assign n77720 = pi16 ? n2856 : ~n2964;
  assign n77721 = pi16 ? n3946 : ~n2964;
  assign n77722 = pi15 ? n77720 : n77721;
  assign n77723 = pi14 ? n77719 : n77722;
  assign n77724 = pi13 ? n77718 : n77723;
  assign n77725 = pi16 ? n2629 : ~n2964;
  assign n77726 = pi14 ? n77725 : n77172;
  assign n77727 = pi15 ? n77113 : n76893;
  assign n77728 = pi15 ? n76893 : n77001;
  assign n77729 = pi14 ? n77727 : n77728;
  assign n77730 = pi13 ? n77726 : n77729;
  assign n77731 = pi12 ? n77724 : n77730;
  assign n77732 = pi11 ? n77714 : n77731;
  assign n77733 = pi16 ? n2756 : ~n3061;
  assign n77734 = pi15 ? n77001 : n77733;
  assign n77735 = pi14 ? n77734 : n76854;
  assign n77736 = pi16 ? n2426 : ~n2840;
  assign n77737 = pi15 ? n76853 : n77736;
  assign n77738 = pi16 ? n3788 : ~n2851;
  assign n77739 = pi15 ? n77736 : n77738;
  assign n77740 = pi14 ? n77737 : n77739;
  assign n77741 = pi13 ? n77735 : n77740;
  assign n77742 = pi16 ? n3788 : ~n3068;
  assign n77743 = pi15 ? n77738 : n77742;
  assign n77744 = pi14 ? n77743 : n77742;
  assign n77745 = pi16 ? n2306 : ~n3068;
  assign n77746 = pi16 ? n2306 : ~n2725;
  assign n77747 = pi14 ? n77745 : n77746;
  assign n77748 = pi13 ? n77744 : n77747;
  assign n77749 = pi12 ? n77741 : n77748;
  assign n77750 = pi16 ? n2320 : ~n2732;
  assign n77751 = pi16 ? n2320 : ~n2617;
  assign n77752 = pi14 ? n77750 : n77751;
  assign n77753 = pi16 ? n1934 : ~n2617;
  assign n77754 = pi16 ? n2300 : ~n2856;
  assign n77755 = pi16 ? n2300 : ~n2624;
  assign n77756 = pi15 ? n77754 : n77755;
  assign n77757 = pi14 ? n77753 : n77756;
  assign n77758 = pi13 ? n77752 : n77757;
  assign n77759 = pi16 ? n2300 : ~n2860;
  assign n77760 = pi15 ? n77755 : n77759;
  assign n77761 = pi16 ? n2530 : ~n4100;
  assign n77762 = pi16 ? n3625 : ~n3946;
  assign n77763 = pi15 ? n77761 : n77762;
  assign n77764 = pi14 ? n77760 : n77763;
  assign n77765 = pi15 ? n77762 : n66060;
  assign n77766 = pi16 ? n3625 : ~n2513;
  assign n77767 = pi16 ? n2654 : ~n2749;
  assign n77768 = pi15 ? n77766 : n77767;
  assign n77769 = pi14 ? n77765 : n77768;
  assign n77770 = pi13 ? n77764 : n77769;
  assign n77771 = pi12 ? n77758 : n77770;
  assign n77772 = pi11 ? n77749 : n77771;
  assign n77773 = pi10 ? n77732 : n77772;
  assign n77774 = pi09 ? n77690 : n77773;
  assign n77775 = pi08 ? n77677 : n77774;
  assign n77776 = pi17 ? n2355 : ~n3050;
  assign n77777 = pi16 ? n32 : n77776;
  assign n77778 = pi15 ? n32 : n77777;
  assign n77779 = pi17 ? n4023 : ~n3050;
  assign n77780 = pi16 ? n32 : n77779;
  assign n77781 = pi17 ? n1120 : ~n3050;
  assign n77782 = pi16 ? n32 : n77781;
  assign n77783 = pi15 ? n77780 : n77782;
  assign n77784 = pi14 ? n77778 : n77783;
  assign n77785 = pi13 ? n32 : n77784;
  assign n77786 = pi12 ? n32 : n77785;
  assign n77787 = pi11 ? n32 : n77786;
  assign n77788 = pi10 ? n32 : n77787;
  assign n77789 = pi17 ? n4034 : ~n3050;
  assign n77790 = pi16 ? n32 : n77789;
  assign n77791 = pi17 ? n4037 : ~n3050;
  assign n77792 = pi16 ? n32 : n77791;
  assign n77793 = pi15 ? n77790 : n77792;
  assign n77794 = pi17 ? n4041 : ~n2952;
  assign n77795 = pi16 ? n32 : n77794;
  assign n77796 = pi15 ? n77795 : n77596;
  assign n77797 = pi14 ? n77793 : n77796;
  assign n77798 = pi17 ? n1028 : ~n2952;
  assign n77799 = pi16 ? n32 : n77798;
  assign n77800 = pi15 ? n77598 : n77799;
  assign n77801 = pi17 ? n3719 : ~n2952;
  assign n77802 = pi16 ? n32 : n77801;
  assign n77803 = pi15 ? n77802 : n77699;
  assign n77804 = pi14 ? n77800 : n77803;
  assign n77805 = pi13 ? n77797 : n77804;
  assign n77806 = pi16 ? n3438 : ~n2953;
  assign n77807 = pi16 ? n3729 : ~n2953;
  assign n77808 = pi15 ? n77806 : n77807;
  assign n77809 = pi16 ? n3165 : ~n2953;
  assign n77810 = pi15 ? n77809 : n77495;
  assign n77811 = pi14 ? n77808 : n77810;
  assign n77812 = pi16 ? n3183 : ~n2953;
  assign n77813 = pi15 ? n77611 : n77812;
  assign n77814 = pi14 ? n77610 : n77813;
  assign n77815 = pi13 ? n77811 : n77814;
  assign n77816 = pi12 ? n77805 : n77815;
  assign n77817 = pi16 ? n3061 : ~n3176;
  assign n77818 = pi15 ? n77812 : n77817;
  assign n77819 = pi15 ? n77817 : n77306;
  assign n77820 = pi14 ? n77818 : n77819;
  assign n77821 = pi16 ? n2725 : ~n2958;
  assign n77822 = pi14 ? n77310 : n77821;
  assign n77823 = pi13 ? n77820 : n77822;
  assign n77824 = pi15 ? n77716 : n77412;
  assign n77825 = pi16 ? n4100 : ~n2964;
  assign n77826 = pi15 ? n77238 : n77825;
  assign n77827 = pi14 ? n77824 : n77826;
  assign n77828 = pi16 ? n4100 : ~n3183;
  assign n77829 = pi16 ? n4100 : ~n2832;
  assign n77830 = pi15 ? n77828 : n77829;
  assign n77831 = pi16 ? n3946 : ~n2832;
  assign n77832 = pi14 ? n77830 : n77831;
  assign n77833 = pi13 ? n77827 : n77832;
  assign n77834 = pi12 ? n77823 : n77833;
  assign n77835 = pi11 ? n77816 : n77834;
  assign n77836 = pi16 ? n2749 : ~n3061;
  assign n77837 = pi15 ? n76891 : n77836;
  assign n77838 = pi14 ? n76891 : n77837;
  assign n77839 = pi16 ? n2749 : ~n2840;
  assign n77840 = pi15 ? n77836 : n77839;
  assign n77841 = pi16 ? n2409 : ~n2840;
  assign n77842 = pi16 ? n2409 : ~n2851;
  assign n77843 = pi15 ? n77841 : n77842;
  assign n77844 = pi14 ? n77840 : n77843;
  assign n77845 = pi13 ? n77838 : n77844;
  assign n77846 = pi16 ? n2120 : ~n2851;
  assign n77847 = pi15 ? n77842 : n77846;
  assign n77848 = pi14 ? n77842 : n77847;
  assign n77849 = pi16 ? n2120 : ~n3068;
  assign n77850 = pi16 ? n2120 : ~n2725;
  assign n77851 = pi14 ? n77849 : n77850;
  assign n77852 = pi13 ? n77848 : n77851;
  assign n77853 = pi12 ? n77845 : n77852;
  assign n77854 = pi16 ? n3625 : ~n2732;
  assign n77855 = pi16 ? n3625 : ~n2745;
  assign n77856 = pi14 ? n77854 : n77855;
  assign n77857 = pi16 ? n2426 : ~n2617;
  assign n77858 = pi16 ? n2120 : ~n2856;
  assign n77859 = pi16 ? n2426 : ~n2624;
  assign n77860 = pi15 ? n77858 : n77859;
  assign n77861 = pi14 ? n77857 : n77860;
  assign n77862 = pi13 ? n77856 : n77861;
  assign n77863 = pi16 ? n2120 : ~n2624;
  assign n77864 = pi16 ? n2120 : ~n2860;
  assign n77865 = pi15 ? n77863 : n77864;
  assign n77866 = pi16 ? n2293 : ~n4100;
  assign n77867 = pi15 ? n66183 : n77866;
  assign n77868 = pi14 ? n77865 : n77867;
  assign n77869 = pi16 ? n2293 : ~n2513;
  assign n77870 = pi16 ? n2293 : ~n2749;
  assign n77871 = pi15 ? n77869 : n77870;
  assign n77872 = pi14 ? n66193 : n77871;
  assign n77873 = pi13 ? n77868 : n77872;
  assign n77874 = pi12 ? n77862 : n77873;
  assign n77875 = pi11 ? n77853 : n77874;
  assign n77876 = pi10 ? n77835 : n77875;
  assign n77877 = pi09 ? n77788 : n77876;
  assign n77878 = pi17 ? n2461 : ~n3050;
  assign n77879 = pi16 ? n32 : n77878;
  assign n77880 = pi15 ? n32 : n77879;
  assign n77881 = pi17 ? n4167 : ~n3050;
  assign n77882 = pi16 ? n32 : n77881;
  assign n77883 = pi17 ? n1215 : ~n3050;
  assign n77884 = pi16 ? n32 : n77883;
  assign n77885 = pi15 ? n77882 : n77884;
  assign n77886 = pi14 ? n77880 : n77885;
  assign n77887 = pi13 ? n32 : n77886;
  assign n77888 = pi12 ? n32 : n77887;
  assign n77889 = pi11 ? n32 : n77888;
  assign n77890 = pi10 ? n32 : n77889;
  assign n77891 = pi15 ? n77777 : n77792;
  assign n77892 = pi17 ? n1605 : ~n2952;
  assign n77893 = pi16 ? n32 : n77892;
  assign n77894 = pi15 ? n77893 : n77684;
  assign n77895 = pi14 ? n77891 : n77894;
  assign n77896 = pi17 ? n1726 : ~n3050;
  assign n77897 = pi16 ? n32 : n77896;
  assign n77898 = pi15 ? n77692 : n77897;
  assign n77899 = pi17 ? n4041 : ~n3050;
  assign n77900 = pi16 ? n32 : n77899;
  assign n77901 = pi17 ? n3719 : ~n3050;
  assign n77902 = pi16 ? n32 : n77901;
  assign n77903 = pi15 ? n77900 : n77902;
  assign n77904 = pi14 ? n77898 : n77903;
  assign n77905 = pi13 ? n77895 : n77904;
  assign n77906 = pi16 ? n32 : ~n3051;
  assign n77907 = pi16 ? n3570 : ~n3051;
  assign n77908 = pi15 ? n77906 : n77907;
  assign n77909 = pi16 ? n3283 : ~n3051;
  assign n77910 = pi15 ? n77909 : n77699;
  assign n77911 = pi14 ? n77908 : n77910;
  assign n77912 = pi15 ? n77700 : n77704;
  assign n77913 = pi15 ? n77705 : n77707;
  assign n77914 = pi14 ? n77912 : n77913;
  assign n77915 = pi13 ? n77911 : n77914;
  assign n77916 = pi12 ? n77905 : n77915;
  assign n77917 = pi15 ? n77707 : n77503;
  assign n77918 = pi15 ? n77503 : n77406;
  assign n77919 = pi14 ? n77917 : n77918;
  assign n77920 = pi16 ? n2832 : ~n2958;
  assign n77921 = pi14 ? n77231 : n77920;
  assign n77922 = pi13 ? n77919 : n77921;
  assign n77923 = pi15 ? n77817 : n77504;
  assign n77924 = pi16 ? n4246 : ~n2958;
  assign n77925 = pi15 ? n77308 : n77924;
  assign n77926 = pi14 ? n77923 : n77925;
  assign n77927 = pi16 ? n4246 : ~n3183;
  assign n77928 = pi15 ? n76989 : n76991;
  assign n77929 = pi14 ? n77927 : n77928;
  assign n77930 = pi13 ? n77926 : n77929;
  assign n77931 = pi12 ? n77922 : n77930;
  assign n77932 = pi11 ? n77916 : n77931;
  assign n77933 = pi16 ? n2860 : ~n2832;
  assign n77934 = pi15 ? n76937 : n77933;
  assign n77935 = pi14 ? n76937 : n77934;
  assign n77936 = pi16 ? n3946 : ~n2837;
  assign n77937 = pi15 ? n77933 : n77936;
  assign n77938 = pi16 ? n3946 : ~n2840;
  assign n77939 = pi15 ? n77936 : n77938;
  assign n77940 = pi14 ? n77937 : n77939;
  assign n77941 = pi13 ? n77935 : n77940;
  assign n77942 = pi16 ? n3946 : ~n2851;
  assign n77943 = pi15 ? n77938 : n77942;
  assign n77944 = pi16 ? n2756 : ~n2851;
  assign n77945 = pi15 ? n77942 : n77944;
  assign n77946 = pi14 ? n77943 : n77945;
  assign n77947 = pi16 ? n2756 : ~n3068;
  assign n77948 = pi15 ? n77944 : n77947;
  assign n77949 = pi16 ? n2756 : ~n4246;
  assign n77950 = pi14 ? n77948 : n77949;
  assign n77951 = pi13 ? n77946 : n77950;
  assign n77952 = pi12 ? n77941 : n77951;
  assign n77953 = pi16 ? n2293 : ~n2725;
  assign n77954 = pi16 ? n2293 : ~n2732;
  assign n77955 = pi15 ? n77953 : n77954;
  assign n77956 = pi16 ? n2293 : ~n2745;
  assign n77957 = pi14 ? n77955 : n77956;
  assign n77958 = pi16 ? n3769 : ~n2617;
  assign n77959 = pi15 ? n63613 : n77958;
  assign n77960 = pi16 ? n2749 : ~n2856;
  assign n77961 = pi16 ? n3769 : ~n2856;
  assign n77962 = pi15 ? n77960 : n77961;
  assign n77963 = pi14 ? n77959 : n77962;
  assign n77964 = pi13 ? n77957 : n77963;
  assign n77965 = pi16 ? n2749 : ~n2624;
  assign n77966 = pi16 ? n2749 : ~n2860;
  assign n77967 = pi15 ? n77965 : n77966;
  assign n77968 = pi15 ? n66307 : n66311;
  assign n77969 = pi14 ? n77967 : n77968;
  assign n77970 = pi16 ? n2513 : ~n2513;
  assign n77971 = pi16 ? n4100 : ~n2513;
  assign n77972 = pi15 ? n77970 : n77971;
  assign n77973 = pi14 ? n66313 : n77972;
  assign n77974 = pi13 ? n77969 : n77973;
  assign n77975 = pi12 ? n77964 : n77974;
  assign n77976 = pi11 ? n77952 : n77975;
  assign n77977 = pi10 ? n77932 : n77976;
  assign n77978 = pi09 ? n77890 : n77977;
  assign n77979 = pi08 ? n77877 : n77978;
  assign n77980 = pi07 ? n77775 : n77979;
  assign n77981 = pi17 ? n1480 : ~n2959;
  assign n77982 = pi16 ? n32 : n77981;
  assign n77983 = pi15 ? n32 : n77982;
  assign n77984 = pi17 ? n4341 : ~n2959;
  assign n77985 = pi16 ? n32 : n77984;
  assign n77986 = pi17 ? n1989 : ~n2959;
  assign n77987 = pi16 ? n32 : n77986;
  assign n77988 = pi15 ? n77985 : n77987;
  assign n77989 = pi14 ? n77983 : n77988;
  assign n77990 = pi13 ? n32 : n77989;
  assign n77991 = pi12 ? n32 : n77990;
  assign n77992 = pi11 ? n32 : n77991;
  assign n77993 = pi10 ? n32 : n77992;
  assign n77994 = pi17 ? n2461 : ~n2959;
  assign n77995 = pi16 ? n32 : n77994;
  assign n77996 = pi17 ? n2355 : ~n2959;
  assign n77997 = pi16 ? n32 : n77996;
  assign n77998 = pi15 ? n77995 : n77997;
  assign n77999 = pi14 ? n77998 : n77783;
  assign n78000 = pi17 ? n1219 : ~n3050;
  assign n78001 = pi16 ? n32 : n78000;
  assign n78002 = pi15 ? n77790 : n78001;
  assign n78003 = pi17 ? n1605 : ~n3050;
  assign n78004 = pi16 ? n32 : n78003;
  assign n78005 = pi15 ? n78004 : n77900;
  assign n78006 = pi14 ? n78002 : n78005;
  assign n78007 = pi13 ? n77999 : n78006;
  assign n78008 = pi17 ? n2005 : ~n3050;
  assign n78009 = pi16 ? n32 : n78008;
  assign n78010 = pi17 ? n3715 : ~n3050;
  assign n78011 = pi16 ? n32 : n78010;
  assign n78012 = pi15 ? n78009 : n78011;
  assign n78013 = pi17 ? n1028 : ~n3050;
  assign n78014 = pi16 ? n32 : n78013;
  assign n78015 = pi15 ? n78014 : n77802;
  assign n78016 = pi14 ? n78012 : n78015;
  assign n78017 = pi15 ? n77699 : n77806;
  assign n78018 = pi16 ? n3729 : ~n3051;
  assign n78019 = pi16 ? n3165 : ~n3051;
  assign n78020 = pi15 ? n78018 : n78019;
  assign n78021 = pi14 ? n78017 : n78020;
  assign n78022 = pi13 ? n78016 : n78021;
  assign n78023 = pi12 ? n78007 : n78022;
  assign n78024 = pi16 ? n3047 : ~n3051;
  assign n78025 = pi15 ? n78024 : n77700;
  assign n78026 = pi14 ? n78025 : n77912;
  assign n78027 = pi16 ? n3051 : ~n3176;
  assign n78028 = pi14 ? n78027 : n77500;
  assign n78029 = pi13 ? n78026 : n78028;
  assign n78030 = pi15 ? n77406 : n77408;
  assign n78031 = pi14 ? n77610 : n78030;
  assign n78032 = pi16 ? n3183 : ~n3183;
  assign n78033 = pi16 ? n3061 : ~n3183;
  assign n78034 = pi15 ? n77040 : n78033;
  assign n78035 = pi14 ? n78032 : n78034;
  assign n78036 = pi13 ? n78031 : n78035;
  assign n78037 = pi12 ? n78029 : n78036;
  assign n78038 = pi11 ? n78023 : n78037;
  assign n78039 = pi16 ? n3068 : ~n2832;
  assign n78040 = pi15 ? n77050 : n78039;
  assign n78041 = pi14 ? n77050 : n78040;
  assign n78042 = pi16 ? n4246 : ~n2832;
  assign n78043 = pi16 ? n2617 : ~n2837;
  assign n78044 = pi15 ? n78042 : n78043;
  assign n78045 = pi16 ? n2617 : ~n2840;
  assign n78046 = pi15 ? n78043 : n78045;
  assign n78047 = pi14 ? n78044 : n78046;
  assign n78048 = pi13 ? n78041 : n78047;
  assign n78049 = pi16 ? n2624 : ~n2840;
  assign n78050 = pi16 ? n2624 : ~n2851;
  assign n78051 = pi15 ? n78049 : n78050;
  assign n78052 = pi14 ? n78045 : n78051;
  assign n78053 = pi16 ? n2624 : ~n3068;
  assign n78054 = pi15 ? n78050 : n78053;
  assign n78055 = pi16 ? n2624 : ~n4246;
  assign n78056 = pi14 ? n78054 : n78055;
  assign n78057 = pi13 ? n78052 : n78056;
  assign n78058 = pi12 ? n78048 : n78057;
  assign n78059 = pi16 ? n2513 : ~n2725;
  assign n78060 = pi16 ? n2513 : ~n2732;
  assign n78061 = pi16 ? n2513 : ~n2745;
  assign n78062 = pi15 ? n78060 : n78061;
  assign n78063 = pi14 ? n78059 : n78062;
  assign n78064 = pi15 ? n63611 : n63422;
  assign n78065 = pi14 ? n78064 : n63534;
  assign n78066 = pi13 ? n78063 : n78065;
  assign n78067 = pi16 ? n4100 : ~n2624;
  assign n78068 = pi15 ? n78067 : n66456;
  assign n78069 = pi14 ? n62285 : n78068;
  assign n78070 = pi16 ? n2745 : ~n3946;
  assign n78071 = pi15 ? n66456 : n78070;
  assign n78072 = pi16 ? n2745 : ~n2629;
  assign n78073 = pi16 ? n2745 : ~n2513;
  assign n78074 = pi15 ? n78072 : n78073;
  assign n78075 = pi14 ? n78071 : n78074;
  assign n78076 = pi13 ? n78069 : n78075;
  assign n78077 = pi12 ? n78066 : n78076;
  assign n78078 = pi11 ? n78058 : n78077;
  assign n78079 = pi10 ? n78038 : n78078;
  assign n78080 = pi09 ? n77993 : n78079;
  assign n78081 = pi17 ? n2159 : ~n2959;
  assign n78082 = pi16 ? n32 : n78081;
  assign n78083 = pi15 ? n32 : n78082;
  assign n78084 = pi17 ? n4497 : ~n2959;
  assign n78085 = pi16 ? n32 : n78084;
  assign n78086 = pi17 ? n1472 : ~n2959;
  assign n78087 = pi16 ? n32 : n78086;
  assign n78088 = pi15 ? n78085 : n78087;
  assign n78089 = pi14 ? n78083 : n78088;
  assign n78090 = pi13 ? n32 : n78089;
  assign n78091 = pi12 ? n32 : n78090;
  assign n78092 = pi11 ? n32 : n78091;
  assign n78093 = pi10 ? n32 : n78092;
  assign n78094 = pi15 ? n77982 : n77995;
  assign n78095 = pi14 ? n78094 : n77885;
  assign n78096 = pi17 ? n4515 : ~n3050;
  assign n78097 = pi16 ? n32 : n78096;
  assign n78098 = pi17 ? n4023 : ~n2959;
  assign n78099 = pi16 ? n32 : n78098;
  assign n78100 = pi15 ? n78097 : n78099;
  assign n78101 = pi17 ? n1605 : ~n2959;
  assign n78102 = pi16 ? n32 : n78101;
  assign n78103 = pi14 ? n78100 : n78102;
  assign n78104 = pi13 ? n78095 : n78103;
  assign n78105 = pi17 ? n1227 : ~n2959;
  assign n78106 = pi16 ? n32 : n78105;
  assign n78107 = pi17 ? n3553 : ~n2959;
  assign n78108 = pi16 ? n32 : n78107;
  assign n78109 = pi15 ? n78106 : n78108;
  assign n78110 = pi17 ? n1726 : ~n2959;
  assign n78111 = pi16 ? n32 : n78110;
  assign n78112 = pi15 ? n78111 : n77900;
  assign n78113 = pi14 ? n78109 : n78112;
  assign n78114 = pi15 ? n77902 : n77906;
  assign n78115 = pi15 ? n77907 : n77909;
  assign n78116 = pi14 ? n78114 : n78115;
  assign n78117 = pi13 ? n78113 : n78116;
  assign n78118 = pi12 ? n78104 : n78117;
  assign n78119 = pi16 ? n3156 : ~n3051;
  assign n78120 = pi15 ? n78119 : n77699;
  assign n78121 = pi14 ? n78120 : n78017;
  assign n78122 = pi16 ? n3161 : ~n3176;
  assign n78123 = pi15 ? n78122 : n77403;
  assign n78124 = pi14 ? n78123 : n77403;
  assign n78125 = pi13 ? n78121 : n78124;
  assign n78126 = pi16 ? n4578 : ~n2953;
  assign n78127 = pi15 ? n77700 : n78126;
  assign n78128 = pi16 ? n4578 : ~n3176;
  assign n78129 = pi15 ? n78128 : n78027;
  assign n78130 = pi14 ? n78127 : n78129;
  assign n78131 = pi14 ? n77157 : n77097;
  assign n78132 = pi13 ? n78130 : n78131;
  assign n78133 = pi12 ? n78125 : n78132;
  assign n78134 = pi11 ? n78118 : n78133;
  assign n78135 = pi16 ? n2958 : ~n3183;
  assign n78136 = pi16 ? n2964 : ~n3183;
  assign n78137 = pi15 ? n78135 : n78136;
  assign n78138 = pi14 ? n78135 : n78137;
  assign n78139 = pi16 ? n3183 : ~n2832;
  assign n78140 = pi16 ? n2840 : ~n3061;
  assign n78141 = pi15 ? n78139 : n78140;
  assign n78142 = pi16 ? n2837 : ~n3061;
  assign n78143 = pi16 ? n2837 : ~n2837;
  assign n78144 = pi15 ? n78142 : n78143;
  assign n78145 = pi14 ? n78141 : n78144;
  assign n78146 = pi13 ? n78138 : n78145;
  assign n78147 = pi16 ? n2837 : ~n2840;
  assign n78148 = pi16 ? n2840 : ~n2840;
  assign n78149 = pi15 ? n78147 : n78148;
  assign n78150 = pi16 ? n2725 : ~n2840;
  assign n78151 = pi14 ? n78149 : n78150;
  assign n78152 = pi16 ? n2725 : ~n2851;
  assign n78153 = pi16 ? n2725 : ~n3068;
  assign n78154 = pi15 ? n78152 : n78153;
  assign n78155 = pi16 ? n2745 : ~n4246;
  assign n78156 = pi15 ? n78153 : n78155;
  assign n78157 = pi14 ? n78154 : n78156;
  assign n78158 = pi13 ? n78151 : n78157;
  assign n78159 = pi12 ? n78146 : n78158;
  assign n78160 = pi16 ? n2745 : ~n2725;
  assign n78161 = pi14 ? n78160 : n63697;
  assign n78162 = pi16 ? n2732 : ~n2732;
  assign n78163 = pi15 ? n78162 : n63404;
  assign n78164 = pi16 ? n3068 : ~n2856;
  assign n78165 = pi15 ? n63404 : n78164;
  assign n78166 = pi14 ? n78163 : n78165;
  assign n78167 = pi13 ? n78161 : n78166;
  assign n78168 = pi16 ? n4246 : ~n2624;
  assign n78169 = pi16 ? n2851 : ~n4100;
  assign n78170 = pi15 ? n78168 : n78169;
  assign n78171 = pi14 ? n49412 : n78170;
  assign n78172 = pi16 ? n2851 : ~n3946;
  assign n78173 = pi15 ? n66579 : n78172;
  assign n78174 = pi16 ? n2837 : ~n2629;
  assign n78175 = pi15 ? n46675 : n78174;
  assign n78176 = pi14 ? n78173 : n78175;
  assign n78177 = pi13 ? n78171 : n78176;
  assign n78178 = pi12 ? n78167 : n78177;
  assign n78179 = pi11 ? n78159 : n78178;
  assign n78180 = pi10 ? n78134 : n78179;
  assign n78181 = pi09 ? n78093 : n78180;
  assign n78182 = pi08 ? n78080 : n78181;
  assign n78183 = pi17 ? n1706 : ~n3587;
  assign n78184 = pi16 ? n32 : n78183;
  assign n78185 = pi15 ? n32 : n78184;
  assign n78186 = pi17 ? n4656 : ~n3587;
  assign n78187 = pi16 ? n32 : n78186;
  assign n78188 = pi17 ? n4659 : ~n3587;
  assign n78189 = pi16 ? n32 : n78188;
  assign n78190 = pi15 ? n78187 : n78189;
  assign n78191 = pi14 ? n78185 : n78190;
  assign n78192 = pi13 ? n32 : n78191;
  assign n78193 = pi12 ? n32 : n78192;
  assign n78194 = pi11 ? n32 : n78193;
  assign n78195 = pi10 ? n32 : n78194;
  assign n78196 = pi17 ? n2159 : ~n3587;
  assign n78197 = pi16 ? n32 : n78196;
  assign n78198 = pi17 ? n1480 : ~n3587;
  assign n78199 = pi16 ? n32 : n78198;
  assign n78200 = pi15 ? n78197 : n78199;
  assign n78201 = pi14 ? n78200 : n77988;
  assign n78202 = pi17 ? n4682 : ~n2959;
  assign n78203 = pi16 ? n32 : n78202;
  assign n78204 = pi17 ? n4167 : ~n2959;
  assign n78205 = pi16 ? n32 : n78204;
  assign n78206 = pi15 ? n78203 : n78205;
  assign n78207 = pi14 ? n78206 : n78099;
  assign n78208 = pi13 ? n78201 : n78207;
  assign n78209 = pi17 ? n1120 : ~n2959;
  assign n78210 = pi16 ? n32 : n78209;
  assign n78211 = pi17 ? n4034 : ~n2959;
  assign n78212 = pi16 ? n32 : n78211;
  assign n78213 = pi15 ? n78210 : n78212;
  assign n78214 = pi15 ? n78001 : n78004;
  assign n78215 = pi14 ? n78213 : n78214;
  assign n78216 = pi17 ? n2005 : ~n2959;
  assign n78217 = pi16 ? n32 : n78216;
  assign n78218 = pi15 ? n77900 : n78217;
  assign n78219 = pi17 ? n3715 : ~n2959;
  assign n78220 = pi16 ? n32 : n78219;
  assign n78221 = pi17 ? n1028 : ~n2959;
  assign n78222 = pi16 ? n32 : n78221;
  assign n78223 = pi15 ? n78220 : n78222;
  assign n78224 = pi14 ? n78218 : n78223;
  assign n78225 = pi13 ? n78215 : n78224;
  assign n78226 = pi12 ? n78208 : n78225;
  assign n78227 = pi17 ? n3719 : ~n2959;
  assign n78228 = pi16 ? n32 : n78227;
  assign n78229 = pi15 ? n78228 : n77902;
  assign n78230 = pi17 ? n3557 : ~n3050;
  assign n78231 = pi16 ? n32 : n78230;
  assign n78232 = pi15 ? n78231 : n77906;
  assign n78233 = pi14 ? n78229 : n78232;
  assign n78234 = pi16 ? n3570 : ~n2953;
  assign n78235 = pi15 ? n78234 : n77697;
  assign n78236 = pi14 ? n78235 : n77697;
  assign n78237 = pi13 ? n78233 : n78236;
  assign n78238 = pi16 ? n4740 : ~n2953;
  assign n78239 = pi15 ? n77699 : n78238;
  assign n78240 = pi14 ? n78239 : n78122;
  assign n78241 = pi16 ? n3161 : ~n2964;
  assign n78242 = pi16 ? n3293 : ~n2964;
  assign n78243 = pi14 ? n78241 : n78242;
  assign n78244 = pi13 ? n78240 : n78243;
  assign n78245 = pi12 ? n78237 : n78244;
  assign n78246 = pi11 ? n78226 : n78245;
  assign n78247 = pi16 ? n3588 : ~n2964;
  assign n78248 = pi16 ? n3588 : ~n3183;
  assign n78249 = pi16 ? n4578 : ~n3183;
  assign n78250 = pi15 ? n78248 : n78249;
  assign n78251 = pi14 ? n78247 : n78250;
  assign n78252 = pi16 ? n4578 : ~n2832;
  assign n78253 = pi16 ? n2953 : ~n3061;
  assign n78254 = pi15 ? n78252 : n78253;
  assign n78255 = pi16 ? n2953 : ~n2837;
  assign n78256 = pi15 ? n78253 : n78255;
  assign n78257 = pi14 ? n78254 : n78256;
  assign n78258 = pi13 ? n78251 : n78257;
  assign n78259 = pi16 ? n3176 : ~n2837;
  assign n78260 = pi15 ? n78255 : n78259;
  assign n78261 = pi16 ? n2832 : ~n2840;
  assign n78262 = pi14 ? n78260 : n78261;
  assign n78263 = pi16 ? n2832 : ~n2851;
  assign n78264 = pi16 ? n3183 : ~n3068;
  assign n78265 = pi15 ? n78263 : n78264;
  assign n78266 = pi16 ? n2832 : ~n3068;
  assign n78267 = pi16 ? n2851 : ~n3068;
  assign n78268 = pi15 ? n78266 : n78267;
  assign n78269 = pi14 ? n78265 : n78268;
  assign n78270 = pi13 ? n78262 : n78269;
  assign n78271 = pi12 ? n78258 : n78270;
  assign n78272 = pi16 ? n2851 : ~n4246;
  assign n78273 = pi16 ? n2851 : ~n2732;
  assign n78274 = pi16 ? n3061 : ~n2732;
  assign n78275 = pi15 ? n78273 : n78274;
  assign n78276 = pi14 ? n78272 : n78275;
  assign n78277 = pi16 ? n2832 : ~n2745;
  assign n78278 = pi15 ? n78274 : n78277;
  assign n78279 = pi16 ? n2832 : ~n2617;
  assign n78280 = pi14 ? n78278 : n78279;
  assign n78281 = pi13 ? n78276 : n78280;
  assign n78282 = pi15 ? n62269 : n66713;
  assign n78283 = pi15 ? n61765 : n47041;
  assign n78284 = pi14 ? n78282 : n78283;
  assign n78285 = pi16 ? n3176 : ~n4100;
  assign n78286 = pi15 ? n78285 : n47041;
  assign n78287 = pi14 ? n78286 : n63968;
  assign n78288 = pi13 ? n78284 : n78287;
  assign n78289 = pi12 ? n78281 : n78288;
  assign n78290 = pi11 ? n78271 : n78289;
  assign n78291 = pi10 ? n78246 : n78290;
  assign n78292 = pi09 ? n78195 : n78291;
  assign n78293 = pi17 ? n4798 : ~n3587;
  assign n78294 = pi16 ? n32 : n78293;
  assign n78295 = pi15 ? n32 : n78294;
  assign n78296 = pi17 ? n1966 : ~n3587;
  assign n78297 = pi16 ? n32 : n78296;
  assign n78298 = pi17 ? n4804 : ~n3587;
  assign n78299 = pi16 ? n32 : n78298;
  assign n78300 = pi15 ? n78297 : n78299;
  assign n78301 = pi14 ? n78295 : n78300;
  assign n78302 = pi13 ? n32 : n78301;
  assign n78303 = pi12 ? n32 : n78302;
  assign n78304 = pi11 ? n32 : n78303;
  assign n78305 = pi10 ? n32 : n78304;
  assign n78306 = pi15 ? n78184 : n78197;
  assign n78307 = pi14 ? n78306 : n78088;
  assign n78308 = pi17 ? n4822 : ~n3587;
  assign n78309 = pi16 ? n32 : n78308;
  assign n78310 = pi17 ? n4341 : ~n3587;
  assign n78311 = pi16 ? n32 : n78310;
  assign n78312 = pi15 ? n78309 : n78311;
  assign n78313 = pi17 ? n4167 : ~n3587;
  assign n78314 = pi16 ? n32 : n78313;
  assign n78315 = pi14 ? n78312 : n78314;
  assign n78316 = pi13 ? n78307 : n78315;
  assign n78317 = pi17 ? n1215 : ~n3587;
  assign n78318 = pi16 ? n32 : n78317;
  assign n78319 = pi17 ? n4515 : ~n3587;
  assign n78320 = pi16 ? n32 : n78319;
  assign n78321 = pi15 ? n78318 : n78320;
  assign n78322 = pi17 ? n4023 : ~n3587;
  assign n78323 = pi16 ? n32 : n78322;
  assign n78324 = pi15 ? n78323 : n78102;
  assign n78325 = pi14 ? n78321 : n78324;
  assign n78326 = pi15 ? n78102 : n78106;
  assign n78327 = pi15 ? n78108 : n78111;
  assign n78328 = pi14 ? n78326 : n78327;
  assign n78329 = pi13 ? n78325 : n78328;
  assign n78330 = pi12 ? n78316 : n78329;
  assign n78331 = pi17 ? n4041 : ~n2959;
  assign n78332 = pi16 ? n32 : n78331;
  assign n78333 = pi15 ? n78332 : n77900;
  assign n78334 = pi17 ? n3704 : ~n3050;
  assign n78335 = pi16 ? n32 : n78334;
  assign n78336 = pi15 ? n78335 : n77596;
  assign n78337 = pi14 ? n78333 : n78336;
  assign n78338 = pi17 ? n2008 : ~n2952;
  assign n78339 = pi16 ? n32 : n78338;
  assign n78340 = pi15 ? n77799 : n78339;
  assign n78341 = pi14 ? n77800 : n78340;
  assign n78342 = pi13 ? n78337 : n78341;
  assign n78343 = pi15 ? n78231 : n77694;
  assign n78344 = pi15 ? n78234 : n77493;
  assign n78345 = pi14 ? n78343 : n78344;
  assign n78346 = pi16 ? n3570 : ~n2958;
  assign n78347 = pi16 ? n3438 : ~n2958;
  assign n78348 = pi16 ? n3729 : ~n2964;
  assign n78349 = pi15 ? n78347 : n78348;
  assign n78350 = pi14 ? n78346 : n78349;
  assign n78351 = pi13 ? n78345 : n78350;
  assign n78352 = pi12 ? n78342 : n78351;
  assign n78353 = pi11 ? n78330 : n78352;
  assign n78354 = pi16 ? n3165 : ~n3183;
  assign n78355 = pi15 ? n78348 : n78354;
  assign n78356 = pi14 ? n78348 : n78355;
  assign n78357 = pi16 ? n3165 : ~n2832;
  assign n78358 = pi16 ? n3047 : ~n2832;
  assign n78359 = pi15 ? n78357 : n78358;
  assign n78360 = pi16 ? n3047 : ~n3061;
  assign n78361 = pi16 ? n3047 : ~n2837;
  assign n78362 = pi15 ? n78360 : n78361;
  assign n78363 = pi14 ? n78359 : n78362;
  assign n78364 = pi13 ? n78356 : n78363;
  assign n78365 = pi16 ? n3588 : ~n2837;
  assign n78366 = pi15 ? n78255 : n78365;
  assign n78367 = pi14 ? n78361 : n78366;
  assign n78368 = pi16 ? n3588 : ~n2851;
  assign n78369 = pi16 ? n4578 : ~n3068;
  assign n78370 = pi16 ? n2832 : ~n4246;
  assign n78371 = pi15 ? n78369 : n78370;
  assign n78372 = pi14 ? n78368 : n78371;
  assign n78373 = pi13 ? n78367 : n78372;
  assign n78374 = pi12 ? n78364 : n78373;
  assign n78375 = pi16 ? n2958 : ~n4246;
  assign n78376 = pi16 ? n3176 : ~n2732;
  assign n78377 = pi15 ? n63823 : n78376;
  assign n78378 = pi14 ? n78375 : n78377;
  assign n78379 = pi16 ? n3176 : ~n2745;
  assign n78380 = pi15 ? n78376 : n78379;
  assign n78381 = pi16 ? n4578 : ~n2745;
  assign n78382 = pi15 ? n78379 : n78381;
  assign n78383 = pi14 ? n78380 : n78382;
  assign n78384 = pi13 ? n78378 : n78383;
  assign n78385 = pi16 ? n4578 : ~n2617;
  assign n78386 = pi15 ? n78385 : n66838;
  assign n78387 = pi16 ? n3588 : ~n2624;
  assign n78388 = pi16 ? n3588 : ~n2860;
  assign n78389 = pi15 ? n78387 : n78388;
  assign n78390 = pi14 ? n78386 : n78389;
  assign n78391 = pi16 ? n3165 : ~n4100;
  assign n78392 = pi15 ? n78388 : n78391;
  assign n78393 = pi16 ? n3047 : ~n3946;
  assign n78394 = pi16 ? n3047 : ~n2629;
  assign n78395 = pi15 ? n78393 : n78394;
  assign n78396 = pi14 ? n78392 : n78395;
  assign n78397 = pi13 ? n78390 : n78396;
  assign n78398 = pi12 ? n78384 : n78397;
  assign n78399 = pi11 ? n78374 : n78398;
  assign n78400 = pi10 ? n78353 : n78399;
  assign n78401 = pi09 ? n78305 : n78400;
  assign n78402 = pi08 ? n78292 : n78401;
  assign n78403 = pi07 ? n78182 : n78402;
  assign n78404 = pi06 ? n77980 : n78403;
  assign n78405 = pi17 ? n1971 : ~n3292;
  assign n78406 = pi16 ? n32 : n78405;
  assign n78407 = pi15 ? n32 : n78406;
  assign n78408 = pi17 ? n930 : ~n3292;
  assign n78409 = pi16 ? n32 : n78408;
  assign n78410 = pi17 ? n1134 : ~n3292;
  assign n78411 = pi16 ? n32 : n78410;
  assign n78412 = pi15 ? n78409 : n78411;
  assign n78413 = pi14 ? n78407 : n78412;
  assign n78414 = pi13 ? n32 : n78413;
  assign n78415 = pi12 ? n32 : n78414;
  assign n78416 = pi11 ? n32 : n78415;
  assign n78417 = pi10 ? n32 : n78416;
  assign n78418 = pi17 ? n1706 : ~n3292;
  assign n78419 = pi16 ? n32 : n78418;
  assign n78420 = pi17 ? n1700 : ~n3587;
  assign n78421 = pi16 ? n32 : n78420;
  assign n78422 = pi15 ? n78187 : n78421;
  assign n78423 = pi14 ? n78419 : n78422;
  assign n78424 = pi17 ? n4497 : ~n3587;
  assign n78425 = pi16 ? n32 : n78424;
  assign n78426 = pi15 ? n78197 : n78425;
  assign n78427 = pi14 ? n78426 : n78311;
  assign n78428 = pi13 ? n78423 : n78427;
  assign n78429 = pi17 ? n1989 : ~n3587;
  assign n78430 = pi16 ? n32 : n78429;
  assign n78431 = pi17 ? n4682 : ~n3587;
  assign n78432 = pi16 ? n32 : n78431;
  assign n78433 = pi15 ? n78430 : n78432;
  assign n78434 = pi15 ? n78314 : n78099;
  assign n78435 = pi14 ? n78433 : n78434;
  assign n78436 = pi17 ? n1120 : ~n3587;
  assign n78437 = pi16 ? n32 : n78436;
  assign n78438 = pi15 ? n78099 : n78437;
  assign n78439 = pi17 ? n4034 : ~n3587;
  assign n78440 = pi16 ? n32 : n78439;
  assign n78441 = pi17 ? n1219 : ~n3587;
  assign n78442 = pi16 ? n32 : n78441;
  assign n78443 = pi15 ? n78440 : n78442;
  assign n78444 = pi14 ? n78438 : n78443;
  assign n78445 = pi13 ? n78435 : n78444;
  assign n78446 = pi12 ? n78428 : n78445;
  assign n78447 = pi17 ? n1605 : ~n3587;
  assign n78448 = pi16 ? n32 : n78447;
  assign n78449 = pi15 ? n78448 : n78102;
  assign n78450 = pi17 ? n3855 : ~n2959;
  assign n78451 = pi16 ? n32 : n78450;
  assign n78452 = pi17 ? n1227 : ~n3050;
  assign n78453 = pi16 ? n32 : n78452;
  assign n78454 = pi15 ? n78451 : n78453;
  assign n78455 = pi14 ? n78449 : n78454;
  assign n78456 = pi17 ? n3553 : ~n3050;
  assign n78457 = pi16 ? n32 : n78456;
  assign n78458 = pi15 ? n78457 : n77897;
  assign n78459 = pi17 ? n1500 : ~n3050;
  assign n78460 = pi16 ? n32 : n78459;
  assign n78461 = pi15 ? n77897 : n78460;
  assign n78462 = pi14 ? n78458 : n78461;
  assign n78463 = pi13 ? n78455 : n78462;
  assign n78464 = pi17 ? n3715 : ~n3175;
  assign n78465 = pi16 ? n32 : n78464;
  assign n78466 = pi15 ? n77598 : n78465;
  assign n78467 = pi14 ? n78336 : n78466;
  assign n78468 = pi17 ? n3719 : ~n2726;
  assign n78469 = pi16 ? n32 : n78468;
  assign n78470 = pi17 ? n2008 : ~n2726;
  assign n78471 = pi16 ? n32 : n78470;
  assign n78472 = pi17 ? n3557 : ~n2726;
  assign n78473 = pi16 ? n32 : n78472;
  assign n78474 = pi15 ? n78471 : n78473;
  assign n78475 = pi14 ? n78469 : n78474;
  assign n78476 = pi13 ? n78467 : n78475;
  assign n78477 = pi12 ? n78463 : n78476;
  assign n78478 = pi11 ? n78446 : n78477;
  assign n78479 = pi17 ? n3557 : ~n2963;
  assign n78480 = pi16 ? n32 : n78479;
  assign n78481 = pi15 ? n78473 : n78480;
  assign n78482 = pi16 ? n3283 : ~n3183;
  assign n78483 = pi15 ? n78480 : n78482;
  assign n78484 = pi14 ? n78481 : n78483;
  assign n78485 = pi16 ? n3156 : ~n2832;
  assign n78486 = pi16 ? n3156 : ~n3061;
  assign n78487 = pi15 ? n78485 : n78486;
  assign n78488 = pi14 ? n78485 : n78487;
  assign n78489 = pi13 ? n78484 : n78488;
  assign n78490 = pi16 ? n3729 : ~n3061;
  assign n78491 = pi16 ? n3729 : ~n2837;
  assign n78492 = pi15 ? n78490 : n78491;
  assign n78493 = pi16 ? n4740 : ~n2837;
  assign n78494 = pi14 ? n78492 : n78493;
  assign n78495 = pi16 ? n4740 : ~n2840;
  assign n78496 = pi16 ? n4740 : ~n2851;
  assign n78497 = pi15 ? n78495 : n78496;
  assign n78498 = pi16 ? n3588 : ~n3068;
  assign n78499 = pi15 ? n78496 : n78498;
  assign n78500 = pi14 ? n78497 : n78499;
  assign n78501 = pi13 ? n78494 : n78500;
  assign n78502 = pi12 ? n78489 : n78501;
  assign n78503 = pi16 ? n3588 : ~n4246;
  assign n78504 = pi15 ? n78498 : n78503;
  assign n78505 = pi14 ? n78504 : n63810;
  assign n78506 = pi16 ? n3165 : ~n2745;
  assign n78507 = pi15 ? n63810 : n78506;
  assign n78508 = pi16 ? n3161 : ~n2617;
  assign n78509 = pi15 ? n78506 : n78508;
  assign n78510 = pi14 ? n78507 : n78509;
  assign n78511 = pi13 ? n78505 : n78510;
  assign n78512 = pi16 ? n3161 : ~n2856;
  assign n78513 = pi16 ? n3438 : ~n2624;
  assign n78514 = pi16 ? n3438 : ~n2860;
  assign n78515 = pi15 ? n78513 : n78514;
  assign n78516 = pi14 ? n78512 : n78515;
  assign n78517 = pi16 ? n3438 : ~n4100;
  assign n78518 = pi16 ? n3156 : ~n4100;
  assign n78519 = pi15 ? n78517 : n78518;
  assign n78520 = pi16 ? n3438 : ~n3946;
  assign n78521 = pi15 ? n78520 : n49846;
  assign n78522 = pi14 ? n78519 : n78521;
  assign n78523 = pi13 ? n78516 : n78522;
  assign n78524 = pi12 ? n78511 : n78523;
  assign n78525 = pi11 ? n78502 : n78524;
  assign n78526 = pi10 ? n78478 : n78525;
  assign n78527 = pi09 ? n78417 : n78526;
  assign n78528 = pi17 ? n1593 : ~n3292;
  assign n78529 = pi16 ? n32 : n78528;
  assign n78530 = pi15 ? n32 : n78529;
  assign n78531 = pi17 ? n1470 : ~n3292;
  assign n78532 = pi16 ? n32 : n78531;
  assign n78533 = pi14 ? n78530 : n78532;
  assign n78534 = pi13 ? n32 : n78533;
  assign n78535 = pi12 ? n32 : n78534;
  assign n78536 = pi11 ? n32 : n78535;
  assign n78537 = pi10 ? n32 : n78536;
  assign n78538 = pi14 ? n78411 : n78300;
  assign n78539 = pi17 ? n4656 : ~n3292;
  assign n78540 = pi16 ? n32 : n78539;
  assign n78541 = pi15 ? n78419 : n78540;
  assign n78542 = pi17 ? n4497 : ~n3292;
  assign n78543 = pi16 ? n32 : n78542;
  assign n78544 = pi14 ? n78541 : n78543;
  assign n78545 = pi13 ? n78538 : n78544;
  assign n78546 = pi17 ? n1472 : ~n3292;
  assign n78547 = pi16 ? n32 : n78546;
  assign n78548 = pi17 ? n4822 : ~n3292;
  assign n78549 = pi16 ? n32 : n78548;
  assign n78550 = pi15 ? n78547 : n78549;
  assign n78551 = pi17 ? n4341 : ~n3292;
  assign n78552 = pi16 ? n32 : n78551;
  assign n78553 = pi15 ? n78552 : n78314;
  assign n78554 = pi14 ? n78550 : n78553;
  assign n78555 = pi15 ? n78314 : n78318;
  assign n78556 = pi15 ? n78320 : n78323;
  assign n78557 = pi14 ? n78555 : n78556;
  assign n78558 = pi13 ? n78554 : n78557;
  assign n78559 = pi12 ? n78545 : n78558;
  assign n78560 = pi15 ? n78323 : n78099;
  assign n78561 = pi15 ? n78099 : n77782;
  assign n78562 = pi14 ? n78560 : n78561;
  assign n78563 = pi15 ? n77792 : n78004;
  assign n78564 = pi14 ? n77793 : n78563;
  assign n78565 = pi13 ? n78562 : n78564;
  assign n78566 = pi15 ? n78457 : n77692;
  assign n78567 = pi14 ? n78454 : n78566;
  assign n78568 = pi17 ? n4041 : ~n3175;
  assign n78569 = pi16 ? n32 : n78568;
  assign n78570 = pi17 ? n1500 : ~n2726;
  assign n78571 = pi16 ? n32 : n78570;
  assign n78572 = pi17 ? n3704 : ~n2726;
  assign n78573 = pi16 ? n32 : n78572;
  assign n78574 = pi15 ? n78571 : n78573;
  assign n78575 = pi14 ? n78569 : n78574;
  assign n78576 = pi13 ? n78567 : n78575;
  assign n78577 = pi12 ? n78565 : n78576;
  assign n78578 = pi11 ? n78559 : n78577;
  assign n78579 = pi17 ? n3715 : ~n2726;
  assign n78580 = pi16 ? n32 : n78579;
  assign n78581 = pi15 ? n78573 : n78580;
  assign n78582 = pi17 ? n1028 : ~n2726;
  assign n78583 = pi16 ? n32 : n78582;
  assign n78584 = pi15 ? n78580 : n78583;
  assign n78585 = pi14 ? n78581 : n78584;
  assign n78586 = pi17 ? n3719 : ~n3182;
  assign n78587 = pi16 ? n32 : n78586;
  assign n78588 = pi17 ? n3719 : ~n2831;
  assign n78589 = pi16 ? n32 : n78588;
  assign n78590 = pi17 ? n3719 : ~n2733;
  assign n78591 = pi16 ? n32 : n78590;
  assign n78592 = pi15 ? n78589 : n78591;
  assign n78593 = pi14 ? n78587 : n78592;
  assign n78594 = pi13 ? n78585 : n78593;
  assign n78595 = pi17 ? n3557 : ~n2733;
  assign n78596 = pi16 ? n32 : n78595;
  assign n78597 = pi16 ? n3283 : ~n3061;
  assign n78598 = pi15 ? n78596 : n78597;
  assign n78599 = pi16 ? n32 : ~n2837;
  assign n78600 = pi16 ? n3283 : ~n2837;
  assign n78601 = pi15 ? n78599 : n78600;
  assign n78602 = pi14 ? n78598 : n78601;
  assign n78603 = pi16 ? n3283 : ~n2840;
  assign n78604 = pi15 ? n78599 : n78603;
  assign n78605 = pi16 ? n3729 : ~n2851;
  assign n78606 = pi15 ? n78603 : n78605;
  assign n78607 = pi14 ? n78604 : n78606;
  assign n78608 = pi13 ? n78602 : n78607;
  assign n78609 = pi12 ? n78594 : n78608;
  assign n78610 = pi16 ? n3438 : ~n3068;
  assign n78611 = pi16 ? n3438 : ~n4246;
  assign n78612 = pi15 ? n78610 : n78611;
  assign n78613 = pi16 ? n3156 : ~n2725;
  assign n78614 = pi14 ? n78612 : n78613;
  assign n78615 = pi16 ? n3156 : ~n2732;
  assign n78616 = pi16 ? n3570 : ~n2732;
  assign n78617 = pi15 ? n78615 : n78616;
  assign n78618 = pi16 ? n3156 : ~n2745;
  assign n78619 = pi16 ? n3570 : ~n2745;
  assign n78620 = pi15 ? n78618 : n78619;
  assign n78621 = pi14 ? n78617 : n78620;
  assign n78622 = pi13 ? n78614 : n78621;
  assign n78623 = pi16 ? n32 : ~n2617;
  assign n78624 = pi17 ? n3557 : ~n2855;
  assign n78625 = pi16 ? n32 : n78624;
  assign n78626 = pi14 ? n78623 : n78625;
  assign n78627 = pi17 ? n3557 : ~n2750;
  assign n78628 = pi16 ? n32 : n78627;
  assign n78629 = pi17 ? n3719 : ~n4099;
  assign n78630 = pi16 ? n32 : n78629;
  assign n78631 = pi15 ? n78628 : n78630;
  assign n78632 = pi17 ? n1028 : ~n2618;
  assign n78633 = pi16 ? n32 : n78632;
  assign n78634 = pi17 ? n1028 : ~n2628;
  assign n78635 = pi16 ? n32 : n78634;
  assign n78636 = pi15 ? n78633 : n78635;
  assign n78637 = pi14 ? n78631 : n78636;
  assign n78638 = pi13 ? n78626 : n78637;
  assign n78639 = pi12 ? n78622 : n78638;
  assign n78640 = pi11 ? n78609 : n78639;
  assign n78641 = pi10 ? n78578 : n78640;
  assign n78642 = pi09 ? n78537 : n78641;
  assign n78643 = pi08 ? n78527 : n78642;
  assign n78644 = pi17 ? n1833 : ~n3046;
  assign n78645 = pi16 ? n32 : n78644;
  assign n78646 = pi15 ? n32 : n78645;
  assign n78647 = pi17 ? n2143 : ~n3046;
  assign n78648 = pi16 ? n32 : n78647;
  assign n78649 = pi17 ? n1322 : ~n3046;
  assign n78650 = pi16 ? n32 : n78649;
  assign n78651 = pi15 ? n78648 : n78650;
  assign n78652 = pi14 ? n78646 : n78651;
  assign n78653 = pi13 ? n32 : n78652;
  assign n78654 = pi12 ? n32 : n78653;
  assign n78655 = pi11 ? n32 : n78654;
  assign n78656 = pi10 ? n32 : n78655;
  assign n78657 = pi17 ? n1971 : ~n3046;
  assign n78658 = pi16 ? n32 : n78657;
  assign n78659 = pi17 ? n1213 : ~n3046;
  assign n78660 = pi16 ? n32 : n78659;
  assign n78661 = pi15 ? n78660 : n78411;
  assign n78662 = pi14 ? n78658 : n78661;
  assign n78663 = pi17 ? n1232 : ~n3292;
  assign n78664 = pi16 ? n32 : n78663;
  assign n78665 = pi15 ? n78664 : n78540;
  assign n78666 = pi14 ? n78665 : n78540;
  assign n78667 = pi13 ? n78662 : n78666;
  assign n78668 = pi17 ? n1700 : ~n3292;
  assign n78669 = pi16 ? n32 : n78668;
  assign n78670 = pi17 ? n2159 : ~n3292;
  assign n78671 = pi16 ? n32 : n78670;
  assign n78672 = pi15 ? n78669 : n78671;
  assign n78673 = pi15 ? n78543 : n78311;
  assign n78674 = pi14 ? n78672 : n78673;
  assign n78675 = pi17 ? n1989 : ~n3292;
  assign n78676 = pi16 ? n32 : n78675;
  assign n78677 = pi15 ? n78311 : n78676;
  assign n78678 = pi17 ? n4682 : ~n3292;
  assign n78679 = pi16 ? n32 : n78678;
  assign n78680 = pi17 ? n4167 : ~n3292;
  assign n78681 = pi16 ? n32 : n78680;
  assign n78682 = pi15 ? n78679 : n78681;
  assign n78683 = pi14 ? n78677 : n78682;
  assign n78684 = pi13 ? n78674 : n78683;
  assign n78685 = pi12 ? n78667 : n78684;
  assign n78686 = pi15 ? n78681 : n78314;
  assign n78687 = pi17 ? n1215 : ~n2959;
  assign n78688 = pi16 ? n32 : n78687;
  assign n78689 = pi15 ? n78314 : n78688;
  assign n78690 = pi14 ? n78686 : n78689;
  assign n78691 = pi13 ? n78690 : n77997;
  assign n78692 = pi15 ? n78001 : n77583;
  assign n78693 = pi14 ? n78561 : n78692;
  assign n78694 = pi17 ? n4037 : ~n3175;
  assign n78695 = pi16 ? n32 : n78694;
  assign n78696 = pi17 ? n1605 : ~n3175;
  assign n78697 = pi16 ? n32 : n78696;
  assign n78698 = pi17 ? n3855 : ~n3175;
  assign n78699 = pi16 ? n32 : n78698;
  assign n78700 = pi15 ? n78697 : n78699;
  assign n78701 = pi14 ? n78695 : n78700;
  assign n78702 = pi13 ? n78693 : n78701;
  assign n78703 = pi12 ? n78691 : n78702;
  assign n78704 = pi11 ? n78685 : n78703;
  assign n78705 = pi17 ? n3553 : ~n2726;
  assign n78706 = pi16 ? n32 : n78705;
  assign n78707 = pi15 ? n78699 : n78706;
  assign n78708 = pi17 ? n1726 : ~n2726;
  assign n78709 = pi16 ? n32 : n78708;
  assign n78710 = pi15 ? n78706 : n78709;
  assign n78711 = pi14 ? n78707 : n78710;
  assign n78712 = pi17 ? n4041 : ~n2963;
  assign n78713 = pi16 ? n32 : n78712;
  assign n78714 = pi17 ? n4041 : ~n3182;
  assign n78715 = pi16 ? n32 : n78714;
  assign n78716 = pi15 ? n78713 : n78715;
  assign n78717 = pi17 ? n3704 : ~n3182;
  assign n78718 = pi16 ? n32 : n78717;
  assign n78719 = pi17 ? n3704 : ~n2831;
  assign n78720 = pi16 ? n32 : n78719;
  assign n78721 = pi15 ? n78718 : n78720;
  assign n78722 = pi14 ? n78716 : n78721;
  assign n78723 = pi13 ? n78711 : n78722;
  assign n78724 = pi17 ? n1028 : ~n2733;
  assign n78725 = pi16 ? n32 : n78724;
  assign n78726 = pi15 ? n78720 : n78725;
  assign n78727 = pi17 ? n2005 : ~n2836;
  assign n78728 = pi16 ? n32 : n78727;
  assign n78729 = pi17 ? n1028 : ~n2836;
  assign n78730 = pi16 ? n32 : n78729;
  assign n78731 = pi15 ? n78728 : n78730;
  assign n78732 = pi14 ? n78726 : n78731;
  assign n78733 = pi17 ? n1028 : ~n2839;
  assign n78734 = pi16 ? n32 : n78733;
  assign n78735 = pi15 ? n78728 : n78734;
  assign n78736 = pi17 ? n3557 : ~n2839;
  assign n78737 = pi16 ? n32 : n78736;
  assign n78738 = pi17 ? n3557 : ~n2850;
  assign n78739 = pi16 ? n32 : n78738;
  assign n78740 = pi15 ? n78737 : n78739;
  assign n78741 = pi14 ? n78735 : n78740;
  assign n78742 = pi13 ? n78732 : n78741;
  assign n78743 = pi12 ? n78723 : n78742;
  assign n78744 = pi17 ? n3557 : ~n3067;
  assign n78745 = pi16 ? n32 : n78744;
  assign n78746 = pi17 ? n3719 : ~n2724;
  assign n78747 = pi16 ? n32 : n78746;
  assign n78748 = pi17 ? n3715 : ~n2724;
  assign n78749 = pi16 ? n32 : n78748;
  assign n78750 = pi15 ? n78747 : n78749;
  assign n78751 = pi14 ? n78745 : n78750;
  assign n78752 = pi17 ? n3715 : ~n2731;
  assign n78753 = pi16 ? n32 : n78752;
  assign n78754 = pi17 ? n3715 : ~n2736;
  assign n78755 = pi16 ? n32 : n78754;
  assign n78756 = pi15 ? n78753 : n78755;
  assign n78757 = pi14 ? n78753 : n78756;
  assign n78758 = pi13 ? n78751 : n78757;
  assign n78759 = pi17 ? n3715 : ~n2616;
  assign n78760 = pi16 ? n32 : n78759;
  assign n78761 = pi15 ? n78755 : n78760;
  assign n78762 = pi17 ? n3704 : ~n2855;
  assign n78763 = pi16 ? n32 : n78762;
  assign n78764 = pi17 ? n4041 : ~n2855;
  assign n78765 = pi16 ? n32 : n78764;
  assign n78766 = pi15 ? n78763 : n78765;
  assign n78767 = pi14 ? n78761 : n78766;
  assign n78768 = pi17 ? n3704 : ~n2623;
  assign n78769 = pi16 ? n32 : n78768;
  assign n78770 = pi17 ? n4041 : ~n2750;
  assign n78771 = pi16 ? n32 : n78770;
  assign n78772 = pi15 ? n78769 : n78771;
  assign n78773 = pi17 ? n4041 : ~n4099;
  assign n78774 = pi16 ? n32 : n78773;
  assign n78775 = pi17 ? n1500 : ~n2618;
  assign n78776 = pi16 ? n32 : n78775;
  assign n78777 = pi15 ? n78774 : n78776;
  assign n78778 = pi14 ? n78772 : n78777;
  assign n78779 = pi13 ? n78767 : n78778;
  assign n78780 = pi12 ? n78758 : n78779;
  assign n78781 = pi11 ? n78743 : n78780;
  assign n78782 = pi10 ? n78704 : n78781;
  assign n78783 = pi09 ? n78656 : n78782;
  assign n78784 = pi17 ? n1943 : ~n3046;
  assign n78785 = pi16 ? n32 : n78784;
  assign n78786 = pi15 ? n32 : n78785;
  assign n78787 = pi17 ? n2325 : ~n3046;
  assign n78788 = pi16 ? n32 : n78787;
  assign n78789 = pi17 ? n1682 : ~n3046;
  assign n78790 = pi16 ? n32 : n78789;
  assign n78791 = pi15 ? n78788 : n78790;
  assign n78792 = pi14 ? n78786 : n78791;
  assign n78793 = pi13 ? n32 : n78792;
  assign n78794 = pi12 ? n32 : n78793;
  assign n78795 = pi11 ? n32 : n78794;
  assign n78796 = pi10 ? n32 : n78795;
  assign n78797 = pi17 ? n1842 : ~n3046;
  assign n78798 = pi16 ? n32 : n78797;
  assign n78799 = pi17 ? n1478 : ~n3292;
  assign n78800 = pi16 ? n32 : n78799;
  assign n78801 = pi15 ? n78798 : n78800;
  assign n78802 = pi14 ? n78650 : n78801;
  assign n78803 = pi17 ? n1478 : ~n3046;
  assign n78804 = pi16 ? n32 : n78803;
  assign n78805 = pi17 ? n1232 : ~n3046;
  assign n78806 = pi16 ? n32 : n78805;
  assign n78807 = pi15 ? n78804 : n78806;
  assign n78808 = pi17 ? n1966 : ~n3046;
  assign n78809 = pi16 ? n32 : n78808;
  assign n78810 = pi15 ? n78806 : n78809;
  assign n78811 = pi14 ? n78807 : n78810;
  assign n78812 = pi13 ? n78802 : n78811;
  assign n78813 = pi17 ? n4804 : ~n3046;
  assign n78814 = pi16 ? n32 : n78813;
  assign n78815 = pi17 ? n1706 : ~n3046;
  assign n78816 = pi16 ? n32 : n78815;
  assign n78817 = pi15 ? n78814 : n78816;
  assign n78818 = pi17 ? n4656 : ~n3046;
  assign n78819 = pi16 ? n32 : n78818;
  assign n78820 = pi15 ? n78819 : n78543;
  assign n78821 = pi14 ? n78817 : n78820;
  assign n78822 = pi15 ? n78543 : n78547;
  assign n78823 = pi15 ? n78549 : n78552;
  assign n78824 = pi14 ? n78822 : n78823;
  assign n78825 = pi13 ? n78821 : n78824;
  assign n78826 = pi12 ? n78812 : n78825;
  assign n78827 = pi15 ? n78552 : n78311;
  assign n78828 = pi15 ? n78311 : n77987;
  assign n78829 = pi14 ? n78827 : n78828;
  assign n78830 = pi13 ? n78829 : n77995;
  assign n78831 = pi17 ? n5541 : ~n2959;
  assign n78832 = pi16 ? n32 : n78831;
  assign n78833 = pi15 ? n78314 : n78832;
  assign n78834 = pi14 ? n78833 : n78832;
  assign n78835 = pi17 ? n5541 : ~n2952;
  assign n78836 = pi16 ? n32 : n78835;
  assign n78837 = pi17 ? n2355 : ~n3175;
  assign n78838 = pi16 ? n32 : n78837;
  assign n78839 = pi17 ? n1120 : ~n3175;
  assign n78840 = pi16 ? n32 : n78839;
  assign n78841 = pi15 ? n78838 : n78840;
  assign n78842 = pi14 ? n78836 : n78841;
  assign n78843 = pi13 ? n78834 : n78842;
  assign n78844 = pi12 ? n78830 : n78843;
  assign n78845 = pi11 ? n78826 : n78844;
  assign n78846 = pi17 ? n4034 : ~n3175;
  assign n78847 = pi16 ? n32 : n78846;
  assign n78848 = pi15 ? n78840 : n78847;
  assign n78849 = pi17 ? n4034 : ~n2726;
  assign n78850 = pi16 ? n32 : n78849;
  assign n78851 = pi17 ? n1219 : ~n2726;
  assign n78852 = pi16 ? n32 : n78851;
  assign n78853 = pi15 ? n78850 : n78852;
  assign n78854 = pi14 ? n78848 : n78853;
  assign n78855 = pi17 ? n4037 : ~n2726;
  assign n78856 = pi16 ? n32 : n78855;
  assign n78857 = pi17 ? n4037 : ~n2963;
  assign n78858 = pi16 ? n32 : n78857;
  assign n78859 = pi15 ? n78856 : n78858;
  assign n78860 = pi17 ? n3855 : ~n2963;
  assign n78861 = pi16 ? n32 : n78860;
  assign n78862 = pi17 ? n3855 : ~n3182;
  assign n78863 = pi16 ? n32 : n78862;
  assign n78864 = pi15 ? n78861 : n78863;
  assign n78865 = pi14 ? n78859 : n78864;
  assign n78866 = pi13 ? n78854 : n78865;
  assign n78867 = pi17 ? n3855 : ~n2831;
  assign n78868 = pi16 ? n32 : n78867;
  assign n78869 = pi17 ? n1726 : ~n2733;
  assign n78870 = pi16 ? n32 : n78869;
  assign n78871 = pi15 ? n78868 : n78870;
  assign n78872 = pi17 ? n1227 : ~n2733;
  assign n78873 = pi16 ? n32 : n78872;
  assign n78874 = pi15 ? n78873 : n78870;
  assign n78875 = pi14 ? n78871 : n78874;
  assign n78876 = pi17 ? n1726 : ~n2836;
  assign n78877 = pi16 ? n32 : n78876;
  assign n78878 = pi17 ? n1726 : ~n2839;
  assign n78879 = pi16 ? n32 : n78878;
  assign n78880 = pi15 ? n78877 : n78879;
  assign n78881 = pi17 ? n3715 : ~n2839;
  assign n78882 = pi16 ? n32 : n78881;
  assign n78883 = pi17 ? n3704 : ~n2839;
  assign n78884 = pi16 ? n32 : n78883;
  assign n78885 = pi15 ? n78882 : n78884;
  assign n78886 = pi14 ? n78880 : n78885;
  assign n78887 = pi13 ? n78875 : n78886;
  assign n78888 = pi12 ? n78866 : n78887;
  assign n78889 = pi17 ? n3704 : ~n2850;
  assign n78890 = pi16 ? n32 : n78889;
  assign n78891 = pi17 ? n4041 : ~n3067;
  assign n78892 = pi16 ? n32 : n78891;
  assign n78893 = pi14 ? n78890 : n78892;
  assign n78894 = pi17 ? n4041 : ~n2724;
  assign n78895 = pi16 ? n32 : n78894;
  assign n78896 = pi17 ? n4041 : ~n2731;
  assign n78897 = pi16 ? n32 : n78896;
  assign n78898 = pi15 ? n78895 : n78897;
  assign n78899 = pi17 ? n3553 : ~n2736;
  assign n78900 = pi16 ? n32 : n78899;
  assign n78901 = pi15 ? n78897 : n78900;
  assign n78902 = pi14 ? n78898 : n78901;
  assign n78903 = pi13 ? n78893 : n78902;
  assign n78904 = pi15 ? n78900 : n67410;
  assign n78905 = pi17 ? n3855 : ~n2616;
  assign n78906 = pi16 ? n32 : n78905;
  assign n78907 = pi17 ? n3855 : ~n2855;
  assign n78908 = pi16 ? n32 : n78907;
  assign n78909 = pi15 ? n78906 : n78908;
  assign n78910 = pi14 ? n78904 : n78909;
  assign n78911 = pi17 ? n4037 : ~n2750;
  assign n78912 = pi16 ? n32 : n78911;
  assign n78913 = pi15 ? n78908 : n78912;
  assign n78914 = pi17 ? n4037 : ~n4099;
  assign n78915 = pi16 ? n32 : n78914;
  assign n78916 = pi17 ? n1605 : ~n2618;
  assign n78917 = pi16 ? n32 : n78916;
  assign n78918 = pi15 ? n78915 : n78917;
  assign n78919 = pi14 ? n78913 : n78918;
  assign n78920 = pi13 ? n78910 : n78919;
  assign n78921 = pi12 ? n78903 : n78920;
  assign n78922 = pi11 ? n78888 : n78921;
  assign n78923 = pi10 ? n78845 : n78922;
  assign n78924 = pi09 ? n78796 : n78923;
  assign n78925 = pi08 ? n78783 : n78924;
  assign n78926 = pi07 ? n78643 : n78925;
  assign n78927 = pi17 ? n3337 : ~n3164;
  assign n78928 = pi16 ? n32 : n78927;
  assign n78929 = pi15 ? n32 : n78928;
  assign n78930 = pi17 ? n1814 : ~n3164;
  assign n78931 = pi16 ? n32 : n78930;
  assign n78932 = pi14 ? n78929 : n78931;
  assign n78933 = pi13 ? n32 : n78932;
  assign n78934 = pi12 ? n32 : n78933;
  assign n78935 = pi11 ? n32 : n78934;
  assign n78936 = pi10 ? n32 : n78935;
  assign n78937 = pi17 ? n1682 : ~n3164;
  assign n78938 = pi16 ? n32 : n78937;
  assign n78939 = pi17 ? n1576 : ~n3164;
  assign n78940 = pi16 ? n32 : n78939;
  assign n78941 = pi15 ? n78938 : n78940;
  assign n78942 = pi17 ? n2143 : ~n3164;
  assign n78943 = pi16 ? n32 : n78942;
  assign n78944 = pi17 ? n1580 : ~n3046;
  assign n78945 = pi16 ? n32 : n78944;
  assign n78946 = pi15 ? n78943 : n78945;
  assign n78947 = pi14 ? n78941 : n78946;
  assign n78948 = pi17 ? n1593 : ~n3046;
  assign n78949 = pi16 ? n32 : n78948;
  assign n78950 = pi15 ? n78949 : n78660;
  assign n78951 = pi14 ? n78950 : n78660;
  assign n78952 = pi13 ? n78947 : n78951;
  assign n78953 = pi17 ? n1134 : ~n3046;
  assign n78954 = pi16 ? n32 : n78953;
  assign n78955 = pi15 ? n78954 : n78806;
  assign n78956 = pi15 ? n78819 : n78540;
  assign n78957 = pi14 ? n78955 : n78956;
  assign n78958 = pi17 ? n1700 : ~n3046;
  assign n78959 = pi16 ? n32 : n78958;
  assign n78960 = pi15 ? n78540 : n78959;
  assign n78961 = pi17 ? n2159 : ~n3046;
  assign n78962 = pi16 ? n32 : n78961;
  assign n78963 = pi17 ? n4497 : ~n3046;
  assign n78964 = pi16 ? n32 : n78963;
  assign n78965 = pi15 ? n78962 : n78964;
  assign n78966 = pi14 ? n78960 : n78965;
  assign n78967 = pi13 ? n78957 : n78966;
  assign n78968 = pi12 ? n78952 : n78967;
  assign n78969 = pi15 ? n78964 : n78543;
  assign n78970 = pi17 ? n1472 : ~n3587;
  assign n78971 = pi16 ? n32 : n78970;
  assign n78972 = pi15 ? n78543 : n78971;
  assign n78973 = pi14 ? n78969 : n78972;
  assign n78974 = pi13 ? n78973 : n78199;
  assign n78975 = pi17 ? n5765 : ~n2959;
  assign n78976 = pi16 ? n32 : n78975;
  assign n78977 = pi15 ? n78311 : n78976;
  assign n78978 = pi14 ? n78977 : n78976;
  assign n78979 = pi17 ? n5765 : ~n3050;
  assign n78980 = pi16 ? n32 : n78979;
  assign n78981 = pi17 ? n5765 : ~n2952;
  assign n78982 = pi16 ? n32 : n78981;
  assign n78983 = pi15 ? n78980 : n78982;
  assign n78984 = pi17 ? n4515 : ~n2952;
  assign n78985 = pi16 ? n32 : n78984;
  assign n78986 = pi14 ? n78983 : n78985;
  assign n78987 = pi13 ? n78978 : n78986;
  assign n78988 = pi12 ? n78974 : n78987;
  assign n78989 = pi11 ? n78968 : n78988;
  assign n78990 = pi17 ? n4515 : ~n3175;
  assign n78991 = pi16 ? n32 : n78990;
  assign n78992 = pi15 ? n78985 : n78991;
  assign n78993 = pi17 ? n4515 : ~n2726;
  assign n78994 = pi16 ? n32 : n78993;
  assign n78995 = pi17 ? n2465 : ~n2726;
  assign n78996 = pi16 ? n32 : n78995;
  assign n78997 = pi15 ? n78994 : n78996;
  assign n78998 = pi14 ? n78992 : n78997;
  assign n78999 = pi17 ? n2355 : ~n2963;
  assign n79000 = pi16 ? n32 : n78999;
  assign n79001 = pi17 ? n4023 : ~n2963;
  assign n79002 = pi16 ? n32 : n79001;
  assign n79003 = pi17 ? n4023 : ~n3182;
  assign n79004 = pi16 ? n32 : n79003;
  assign n79005 = pi15 ? n79002 : n79004;
  assign n79006 = pi14 ? n79000 : n79005;
  assign n79007 = pi13 ? n78998 : n79006;
  assign n79008 = pi17 ? n4023 : ~n2831;
  assign n79009 = pi16 ? n32 : n79008;
  assign n79010 = pi17 ? n1219 : ~n2733;
  assign n79011 = pi16 ? n32 : n79010;
  assign n79012 = pi15 ? n79009 : n79011;
  assign n79013 = pi17 ? n1120 : ~n2733;
  assign n79014 = pi16 ? n32 : n79013;
  assign n79015 = pi15 ? n79014 : n79011;
  assign n79016 = pi14 ? n79012 : n79015;
  assign n79017 = pi17 ? n1219 : ~n2836;
  assign n79018 = pi16 ? n32 : n79017;
  assign n79019 = pi17 ? n1227 : ~n2836;
  assign n79020 = pi16 ? n32 : n79019;
  assign n79021 = pi17 ? n3855 : ~n2839;
  assign n79022 = pi16 ? n32 : n79021;
  assign n79023 = pi15 ? n79020 : n79022;
  assign n79024 = pi14 ? n79018 : n79023;
  assign n79025 = pi13 ? n79016 : n79024;
  assign n79026 = pi12 ? n79007 : n79025;
  assign n79027 = pi17 ? n3855 : ~n2850;
  assign n79028 = pi16 ? n32 : n79027;
  assign n79029 = pi15 ? n79022 : n79028;
  assign n79030 = pi17 ? n4037 : ~n3067;
  assign n79031 = pi16 ? n32 : n79030;
  assign n79032 = pi14 ? n79029 : n79031;
  assign n79033 = pi17 ? n4037 : ~n4245;
  assign n79034 = pi16 ? n32 : n79033;
  assign n79035 = pi17 ? n4037 : ~n2724;
  assign n79036 = pi16 ? n32 : n79035;
  assign n79037 = pi17 ? n4034 : ~n2731;
  assign n79038 = pi16 ? n32 : n79037;
  assign n79039 = pi15 ? n79036 : n79038;
  assign n79040 = pi14 ? n79034 : n79039;
  assign n79041 = pi13 ? n79032 : n79040;
  assign n79042 = pi17 ? n4034 : ~n2616;
  assign n79043 = pi16 ? n32 : n79042;
  assign n79044 = pi15 ? n79038 : n79043;
  assign n79045 = pi17 ? n4023 : ~n2855;
  assign n79046 = pi16 ? n32 : n79045;
  assign n79047 = pi14 ? n79044 : n79046;
  assign n79048 = pi17 ? n4023 : ~n2623;
  assign n79049 = pi16 ? n32 : n79048;
  assign n79050 = pi15 ? n79049 : n5838;
  assign n79051 = pi17 ? n5541 : ~n4099;
  assign n79052 = pi16 ? n32 : n79051;
  assign n79053 = pi17 ? n2355 : ~n2618;
  assign n79054 = pi16 ? n32 : n79053;
  assign n79055 = pi15 ? n79052 : n79054;
  assign n79056 = pi14 ? n79050 : n79055;
  assign n79057 = pi13 ? n79047 : n79056;
  assign n79058 = pi12 ? n79041 : n79057;
  assign n79059 = pi11 ? n79026 : n79058;
  assign n79060 = pi10 ? n78989 : n79059;
  assign n79061 = pi09 ? n78936 : n79060;
  assign n79062 = pi17 ? n2305 : ~n3164;
  assign n79063 = pi16 ? n32 : n79062;
  assign n79064 = pi15 ? n32 : n79063;
  assign n79065 = pi17 ? n1933 : ~n3164;
  assign n79066 = pi16 ? n32 : n79065;
  assign n79067 = pi15 ? n79066 : n78931;
  assign n79068 = pi14 ? n79064 : n79067;
  assign n79069 = pi13 ? n32 : n79068;
  assign n79070 = pi12 ? n32 : n79069;
  assign n79071 = pi11 ? n32 : n79070;
  assign n79072 = pi10 ? n32 : n79071;
  assign n79073 = pi17 ? n2136 : ~n3164;
  assign n79074 = pi16 ? n32 : n79073;
  assign n79075 = pi15 ? n78931 : n79074;
  assign n79076 = pi17 ? n2325 : ~n3164;
  assign n79077 = pi16 ? n32 : n79076;
  assign n79078 = pi17 ? n3351 : ~n3046;
  assign n79079 = pi16 ? n32 : n79078;
  assign n79080 = pi15 ? n79077 : n79079;
  assign n79081 = pi14 ? n79075 : n79080;
  assign n79082 = pi17 ? n1593 : ~n3164;
  assign n79083 = pi16 ? n32 : n79082;
  assign n79084 = pi15 ? n78940 : n79083;
  assign n79085 = pi17 ? n1842 : ~n3164;
  assign n79086 = pi16 ? n32 : n79085;
  assign n79087 = pi15 ? n79083 : n79086;
  assign n79088 = pi14 ? n79084 : n79087;
  assign n79089 = pi13 ? n79081 : n79088;
  assign n79090 = pi17 ? n1478 : ~n3164;
  assign n79091 = pi16 ? n32 : n79090;
  assign n79092 = pi17 ? n1232 : ~n3164;
  assign n79093 = pi16 ? n32 : n79092;
  assign n79094 = pi15 ? n79093 : n78806;
  assign n79095 = pi14 ? n79091 : n79094;
  assign n79096 = pi15 ? n78809 : n78814;
  assign n79097 = pi15 ? n78816 : n78819;
  assign n79098 = pi14 ? n79096 : n79097;
  assign n79099 = pi13 ? n79095 : n79098;
  assign n79100 = pi12 ? n79089 : n79099;
  assign n79101 = pi15 ? n78540 : n78189;
  assign n79102 = pi14 ? n78956 : n79101;
  assign n79103 = pi13 ? n79102 : n78197;
  assign n79104 = pi17 ? n5930 : ~n3587;
  assign n79105 = pi16 ? n32 : n79104;
  assign n79106 = pi15 ? n78543 : n79105;
  assign n79107 = pi17 ? n5930 : ~n2959;
  assign n79108 = pi16 ? n32 : n79107;
  assign n79109 = pi14 ? n79106 : n79108;
  assign n79110 = pi17 ? n5930 : ~n3050;
  assign n79111 = pi16 ? n32 : n79110;
  assign n79112 = pi17 ? n4682 : ~n3050;
  assign n79113 = pi16 ? n32 : n79112;
  assign n79114 = pi14 ? n79111 : n79113;
  assign n79115 = pi13 ? n79109 : n79114;
  assign n79116 = pi12 ? n79103 : n79115;
  assign n79117 = pi11 ? n79100 : n79116;
  assign n79118 = pi17 ? n4682 : ~n2952;
  assign n79119 = pi16 ? n32 : n79118;
  assign n79120 = pi17 ? n4682 : ~n3175;
  assign n79121 = pi16 ? n32 : n79120;
  assign n79122 = pi15 ? n79119 : n79121;
  assign n79123 = pi17 ? n4167 : ~n3175;
  assign n79124 = pi16 ? n32 : n79123;
  assign n79125 = pi15 ? n79121 : n79124;
  assign n79126 = pi14 ? n79122 : n79125;
  assign n79127 = pi17 ? n4167 : ~n2963;
  assign n79128 = pi16 ? n32 : n79127;
  assign n79129 = pi17 ? n4167 : ~n3182;
  assign n79130 = pi16 ? n32 : n79129;
  assign n79131 = pi15 ? n79128 : n79130;
  assign n79132 = pi14 ? n79128 : n79131;
  assign n79133 = pi13 ? n79126 : n79132;
  assign n79134 = pi17 ? n2465 : ~n3182;
  assign n79135 = pi16 ? n32 : n79134;
  assign n79136 = pi15 ? n79130 : n79135;
  assign n79137 = pi17 ? n4515 : ~n3182;
  assign n79138 = pi16 ? n32 : n79137;
  assign n79139 = pi15 ? n79138 : n79135;
  assign n79140 = pi14 ? n79136 : n79139;
  assign n79141 = pi17 ? n2465 : ~n2836;
  assign n79142 = pi16 ? n32 : n79141;
  assign n79143 = pi17 ? n1120 : ~n2836;
  assign n79144 = pi16 ? n32 : n79143;
  assign n79145 = pi17 ? n1120 : ~n2839;
  assign n79146 = pi16 ? n32 : n79145;
  assign n79147 = pi15 ? n79144 : n79146;
  assign n79148 = pi14 ? n79142 : n79147;
  assign n79149 = pi13 ? n79140 : n79148;
  assign n79150 = pi12 ? n79133 : n79149;
  assign n79151 = pi17 ? n4023 : ~n2839;
  assign n79152 = pi16 ? n32 : n79151;
  assign n79153 = pi17 ? n4023 : ~n2850;
  assign n79154 = pi16 ? n32 : n79153;
  assign n79155 = pi15 ? n79152 : n79154;
  assign n79156 = pi17 ? n5541 : ~n3067;
  assign n79157 = pi16 ? n32 : n79156;
  assign n79158 = pi14 ? n79155 : n79157;
  assign n79159 = pi17 ? n5541 : ~n4245;
  assign n79160 = pi16 ? n32 : n79159;
  assign n79161 = pi17 ? n5541 : ~n2724;
  assign n79162 = pi16 ? n32 : n79161;
  assign n79163 = pi17 ? n2465 : ~n2731;
  assign n79164 = pi16 ? n32 : n79163;
  assign n79165 = pi15 ? n79162 : n79164;
  assign n79166 = pi14 ? n79160 : n79165;
  assign n79167 = pi13 ? n79158 : n79166;
  assign n79168 = pi17 ? n4515 : ~n2731;
  assign n79169 = pi16 ? n32 : n79168;
  assign n79170 = pi17 ? n4515 : ~n2616;
  assign n79171 = pi16 ? n32 : n79170;
  assign n79172 = pi15 ? n79169 : n79171;
  assign n79173 = pi17 ? n4167 : ~n2855;
  assign n79174 = pi16 ? n32 : n79173;
  assign n79175 = pi14 ? n79172 : n79174;
  assign n79176 = pi17 ? n5765 : ~n4099;
  assign n79177 = pi16 ? n32 : n79176;
  assign n79178 = pi17 ? n2461 : ~n2618;
  assign n79179 = pi16 ? n32 : n79178;
  assign n79180 = pi15 ? n79177 : n79179;
  assign n79181 = pi14 ? n6005 : n79180;
  assign n79182 = pi13 ? n79175 : n79181;
  assign n79183 = pi12 ? n79167 : n79182;
  assign n79184 = pi11 ? n79150 : n79183;
  assign n79185 = pi10 ? n79117 : n79184;
  assign n79186 = pi09 ? n79072 : n79185;
  assign n79187 = pi08 ? n79061 : n79186;
  assign n79188 = pi17 ? n2531 : ~n3160;
  assign n79189 = pi16 ? n32 : n79188;
  assign n79190 = pi15 ? n32 : n79189;
  assign n79191 = pi17 ? n1933 : ~n3160;
  assign n79192 = pi16 ? n32 : n79191;
  assign n79193 = pi14 ? n79190 : n79192;
  assign n79194 = pi13 ? n32 : n79193;
  assign n79195 = pi12 ? n32 : n79194;
  assign n79196 = pi11 ? n32 : n79195;
  assign n79197 = pi10 ? n32 : n79196;
  assign n79198 = pi17 ? n2319 : ~n3160;
  assign n79199 = pi16 ? n32 : n79198;
  assign n79200 = pi17 ? n2537 : ~n3160;
  assign n79201 = pi16 ? n32 : n79200;
  assign n79202 = pi15 ? n79199 : n79201;
  assign n79203 = pi17 ? n1807 : ~n3160;
  assign n79204 = pi16 ? n32 : n79203;
  assign n79205 = pi15 ? n79204 : n79074;
  assign n79206 = pi14 ? n79202 : n79205;
  assign n79207 = pi15 ? n79074 : n78940;
  assign n79208 = pi17 ? n1833 : ~n3164;
  assign n79209 = pi16 ? n32 : n79208;
  assign n79210 = pi15 ? n79209 : n78943;
  assign n79211 = pi14 ? n79207 : n79210;
  assign n79212 = pi13 ? n79206 : n79211;
  assign n79213 = pi17 ? n1580 : ~n3164;
  assign n79214 = pi16 ? n32 : n79213;
  assign n79215 = pi15 ? n79214 : n79083;
  assign n79216 = pi17 ? n1213 : ~n3164;
  assign n79217 = pi16 ? n32 : n79216;
  assign n79218 = pi15 ? n79217 : n78660;
  assign n79219 = pi14 ? n79215 : n79218;
  assign n79220 = pi17 ? n1134 : ~n3164;
  assign n79221 = pi16 ? n32 : n79220;
  assign n79222 = pi15 ? n78660 : n79221;
  assign n79223 = pi14 ? n79222 : n79093;
  assign n79224 = pi13 ? n79219 : n79223;
  assign n79225 = pi12 ? n79212 : n79224;
  assign n79226 = pi15 ? n79093 : n78809;
  assign n79227 = pi14 ? n79226 : n79096;
  assign n79228 = pi13 ? n79227 : n78419;
  assign n79229 = pi17 ? n1978 : ~n3292;
  assign n79230 = pi16 ? n32 : n79229;
  assign n79231 = pi15 ? n79230 : n78189;
  assign n79232 = pi17 ? n4659 : ~n2959;
  assign n79233 = pi16 ? n32 : n79232;
  assign n79234 = pi14 ? n79231 : n79233;
  assign n79235 = pi17 ? n4659 : ~n3050;
  assign n79236 = pi16 ? n32 : n79235;
  assign n79237 = pi17 ? n4822 : ~n3050;
  assign n79238 = pi16 ? n32 : n79237;
  assign n79239 = pi14 ? n79236 : n79238;
  assign n79240 = pi13 ? n79234 : n79239;
  assign n79241 = pi12 ? n79228 : n79240;
  assign n79242 = pi11 ? n79225 : n79241;
  assign n79243 = pi17 ? n4822 : ~n2952;
  assign n79244 = pi16 ? n32 : n79243;
  assign n79245 = pi17 ? n4822 : ~n3175;
  assign n79246 = pi16 ? n32 : n79245;
  assign n79247 = pi15 ? n79244 : n79246;
  assign n79248 = pi17 ? n4341 : ~n3175;
  assign n79249 = pi16 ? n32 : n79248;
  assign n79250 = pi15 ? n79246 : n79249;
  assign n79251 = pi14 ? n79247 : n79250;
  assign n79252 = pi17 ? n4341 : ~n2726;
  assign n79253 = pi16 ? n32 : n79252;
  assign n79254 = pi17 ? n4341 : ~n2963;
  assign n79255 = pi16 ? n32 : n79254;
  assign n79256 = pi15 ? n79253 : n79255;
  assign n79257 = pi14 ? n79253 : n79256;
  assign n79258 = pi13 ? n79251 : n79257;
  assign n79259 = pi17 ? n1718 : ~n2963;
  assign n79260 = pi16 ? n32 : n79259;
  assign n79261 = pi17 ? n5765 : ~n3182;
  assign n79262 = pi16 ? n32 : n79261;
  assign n79263 = pi15 ? n79260 : n79262;
  assign n79264 = pi17 ? n1718 : ~n3182;
  assign n79265 = pi16 ? n32 : n79264;
  assign n79266 = pi15 ? n79265 : n79262;
  assign n79267 = pi14 ? n79263 : n79266;
  assign n79268 = pi17 ? n1718 : ~n2831;
  assign n79269 = pi16 ? n32 : n79268;
  assign n79270 = pi17 ? n1215 : ~n2733;
  assign n79271 = pi16 ? n32 : n79270;
  assign n79272 = pi17 ? n4167 : ~n2836;
  assign n79273 = pi16 ? n32 : n79272;
  assign n79274 = pi15 ? n79271 : n79273;
  assign n79275 = pi14 ? n79269 : n79274;
  assign n79276 = pi13 ? n79267 : n79275;
  assign n79277 = pi12 ? n79258 : n79276;
  assign n79278 = pi17 ? n4167 : ~n2850;
  assign n79279 = pi16 ? n32 : n79278;
  assign n79280 = pi15 ? n79273 : n79279;
  assign n79281 = pi17 ? n2461 : ~n3067;
  assign n79282 = pi16 ? n32 : n79281;
  assign n79283 = pi17 ? n5765 : ~n3067;
  assign n79284 = pi16 ? n32 : n79283;
  assign n79285 = pi15 ? n79282 : n79284;
  assign n79286 = pi14 ? n79280 : n79285;
  assign n79287 = pi17 ? n5765 : ~n4245;
  assign n79288 = pi16 ? n32 : n79287;
  assign n79289 = pi17 ? n5765 : ~n2724;
  assign n79290 = pi16 ? n32 : n79289;
  assign n79291 = pi17 ? n4682 : ~n2731;
  assign n79292 = pi16 ? n32 : n79291;
  assign n79293 = pi15 ? n79290 : n79292;
  assign n79294 = pi14 ? n79288 : n79293;
  assign n79295 = pi13 ? n79286 : n79294;
  assign n79296 = pi17 ? n4682 : ~n2616;
  assign n79297 = pi16 ? n32 : n79296;
  assign n79298 = pi15 ? n79292 : n79297;
  assign n79299 = pi17 ? n1989 : ~n2855;
  assign n79300 = pi16 ? n32 : n79299;
  assign n79301 = pi15 ? n79300 : n6257;
  assign n79302 = pi14 ? n79298 : n79301;
  assign n79303 = pi17 ? n5930 : ~n4099;
  assign n79304 = pi16 ? n32 : n79303;
  assign n79305 = pi17 ? n1480 : ~n2618;
  assign n79306 = pi16 ? n32 : n79305;
  assign n79307 = pi15 ? n79304 : n79306;
  assign n79308 = pi14 ? n6264 : n79307;
  assign n79309 = pi13 ? n79302 : n79308;
  assign n79310 = pi12 ? n79295 : n79309;
  assign n79311 = pi11 ? n79277 : n79310;
  assign n79312 = pi10 ? n79242 : n79311;
  assign n79313 = pi09 ? n79197 : n79312;
  assign n79314 = pi17 ? n2408 : ~n3160;
  assign n79315 = pi16 ? n32 : n79314;
  assign n79316 = pi15 ? n32 : n79315;
  assign n79317 = pi14 ? n79316 : n79189;
  assign n79318 = pi13 ? n32 : n79317;
  assign n79319 = pi12 ? n32 : n79318;
  assign n79320 = pi11 ? n32 : n79319;
  assign n79321 = pi10 ? n32 : n79320;
  assign n79322 = pi17 ? n2299 : ~n3160;
  assign n79323 = pi16 ? n32 : n79322;
  assign n79324 = pi17 ? n2410 : ~n3160;
  assign n79325 = pi16 ? n32 : n79324;
  assign n79326 = pi15 ? n79323 : n79325;
  assign n79327 = pi17 ? n2319 : ~n3164;
  assign n79328 = pi16 ? n32 : n79327;
  assign n79329 = pi15 ? n79192 : n79328;
  assign n79330 = pi14 ? n79326 : n79329;
  assign n79331 = pi17 ? n2136 : ~n3160;
  assign n79332 = pi16 ? n32 : n79331;
  assign n79333 = pi17 ? n1943 : ~n3160;
  assign n79334 = pi16 ? n32 : n79333;
  assign n79335 = pi17 ? n2325 : ~n3160;
  assign n79336 = pi16 ? n32 : n79335;
  assign n79337 = pi15 ? n79334 : n79336;
  assign n79338 = pi14 ? n79332 : n79337;
  assign n79339 = pi13 ? n79330 : n79338;
  assign n79340 = pi17 ? n3351 : ~n3160;
  assign n79341 = pi16 ? n32 : n79340;
  assign n79342 = pi17 ? n1576 : ~n3160;
  assign n79343 = pi16 ? n32 : n79342;
  assign n79344 = pi15 ? n79341 : n79343;
  assign n79345 = pi17 ? n1593 : ~n3160;
  assign n79346 = pi16 ? n32 : n79345;
  assign n79347 = pi15 ? n79346 : n79083;
  assign n79348 = pi14 ? n79344 : n79347;
  assign n79349 = pi15 ? n79086 : n79091;
  assign n79350 = pi15 ? n79091 : n79217;
  assign n79351 = pi14 ? n79349 : n79350;
  assign n79352 = pi13 ? n79348 : n79351;
  assign n79353 = pi12 ? n79339 : n79352;
  assign n79354 = pi17 ? n930 : ~n3046;
  assign n79355 = pi16 ? n32 : n79354;
  assign n79356 = pi15 ? n79355 : n78954;
  assign n79357 = pi14 ? n79218 : n79356;
  assign n79358 = pi17 ? n4798 : ~n3046;
  assign n79359 = pi16 ? n32 : n79358;
  assign n79360 = pi14 ? n78954 : n79359;
  assign n79361 = pi13 ? n79357 : n79360;
  assign n79362 = pi17 ? n1966 : ~n3292;
  assign n79363 = pi16 ? n32 : n79362;
  assign n79364 = pi15 ? n79363 : n78299;
  assign n79365 = pi14 ? n79364 : n78299;
  assign n79366 = pi17 ? n4804 : ~n3050;
  assign n79367 = pi16 ? n32 : n79366;
  assign n79368 = pi17 ? n1700 : ~n3050;
  assign n79369 = pi16 ? n32 : n79368;
  assign n79370 = pi15 ? n79367 : n79369;
  assign n79371 = pi17 ? n6439 : ~n3050;
  assign n79372 = pi16 ? n32 : n79371;
  assign n79373 = pi14 ? n79370 : n79372;
  assign n79374 = pi13 ? n79365 : n79373;
  assign n79375 = pi12 ? n79361 : n79374;
  assign n79376 = pi11 ? n79353 : n79375;
  assign n79377 = pi17 ? n6439 : ~n2959;
  assign n79378 = pi16 ? n32 : n79377;
  assign n79379 = pi15 ? n79378 : n79372;
  assign n79380 = pi17 ? n4497 : ~n3050;
  assign n79381 = pi16 ? n32 : n79380;
  assign n79382 = pi15 ? n79372 : n79381;
  assign n79383 = pi14 ? n79379 : n79382;
  assign n79384 = pi17 ? n4497 : ~n2726;
  assign n79385 = pi16 ? n32 : n79384;
  assign n79386 = pi17 ? n4497 : ~n2963;
  assign n79387 = pi16 ? n32 : n79386;
  assign n79388 = pi15 ? n79385 : n79387;
  assign n79389 = pi14 ? n79385 : n79388;
  assign n79390 = pi13 ? n79383 : n79389;
  assign n79391 = pi17 ? n1984 : ~n2963;
  assign n79392 = pi16 ? n32 : n79391;
  assign n79393 = pi17 ? n1984 : ~n3182;
  assign n79394 = pi16 ? n32 : n79393;
  assign n79395 = pi15 ? n79392 : n79394;
  assign n79396 = pi14 ? n79395 : n79394;
  assign n79397 = pi17 ? n1984 : ~n2831;
  assign n79398 = pi16 ? n32 : n79397;
  assign n79399 = pi17 ? n1989 : ~n2831;
  assign n79400 = pi16 ? n32 : n79399;
  assign n79401 = pi15 ? n79398 : n79400;
  assign n79402 = pi17 ? n1989 : ~n2733;
  assign n79403 = pi16 ? n32 : n79402;
  assign n79404 = pi17 ? n1989 : ~n2836;
  assign n79405 = pi16 ? n32 : n79404;
  assign n79406 = pi15 ? n79403 : n79405;
  assign n79407 = pi14 ? n79401 : n79406;
  assign n79408 = pi13 ? n79396 : n79407;
  assign n79409 = pi12 ? n79390 : n79408;
  assign n79410 = pi17 ? n4341 : ~n2836;
  assign n79411 = pi16 ? n32 : n79410;
  assign n79412 = pi17 ? n4341 : ~n2850;
  assign n79413 = pi16 ? n32 : n79412;
  assign n79414 = pi15 ? n79411 : n79413;
  assign n79415 = pi17 ? n5930 : ~n3067;
  assign n79416 = pi16 ? n32 : n79415;
  assign n79417 = pi14 ? n79414 : n79416;
  assign n79418 = pi17 ? n5930 : ~n4245;
  assign n79419 = pi16 ? n32 : n79418;
  assign n79420 = pi17 ? n5930 : ~n2724;
  assign n79421 = pi16 ? n32 : n79420;
  assign n79422 = pi17 ? n1984 : ~n2731;
  assign n79423 = pi16 ? n32 : n79422;
  assign n79424 = pi15 ? n79421 : n79423;
  assign n79425 = pi14 ? n79419 : n79424;
  assign n79426 = pi13 ? n79417 : n79425;
  assign n79427 = pi17 ? n4822 : ~n2731;
  assign n79428 = pi16 ? n32 : n79427;
  assign n79429 = pi17 ? n4822 : ~n2616;
  assign n79430 = pi16 ? n32 : n79429;
  assign n79431 = pi15 ? n79428 : n79430;
  assign n79432 = pi14 ? n79431 : n6497;
  assign n79433 = pi17 ? n4497 : ~n2623;
  assign n79434 = pi16 ? n32 : n79433;
  assign n79435 = pi17 ? n2159 : ~n2623;
  assign n79436 = pi16 ? n32 : n79435;
  assign n79437 = pi15 ? n79434 : n79436;
  assign n79438 = pi17 ? n4659 : ~n4099;
  assign n79439 = pi16 ? n32 : n79438;
  assign n79440 = pi17 ? n2159 : ~n2618;
  assign n79441 = pi16 ? n32 : n79440;
  assign n79442 = pi15 ? n79439 : n79441;
  assign n79443 = pi14 ? n79437 : n79442;
  assign n79444 = pi13 ? n79432 : n79443;
  assign n79445 = pi12 ? n79426 : n79444;
  assign n79446 = pi11 ? n79409 : n79445;
  assign n79447 = pi10 ? n79376 : n79446;
  assign n79448 = pi09 ? n79321 : n79447;
  assign n79449 = pi08 ? n79313 : n79448;
  assign n79450 = pi07 ? n79187 : n79449;
  assign n79451 = pi06 ? n78926 : n79450;
  assign n79452 = pi05 ? n78404 : n79451;
  assign n79453 = pi04 ? n77581 : n79452;
  assign n79454 = pi03 ? n76650 : n79453;
  assign n79455 = pi02 ? n75738 : n79454;
  assign n79456 = pi01 ? n32 : n79455;
  assign n79457 = pi17 ? n2414 : ~n4111;
  assign n79458 = pi16 ? n32 : n79457;
  assign n79459 = pi15 ? n32 : n79458;
  assign n79460 = pi17 ? n2119 : ~n4111;
  assign n79461 = pi16 ? n32 : n79460;
  assign n79462 = pi15 ? n79458 : n79461;
  assign n79463 = pi14 ? n79459 : n79462;
  assign n79464 = pi13 ? n32 : n79463;
  assign n79465 = pi12 ? n32 : n79464;
  assign n79466 = pi11 ? n32 : n79465;
  assign n79467 = pi10 ? n32 : n79466;
  assign n79468 = pi17 ? n2425 : ~n4111;
  assign n79469 = pi16 ? n32 : n79468;
  assign n79470 = pi17 ? n2531 : ~n4111;
  assign n79471 = pi16 ? n32 : n79470;
  assign n79472 = pi15 ? n79469 : n79471;
  assign n79473 = pi17 ? n2299 : ~n4111;
  assign n79474 = pi16 ? n32 : n79473;
  assign n79475 = pi15 ? n79474 : n79199;
  assign n79476 = pi14 ? n79472 : n79475;
  assign n79477 = pi17 ? n3337 : ~n3160;
  assign n79478 = pi16 ? n32 : n79477;
  assign n79479 = pi15 ? n79478 : n79204;
  assign n79480 = pi14 ? n79202 : n79479;
  assign n79481 = pi13 ? n79476 : n79480;
  assign n79482 = pi15 ? n79343 : n79209;
  assign n79483 = pi14 ? n79332 : n79482;
  assign n79484 = pi17 ? n1580 : ~n3160;
  assign n79485 = pi16 ? n32 : n79484;
  assign n79486 = pi15 ? n78943 : n79485;
  assign n79487 = pi14 ? n79486 : n79346;
  assign n79488 = pi13 ? n79483 : n79487;
  assign n79489 = pi12 ? n79481 : n79488;
  assign n79490 = pi15 ? n79346 : n79086;
  assign n79491 = pi17 ? n1470 : ~n3046;
  assign n79492 = pi16 ? n32 : n79491;
  assign n79493 = pi14 ? n79490 : n79492;
  assign n79494 = pi15 ? n78658 : n78660;
  assign n79495 = pi14 ? n78658 : n79494;
  assign n79496 = pi13 ? n79493 : n79495;
  assign n79497 = pi17 ? n930 : ~n3587;
  assign n79498 = pi16 ? n32 : n79497;
  assign n79499 = pi15 ? n78409 : n79498;
  assign n79500 = pi17 ? n1697 : ~n3587;
  assign n79501 = pi16 ? n32 : n79500;
  assign n79502 = pi15 ? n79498 : n79501;
  assign n79503 = pi14 ? n79499 : n79502;
  assign n79504 = pi17 ? n1697 : ~n2959;
  assign n79505 = pi16 ? n32 : n79504;
  assign n79506 = pi17 ? n4798 : ~n2959;
  assign n79507 = pi16 ? n32 : n79506;
  assign n79508 = pi14 ? n79505 : n79507;
  assign n79509 = pi13 ? n79503 : n79508;
  assign n79510 = pi12 ? n79496 : n79509;
  assign n79511 = pi11 ? n79489 : n79510;
  assign n79512 = pi17 ? n4798 : ~n3050;
  assign n79513 = pi16 ? n32 : n79512;
  assign n79514 = pi15 ? n79507 : n79513;
  assign n79515 = pi17 ? n1706 : ~n3050;
  assign n79516 = pi16 ? n32 : n79515;
  assign n79517 = pi17 ? n4656 : ~n3050;
  assign n79518 = pi16 ? n32 : n79517;
  assign n79519 = pi15 ? n79516 : n79518;
  assign n79520 = pi14 ? n79514 : n79519;
  assign n79521 = pi17 ? n4656 : ~n2952;
  assign n79522 = pi16 ? n32 : n79521;
  assign n79523 = pi17 ? n4656 : ~n3175;
  assign n79524 = pi16 ? n32 : n79523;
  assign n79525 = pi17 ? n4656 : ~n2726;
  assign n79526 = pi16 ? n32 : n79525;
  assign n79527 = pi15 ? n79524 : n79526;
  assign n79528 = pi14 ? n79522 : n79527;
  assign n79529 = pi13 ? n79520 : n79528;
  assign n79530 = pi17 ? n1978 : ~n2726;
  assign n79531 = pi16 ? n32 : n79530;
  assign n79532 = pi17 ? n4659 : ~n3182;
  assign n79533 = pi16 ? n32 : n79532;
  assign n79534 = pi15 ? n79531 : n79533;
  assign n79535 = pi17 ? n1978 : ~n3182;
  assign n79536 = pi16 ? n32 : n79535;
  assign n79537 = pi15 ? n79536 : n79533;
  assign n79538 = pi14 ? n79534 : n79537;
  assign n79539 = pi17 ? n1978 : ~n2831;
  assign n79540 = pi16 ? n32 : n79539;
  assign n79541 = pi17 ? n1472 : ~n2831;
  assign n79542 = pi16 ? n32 : n79541;
  assign n79543 = pi15 ? n79540 : n79542;
  assign n79544 = pi17 ? n4497 : ~n2836;
  assign n79545 = pi16 ? n32 : n79544;
  assign n79546 = pi15 ? n6682 : n79545;
  assign n79547 = pi14 ? n79543 : n79546;
  assign n79548 = pi13 ? n79538 : n79547;
  assign n79549 = pi12 ? n79529 : n79548;
  assign n79550 = pi17 ? n4497 : ~n2850;
  assign n79551 = pi16 ? n32 : n79550;
  assign n79552 = pi15 ? n79545 : n79551;
  assign n79553 = pi14 ? n79552 : n6701;
  assign n79554 = pi17 ? n2159 : ~n4245;
  assign n79555 = pi16 ? n32 : n79554;
  assign n79556 = pi17 ? n4659 : ~n4245;
  assign n79557 = pi16 ? n32 : n79556;
  assign n79558 = pi15 ? n79555 : n79557;
  assign n79559 = pi17 ? n4659 : ~n2724;
  assign n79560 = pi16 ? n32 : n79559;
  assign n79561 = pi17 ? n6439 : ~n2731;
  assign n79562 = pi16 ? n32 : n79561;
  assign n79563 = pi15 ? n79560 : n79562;
  assign n79564 = pi14 ? n79558 : n79563;
  assign n79565 = pi13 ? n79553 : n79564;
  assign n79566 = pi17 ? n6439 : ~n2616;
  assign n79567 = pi16 ? n32 : n79566;
  assign n79568 = pi15 ? n79562 : n79567;
  assign n79569 = pi17 ? n4656 : ~n2855;
  assign n79570 = pi16 ? n32 : n79569;
  assign n79571 = pi15 ? n6717 : n79570;
  assign n79572 = pi14 ? n79568 : n79571;
  assign n79573 = pi17 ? n4656 : ~n2623;
  assign n79574 = pi16 ? n32 : n79573;
  assign n79575 = pi17 ? n4804 : ~n2623;
  assign n79576 = pi16 ? n32 : n79575;
  assign n79577 = pi15 ? n79574 : n79576;
  assign n79578 = pi17 ? n4804 : ~n4099;
  assign n79579 = pi16 ? n32 : n79578;
  assign n79580 = pi17 ? n1706 : ~n2618;
  assign n79581 = pi16 ? n32 : n79580;
  assign n79582 = pi15 ? n79579 : n79581;
  assign n79583 = pi14 ? n79577 : n79582;
  assign n79584 = pi13 ? n79572 : n79583;
  assign n79585 = pi12 ? n79565 : n79584;
  assign n79586 = pi11 ? n79549 : n79585;
  assign n79587 = pi10 ? n79511 : n79586;
  assign n79588 = pi09 ? n79467 : n79587;
  assign n79589 = pi17 ? n2512 : ~n4111;
  assign n79590 = pi16 ? n32 : n79589;
  assign n79591 = pi15 ? n32 : n79590;
  assign n79592 = pi17 ? n2517 : ~n4111;
  assign n79593 = pi16 ? n32 : n79592;
  assign n79594 = pi15 ? n79590 : n79593;
  assign n79595 = pi14 ? n79591 : n79594;
  assign n79596 = pi13 ? n32 : n79595;
  assign n79597 = pi12 ? n32 : n79596;
  assign n79598 = pi11 ? n32 : n79597;
  assign n79599 = pi10 ? n32 : n79598;
  assign n79600 = pi17 ? n2755 : ~n4111;
  assign n79601 = pi16 ? n32 : n79600;
  assign n79602 = pi17 ? n2408 : ~n4111;
  assign n79603 = pi16 ? n32 : n79602;
  assign n79604 = pi15 ? n79601 : n79603;
  assign n79605 = pi15 ? n79458 : n79323;
  assign n79606 = pi14 ? n79604 : n79605;
  assign n79607 = pi17 ? n2410 : ~n4111;
  assign n79608 = pi16 ? n32 : n79607;
  assign n79609 = pi15 ? n79474 : n79608;
  assign n79610 = pi17 ? n2305 : ~n4111;
  assign n79611 = pi16 ? n32 : n79610;
  assign n79612 = pi17 ? n1933 : ~n4111;
  assign n79613 = pi16 ? n32 : n79612;
  assign n79614 = pi15 ? n79611 : n79613;
  assign n79615 = pi14 ? n79609 : n79614;
  assign n79616 = pi13 ? n79606 : n79615;
  assign n79617 = pi17 ? n2319 : ~n4111;
  assign n79618 = pi16 ? n32 : n79617;
  assign n79619 = pi17 ? n2136 : ~n4111;
  assign n79620 = pi16 ? n32 : n79619;
  assign n79621 = pi15 ? n79618 : n79620;
  assign n79622 = pi17 ? n1943 : ~n4111;
  assign n79623 = pi16 ? n32 : n79622;
  assign n79624 = pi15 ? n79620 : n79623;
  assign n79625 = pi14 ? n79621 : n79624;
  assign n79626 = pi15 ? n79336 : n79341;
  assign n79627 = pi14 ? n79626 : n79343;
  assign n79628 = pi13 ? n79625 : n79627;
  assign n79629 = pi12 ? n79616 : n79628;
  assign n79630 = pi14 ? n79482 : n78648;
  assign n79631 = pi17 ? n1322 : ~n3164;
  assign n79632 = pi16 ? n32 : n79631;
  assign n79633 = pi15 ? n79632 : n79083;
  assign n79634 = pi14 ? n78650 : n79633;
  assign n79635 = pi13 ? n79630 : n79634;
  assign n79636 = pi15 ? n79086 : n78798;
  assign n79637 = pi17 ? n1704 : ~n3046;
  assign n79638 = pi16 ? n32 : n79637;
  assign n79639 = pi14 ? n79636 : n79638;
  assign n79640 = pi17 ? n1704 : ~n2959;
  assign n79641 = pi16 ? n32 : n79640;
  assign n79642 = pi17 ? n1971 : ~n2959;
  assign n79643 = pi16 ? n32 : n79642;
  assign n79644 = pi15 ? n79641 : n79643;
  assign n79645 = pi14 ? n79644 : n79643;
  assign n79646 = pi13 ? n79639 : n79645;
  assign n79647 = pi12 ? n79635 : n79646;
  assign n79648 = pi11 ? n79629 : n79647;
  assign n79649 = pi17 ? n1134 : ~n3050;
  assign n79650 = pi16 ? n32 : n79649;
  assign n79651 = pi15 ? n79643 : n79650;
  assign n79652 = pi17 ? n1232 : ~n3050;
  assign n79653 = pi16 ? n32 : n79652;
  assign n79654 = pi15 ? n79650 : n79653;
  assign n79655 = pi14 ? n79651 : n79654;
  assign n79656 = pi17 ? n1232 : ~n2952;
  assign n79657 = pi16 ? n32 : n79656;
  assign n79658 = pi17 ? n1232 : ~n3175;
  assign n79659 = pi16 ? n32 : n79658;
  assign n79660 = pi17 ? n1966 : ~n2726;
  assign n79661 = pi16 ? n32 : n79660;
  assign n79662 = pi15 ? n79659 : n79661;
  assign n79663 = pi14 ? n79657 : n79662;
  assign n79664 = pi13 ? n79655 : n79663;
  assign n79665 = pi17 ? n1966 : ~n3182;
  assign n79666 = pi16 ? n32 : n79665;
  assign n79667 = pi15 ? n79661 : n79666;
  assign n79668 = pi14 ? n79667 : n79666;
  assign n79669 = pi17 ? n1966 : ~n2831;
  assign n79670 = pi16 ? n32 : n79669;
  assign n79671 = pi17 ? n1700 : ~n2831;
  assign n79672 = pi16 ? n32 : n79671;
  assign n79673 = pi15 ? n79670 : n79672;
  assign n79674 = pi17 ? n1700 : ~n2836;
  assign n79675 = pi16 ? n32 : n79674;
  assign n79676 = pi15 ? n6877 : n79675;
  assign n79677 = pi14 ? n79673 : n79676;
  assign n79678 = pi13 ? n79668 : n79677;
  assign n79679 = pi12 ? n79664 : n79678;
  assign n79680 = pi17 ? n4656 : ~n2836;
  assign n79681 = pi16 ? n32 : n79680;
  assign n79682 = pi17 ? n4656 : ~n2850;
  assign n79683 = pi16 ? n32 : n79682;
  assign n79684 = pi15 ? n79681 : n79683;
  assign n79685 = pi14 ? n79684 : n6894;
  assign n79686 = pi17 ? n4804 : ~n4245;
  assign n79687 = pi16 ? n32 : n79686;
  assign n79688 = pi17 ? n4804 : ~n2724;
  assign n79689 = pi16 ? n32 : n79688;
  assign n79690 = pi17 ? n1966 : ~n2731;
  assign n79691 = pi16 ? n32 : n79690;
  assign n79692 = pi15 ? n79689 : n79691;
  assign n79693 = pi14 ? n79687 : n79692;
  assign n79694 = pi13 ? n79685 : n79693;
  assign n79695 = pi17 ? n4798 : ~n2616;
  assign n79696 = pi16 ? n32 : n79695;
  assign n79697 = pi15 ? n6912 : n79696;
  assign n79698 = pi17 ? n1232 : ~n2623;
  assign n79699 = pi16 ? n32 : n79698;
  assign n79700 = pi15 ? n6917 : n79699;
  assign n79701 = pi14 ? n79697 : n79700;
  assign n79702 = pi17 ? n1134 : ~n2750;
  assign n79703 = pi16 ? n32 : n79702;
  assign n79704 = pi15 ? n79699 : n79703;
  assign n79705 = pi17 ? n930 : ~n4099;
  assign n79706 = pi16 ? n32 : n79705;
  assign n79707 = pi17 ? n1134 : ~n2618;
  assign n79708 = pi16 ? n32 : n79707;
  assign n79709 = pi15 ? n79706 : n79708;
  assign n79710 = pi14 ? n79704 : n79709;
  assign n79711 = pi13 ? n79701 : n79710;
  assign n79712 = pi12 ? n79694 : n79711;
  assign n79713 = pi11 ? n79679 : n79712;
  assign n79714 = pi10 ? n79648 : n79713;
  assign n79715 = pi09 ? n79599 : n79714;
  assign n79716 = pi08 ? n79588 : n79715;
  assign n79717 = pi17 ? n2623 : ~n3728;
  assign n79718 = pi16 ? n32 : n79717;
  assign n79719 = pi15 ? n32 : n79718;
  assign n79720 = pi17 ? n4099 : ~n3728;
  assign n79721 = pi16 ? n32 : n79720;
  assign n79722 = pi15 ? n79718 : n79721;
  assign n79723 = pi14 ? n79719 : n79722;
  assign n79724 = pi13 ? n32 : n79723;
  assign n79725 = pi12 ? n32 : n79724;
  assign n79726 = pi11 ? n32 : n79725;
  assign n79727 = pi10 ? n32 : n79726;
  assign n79728 = pi17 ? n2618 : ~n3728;
  assign n79729 = pi16 ? n32 : n79728;
  assign n79730 = pi17 ? n2512 : ~n3728;
  assign n79731 = pi16 ? n32 : n79730;
  assign n79732 = pi15 ? n79729 : n79731;
  assign n79733 = pi17 ? n2748 : ~n3728;
  assign n79734 = pi16 ? n32 : n79733;
  assign n79735 = pi15 ? n79734 : n79461;
  assign n79736 = pi14 ? n79732 : n79735;
  assign n79737 = pi15 ? n79461 : n79469;
  assign n79738 = pi17 ? n2653 : ~n4111;
  assign n79739 = pi16 ? n32 : n79738;
  assign n79740 = pi15 ? n79739 : n79474;
  assign n79741 = pi14 ? n79737 : n79740;
  assign n79742 = pi13 ? n79736 : n79741;
  assign n79743 = pi15 ? n79474 : n79618;
  assign n79744 = pi17 ? n2537 : ~n4111;
  assign n79745 = pi16 ? n32 : n79744;
  assign n79746 = pi15 ? n79618 : n79745;
  assign n79747 = pi14 ? n79743 : n79746;
  assign n79748 = pi17 ? n3337 : ~n4111;
  assign n79749 = pi16 ? n32 : n79748;
  assign n79750 = pi17 ? n1807 : ~n4111;
  assign n79751 = pi16 ? n32 : n79750;
  assign n79752 = pi15 ? n79749 : n79751;
  assign n79753 = pi14 ? n79752 : n79620;
  assign n79754 = pi13 ? n79747 : n79753;
  assign n79755 = pi12 ? n79742 : n79754;
  assign n79756 = pi17 ? n1943 : ~n3164;
  assign n79757 = pi16 ? n32 : n79756;
  assign n79758 = pi15 ? n79620 : n79757;
  assign n79759 = pi14 ? n79758 : n79077;
  assign n79760 = pi14 ? n78938 : n78941;
  assign n79761 = pi13 ? n79759 : n79760;
  assign n79762 = pi15 ? n79209 : n78645;
  assign n79763 = pi14 ? n79762 : n78945;
  assign n79764 = pi17 ? n1580 : ~n3292;
  assign n79765 = pi16 ? n32 : n79764;
  assign n79766 = pi17 ? n1322 : ~n3292;
  assign n79767 = pi16 ? n32 : n79766;
  assign n79768 = pi15 ? n79765 : n79767;
  assign n79769 = pi17 ? n1322 : ~n3587;
  assign n79770 = pi16 ? n32 : n79769;
  assign n79771 = pi15 ? n79767 : n79770;
  assign n79772 = pi14 ? n79768 : n79771;
  assign n79773 = pi13 ? n79763 : n79772;
  assign n79774 = pi12 ? n79761 : n79773;
  assign n79775 = pi11 ? n79755 : n79774;
  assign n79776 = pi17 ? n1470 : ~n3587;
  assign n79777 = pi16 ? n32 : n79776;
  assign n79778 = pi17 ? n1470 : ~n3050;
  assign n79779 = pi16 ? n32 : n79778;
  assign n79780 = pi17 ? n1478 : ~n3050;
  assign n79781 = pi16 ? n32 : n79780;
  assign n79782 = pi15 ? n79779 : n79781;
  assign n79783 = pi14 ? n79777 : n79782;
  assign n79784 = pi17 ? n1478 : ~n2952;
  assign n79785 = pi16 ? n32 : n79784;
  assign n79786 = pi17 ? n1213 : ~n2726;
  assign n79787 = pi16 ? n32 : n79786;
  assign n79788 = pi15 ? n79785 : n79787;
  assign n79789 = pi14 ? n79785 : n79788;
  assign n79790 = pi13 ? n79783 : n79789;
  assign n79791 = pi17 ? n1213 : ~n3182;
  assign n79792 = pi16 ? n32 : n79791;
  assign n79793 = pi14 ? n79787 : n79792;
  assign n79794 = pi17 ? n1213 : ~n2831;
  assign n79795 = pi16 ? n32 : n79794;
  assign n79796 = pi17 ? n1697 : ~n2831;
  assign n79797 = pi16 ? n32 : n79796;
  assign n79798 = pi15 ? n79795 : n79797;
  assign n79799 = pi17 ? n1232 : ~n2836;
  assign n79800 = pi16 ? n32 : n79799;
  assign n79801 = pi15 ? n7054 : n79800;
  assign n79802 = pi14 ? n79798 : n79801;
  assign n79803 = pi13 ? n79793 : n79802;
  assign n79804 = pi12 ? n79790 : n79803;
  assign n79805 = pi15 ? n79800 : n7066;
  assign n79806 = pi15 ? n6841 : n6611;
  assign n79807 = pi14 ? n79805 : n79806;
  assign n79808 = pi17 ? n1134 : ~n4245;
  assign n79809 = pi16 ? n32 : n79808;
  assign n79810 = pi15 ? n79809 : n7075;
  assign n79811 = pi17 ? n930 : ~n2724;
  assign n79812 = pi16 ? n32 : n79811;
  assign n79813 = pi15 ? n79812 : n7083;
  assign n79814 = pi14 ? n79810 : n79813;
  assign n79815 = pi13 ? n79807 : n79814;
  assign n79816 = pi17 ? n1971 : ~n2616;
  assign n79817 = pi16 ? n32 : n79816;
  assign n79818 = pi15 ? n7083 : n79817;
  assign n79819 = pi17 ? n1478 : ~n2623;
  assign n79820 = pi16 ? n32 : n79819;
  assign n79821 = pi15 ? n7088 : n79820;
  assign n79822 = pi14 ? n79818 : n79821;
  assign n79823 = pi17 ? n1842 : ~n2750;
  assign n79824 = pi16 ? n32 : n79823;
  assign n79825 = pi15 ? n79820 : n79824;
  assign n79826 = pi17 ? n1842 : ~n4099;
  assign n79827 = pi16 ? n32 : n79826;
  assign n79828 = pi15 ? n79827 : n7115;
  assign n79829 = pi14 ? n79825 : n79828;
  assign n79830 = pi13 ? n79822 : n79829;
  assign n79831 = pi12 ? n79815 : n79830;
  assign n79832 = pi11 ? n79804 : n79831;
  assign n79833 = pi10 ? n79775 : n79832;
  assign n79834 = pi09 ? n79727 : n79833;
  assign n79835 = pi17 ? n3067 : ~n3728;
  assign n79836 = pi16 ? n32 : n79835;
  assign n79837 = pi15 ? n32 : n79836;
  assign n79838 = pi17 ? n4245 : ~n3728;
  assign n79839 = pi16 ? n32 : n79838;
  assign n79840 = pi17 ? n2724 : ~n3728;
  assign n79841 = pi16 ? n32 : n79840;
  assign n79842 = pi15 ? n79839 : n79841;
  assign n79843 = pi14 ? n79837 : n79842;
  assign n79844 = pi13 ? n32 : n79843;
  assign n79845 = pi12 ? n32 : n79844;
  assign n79846 = pi11 ? n32 : n79845;
  assign n79847 = pi10 ? n32 : n79846;
  assign n79848 = pi17 ? n2731 : ~n3728;
  assign n79849 = pi16 ? n32 : n79848;
  assign n79850 = pi15 ? n79849 : n79718;
  assign n79851 = pi17 ? n2750 : ~n3728;
  assign n79852 = pi16 ? n32 : n79851;
  assign n79853 = pi17 ? n2748 : ~n4111;
  assign n79854 = pi16 ? n32 : n79853;
  assign n79855 = pi15 ? n79852 : n79854;
  assign n79856 = pi14 ? n79850 : n79855;
  assign n79857 = pi17 ? n2755 : ~n3728;
  assign n79858 = pi16 ? n32 : n79857;
  assign n79859 = pi15 ? n79734 : n79858;
  assign n79860 = pi17 ? n2519 : ~n3728;
  assign n79861 = pi16 ? n32 : n79860;
  assign n79862 = pi17 ? n2414 : ~n3728;
  assign n79863 = pi16 ? n32 : n79862;
  assign n79864 = pi15 ? n79861 : n79863;
  assign n79865 = pi14 ? n79859 : n79864;
  assign n79866 = pi13 ? n79856 : n79865;
  assign n79867 = pi17 ? n2299 : ~n3728;
  assign n79868 = pi16 ? n32 : n79867;
  assign n79869 = pi15 ? n79863 : n79868;
  assign n79870 = pi14 ? n79869 : n79609;
  assign n79871 = pi14 ? n79614 : n79618;
  assign n79872 = pi13 ? n79870 : n79871;
  assign n79873 = pi12 ? n79866 : n79872;
  assign n79874 = pi17 ? n2537 : ~n3164;
  assign n79875 = pi16 ? n32 : n79874;
  assign n79876 = pi15 ? n79199 : n79875;
  assign n79877 = pi14 ? n79876 : n78928;
  assign n79878 = pi14 ? n78931 : n79075;
  assign n79879 = pi13 ? n79877 : n79878;
  assign n79880 = pi15 ? n79757 : n78785;
  assign n79881 = pi17 ? n1677 : ~n3046;
  assign n79882 = pi16 ? n32 : n79881;
  assign n79883 = pi14 ? n79880 : n79882;
  assign n79884 = pi17 ? n1677 : ~n3292;
  assign n79885 = pi16 ? n32 : n79884;
  assign n79886 = pi17 ? n1682 : ~n3292;
  assign n79887 = pi16 ? n32 : n79886;
  assign n79888 = pi15 ? n79885 : n79887;
  assign n79889 = pi17 ? n1682 : ~n3587;
  assign n79890 = pi16 ? n32 : n79889;
  assign n79891 = pi14 ? n79888 : n79890;
  assign n79892 = pi13 ? n79883 : n79891;
  assign n79893 = pi12 ? n79879 : n79892;
  assign n79894 = pi11 ? n79873 : n79893;
  assign n79895 = pi17 ? n1833 : ~n3587;
  assign n79896 = pi16 ? n32 : n79895;
  assign n79897 = pi17 ? n1833 : ~n3050;
  assign n79898 = pi16 ? n32 : n79897;
  assign n79899 = pi15 ? n79896 : n79898;
  assign n79900 = pi17 ? n2143 : ~n3050;
  assign n79901 = pi16 ? n32 : n79900;
  assign n79902 = pi15 ? n79898 : n79901;
  assign n79903 = pi14 ? n79899 : n79902;
  assign n79904 = pi17 ? n2143 : ~n2952;
  assign n79905 = pi16 ? n32 : n79904;
  assign n79906 = pi17 ? n1593 : ~n3175;
  assign n79907 = pi16 ? n32 : n79906;
  assign n79908 = pi17 ? n1593 : ~n2726;
  assign n79909 = pi16 ? n32 : n79908;
  assign n79910 = pi15 ? n79907 : n79909;
  assign n79911 = pi14 ? n79905 : n79910;
  assign n79912 = pi13 ? n79903 : n79911;
  assign n79913 = pi17 ? n1593 : ~n3182;
  assign n79914 = pi16 ? n32 : n79913;
  assign n79915 = pi15 ? n79909 : n79914;
  assign n79916 = pi14 ? n79915 : n79914;
  assign n79917 = pi17 ? n1593 : ~n2831;
  assign n79918 = pi16 ? n32 : n79917;
  assign n79919 = pi17 ? n1704 : ~n2831;
  assign n79920 = pi16 ? n32 : n79919;
  assign n79921 = pi15 ? n79918 : n79920;
  assign n79922 = pi17 ? n1704 : ~n2836;
  assign n79923 = pi16 ? n32 : n79922;
  assign n79924 = pi15 ? n7239 : n79923;
  assign n79925 = pi14 ? n79921 : n79924;
  assign n79926 = pi13 ? n79916 : n79925;
  assign n79927 = pi12 ? n79912 : n79926;
  assign n79928 = pi15 ? n7245 : n7022;
  assign n79929 = pi17 ? n1842 : ~n4245;
  assign n79930 = pi16 ? n32 : n79929;
  assign n79931 = pi15 ? n6812 : n79930;
  assign n79932 = pi14 ? n79928 : n79931;
  assign n79933 = pi15 ? n79930 : n7252;
  assign n79934 = pi17 ? n1593 : ~n2724;
  assign n79935 = pi16 ? n32 : n79934;
  assign n79936 = pi15 ? n79935 : n7261;
  assign n79937 = pi14 ? n79933 : n79936;
  assign n79938 = pi13 ? n79932 : n79937;
  assign n79939 = pi17 ? n1322 : ~n2616;
  assign n79940 = pi16 ? n32 : n79939;
  assign n79941 = pi17 ? n2143 : ~n2623;
  assign n79942 = pi16 ? n32 : n79941;
  assign n79943 = pi15 ? n7271 : n79942;
  assign n79944 = pi14 ? n79940 : n79943;
  assign n79945 = pi17 ? n1833 : ~n2623;
  assign n79946 = pi16 ? n32 : n79945;
  assign n79947 = pi17 ? n1833 : ~n2750;
  assign n79948 = pi16 ? n32 : n79947;
  assign n79949 = pi15 ? n79946 : n79948;
  assign n79950 = pi17 ? n1576 : ~n4099;
  assign n79951 = pi16 ? n32 : n79950;
  assign n79952 = pi15 ? n79951 : n7289;
  assign n79953 = pi14 ? n79949 : n79952;
  assign n79954 = pi13 ? n79944 : n79953;
  assign n79955 = pi12 ? n79938 : n79954;
  assign n79956 = pi11 ? n79927 : n79955;
  assign n79957 = pi10 ? n79894 : n79956;
  assign n79958 = pi09 ? n79847 : n79957;
  assign n79959 = pi08 ? n79834 : n79958;
  assign n79960 = pi07 ? n79716 : n79959;
  assign n79961 = pi17 ? n2733 : ~n2954;
  assign n79962 = pi16 ? n32 : n79961;
  assign n79963 = pi15 ? n32 : n79962;
  assign n79964 = pi17 ? n2836 : ~n2954;
  assign n79965 = pi16 ? n32 : n79964;
  assign n79966 = pi15 ? n79962 : n79965;
  assign n79967 = pi14 ? n79963 : n79966;
  assign n79968 = pi13 ? n32 : n79967;
  assign n79969 = pi12 ? n32 : n79968;
  assign n79970 = pi11 ? n32 : n79969;
  assign n79971 = pi10 ? n32 : n79970;
  assign n79972 = pi17 ? n2839 : ~n2954;
  assign n79973 = pi16 ? n32 : n79972;
  assign n79974 = pi17 ? n3067 : ~n2954;
  assign n79975 = pi16 ? n32 : n79974;
  assign n79976 = pi15 ? n79973 : n79975;
  assign n79977 = pi17 ? n2750 : ~n2954;
  assign n79978 = pi16 ? n32 : n79977;
  assign n79979 = pi14 ? n79976 : n79978;
  assign n79980 = pi15 ? n79852 : n79729;
  assign n79981 = pi17 ? n2628 : ~n3728;
  assign n79982 = pi16 ? n32 : n79981;
  assign n79983 = pi15 ? n79982 : n79734;
  assign n79984 = pi14 ? n79980 : n79983;
  assign n79985 = pi13 ? n79979 : n79984;
  assign n79986 = pi17 ? n2119 : ~n3728;
  assign n79987 = pi16 ? n32 : n79986;
  assign n79988 = pi15 ? n79734 : n79987;
  assign n79989 = pi14 ? n79988 : n79737;
  assign n79990 = pi17 ? n2653 : ~n3728;
  assign n79991 = pi16 ? n32 : n79990;
  assign n79992 = pi15 ? n79991 : n79868;
  assign n79993 = pi14 ? n79992 : n79868;
  assign n79994 = pi13 ? n79989 : n79993;
  assign n79995 = pi12 ? n79985 : n79994;
  assign n79996 = pi15 ? n79868 : n79608;
  assign n79997 = pi14 ? n79996 : n79611;
  assign n79998 = pi15 ? n79613 : n79199;
  assign n79999 = pi14 ? n79613 : n79998;
  assign n80000 = pi13 ? n79997 : n79999;
  assign n80001 = pi17 ? n1807 : ~n3046;
  assign n80002 = pi16 ? n32 : n80001;
  assign n80003 = pi14 ? n79201 : n80002;
  assign n80004 = pi17 ? n1807 : ~n3292;
  assign n80005 = pi16 ? n32 : n80004;
  assign n80006 = pi17 ? n1814 : ~n3292;
  assign n80007 = pi16 ? n32 : n80006;
  assign n80008 = pi15 ? n80005 : n80007;
  assign n80009 = pi17 ? n1814 : ~n3587;
  assign n80010 = pi16 ? n32 : n80009;
  assign n80011 = pi15 ? n80007 : n80010;
  assign n80012 = pi14 ? n80008 : n80011;
  assign n80013 = pi13 ? n80003 : n80012;
  assign n80014 = pi12 ? n80000 : n80013;
  assign n80015 = pi11 ? n79995 : n80014;
  assign n80016 = pi17 ? n3351 : ~n3587;
  assign n80017 = pi16 ? n32 : n80016;
  assign n80018 = pi17 ? n3351 : ~n3050;
  assign n80019 = pi16 ? n32 : n80018;
  assign n80020 = pi17 ? n2123 : ~n3050;
  assign n80021 = pi16 ? n32 : n80020;
  assign n80022 = pi15 ? n80019 : n80021;
  assign n80023 = pi14 ? n80017 : n80022;
  assign n80024 = pi17 ? n2123 : ~n2952;
  assign n80025 = pi16 ? n32 : n80024;
  assign n80026 = pi17 ? n1682 : ~n2952;
  assign n80027 = pi16 ? n32 : n80026;
  assign n80028 = pi17 ? n1682 : ~n2726;
  assign n80029 = pi16 ? n32 : n80028;
  assign n80030 = pi15 ? n80027 : n80029;
  assign n80031 = pi14 ? n80025 : n80030;
  assign n80032 = pi13 ? n80023 : n80031;
  assign n80033 = pi17 ? n1682 : ~n3182;
  assign n80034 = pi16 ? n32 : n80033;
  assign n80035 = pi14 ? n80029 : n80034;
  assign n80036 = pi17 ? n1580 : ~n2831;
  assign n80037 = pi16 ? n32 : n80036;
  assign n80038 = pi17 ? n2143 : ~n2733;
  assign n80039 = pi16 ? n32 : n80038;
  assign n80040 = pi17 ? n2143 : ~n2836;
  assign n80041 = pi16 ? n32 : n80040;
  assign n80042 = pi15 ? n80039 : n80041;
  assign n80043 = pi14 ? n80037 : n80042;
  assign n80044 = pi13 ? n80035 : n80043;
  assign n80045 = pi12 ? n80032 : n80044;
  assign n80046 = pi15 ? n80041 : n7185;
  assign n80047 = pi17 ? n1576 : ~n4245;
  assign n80048 = pi16 ? n32 : n80047;
  assign n80049 = pi15 ? n6568 : n80048;
  assign n80050 = pi14 ? n80046 : n80049;
  assign n80051 = pi17 ? n1576 : ~n2724;
  assign n80052 = pi16 ? n32 : n80051;
  assign n80053 = pi15 ? n80048 : n80052;
  assign n80054 = pi17 ? n1677 : ~n2731;
  assign n80055 = pi16 ? n32 : n80054;
  assign n80056 = pi15 ? n64265 : n80055;
  assign n80057 = pi14 ? n80053 : n80056;
  assign n80058 = pi13 ? n80050 : n80057;
  assign n80059 = pi17 ? n1677 : ~n2616;
  assign n80060 = pi16 ? n32 : n80059;
  assign n80061 = pi17 ? n2123 : ~n2616;
  assign n80062 = pi16 ? n32 : n80061;
  assign n80063 = pi15 ? n80060 : n80062;
  assign n80064 = pi17 ? n2123 : ~n2623;
  assign n80065 = pi16 ? n32 : n80064;
  assign n80066 = pi15 ? n80065 : n7524;
  assign n80067 = pi14 ? n80063 : n80066;
  assign n80068 = pi14 ? n7531 : n7533;
  assign n80069 = pi13 ? n80067 : n80068;
  assign n80070 = pi12 ? n80058 : n80069;
  assign n80071 = pi11 ? n80045 : n80070;
  assign n80072 = pi10 ? n80015 : n80071;
  assign n80073 = pi09 ? n79971 : n80072;
  assign n80074 = pi17 ? n3175 : ~n2954;
  assign n80075 = pi16 ? n32 : n80074;
  assign n80076 = pi15 ? n32 : n80075;
  assign n80077 = pi17 ? n2963 : ~n2954;
  assign n80078 = pi16 ? n32 : n80077;
  assign n80079 = pi15 ? n80075 : n80078;
  assign n80080 = pi14 ? n80076 : n80079;
  assign n80081 = pi13 ? n32 : n80080;
  assign n80082 = pi12 ? n32 : n80081;
  assign n80083 = pi11 ? n32 : n80082;
  assign n80084 = pi10 ? n32 : n80083;
  assign n80085 = pi17 ? n2831 : ~n2954;
  assign n80086 = pi16 ? n32 : n80085;
  assign n80087 = pi15 ? n80086 : n79962;
  assign n80088 = pi17 ? n4245 : ~n2954;
  assign n80089 = pi16 ? n32 : n80088;
  assign n80090 = pi17 ? n4245 : ~n3155;
  assign n80091 = pi16 ? n32 : n80090;
  assign n80092 = pi15 ? n80089 : n80091;
  assign n80093 = pi14 ? n80087 : n80092;
  assign n80094 = pi17 ? n2724 : ~n2954;
  assign n80095 = pi16 ? n32 : n80094;
  assign n80096 = pi17 ? n2731 : ~n2954;
  assign n80097 = pi16 ? n32 : n80096;
  assign n80098 = pi15 ? n80095 : n80097;
  assign n80099 = pi17 ? n2736 : ~n2954;
  assign n80100 = pi16 ? n32 : n80099;
  assign n80101 = pi15 ? n80100 : n79978;
  assign n80102 = pi14 ? n80098 : n80101;
  assign n80103 = pi13 ? n80093 : n80102;
  assign n80104 = pi15 ? n79978 : n79734;
  assign n80105 = pi14 ? n80104 : n79859;
  assign n80106 = pi15 ? n79863 : n79987;
  assign n80107 = pi14 ? n79864 : n80106;
  assign n80108 = pi13 ? n80105 : n80107;
  assign n80109 = pi12 ? n80103 : n80108;
  assign n80110 = pi15 ? n79987 : n79469;
  assign n80111 = pi15 ? n79739 : n79471;
  assign n80112 = pi14 ? n80110 : n80111;
  assign n80113 = pi15 ? n79471 : n79323;
  assign n80114 = pi14 ? n79471 : n80113;
  assign n80115 = pi13 ? n80112 : n80114;
  assign n80116 = pi17 ? n2305 : ~n3046;
  assign n80117 = pi16 ? n32 : n80116;
  assign n80118 = pi14 ? n79325 : n80117;
  assign n80119 = pi17 ? n2305 : ~n3292;
  assign n80120 = pi16 ? n32 : n80119;
  assign n80121 = pi17 ? n1933 : ~n3292;
  assign n80122 = pi16 ? n32 : n80121;
  assign n80123 = pi15 ? n80120 : n80122;
  assign n80124 = pi17 ? n1933 : ~n3587;
  assign n80125 = pi16 ? n32 : n80124;
  assign n80126 = pi15 ? n80122 : n80125;
  assign n80127 = pi14 ? n80123 : n80126;
  assign n80128 = pi13 ? n80118 : n80127;
  assign n80129 = pi12 ? n80115 : n80128;
  assign n80130 = pi11 ? n80109 : n80129;
  assign n80131 = pi17 ? n3337 : ~n3587;
  assign n80132 = pi16 ? n32 : n80131;
  assign n80133 = pi17 ? n2537 : ~n3587;
  assign n80134 = pi16 ? n32 : n80133;
  assign n80135 = pi15 ? n80132 : n80134;
  assign n80136 = pi17 ? n2537 : ~n3050;
  assign n80137 = pi16 ? n32 : n80136;
  assign n80138 = pi17 ? n3337 : ~n3050;
  assign n80139 = pi16 ? n32 : n80138;
  assign n80140 = pi15 ? n80137 : n80139;
  assign n80141 = pi14 ? n80135 : n80140;
  assign n80142 = pi17 ? n3337 : ~n2952;
  assign n80143 = pi16 ? n32 : n80142;
  assign n80144 = pi17 ? n1943 : ~n3175;
  assign n80145 = pi16 ? n32 : n80144;
  assign n80146 = pi17 ? n1943 : ~n2726;
  assign n80147 = pi16 ? n32 : n80146;
  assign n80148 = pi15 ? n80145 : n80147;
  assign n80149 = pi14 ? n80143 : n80148;
  assign n80150 = pi13 ? n80141 : n80149;
  assign n80151 = pi17 ? n1943 : ~n3182;
  assign n80152 = pi16 ? n32 : n80151;
  assign n80153 = pi15 ? n80147 : n80152;
  assign n80154 = pi17 ? n1943 : ~n2831;
  assign n80155 = pi16 ? n32 : n80154;
  assign n80156 = pi15 ? n80152 : n80155;
  assign n80157 = pi14 ? n80153 : n80156;
  assign n80158 = pi17 ? n1677 : ~n2831;
  assign n80159 = pi16 ? n32 : n80158;
  assign n80160 = pi17 ? n3351 : ~n2733;
  assign n80161 = pi16 ? n32 : n80160;
  assign n80162 = pi15 ? n80159 : n80161;
  assign n80163 = pi17 ? n2123 : ~n2836;
  assign n80164 = pi16 ? n32 : n80163;
  assign n80165 = pi15 ? n80161 : n80164;
  assign n80166 = pi14 ? n80162 : n80165;
  assign n80167 = pi13 ? n80157 : n80166;
  assign n80168 = pi12 ? n80150 : n80167;
  assign n80169 = pi17 ? n2123 : ~n2850;
  assign n80170 = pi16 ? n32 : n80169;
  assign n80171 = pi15 ? n80170 : n7699;
  assign n80172 = pi17 ? n3351 : ~n4245;
  assign n80173 = pi16 ? n32 : n80172;
  assign n80174 = pi15 ? n6784 : n80173;
  assign n80175 = pi14 ? n80171 : n80174;
  assign n80176 = pi17 ? n2325 : ~n4245;
  assign n80177 = pi16 ? n32 : n80176;
  assign n80178 = pi17 ? n2136 : ~n2724;
  assign n80179 = pi16 ? n32 : n80178;
  assign n80180 = pi15 ? n80177 : n80179;
  assign n80181 = pi17 ? n2136 : ~n2616;
  assign n80182 = pi16 ? n32 : n80181;
  assign n80183 = pi15 ? n80179 : n80182;
  assign n80184 = pi14 ? n80180 : n80183;
  assign n80185 = pi13 ? n80175 : n80184;
  assign n80186 = pi17 ? n1814 : ~n2616;
  assign n80187 = pi16 ? n32 : n80186;
  assign n80188 = pi15 ? n80182 : n80187;
  assign n80189 = pi17 ? n1814 : ~n2623;
  assign n80190 = pi16 ? n32 : n80189;
  assign n80191 = pi15 ? n80190 : n7725;
  assign n80192 = pi14 ? n80188 : n80191;
  assign n80193 = pi14 ? n7729 : n7731;
  assign n80194 = pi13 ? n80192 : n80193;
  assign n80195 = pi12 ? n80185 : n80194;
  assign n80196 = pi11 ? n80168 : n80195;
  assign n80197 = pi10 ? n80130 : n80196;
  assign n80198 = pi09 ? n80084 : n80197;
  assign n80199 = pi08 ? n80073 : n80198;
  assign n80200 = pi17 ? n3164 : ~n3155;
  assign n80201 = pi16 ? n32 : n80200;
  assign n80202 = pi15 ? n32 : n80201;
  assign n80203 = pi17 ? n3046 : ~n3155;
  assign n80204 = pi16 ? n32 : n80203;
  assign n80205 = pi17 ? n3292 : ~n3155;
  assign n80206 = pi16 ? n32 : n80205;
  assign n80207 = pi15 ? n80204 : n80206;
  assign n80208 = pi14 ? n80202 : n80207;
  assign n80209 = pi13 ? n32 : n80208;
  assign n80210 = pi12 ? n32 : n80209;
  assign n80211 = pi11 ? n32 : n80210;
  assign n80212 = pi10 ? n32 : n80211;
  assign n80213 = pi17 ? n2952 : ~n3155;
  assign n80214 = pi16 ? n32 : n80213;
  assign n80215 = pi17 ? n3175 : ~n3155;
  assign n80216 = pi16 ? n32 : n80215;
  assign n80217 = pi15 ? n80214 : n80216;
  assign n80218 = pi17 ? n2836 : ~n3155;
  assign n80219 = pi16 ? n32 : n80218;
  assign n80220 = pi15 ? n80219 : n79965;
  assign n80221 = pi14 ? n80217 : n80220;
  assign n80222 = pi15 ? n79965 : n79973;
  assign n80223 = pi17 ? n2850 : ~n2954;
  assign n80224 = pi16 ? n32 : n80223;
  assign n80225 = pi15 ? n80224 : n80089;
  assign n80226 = pi14 ? n80222 : n80225;
  assign n80227 = pi13 ? n80221 : n80226;
  assign n80228 = pi15 ? n79978 : n79852;
  assign n80229 = pi14 ? n80228 : n79980;
  assign n80230 = pi14 ? n79983 : n79734;
  assign n80231 = pi13 ? n80229 : n80230;
  assign n80232 = pi12 ? n80227 : n80231;
  assign n80233 = pi15 ? n79734 : n79601;
  assign n80234 = pi17 ? n2519 : ~n4111;
  assign n80235 = pi16 ? n32 : n80234;
  assign n80236 = pi15 ? n80235 : n79603;
  assign n80237 = pi14 ? n80233 : n80236;
  assign n80238 = pi15 ? n79603 : n79458;
  assign n80239 = pi14 ? n80238 : n79462;
  assign n80240 = pi13 ? n80237 : n80239;
  assign n80241 = pi17 ? n2425 : ~n3160;
  assign n80242 = pi16 ? n32 : n80241;
  assign n80243 = pi17 ? n3787 : ~n3160;
  assign n80244 = pi16 ? n32 : n80243;
  assign n80245 = pi15 ? n80242 : n80244;
  assign n80246 = pi17 ? n3787 : ~n3046;
  assign n80247 = pi16 ? n32 : n80246;
  assign n80248 = pi15 ? n80244 : n80247;
  assign n80249 = pi14 ? n80245 : n80248;
  assign n80250 = pi17 ? n3787 : ~n3292;
  assign n80251 = pi16 ? n32 : n80250;
  assign n80252 = pi17 ? n2531 : ~n3292;
  assign n80253 = pi16 ? n32 : n80252;
  assign n80254 = pi15 ? n80251 : n80253;
  assign n80255 = pi14 ? n80254 : n80253;
  assign n80256 = pi13 ? n80249 : n80255;
  assign n80257 = pi12 ? n80240 : n80256;
  assign n80258 = pi11 ? n80232 : n80257;
  assign n80259 = pi17 ? n2299 : ~n3587;
  assign n80260 = pi16 ? n32 : n80259;
  assign n80261 = pi17 ? n2299 : ~n3050;
  assign n80262 = pi16 ? n32 : n80261;
  assign n80263 = pi17 ? n2410 : ~n3050;
  assign n80264 = pi16 ? n32 : n80263;
  assign n80265 = pi15 ? n80262 : n80264;
  assign n80266 = pi14 ? n80260 : n80265;
  assign n80267 = pi17 ? n2410 : ~n2952;
  assign n80268 = pi16 ? n32 : n80267;
  assign n80269 = pi17 ? n2537 : ~n3175;
  assign n80270 = pi16 ? n32 : n80269;
  assign n80271 = pi17 ? n2319 : ~n2726;
  assign n80272 = pi16 ? n32 : n80271;
  assign n80273 = pi15 ? n80270 : n80272;
  assign n80274 = pi14 ? n80268 : n80273;
  assign n80275 = pi13 ? n80266 : n80274;
  assign n80276 = pi17 ? n1933 : ~n3182;
  assign n80277 = pi16 ? n32 : n80276;
  assign n80278 = pi15 ? n80272 : n80277;
  assign n80279 = pi17 ? n2319 : ~n3182;
  assign n80280 = pi16 ? n32 : n80279;
  assign n80281 = pi17 ? n1933 : ~n2831;
  assign n80282 = pi16 ? n32 : n80281;
  assign n80283 = pi15 ? n80280 : n80282;
  assign n80284 = pi14 ? n80278 : n80283;
  assign n80285 = pi17 ? n1807 : ~n2831;
  assign n80286 = pi16 ? n32 : n80285;
  assign n80287 = pi17 ? n1807 : ~n2733;
  assign n80288 = pi16 ? n32 : n80287;
  assign n80289 = pi15 ? n80286 : n80288;
  assign n80290 = pi17 ? n1814 : ~n2836;
  assign n80291 = pi16 ? n32 : n80290;
  assign n80292 = pi15 ? n80288 : n80291;
  assign n80293 = pi14 ? n80289 : n80292;
  assign n80294 = pi13 ? n80284 : n80293;
  assign n80295 = pi12 ? n80275 : n80294;
  assign n80296 = pi17 ? n1814 : ~n2850;
  assign n80297 = pi16 ? n32 : n80296;
  assign n80298 = pi15 ? n80297 : n7904;
  assign n80299 = pi14 ? n80298 : n7909;
  assign n80300 = pi17 ? n2319 : ~n2724;
  assign n80301 = pi16 ? n32 : n80300;
  assign n80302 = pi17 ? n2319 : ~n2616;
  assign n80303 = pi16 ? n32 : n80302;
  assign n80304 = pi14 ? n80301 : n80303;
  assign n80305 = pi13 ? n80299 : n80304;
  assign n80306 = pi17 ? n1933 : ~n2855;
  assign n80307 = pi16 ? n32 : n80306;
  assign n80308 = pi15 ? n80303 : n80307;
  assign n80309 = pi17 ? n2410 : ~n2750;
  assign n80310 = pi16 ? n32 : n80309;
  assign n80311 = pi15 ? n80310 : n7586;
  assign n80312 = pi14 ? n80308 : n80311;
  assign n80313 = pi17 ? n2299 : ~n2628;
  assign n80314 = pi16 ? n32 : n80313;
  assign n80315 = pi15 ? n7586 : n80314;
  assign n80316 = pi14 ? n80315 : n7950;
  assign n80317 = pi13 ? n80312 : n80316;
  assign n80318 = pi12 ? n80305 : n80317;
  assign n80319 = pi11 ? n80295 : n80318;
  assign n80320 = pi10 ? n80258 : n80319;
  assign n80321 = pi09 ? n80212 : n80320;
  assign n80322 = pi17 ? n2954 : ~n3155;
  assign n80323 = pi16 ? n32 : n80322;
  assign n80324 = pi15 ? n32 : n80323;
  assign n80325 = pi17 ? n4111 : ~n3155;
  assign n80326 = pi16 ? n32 : n80325;
  assign n80327 = pi15 ? n80323 : n80326;
  assign n80328 = pi14 ? n80324 : n80327;
  assign n80329 = pi13 ? n32 : n80328;
  assign n80330 = pi12 ? n32 : n80329;
  assign n80331 = pi11 ? n32 : n80330;
  assign n80332 = pi10 ? n32 : n80331;
  assign n80333 = pi17 ? n3160 : ~n3155;
  assign n80334 = pi16 ? n32 : n80333;
  assign n80335 = pi15 ? n80334 : n80201;
  assign n80336 = pi17 ? n2726 : ~n3155;
  assign n80337 = pi16 ? n32 : n80336;
  assign n80338 = pi17 ? n2726 : ~n2954;
  assign n80339 = pi16 ? n32 : n80338;
  assign n80340 = pi15 ? n80337 : n80339;
  assign n80341 = pi14 ? n80335 : n80340;
  assign n80342 = pi17 ? n3182 : ~n3155;
  assign n80343 = pi16 ? n32 : n80342;
  assign n80344 = pi15 ? n80337 : n80343;
  assign n80345 = pi17 ? n2733 : ~n3155;
  assign n80346 = pi16 ? n32 : n80345;
  assign n80347 = pi15 ? n80346 : n80219;
  assign n80348 = pi14 ? n80344 : n80347;
  assign n80349 = pi13 ? n80341 : n80348;
  assign n80350 = pi17 ? n2724 : ~n3155;
  assign n80351 = pi16 ? n32 : n80350;
  assign n80352 = pi17 ? n2731 : ~n3155;
  assign n80353 = pi16 ? n32 : n80352;
  assign n80354 = pi15 ? n80351 : n80353;
  assign n80355 = pi14 ? n80091 : n80354;
  assign n80356 = pi17 ? n2736 : ~n3155;
  assign n80357 = pi16 ? n32 : n80356;
  assign n80358 = pi17 ? n2750 : ~n3155;
  assign n80359 = pi16 ? n32 : n80358;
  assign n80360 = pi15 ? n80357 : n80359;
  assign n80361 = pi14 ? n80360 : n80359;
  assign n80362 = pi13 ? n80355 : n80361;
  assign n80363 = pi12 ? n80349 : n80362;
  assign n80364 = pi17 ? n2618 : ~n2954;
  assign n80365 = pi16 ? n32 : n80364;
  assign n80366 = pi15 ? n79978 : n80365;
  assign n80367 = pi17 ? n2628 : ~n2954;
  assign n80368 = pi16 ? n32 : n80367;
  assign n80369 = pi15 ? n80368 : n79590;
  assign n80370 = pi14 ? n80366 : n80369;
  assign n80371 = pi14 ? n79590 : n79594;
  assign n80372 = pi13 ? n80370 : n80371;
  assign n80373 = pi17 ? n2755 : ~n3160;
  assign n80374 = pi16 ? n32 : n80373;
  assign n80375 = pi17 ? n2292 : ~n3160;
  assign n80376 = pi16 ? n32 : n80375;
  assign n80377 = pi15 ? n80374 : n80376;
  assign n80378 = pi17 ? n2408 : ~n3046;
  assign n80379 = pi16 ? n32 : n80378;
  assign n80380 = pi15 ? n80376 : n80379;
  assign n80381 = pi14 ? n80377 : n80380;
  assign n80382 = pi17 ? n2408 : ~n3292;
  assign n80383 = pi16 ? n32 : n80382;
  assign n80384 = pi17 ? n2414 : ~n3292;
  assign n80385 = pi16 ? n32 : n80384;
  assign n80386 = pi15 ? n80383 : n80385;
  assign n80387 = pi17 ? n2425 : ~n3587;
  assign n80388 = pi16 ? n32 : n80387;
  assign n80389 = pi15 ? n80385 : n80388;
  assign n80390 = pi14 ? n80386 : n80389;
  assign n80391 = pi13 ? n80381 : n80390;
  assign n80392 = pi12 ? n80372 : n80391;
  assign n80393 = pi11 ? n80363 : n80392;
  assign n80394 = pi17 ? n2425 : ~n3050;
  assign n80395 = pi16 ? n32 : n80394;
  assign n80396 = pi17 ? n2653 : ~n3050;
  assign n80397 = pi16 ? n32 : n80396;
  assign n80398 = pi15 ? n80395 : n80397;
  assign n80399 = pi14 ? n80388 : n80398;
  assign n80400 = pi17 ? n2653 : ~n2952;
  assign n80401 = pi16 ? n32 : n80400;
  assign n80402 = pi17 ? n3787 : ~n3175;
  assign n80403 = pi16 ? n32 : n80402;
  assign n80404 = pi17 ? n3787 : ~n2726;
  assign n80405 = pi16 ? n32 : n80404;
  assign n80406 = pi15 ? n80403 : n80405;
  assign n80407 = pi14 ? n80401 : n80406;
  assign n80408 = pi13 ? n80399 : n80407;
  assign n80409 = pi17 ? n3787 : ~n3182;
  assign n80410 = pi16 ? n32 : n80409;
  assign n80411 = pi15 ? n80405 : n80410;
  assign n80412 = pi17 ? n3787 : ~n2831;
  assign n80413 = pi16 ? n32 : n80412;
  assign n80414 = pi15 ? n80410 : n80413;
  assign n80415 = pi14 ? n80411 : n80414;
  assign n80416 = pi17 ? n2305 : ~n2733;
  assign n80417 = pi16 ? n32 : n80416;
  assign n80418 = pi15 ? n80282 : n80417;
  assign n80419 = pi17 ? n2410 : ~n2850;
  assign n80420 = pi16 ? n32 : n80419;
  assign n80421 = pi15 ? n80417 : n80420;
  assign n80422 = pi14 ? n80418 : n80421;
  assign n80423 = pi13 ? n80415 : n80422;
  assign n80424 = pi12 ? n80408 : n80423;
  assign n80425 = pi14 ? n8091 : n8096;
  assign n80426 = pi17 ? n2299 : ~n2724;
  assign n80427 = pi16 ? n32 : n80426;
  assign n80428 = pi17 ? n2531 : ~n2616;
  assign n80429 = pi16 ? n32 : n80428;
  assign n80430 = pi14 ? n80427 : n80429;
  assign n80431 = pi13 ? n80425 : n80430;
  assign n80432 = pi17 ? n2653 : ~n2616;
  assign n80433 = pi16 ? n32 : n80432;
  assign n80434 = pi17 ? n2425 : ~n2855;
  assign n80435 = pi16 ? n32 : n80434;
  assign n80436 = pi15 ? n80433 : n80435;
  assign n80437 = pi17 ? n2653 : ~n2750;
  assign n80438 = pi16 ? n32 : n80437;
  assign n80439 = pi15 ? n80438 : n8121;
  assign n80440 = pi14 ? n80436 : n80439;
  assign n80441 = pi17 ? n2119 : ~n2628;
  assign n80442 = pi16 ? n32 : n80441;
  assign n80443 = pi15 ? n8125 : n80442;
  assign n80444 = pi15 ? n46420 : n8137;
  assign n80445 = pi14 ? n80443 : n80444;
  assign n80446 = pi13 ? n80440 : n80445;
  assign n80447 = pi12 ? n80431 : n80446;
  assign n80448 = pi11 ? n80424 : n80447;
  assign n80449 = pi10 ? n80393 : n80448;
  assign n80450 = pi09 ? n80332 : n80449;
  assign n80451 = pi08 ? n80321 : n80450;
  assign n80452 = pi07 ? n80199 : n80451;
  assign n80453 = pi06 ? n79960 : n80452;
  assign n80454 = pi18 ? n1676 : ~n936;
  assign n80455 = pi17 ? n32 : n80454;
  assign n80456 = pi16 ? n32 : n80455;
  assign n80457 = pi15 ? n32 : n80456;
  assign n80458 = pi17 ? n3569 : ~n3282;
  assign n80459 = pi16 ? n32 : n80458;
  assign n80460 = pi14 ? n80457 : n80459;
  assign n80461 = pi13 ? n32 : n80460;
  assign n80462 = pi12 ? n32 : n80461;
  assign n80463 = pi11 ? n32 : n80462;
  assign n80464 = pi10 ? n32 : n80463;
  assign n80465 = pi17 ? n3282 : ~n3282;
  assign n80466 = pi16 ? n32 : n80465;
  assign n80467 = pi17 ? n3155 : ~n3282;
  assign n80468 = pi16 ? n32 : n80467;
  assign n80469 = pi15 ? n80466 : n80468;
  assign n80470 = pi17 ? n3046 : ~n3282;
  assign n80471 = pi16 ? n32 : n80470;
  assign n80472 = pi15 ? n80471 : n80204;
  assign n80473 = pi14 ? n80469 : n80472;
  assign n80474 = pi17 ? n3587 : ~n3155;
  assign n80475 = pi16 ? n32 : n80474;
  assign n80476 = pi15 ? n80206 : n80475;
  assign n80477 = pi15 ? n80216 : n80337;
  assign n80478 = pi14 ? n80476 : n80477;
  assign n80479 = pi13 ? n80473 : n80478;
  assign n80480 = pi17 ? n2839 : ~n3155;
  assign n80481 = pi16 ? n32 : n80480;
  assign n80482 = pi15 ? n80219 : n80481;
  assign n80483 = pi14 ? n80219 : n80482;
  assign n80484 = pi17 ? n2850 : ~n3155;
  assign n80485 = pi16 ? n32 : n80484;
  assign n80486 = pi15 ? n80485 : n80091;
  assign n80487 = pi14 ? n80486 : n80091;
  assign n80488 = pi13 ? n80483 : n80487;
  assign n80489 = pi12 ? n80479 : n80488;
  assign n80490 = pi17 ? n2623 : ~n4111;
  assign n80491 = pi16 ? n32 : n80490;
  assign n80492 = pi15 ? n80100 : n80491;
  assign n80493 = pi14 ? n80098 : n80492;
  assign n80494 = pi17 ? n4099 : ~n4111;
  assign n80495 = pi16 ? n32 : n80494;
  assign n80496 = pi15 ? n80491 : n80495;
  assign n80497 = pi14 ? n80491 : n80496;
  assign n80498 = pi13 ? n80493 : n80497;
  assign n80499 = pi17 ? n2618 : ~n3160;
  assign n80500 = pi16 ? n32 : n80499;
  assign n80501 = pi17 ? n2628 : ~n3160;
  assign n80502 = pi16 ? n32 : n80501;
  assign n80503 = pi15 ? n80500 : n80502;
  assign n80504 = pi17 ? n2628 : ~n3046;
  assign n80505 = pi16 ? n32 : n80504;
  assign n80506 = pi14 ? n80503 : n80505;
  assign n80507 = pi17 ? n2628 : ~n3292;
  assign n80508 = pi16 ? n32 : n80507;
  assign n80509 = pi17 ? n2748 : ~n3292;
  assign n80510 = pi16 ? n32 : n80509;
  assign n80511 = pi15 ? n80508 : n80510;
  assign n80512 = pi17 ? n2748 : ~n3587;
  assign n80513 = pi16 ? n32 : n80512;
  assign n80514 = pi17 ? n2755 : ~n3587;
  assign n80515 = pi16 ? n32 : n80514;
  assign n80516 = pi15 ? n80513 : n80515;
  assign n80517 = pi14 ? n80511 : n80516;
  assign n80518 = pi13 ? n80506 : n80517;
  assign n80519 = pi12 ? n80498 : n80518;
  assign n80520 = pi11 ? n80489 : n80519;
  assign n80521 = pi17 ? n2519 : ~n3050;
  assign n80522 = pi16 ? n32 : n80521;
  assign n80523 = pi15 ? n80515 : n80522;
  assign n80524 = pi17 ? n2292 : ~n2952;
  assign n80525 = pi16 ? n32 : n80524;
  assign n80526 = pi15 ? n80522 : n80525;
  assign n80527 = pi14 ? n80523 : n80526;
  assign n80528 = pi17 ? n2414 : ~n3175;
  assign n80529 = pi16 ? n32 : n80528;
  assign n80530 = pi15 ? n80525 : n80529;
  assign n80531 = pi15 ? n80529 : n8264;
  assign n80532 = pi14 ? n80530 : n80531;
  assign n80533 = pi13 ? n80527 : n80532;
  assign n80534 = pi17 ? n2414 : ~n3182;
  assign n80535 = pi16 ? n32 : n80534;
  assign n80536 = pi14 ? n80535 : n8284;
  assign n80537 = pi17 ? n3787 : ~n2733;
  assign n80538 = pi16 ? n32 : n80537;
  assign n80539 = pi17 ? n2119 : ~n2733;
  assign n80540 = pi16 ? n32 : n80539;
  assign n80541 = pi15 ? n80538 : n80540;
  assign n80542 = pi17 ? n2119 : ~n2850;
  assign n80543 = pi16 ? n32 : n80542;
  assign n80544 = pi15 ? n80543 : n8295;
  assign n80545 = pi14 ? n80541 : n80544;
  assign n80546 = pi13 ? n80536 : n80545;
  assign n80547 = pi12 ? n80533 : n80546;
  assign n80548 = pi15 ? n8295 : n6964;
  assign n80549 = pi17 ? n2425 : ~n2724;
  assign n80550 = pi16 ? n32 : n80549;
  assign n80551 = pi15 ? n8309 : n80550;
  assign n80552 = pi14 ? n80548 : n80551;
  assign n80553 = pi17 ? n2119 : ~n2616;
  assign n80554 = pi16 ? n32 : n80553;
  assign n80555 = pi15 ? n8309 : n80554;
  assign n80556 = pi14 ? n80555 : n8314;
  assign n80557 = pi13 ? n80552 : n80556;
  assign n80558 = pi17 ? n2519 : ~n2618;
  assign n80559 = pi16 ? n32 : n80558;
  assign n80560 = pi15 ? n8321 : n80559;
  assign n80561 = pi14 ? n8322 : n80560;
  assign n80562 = pi17 ? n2748 : ~n2628;
  assign n80563 = pi16 ? n32 : n80562;
  assign n80564 = pi15 ? n35097 : n80563;
  assign n80565 = pi14 ? n80564 : n8334;
  assign n80566 = pi13 ? n80561 : n80565;
  assign n80567 = pi12 ? n80557 : n80566;
  assign n80568 = pi11 ? n80547 : n80567;
  assign n80569 = pi10 ? n80520 : n80568;
  assign n80570 = pi09 ? n80464 : n80569;
  assign n80571 = pi18 ? n3350 : ~n936;
  assign n80572 = pi17 ? n32 : n80571;
  assign n80573 = pi16 ? n32 : n80572;
  assign n80574 = pi15 ? n32 : n80573;
  assign n80575 = pi14 ? n80574 : n80573;
  assign n80576 = pi13 ? n32 : n80575;
  assign n80577 = pi12 ? n32 : n80576;
  assign n80578 = pi11 ? n32 : n80577;
  assign n80579 = pi10 ? n32 : n80578;
  assign n80580 = pi18 ? n618 : ~n936;
  assign n80581 = pi17 ? n32 : n80580;
  assign n80582 = pi16 ? n32 : n80581;
  assign n80583 = pi15 ? n80582 : n80468;
  assign n80584 = pi17 ? n3728 : ~n3155;
  assign n80585 = pi16 ? n32 : n80584;
  assign n80586 = pi15 ? n80323 : n80585;
  assign n80587 = pi14 ? n80583 : n80586;
  assign n80588 = pi15 ? n80585 : n80334;
  assign n80589 = pi15 ? n80201 : n80204;
  assign n80590 = pi14 ? n80588 : n80589;
  assign n80591 = pi13 ? n80587 : n80590;
  assign n80592 = pi14 ? n80337 : n80344;
  assign n80593 = pi14 ? n80347 : n80219;
  assign n80594 = pi13 ? n80592 : n80593;
  assign n80595 = pi12 ? n80591 : n80594;
  assign n80596 = pi15 ? n80219 : n79973;
  assign n80597 = pi17 ? n3067 : ~n4111;
  assign n80598 = pi16 ? n32 : n80597;
  assign n80599 = pi15 ? n80224 : n80598;
  assign n80600 = pi14 ? n80596 : n80599;
  assign n80601 = pi17 ? n4245 : ~n4111;
  assign n80602 = pi16 ? n32 : n80601;
  assign n80603 = pi17 ? n2724 : ~n4111;
  assign n80604 = pi16 ? n32 : n80603;
  assign n80605 = pi15 ? n80602 : n80604;
  assign n80606 = pi14 ? n80598 : n80605;
  assign n80607 = pi13 ? n80600 : n80606;
  assign n80608 = pi17 ? n2731 : ~n3160;
  assign n80609 = pi16 ? n32 : n80608;
  assign n80610 = pi17 ? n2855 : ~n3160;
  assign n80611 = pi16 ? n32 : n80610;
  assign n80612 = pi15 ? n80609 : n80611;
  assign n80613 = pi17 ? n2855 : ~n3046;
  assign n80614 = pi16 ? n32 : n80613;
  assign n80615 = pi14 ? n80612 : n80614;
  assign n80616 = pi17 ? n2855 : ~n3292;
  assign n80617 = pi16 ? n32 : n80616;
  assign n80618 = pi17 ? n2750 : ~n3292;
  assign n80619 = pi16 ? n32 : n80618;
  assign n80620 = pi15 ? n80617 : n80619;
  assign n80621 = pi17 ? n2750 : ~n3587;
  assign n80622 = pi16 ? n32 : n80621;
  assign n80623 = pi17 ? n4099 : ~n3587;
  assign n80624 = pi16 ? n32 : n80623;
  assign n80625 = pi15 ? n80622 : n80624;
  assign n80626 = pi14 ? n80620 : n80625;
  assign n80627 = pi13 ? n80615 : n80626;
  assign n80628 = pi12 ? n80607 : n80627;
  assign n80629 = pi11 ? n80595 : n80628;
  assign n80630 = pi17 ? n4099 : ~n3050;
  assign n80631 = pi16 ? n32 : n80630;
  assign n80632 = pi15 ? n80624 : n80631;
  assign n80633 = pi17 ? n2628 : ~n2952;
  assign n80634 = pi16 ? n32 : n80633;
  assign n80635 = pi15 ? n80631 : n80634;
  assign n80636 = pi14 ? n80632 : n80635;
  assign n80637 = pi15 ? n80634 : n8447;
  assign n80638 = pi17 ? n2748 : ~n3175;
  assign n80639 = pi16 ? n32 : n80638;
  assign n80640 = pi17 ? n2517 : ~n2726;
  assign n80641 = pi16 ? n32 : n80640;
  assign n80642 = pi15 ? n80639 : n80641;
  assign n80643 = pi14 ? n80637 : n80642;
  assign n80644 = pi13 ? n80636 : n80643;
  assign n80645 = pi17 ? n2517 : ~n3182;
  assign n80646 = pi16 ? n32 : n80645;
  assign n80647 = pi17 ? n2519 : ~n2831;
  assign n80648 = pi16 ? n32 : n80647;
  assign n80649 = pi15 ? n8460 : n80648;
  assign n80650 = pi14 ? n80646 : n80649;
  assign n80651 = pi17 ? n2519 : ~n2733;
  assign n80652 = pi16 ? n32 : n80651;
  assign n80653 = pi17 ? n2519 : ~n2850;
  assign n80654 = pi16 ? n32 : n80653;
  assign n80655 = pi15 ? n80654 : n8466;
  assign n80656 = pi14 ? n80652 : n80655;
  assign n80657 = pi13 ? n80650 : n80656;
  assign n80658 = pi12 ? n80644 : n80657;
  assign n80659 = pi15 ? n80654 : n7781;
  assign n80660 = pi14 ? n80659 : n69306;
  assign n80661 = pi15 ? n8480 : n8485;
  assign n80662 = pi14 ? n80661 : n8485;
  assign n80663 = pi13 ? n80660 : n80662;
  assign n80664 = pi17 ? n2748 : ~n2750;
  assign n80665 = pi16 ? n32 : n80664;
  assign n80666 = pi17 ? n4099 : ~n2618;
  assign n80667 = pi16 ? n32 : n80666;
  assign n80668 = pi15 ? n80665 : n80667;
  assign n80669 = pi14 ? n8489 : n80668;
  assign n80670 = pi17 ? n4099 : ~n2517;
  assign n80671 = pi16 ? n32 : n80670;
  assign n80672 = pi15 ? n8493 : n80671;
  assign n80673 = pi14 ? n8497 : n80672;
  assign n80674 = pi13 ? n80669 : n80673;
  assign n80675 = pi12 ? n80663 : n80674;
  assign n80676 = pi11 ? n80658 : n80675;
  assign n80677 = pi10 ? n80629 : n80676;
  assign n80678 = pi09 ? n80579 : n80677;
  assign n80679 = pi08 ? n80570 : n80678;
  assign n80680 = pi18 ? n1813 : ~n936;
  assign n80681 = pi17 ? n32 : n80680;
  assign n80682 = pi16 ? n32 : n80681;
  assign n80683 = pi15 ? n32 : n80682;
  assign n80684 = pi18 ? n1813 : ~n1575;
  assign n80685 = pi17 ? n32 : n80684;
  assign n80686 = pi16 ? n32 : n80685;
  assign n80687 = pi18 ? n814 : ~n1575;
  assign n80688 = pi17 ? n32 : n80687;
  assign n80689 = pi16 ? n32 : n80688;
  assign n80690 = pi15 ? n80686 : n80689;
  assign n80691 = pi14 ? n80683 : n80690;
  assign n80692 = pi13 ? n32 : n80691;
  assign n80693 = pi12 ? n32 : n80692;
  assign n80694 = pi11 ? n32 : n80693;
  assign n80695 = pi10 ? n32 : n80694;
  assign n80696 = pi18 ? n1676 : ~n1575;
  assign n80697 = pi17 ? n32 : n80696;
  assign n80698 = pi16 ? n32 : n80697;
  assign n80699 = pi15 ? n80689 : n80698;
  assign n80700 = pi17 ? n32 : ~n3569;
  assign n80701 = pi16 ? n32 : n80700;
  assign n80702 = pi14 ? n80699 : n80701;
  assign n80703 = pi17 ? n3282 : ~n3569;
  assign n80704 = pi16 ? n32 : n80703;
  assign n80705 = pi17 ? n3155 : ~n3569;
  assign n80706 = pi16 ? n32 : n80705;
  assign n80707 = pi17 ? n2954 : ~n3569;
  assign n80708 = pi16 ? n32 : n80707;
  assign n80709 = pi15 ? n80706 : n80708;
  assign n80710 = pi14 ? n80704 : n80709;
  assign n80711 = pi13 ? n80702 : n80710;
  assign n80712 = pi17 ? n3046 : ~n3569;
  assign n80713 = pi16 ? n32 : n80712;
  assign n80714 = pi17 ? n3292 : ~n3569;
  assign n80715 = pi16 ? n32 : n80714;
  assign n80716 = pi17 ? n3587 : ~n3569;
  assign n80717 = pi16 ? n32 : n80716;
  assign n80718 = pi15 ? n80715 : n80717;
  assign n80719 = pi14 ? n80713 : n80718;
  assign n80720 = pi14 ? n80477 : n80337;
  assign n80721 = pi13 ? n80719 : n80720;
  assign n80722 = pi12 ? n80711 : n80721;
  assign n80723 = pi17 ? n3182 : ~n2954;
  assign n80724 = pi16 ? n32 : n80723;
  assign n80725 = pi15 ? n80337 : n80724;
  assign n80726 = pi17 ? n2733 : ~n4111;
  assign n80727 = pi16 ? n32 : n80726;
  assign n80728 = pi15 ? n79962 : n80727;
  assign n80729 = pi14 ? n80725 : n80728;
  assign n80730 = pi17 ? n2836 : ~n3160;
  assign n80731 = pi16 ? n32 : n80730;
  assign n80732 = pi15 ? n80727 : n80731;
  assign n80733 = pi14 ? n80727 : n80732;
  assign n80734 = pi13 ? n80729 : n80733;
  assign n80735 = pi17 ? n2839 : ~n3160;
  assign n80736 = pi16 ? n32 : n80735;
  assign n80737 = pi17 ? n2850 : ~n3160;
  assign n80738 = pi16 ? n32 : n80737;
  assign n80739 = pi15 ? n80736 : n80738;
  assign n80740 = pi17 ? n2850 : ~n3046;
  assign n80741 = pi16 ? n32 : n80740;
  assign n80742 = pi14 ? n80739 : n80741;
  assign n80743 = pi17 ? n3067 : ~n3292;
  assign n80744 = pi16 ? n32 : n80743;
  assign n80745 = pi17 ? n4245 : ~n3292;
  assign n80746 = pi16 ? n32 : n80745;
  assign n80747 = pi15 ? n80744 : n80746;
  assign n80748 = pi17 ? n4245 : ~n3587;
  assign n80749 = pi16 ? n32 : n80748;
  assign n80750 = pi17 ? n2736 : ~n3587;
  assign n80751 = pi16 ? n32 : n80750;
  assign n80752 = pi15 ? n80749 : n80751;
  assign n80753 = pi14 ? n80747 : n80752;
  assign n80754 = pi13 ? n80742 : n80753;
  assign n80755 = pi12 ? n80734 : n80754;
  assign n80756 = pi11 ? n80722 : n80755;
  assign n80757 = pi17 ? n2736 : ~n3050;
  assign n80758 = pi16 ? n32 : n80757;
  assign n80759 = pi15 ? n80751 : n80758;
  assign n80760 = pi17 ? n2855 : ~n2952;
  assign n80761 = pi16 ? n32 : n80760;
  assign n80762 = pi15 ? n80758 : n80761;
  assign n80763 = pi14 ? n80759 : n80762;
  assign n80764 = pi17 ? n2623 : ~n3175;
  assign n80765 = pi16 ? n32 : n80764;
  assign n80766 = pi15 ? n80761 : n80765;
  assign n80767 = pi17 ? n2623 : ~n3182;
  assign n80768 = pi16 ? n32 : n80767;
  assign n80769 = pi15 ? n80765 : n80768;
  assign n80770 = pi14 ? n80766 : n80769;
  assign n80771 = pi13 ? n80763 : n80770;
  assign n80772 = pi17 ? n2750 : ~n3182;
  assign n80773 = pi16 ? n32 : n80772;
  assign n80774 = pi15 ? n80768 : n80773;
  assign n80775 = pi17 ? n2750 : ~n2831;
  assign n80776 = pi16 ? n32 : n80775;
  assign n80777 = pi17 ? n2512 : ~n2733;
  assign n80778 = pi16 ? n32 : n80777;
  assign n80779 = pi15 ? n80776 : n80778;
  assign n80780 = pi14 ? n80774 : n80779;
  assign n80781 = pi17 ? n2628 : ~n2733;
  assign n80782 = pi16 ? n32 : n80781;
  assign n80783 = pi15 ? n80778 : n80782;
  assign n80784 = pi17 ? n2628 : ~n2850;
  assign n80785 = pi16 ? n32 : n80784;
  assign n80786 = pi17 ? n2618 : ~n2850;
  assign n80787 = pi16 ? n32 : n80786;
  assign n80788 = pi15 ? n80785 : n80787;
  assign n80789 = pi14 ? n80783 : n80788;
  assign n80790 = pi13 ? n80780 : n80789;
  assign n80791 = pi12 ? n80771 : n80790;
  assign n80792 = pi17 ? n4099 : ~n2850;
  assign n80793 = pi16 ? n32 : n80792;
  assign n80794 = pi15 ? n80793 : n6949;
  assign n80795 = pi14 ? n80794 : n8672;
  assign n80796 = pi14 ? n8686 : n8688;
  assign n80797 = pi13 ? n80795 : n80796;
  assign n80798 = pi17 ? n2855 : ~n2623;
  assign n80799 = pi16 ? n32 : n80798;
  assign n80800 = pi17 ? n2616 : ~n2750;
  assign n80801 = pi16 ? n32 : n80800;
  assign n80802 = pi15 ? n80799 : n80801;
  assign n80803 = pi17 ? n2855 : ~n2618;
  assign n80804 = pi16 ? n32 : n80803;
  assign n80805 = pi17 ? n2616 : ~n2618;
  assign n80806 = pi16 ? n32 : n80805;
  assign n80807 = pi15 ? n80804 : n80806;
  assign n80808 = pi14 ? n80802 : n80807;
  assign n80809 = pi17 ? n2736 : ~n2628;
  assign n80810 = pi16 ? n32 : n80809;
  assign n80811 = pi15 ? n8707 : n80810;
  assign n80812 = pi15 ? n8709 : n8716;
  assign n80813 = pi14 ? n80811 : n80812;
  assign n80814 = pi13 ? n80808 : n80813;
  assign n80815 = pi12 ? n80797 : n80814;
  assign n80816 = pi11 ? n80791 : n80815;
  assign n80817 = pi10 ? n80756 : n80816;
  assign n80818 = pi09 ? n80695 : n80817;
  assign n80819 = pi18 ? n2298 : ~n936;
  assign n80820 = pi17 ? n32 : n80819;
  assign n80821 = pi16 ? n32 : n80820;
  assign n80822 = pi15 ? n32 : n80821;
  assign n80823 = pi18 ? n430 : ~n1575;
  assign n80824 = pi17 ? n32 : n80823;
  assign n80825 = pi16 ? n32 : n80824;
  assign n80826 = pi14 ? n80822 : n80825;
  assign n80827 = pi13 ? n32 : n80826;
  assign n80828 = pi12 ? n32 : n80827;
  assign n80829 = pi11 ? n32 : n80828;
  assign n80830 = pi10 ? n32 : n80829;
  assign n80831 = pi18 ? n2304 : ~n1575;
  assign n80832 = pi17 ? n32 : n80831;
  assign n80833 = pi16 ? n32 : n80832;
  assign n80834 = pi18 ? n1942 : ~n1575;
  assign n80835 = pi17 ? n32 : n80834;
  assign n80836 = pi16 ? n32 : n80835;
  assign n80837 = pi15 ? n80833 : n80836;
  assign n80838 = pi18 ? n237 : ~n1575;
  assign n80839 = pi17 ? n32 : n80838;
  assign n80840 = pi16 ? n32 : n80839;
  assign n80841 = pi18 ? n618 : ~n1575;
  assign n80842 = pi17 ? n32 : n80841;
  assign n80843 = pi16 ? n32 : n80842;
  assign n80844 = pi15 ? n80840 : n80843;
  assign n80845 = pi14 ? n80837 : n80844;
  assign n80846 = pi15 ? n80698 : n80708;
  assign n80847 = pi14 ? n80843 : n80846;
  assign n80848 = pi13 ? n80845 : n80847;
  assign n80849 = pi17 ? n3728 : ~n3569;
  assign n80850 = pi16 ? n32 : n80849;
  assign n80851 = pi15 ? n80708 : n80850;
  assign n80852 = pi17 ? n3160 : ~n3569;
  assign n80853 = pi16 ? n32 : n80852;
  assign n80854 = pi15 ? n80850 : n80853;
  assign n80855 = pi14 ? n80851 : n80854;
  assign n80856 = pi14 ? n80589 : n80204;
  assign n80857 = pi13 ? n80855 : n80856;
  assign n80858 = pi12 ? n80848 : n80857;
  assign n80859 = pi17 ? n3587 : ~n2954;
  assign n80860 = pi16 ? n32 : n80859;
  assign n80861 = pi15 ? n80206 : n80860;
  assign n80862 = pi17 ? n3175 : ~n4111;
  assign n80863 = pi16 ? n32 : n80862;
  assign n80864 = pi15 ? n80075 : n80863;
  assign n80865 = pi14 ? n80861 : n80864;
  assign n80866 = pi17 ? n2963 : ~n3160;
  assign n80867 = pi16 ? n32 : n80866;
  assign n80868 = pi15 ? n80863 : n80867;
  assign n80869 = pi14 ? n80863 : n80868;
  assign n80870 = pi13 ? n80865 : n80869;
  assign n80871 = pi17 ? n2831 : ~n3160;
  assign n80872 = pi16 ? n32 : n80871;
  assign n80873 = pi17 ? n2831 : ~n3046;
  assign n80874 = pi16 ? n32 : n80873;
  assign n80875 = pi14 ? n80872 : n80874;
  assign n80876 = pi17 ? n2831 : ~n3292;
  assign n80877 = pi16 ? n32 : n80876;
  assign n80878 = pi17 ? n2733 : ~n3292;
  assign n80879 = pi16 ? n32 : n80878;
  assign n80880 = pi15 ? n80877 : n80879;
  assign n80881 = pi17 ? n2733 : ~n3587;
  assign n80882 = pi16 ? n32 : n80881;
  assign n80883 = pi17 ? n2836 : ~n3587;
  assign n80884 = pi16 ? n32 : n80883;
  assign n80885 = pi15 ? n80882 : n80884;
  assign n80886 = pi14 ? n80880 : n80885;
  assign n80887 = pi13 ? n80875 : n80886;
  assign n80888 = pi12 ? n80870 : n80887;
  assign n80889 = pi11 ? n80858 : n80888;
  assign n80890 = pi17 ? n2836 : ~n3050;
  assign n80891 = pi16 ? n32 : n80890;
  assign n80892 = pi15 ? n80884 : n80891;
  assign n80893 = pi17 ? n2839 : ~n3050;
  assign n80894 = pi16 ? n32 : n80893;
  assign n80895 = pi17 ? n2850 : ~n2952;
  assign n80896 = pi16 ? n32 : n80895;
  assign n80897 = pi15 ? n80894 : n80896;
  assign n80898 = pi14 ? n80892 : n80897;
  assign n80899 = pi17 ? n2724 : ~n3175;
  assign n80900 = pi16 ? n32 : n80899;
  assign n80901 = pi15 ? n80896 : n80900;
  assign n80902 = pi17 ? n2724 : ~n3182;
  assign n80903 = pi16 ? n32 : n80902;
  assign n80904 = pi15 ? n80900 : n80903;
  assign n80905 = pi14 ? n80901 : n80904;
  assign n80906 = pi13 ? n80898 : n80905;
  assign n80907 = pi17 ? n2731 : ~n3182;
  assign n80908 = pi16 ? n32 : n80907;
  assign n80909 = pi15 ? n80903 : n80908;
  assign n80910 = pi17 ? n2731 : ~n2831;
  assign n80911 = pi16 ? n32 : n80910;
  assign n80912 = pi17 ? n2623 : ~n2733;
  assign n80913 = pi16 ? n32 : n80912;
  assign n80914 = pi15 ? n80911 : n80913;
  assign n80915 = pi14 ? n80909 : n80914;
  assign n80916 = pi17 ? n2736 : ~n2839;
  assign n80917 = pi16 ? n32 : n80916;
  assign n80918 = pi15 ? n80913 : n80917;
  assign n80919 = pi17 ? n2736 : ~n2850;
  assign n80920 = pi16 ? n32 : n80919;
  assign n80921 = pi17 ? n2616 : ~n2850;
  assign n80922 = pi16 ? n32 : n80921;
  assign n80923 = pi15 ? n80920 : n80922;
  assign n80924 = pi14 ? n80918 : n80923;
  assign n80925 = pi13 ? n80915 : n80924;
  assign n80926 = pi12 ? n80906 : n80925;
  assign n80927 = pi15 ? n80922 : n8871;
  assign n80928 = pi14 ? n80927 : n69504;
  assign n80929 = pi14 ? n8883 : n8889;
  assign n80930 = pi13 ? n80928 : n80929;
  assign n80931 = pi17 ? n4245 : ~n2623;
  assign n80932 = pi16 ? n32 : n80931;
  assign n80933 = pi15 ? n80932 : n8894;
  assign n80934 = pi17 ? n4245 : ~n2618;
  assign n80935 = pi16 ? n32 : n80934;
  assign n80936 = pi17 ? n3067 : ~n2618;
  assign n80937 = pi16 ? n32 : n80936;
  assign n80938 = pi15 ? n80935 : n80937;
  assign n80939 = pi14 ? n80933 : n80938;
  assign n80940 = pi17 ? n3067 : ~n2628;
  assign n80941 = pi16 ? n32 : n80940;
  assign n80942 = pi15 ? n80941 : n8905;
  assign n80943 = pi14 ? n80942 : n8913;
  assign n80944 = pi13 ? n80939 : n80943;
  assign n80945 = pi12 ? n80930 : n80944;
  assign n80946 = pi11 ? n80926 : n80945;
  assign n80947 = pi10 ? n80889 : n80946;
  assign n80948 = pi09 ? n80830 : n80947;
  assign n80949 = pi08 ? n80818 : n80948;
  assign n80950 = pi07 ? n80679 : n80949;
  assign n80951 = pi18 ? n418 : ~n936;
  assign n80952 = pi17 ? n32 : n80951;
  assign n80953 = pi16 ? n32 : n80952;
  assign n80954 = pi15 ? n32 : n80953;
  assign n80955 = pi18 ? n418 : ~n1575;
  assign n80956 = pi17 ? n32 : n80955;
  assign n80957 = pi16 ? n32 : n80956;
  assign n80958 = pi14 ? n80954 : n80957;
  assign n80959 = pi13 ? n32 : n80958;
  assign n80960 = pi12 ? n32 : n80959;
  assign n80961 = pi11 ? n32 : n80960;
  assign n80962 = pi10 ? n32 : n80961;
  assign n80963 = pi18 ? n3786 : ~n1575;
  assign n80964 = pi17 ? n32 : n80963;
  assign n80965 = pi16 ? n32 : n80964;
  assign n80966 = pi15 ? n80965 : n80686;
  assign n80967 = pi14 ? n80966 : n80689;
  assign n80968 = pi15 ? n80689 : n80836;
  assign n80969 = pi15 ? n80836 : n80701;
  assign n80970 = pi14 ? n80968 : n80969;
  assign n80971 = pi13 ? n80967 : n80970;
  assign n80972 = pi14 ? n80701 : n80704;
  assign n80973 = pi17 ? n3155 : ~n3155;
  assign n80974 = pi16 ? n32 : n80973;
  assign n80975 = pi15 ? n80974 : n80323;
  assign n80976 = pi14 ? n80975 : n80586;
  assign n80977 = pi13 ? n80972 : n80976;
  assign n80978 = pi12 ? n80971 : n80977;
  assign n80979 = pi17 ? n3160 : ~n2954;
  assign n80980 = pi16 ? n32 : n80979;
  assign n80981 = pi15 ? n80585 : n80980;
  assign n80982 = pi17 ? n3164 : ~n2954;
  assign n80983 = pi16 ? n32 : n80982;
  assign n80984 = pi17 ? n3164 : ~n4111;
  assign n80985 = pi16 ? n32 : n80984;
  assign n80986 = pi15 ? n80983 : n80985;
  assign n80987 = pi14 ? n80981 : n80986;
  assign n80988 = pi17 ? n3046 : ~n4111;
  assign n80989 = pi16 ? n32 : n80988;
  assign n80990 = pi17 ? n3292 : ~n3160;
  assign n80991 = pi16 ? n32 : n80990;
  assign n80992 = pi15 ? n80989 : n80991;
  assign n80993 = pi14 ? n80985 : n80992;
  assign n80994 = pi13 ? n80987 : n80993;
  assign n80995 = pi17 ? n2952 : ~n3160;
  assign n80996 = pi16 ? n32 : n80995;
  assign n80997 = pi17 ? n2952 : ~n3046;
  assign n80998 = pi16 ? n32 : n80997;
  assign n80999 = pi14 ? n80996 : n80998;
  assign n81000 = pi17 ? n2952 : ~n3292;
  assign n81001 = pi16 ? n32 : n81000;
  assign n81002 = pi17 ? n2726 : ~n3292;
  assign n81003 = pi16 ? n32 : n81002;
  assign n81004 = pi15 ? n81001 : n81003;
  assign n81005 = pi17 ? n2963 : ~n3587;
  assign n81006 = pi16 ? n32 : n81005;
  assign n81007 = pi14 ? n81004 : n81006;
  assign n81008 = pi13 ? n80999 : n81007;
  assign n81009 = pi12 ? n80994 : n81008;
  assign n81010 = pi11 ? n80978 : n81009;
  assign n81011 = pi17 ? n2963 : ~n3050;
  assign n81012 = pi16 ? n32 : n81011;
  assign n81013 = pi15 ? n81006 : n81012;
  assign n81014 = pi17 ? n3182 : ~n2952;
  assign n81015 = pi16 ? n32 : n81014;
  assign n81016 = pi15 ? n81012 : n81015;
  assign n81017 = pi14 ? n81013 : n81016;
  assign n81018 = pi17 ? n2831 : ~n3175;
  assign n81019 = pi16 ? n32 : n81018;
  assign n81020 = pi15 ? n81015 : n81019;
  assign n81021 = pi17 ? n2831 : ~n3182;
  assign n81022 = pi16 ? n32 : n81021;
  assign n81023 = pi15 ? n9100 : n81022;
  assign n81024 = pi14 ? n81020 : n81023;
  assign n81025 = pi13 ? n81017 : n81024;
  assign n81026 = pi17 ? n2839 : ~n3182;
  assign n81027 = pi16 ? n32 : n81026;
  assign n81028 = pi17 ? n2733 : ~n3182;
  assign n81029 = pi16 ? n32 : n81028;
  assign n81030 = pi15 ? n81027 : n81029;
  assign n81031 = pi17 ? n2733 : ~n2831;
  assign n81032 = pi16 ? n32 : n81031;
  assign n81033 = pi15 ? n81032 : n9121;
  assign n81034 = pi14 ? n81030 : n81033;
  assign n81035 = pi17 ? n2850 : ~n2839;
  assign n81036 = pi16 ? n32 : n81035;
  assign n81037 = pi15 ? n9121 : n81036;
  assign n81038 = pi17 ? n2850 : ~n2850;
  assign n81039 = pi16 ? n32 : n81038;
  assign n81040 = pi17 ? n3067 : ~n2850;
  assign n81041 = pi16 ? n32 : n81040;
  assign n81042 = pi15 ? n81039 : n81041;
  assign n81043 = pi14 ? n81037 : n81042;
  assign n81044 = pi13 ? n81034 : n81043;
  assign n81045 = pi12 ? n81025 : n81044;
  assign n81046 = pi15 ? n81041 : n50986;
  assign n81047 = pi14 ? n81046 : n9142;
  assign n81048 = pi17 ? n2836 : ~n2616;
  assign n81049 = pi16 ? n32 : n81048;
  assign n81050 = pi15 ? n9145 : n81049;
  assign n81051 = pi14 ? n81050 : n9152;
  assign n81052 = pi13 ? n81047 : n81051;
  assign n81053 = pi17 ? n2733 : ~n2623;
  assign n81054 = pi16 ? n32 : n81053;
  assign n81055 = pi15 ? n81054 : n9157;
  assign n81056 = pi14 ? n81055 : n9162;
  assign n81057 = pi17 ? n2726 : ~n2517;
  assign n81058 = pi16 ? n32 : n81057;
  assign n81059 = pi15 ? n81058 : n9177;
  assign n81060 = pi14 ? n9168 : n81059;
  assign n81061 = pi13 ? n81056 : n81060;
  assign n81062 = pi12 ? n81052 : n81061;
  assign n81063 = pi11 ? n81045 : n81062;
  assign n81064 = pi10 ? n81010 : n81063;
  assign n81065 = pi09 ? n80962 : n81064;
  assign n81066 = pi18 ? n797 : ~n936;
  assign n81067 = pi17 ? n32 : n81066;
  assign n81068 = pi16 ? n32 : n81067;
  assign n81069 = pi15 ? n32 : n81068;
  assign n81070 = pi18 ? n797 : ~n1575;
  assign n81071 = pi17 ? n32 : n81070;
  assign n81072 = pi16 ? n32 : n81071;
  assign n81073 = pi14 ? n81069 : n81072;
  assign n81074 = pi13 ? n32 : n81073;
  assign n81075 = pi12 ? n32 : n81074;
  assign n81076 = pi11 ? n32 : n81075;
  assign n81077 = pi10 ? n32 : n81076;
  assign n81078 = pi18 ? n605 : ~n1575;
  assign n81079 = pi17 ? n32 : n81078;
  assign n81080 = pi16 ? n32 : n81079;
  assign n81081 = pi15 ? n81080 : n80825;
  assign n81082 = pi14 ? n81081 : n80825;
  assign n81083 = pi18 ? n344 : ~n1575;
  assign n81084 = pi17 ? n32 : n81083;
  assign n81085 = pi16 ? n32 : n81084;
  assign n81086 = pi15 ? n81085 : n80840;
  assign n81087 = pi14 ? n80833 : n81086;
  assign n81088 = pi13 ? n81082 : n81087;
  assign n81089 = pi14 ? n80844 : n80843;
  assign n81090 = pi18 ? n1676 : ~n2142;
  assign n81091 = pi17 ? n32 : n81090;
  assign n81092 = pi16 ? n32 : n81091;
  assign n81093 = pi17 ? n32 : ~n3155;
  assign n81094 = pi16 ? n32 : n81093;
  assign n81095 = pi15 ? n81092 : n81094;
  assign n81096 = pi14 ? n81095 : n81094;
  assign n81097 = pi13 ? n81089 : n81096;
  assign n81098 = pi12 ? n81088 : n81097;
  assign n81099 = pi17 ? n3282 : ~n2954;
  assign n81100 = pi16 ? n32 : n81099;
  assign n81101 = pi17 ? n3155 : ~n2954;
  assign n81102 = pi16 ? n32 : n81101;
  assign n81103 = pi17 ? n3155 : ~n4111;
  assign n81104 = pi16 ? n32 : n81103;
  assign n81105 = pi15 ? n81102 : n81104;
  assign n81106 = pi14 ? n81100 : n81105;
  assign n81107 = pi17 ? n2954 : ~n4111;
  assign n81108 = pi16 ? n32 : n81107;
  assign n81109 = pi15 ? n81104 : n81108;
  assign n81110 = pi17 ? n4111 : ~n3160;
  assign n81111 = pi16 ? n32 : n81110;
  assign n81112 = pi15 ? n81108 : n81111;
  assign n81113 = pi14 ? n81109 : n81112;
  assign n81114 = pi13 ? n81106 : n81113;
  assign n81115 = pi17 ? n3160 : ~n3160;
  assign n81116 = pi16 ? n32 : n81115;
  assign n81117 = pi17 ? n3160 : ~n3046;
  assign n81118 = pi16 ? n32 : n81117;
  assign n81119 = pi14 ? n81116 : n81118;
  assign n81120 = pi17 ? n3164 : ~n3292;
  assign n81121 = pi16 ? n32 : n81120;
  assign n81122 = pi17 ? n3046 : ~n3292;
  assign n81123 = pi16 ? n32 : n81122;
  assign n81124 = pi15 ? n81121 : n81123;
  assign n81125 = pi17 ? n2959 : ~n3587;
  assign n81126 = pi16 ? n32 : n81125;
  assign n81127 = pi14 ? n81124 : n81126;
  assign n81128 = pi13 ? n81119 : n81127;
  assign n81129 = pi12 ? n81114 : n81128;
  assign n81130 = pi11 ? n81098 : n81129;
  assign n81131 = pi17 ? n2959 : ~n3050;
  assign n81132 = pi16 ? n32 : n81131;
  assign n81133 = pi17 ? n2952 : ~n2952;
  assign n81134 = pi16 ? n32 : n81133;
  assign n81135 = pi15 ? n81132 : n81134;
  assign n81136 = pi14 ? n81132 : n81135;
  assign n81137 = pi17 ? n3175 : ~n3175;
  assign n81138 = pi16 ? n32 : n81137;
  assign n81139 = pi17 ? n3175 : ~n3182;
  assign n81140 = pi16 ? n32 : n81139;
  assign n81141 = pi15 ? n81138 : n81140;
  assign n81142 = pi14 ? n81138 : n81141;
  assign n81143 = pi13 ? n81136 : n81142;
  assign n81144 = pi17 ? n3175 : ~n2831;
  assign n81145 = pi16 ? n32 : n81144;
  assign n81146 = pi15 ? n81145 : n9381;
  assign n81147 = pi14 ? n81140 : n81146;
  assign n81148 = pi17 ? n2831 : ~n2839;
  assign n81149 = pi16 ? n32 : n81148;
  assign n81150 = pi15 ? n9381 : n81149;
  assign n81151 = pi15 ? n9388 : n9396;
  assign n81152 = pi14 ? n81150 : n81151;
  assign n81153 = pi13 ? n81147 : n81152;
  assign n81154 = pi12 ? n81143 : n81153;
  assign n81155 = pi17 ? n2963 : ~n4245;
  assign n81156 = pi16 ? n32 : n81155;
  assign n81157 = pi15 ? n9396 : n81156;
  assign n81158 = pi14 ? n81157 : n9400;
  assign n81159 = pi17 ? n2726 : ~n2616;
  assign n81160 = pi16 ? n32 : n81159;
  assign n81161 = pi15 ? n9403 : n81160;
  assign n81162 = pi15 ? n81160 : n9415;
  assign n81163 = pi14 ? n81161 : n81162;
  assign n81164 = pi13 ? n81158 : n81163;
  assign n81165 = pi17 ? n3046 : ~n2517;
  assign n81166 = pi16 ? n32 : n81165;
  assign n81167 = pi15 ? n81166 : n9435;
  assign n81168 = pi14 ? n9424 : n81167;
  assign n81169 = pi13 ? n9422 : n81168;
  assign n81170 = pi12 ? n81164 : n81169;
  assign n81171 = pi11 ? n81154 : n81170;
  assign n81172 = pi10 ? n81130 : n81171;
  assign n81173 = pi09 ? n81077 : n81172;
  assign n81174 = pi08 ? n81065 : n81173;
  assign n81175 = pi18 ? n2627 : ~n936;
  assign n81176 = pi17 ? n32 : n81175;
  assign n81177 = pi16 ? n32 : n81176;
  assign n81178 = pi15 ? n32 : n81177;
  assign n81179 = pi18 ? n2627 : ~n1575;
  assign n81180 = pi17 ? n32 : n81179;
  assign n81181 = pi16 ? n32 : n81180;
  assign n81182 = pi15 ? n81181 : n81080;
  assign n81183 = pi14 ? n81178 : n81182;
  assign n81184 = pi13 ? n32 : n81183;
  assign n81185 = pi12 ? n32 : n81184;
  assign n81186 = pi11 ? n32 : n81185;
  assign n81187 = pi10 ? n32 : n81186;
  assign n81188 = pi18 ? n2424 : ~n1575;
  assign n81189 = pi17 ? n32 : n81188;
  assign n81190 = pi16 ? n32 : n81189;
  assign n81191 = pi15 ? n81190 : n80957;
  assign n81192 = pi15 ? n80957 : n80965;
  assign n81193 = pi14 ? n81191 : n81192;
  assign n81194 = pi18 ? n532 : ~n1575;
  assign n81195 = pi17 ? n32 : n81194;
  assign n81196 = pi16 ? n32 : n81195;
  assign n81197 = pi15 ? n81196 : n80686;
  assign n81198 = pi14 ? n80965 : n81197;
  assign n81199 = pi13 ? n81193 : n81198;
  assign n81200 = pi14 ? n80689 : n80968;
  assign n81201 = pi18 ? n1942 : ~n2142;
  assign n81202 = pi17 ? n32 : n81201;
  assign n81203 = pi16 ? n32 : n81202;
  assign n81204 = pi18 ? n237 : ~n2142;
  assign n81205 = pi17 ? n32 : n81204;
  assign n81206 = pi16 ? n32 : n81205;
  assign n81207 = pi15 ? n81203 : n81206;
  assign n81208 = pi18 ? n618 : ~n2142;
  assign n81209 = pi17 ? n32 : n81208;
  assign n81210 = pi16 ? n32 : n81209;
  assign n81211 = pi15 ? n81206 : n81210;
  assign n81212 = pi14 ? n81207 : n81211;
  assign n81213 = pi13 ? n81200 : n81212;
  assign n81214 = pi12 ? n81199 : n81213;
  assign n81215 = pi18 ? n618 : ~n863;
  assign n81216 = pi17 ? n32 : n81215;
  assign n81217 = pi16 ? n32 : n81216;
  assign n81218 = pi18 ? n1676 : ~n863;
  assign n81219 = pi17 ? n32 : n81218;
  assign n81220 = pi16 ? n32 : n81219;
  assign n81221 = pi18 ? n1676 : ~n1592;
  assign n81222 = pi17 ? n32 : n81221;
  assign n81223 = pi16 ? n32 : n81222;
  assign n81224 = pi15 ? n81220 : n81223;
  assign n81225 = pi14 ? n81217 : n81224;
  assign n81226 = pi17 ? n3569 : ~n4111;
  assign n81227 = pi16 ? n32 : n81226;
  assign n81228 = pi17 ? n3569 : ~n3160;
  assign n81229 = pi16 ? n32 : n81228;
  assign n81230 = pi15 ? n81227 : n81229;
  assign n81231 = pi14 ? n81223 : n81230;
  assign n81232 = pi13 ? n81225 : n81231;
  assign n81233 = pi17 ? n3282 : ~n3160;
  assign n81234 = pi16 ? n32 : n81233;
  assign n81235 = pi17 ? n3282 : ~n3046;
  assign n81236 = pi16 ? n32 : n81235;
  assign n81237 = pi17 ? n3155 : ~n3046;
  assign n81238 = pi16 ? n32 : n81237;
  assign n81239 = pi15 ? n81236 : n81238;
  assign n81240 = pi14 ? n81234 : n81239;
  assign n81241 = pi17 ? n3155 : ~n3292;
  assign n81242 = pi16 ? n32 : n81241;
  assign n81243 = pi17 ? n3728 : ~n3292;
  assign n81244 = pi16 ? n32 : n81243;
  assign n81245 = pi15 ? n81242 : n81244;
  assign n81246 = pi17 ? n3728 : ~n3587;
  assign n81247 = pi16 ? n32 : n81246;
  assign n81248 = pi14 ? n81245 : n81247;
  assign n81249 = pi13 ? n81240 : n81248;
  assign n81250 = pi12 ? n81232 : n81249;
  assign n81251 = pi11 ? n81214 : n81250;
  assign n81252 = pi17 ? n3728 : ~n3050;
  assign n81253 = pi16 ? n32 : n81252;
  assign n81254 = pi17 ? n4111 : ~n3050;
  assign n81255 = pi16 ? n32 : n81254;
  assign n81256 = pi17 ? n3160 : ~n2952;
  assign n81257 = pi16 ? n32 : n81256;
  assign n81258 = pi15 ? n81255 : n81257;
  assign n81259 = pi14 ? n81253 : n81258;
  assign n81260 = pi17 ? n3292 : ~n3175;
  assign n81261 = pi16 ? n32 : n81260;
  assign n81262 = pi17 ? n3292 : ~n2963;
  assign n81263 = pi16 ? n32 : n81262;
  assign n81264 = pi17 ? n3292 : ~n3182;
  assign n81265 = pi16 ? n32 : n81264;
  assign n81266 = pi15 ? n81263 : n81265;
  assign n81267 = pi14 ? n81261 : n81266;
  assign n81268 = pi13 ? n81259 : n81267;
  assign n81269 = pi17 ? n3587 : ~n3182;
  assign n81270 = pi16 ? n32 : n81269;
  assign n81271 = pi15 ? n81265 : n81270;
  assign n81272 = pi17 ? n3175 : ~n2733;
  assign n81273 = pi16 ? n32 : n81272;
  assign n81274 = pi14 ? n81271 : n81273;
  assign n81275 = pi17 ? n2959 : ~n2839;
  assign n81276 = pi16 ? n32 : n81275;
  assign n81277 = pi17 ? n3587 : ~n2850;
  assign n81278 = pi16 ? n32 : n81277;
  assign n81279 = pi15 ? n81278 : n9678;
  assign n81280 = pi14 ? n81276 : n81279;
  assign n81281 = pi13 ? n81274 : n81280;
  assign n81282 = pi12 ? n81268 : n81281;
  assign n81283 = pi17 ? n2959 : ~n4245;
  assign n81284 = pi16 ? n32 : n81283;
  assign n81285 = pi15 ? n9678 : n81284;
  assign n81286 = pi14 ? n81285 : n9682;
  assign n81287 = pi15 ? n9681 : n9688;
  assign n81288 = pi14 ? n81287 : n9691;
  assign n81289 = pi13 ? n81286 : n81288;
  assign n81290 = pi15 ? n9690 : n9698;
  assign n81291 = pi14 ? n81290 : n9698;
  assign n81292 = pi13 ? n81291 : n9711;
  assign n81293 = pi12 ? n81289 : n81292;
  assign n81294 = pi11 ? n81282 : n81293;
  assign n81295 = pi10 ? n81251 : n81294;
  assign n81296 = pi09 ? n81187 : n81295;
  assign n81297 = pi18 ? n1750 : ~n936;
  assign n81298 = pi17 ? n32 : n81297;
  assign n81299 = pi16 ? n32 : n81298;
  assign n81300 = pi15 ? n32 : n81299;
  assign n81301 = pi18 ? n2622 : ~n1575;
  assign n81302 = pi17 ? n32 : n81301;
  assign n81303 = pi16 ? n32 : n81302;
  assign n81304 = pi18 ? n323 : ~n1575;
  assign n81305 = pi17 ? n32 : n81304;
  assign n81306 = pi16 ? n32 : n81305;
  assign n81307 = pi15 ? n81303 : n81306;
  assign n81308 = pi14 ? n81300 : n81307;
  assign n81309 = pi13 ? n32 : n81308;
  assign n81310 = pi12 ? n32 : n81309;
  assign n81311 = pi11 ? n32 : n81310;
  assign n81312 = pi10 ? n32 : n81311;
  assign n81313 = pi18 ? n2291 : ~n1575;
  assign n81314 = pi17 ? n32 : n81313;
  assign n81315 = pi16 ? n32 : n81314;
  assign n81316 = pi15 ? n81315 : n81072;
  assign n81317 = pi18 ? n2413 : ~n1575;
  assign n81318 = pi17 ? n32 : n81317;
  assign n81319 = pi16 ? n32 : n81318;
  assign n81320 = pi15 ? n81072 : n81319;
  assign n81321 = pi14 ? n81316 : n81320;
  assign n81322 = pi15 ? n81190 : n80825;
  assign n81323 = pi14 ? n81319 : n81322;
  assign n81324 = pi13 ? n81321 : n81323;
  assign n81325 = pi14 ? n80825 : n80833;
  assign n81326 = pi18 ? n344 : ~n2142;
  assign n81327 = pi17 ? n32 : n81326;
  assign n81328 = pi16 ? n32 : n81327;
  assign n81329 = pi18 ? n1813 : ~n2142;
  assign n81330 = pi17 ? n32 : n81329;
  assign n81331 = pi16 ? n32 : n81330;
  assign n81332 = pi15 ? n81328 : n81331;
  assign n81333 = pi18 ? n814 : ~n2142;
  assign n81334 = pi17 ? n32 : n81333;
  assign n81335 = pi16 ? n32 : n81334;
  assign n81336 = pi14 ? n81332 : n81335;
  assign n81337 = pi13 ? n81325 : n81336;
  assign n81338 = pi12 ? n81324 : n81337;
  assign n81339 = pi18 ? n814 : ~n863;
  assign n81340 = pi17 ? n32 : n81339;
  assign n81341 = pi16 ? n32 : n81340;
  assign n81342 = pi18 ? n1942 : ~n863;
  assign n81343 = pi17 ? n32 : n81342;
  assign n81344 = pi16 ? n32 : n81343;
  assign n81345 = pi15 ? n81341 : n81344;
  assign n81346 = pi18 ? n1942 : ~n1592;
  assign n81347 = pi17 ? n32 : n81346;
  assign n81348 = pi16 ? n32 : n81347;
  assign n81349 = pi15 ? n81344 : n81348;
  assign n81350 = pi14 ? n81345 : n81349;
  assign n81351 = pi18 ? n3350 : ~n1592;
  assign n81352 = pi17 ? n32 : n81351;
  assign n81353 = pi16 ? n32 : n81352;
  assign n81354 = pi15 ? n81348 : n81353;
  assign n81355 = pi18 ? n3350 : ~n1841;
  assign n81356 = pi17 ? n32 : n81355;
  assign n81357 = pi16 ? n32 : n81356;
  assign n81358 = pi15 ? n81353 : n81357;
  assign n81359 = pi14 ? n81354 : n81358;
  assign n81360 = pi13 ? n81350 : n81359;
  assign n81361 = pi18 ? n618 : ~n1841;
  assign n81362 = pi17 ? n32 : n81361;
  assign n81363 = pi16 ? n32 : n81362;
  assign n81364 = pi18 ? n618 : ~n1477;
  assign n81365 = pi17 ? n32 : n81364;
  assign n81366 = pi16 ? n32 : n81365;
  assign n81367 = pi14 ? n81363 : n81366;
  assign n81368 = pi17 ? n32 : ~n3292;
  assign n81369 = pi16 ? n32 : n81368;
  assign n81370 = pi17 ? n32 : ~n3587;
  assign n81371 = pi16 ? n32 : n81370;
  assign n81372 = pi14 ? n81369 : n81371;
  assign n81373 = pi13 ? n81367 : n81372;
  assign n81374 = pi12 ? n81360 : n81373;
  assign n81375 = pi11 ? n81338 : n81374;
  assign n81376 = pi17 ? n32 : ~n3050;
  assign n81377 = pi16 ? n32 : n81376;
  assign n81378 = pi17 ? n3569 : ~n3050;
  assign n81379 = pi16 ? n32 : n81378;
  assign n81380 = pi15 ? n81377 : n81379;
  assign n81381 = pi17 ? n4111 : ~n2952;
  assign n81382 = pi16 ? n32 : n81381;
  assign n81383 = pi15 ? n81379 : n81382;
  assign n81384 = pi14 ? n81380 : n81383;
  assign n81385 = pi17 ? n3155 : ~n3175;
  assign n81386 = pi16 ? n32 : n81385;
  assign n81387 = pi17 ? n4111 : ~n3175;
  assign n81388 = pi16 ? n32 : n81387;
  assign n81389 = pi15 ? n81386 : n81388;
  assign n81390 = pi17 ? n3155 : ~n2963;
  assign n81391 = pi16 ? n32 : n81390;
  assign n81392 = pi17 ? n3155 : ~n3182;
  assign n81393 = pi16 ? n32 : n81392;
  assign n81394 = pi15 ? n81391 : n81393;
  assign n81395 = pi14 ? n81389 : n81394;
  assign n81396 = pi13 ? n81384 : n81395;
  assign n81397 = pi17 ? n2954 : ~n3182;
  assign n81398 = pi16 ? n32 : n81397;
  assign n81399 = pi17 ? n3164 : ~n2733;
  assign n81400 = pi16 ? n32 : n81399;
  assign n81401 = pi14 ? n81398 : n81400;
  assign n81402 = pi17 ? n3160 : ~n2839;
  assign n81403 = pi16 ? n32 : n81402;
  assign n81404 = pi17 ? n3160 : ~n2850;
  assign n81405 = pi16 ? n32 : n81404;
  assign n81406 = pi17 ? n3164 : ~n2850;
  assign n81407 = pi16 ? n32 : n81406;
  assign n81408 = pi15 ? n81405 : n81407;
  assign n81409 = pi14 ? n81403 : n81408;
  assign n81410 = pi13 ? n81401 : n81409;
  assign n81411 = pi12 ? n81396 : n81410;
  assign n81412 = pi14 ? n9949 : n9955;
  assign n81413 = pi15 ? n9958 : n9965;
  assign n81414 = pi14 ? n9959 : n81413;
  assign n81415 = pi13 ? n81412 : n81414;
  assign n81416 = pi17 ? n2954 : ~n4099;
  assign n81417 = pi16 ? n32 : n81416;
  assign n81418 = pi15 ? n81417 : n9970;
  assign n81419 = pi17 ? n3569 : ~n2618;
  assign n81420 = pi16 ? n32 : n81419;
  assign n81421 = pi14 ? n81418 : n81420;
  assign n81422 = pi13 ? n81421 : n9988;
  assign n81423 = pi12 ? n81415 : n81422;
  assign n81424 = pi11 ? n81411 : n81423;
  assign n81425 = pi10 ? n81375 : n81424;
  assign n81426 = pi09 ? n81312 : n81425;
  assign n81427 = pi08 ? n81296 : n81426;
  assign n81428 = pi07 ? n81174 : n81427;
  assign n81429 = pi06 ? n80950 : n81428;
  assign n81430 = pi05 ? n80453 : n81429;
  assign n81431 = pi18 ? n962 : ~n936;
  assign n81432 = pi17 ? n32 : n81431;
  assign n81433 = pi16 ? n32 : n81432;
  assign n81434 = pi15 ? n32 : n81433;
  assign n81435 = pi18 ? n2730 : ~n1575;
  assign n81436 = pi17 ? n32 : n81435;
  assign n81437 = pi16 ? n32 : n81436;
  assign n81438 = pi18 ? n702 : ~n1575;
  assign n81439 = pi17 ? n32 : n81438;
  assign n81440 = pi16 ? n32 : n81439;
  assign n81441 = pi15 ? n81437 : n81440;
  assign n81442 = pi14 ? n81434 : n81441;
  assign n81443 = pi13 ? n32 : n81442;
  assign n81444 = pi12 ? n32 : n81443;
  assign n81445 = pi11 ? n32 : n81444;
  assign n81446 = pi10 ? n32 : n81445;
  assign n81447 = pi18 ? n4098 : ~n1575;
  assign n81448 = pi17 ? n32 : n81447;
  assign n81449 = pi16 ? n32 : n81448;
  assign n81450 = pi18 ? n595 : ~n1575;
  assign n81451 = pi17 ? n32 : n81450;
  assign n81452 = pi16 ? n32 : n81451;
  assign n81453 = pi15 ? n81449 : n81452;
  assign n81454 = pi15 ? n81452 : n81181;
  assign n81455 = pi14 ? n81453 : n81454;
  assign n81456 = pi18 ? n508 : ~n1575;
  assign n81457 = pi17 ? n32 : n81456;
  assign n81458 = pi16 ? n32 : n81457;
  assign n81459 = pi14 ? n81458 : n81191;
  assign n81460 = pi13 ? n81455 : n81459;
  assign n81461 = pi14 ? n80957 : n80965;
  assign n81462 = pi18 ? n532 : ~n2142;
  assign n81463 = pi17 ? n32 : n81462;
  assign n81464 = pi16 ? n32 : n81463;
  assign n81465 = pi18 ? n2298 : ~n2142;
  assign n81466 = pi17 ? n32 : n81465;
  assign n81467 = pi16 ? n32 : n81466;
  assign n81468 = pi15 ? n81464 : n81467;
  assign n81469 = pi18 ? n430 : ~n2142;
  assign n81470 = pi17 ? n32 : n81469;
  assign n81471 = pi16 ? n32 : n81470;
  assign n81472 = pi14 ? n81468 : n81471;
  assign n81473 = pi13 ? n81461 : n81472;
  assign n81474 = pi12 ? n81460 : n81473;
  assign n81475 = pi18 ? n430 : ~n863;
  assign n81476 = pi17 ? n32 : n81475;
  assign n81477 = pi16 ? n32 : n81476;
  assign n81478 = pi18 ? n2304 : ~n863;
  assign n81479 = pi17 ? n32 : n81478;
  assign n81480 = pi16 ? n32 : n81479;
  assign n81481 = pi15 ? n81477 : n81480;
  assign n81482 = pi18 ? n344 : ~n1592;
  assign n81483 = pi17 ? n32 : n81482;
  assign n81484 = pi16 ? n32 : n81483;
  assign n81485 = pi15 ? n81480 : n81484;
  assign n81486 = pi14 ? n81481 : n81485;
  assign n81487 = pi18 ? n350 : ~n1592;
  assign n81488 = pi17 ? n32 : n81487;
  assign n81489 = pi16 ? n32 : n81488;
  assign n81490 = pi18 ? n1813 : ~n1592;
  assign n81491 = pi17 ? n32 : n81490;
  assign n81492 = pi16 ? n32 : n81491;
  assign n81493 = pi15 ? n81489 : n81492;
  assign n81494 = pi18 ? n1813 : ~n1841;
  assign n81495 = pi17 ? n32 : n81494;
  assign n81496 = pi16 ? n32 : n81495;
  assign n81497 = pi15 ? n81492 : n81496;
  assign n81498 = pi14 ? n81493 : n81497;
  assign n81499 = pi13 ? n81486 : n81498;
  assign n81500 = pi18 ? n814 : ~n1841;
  assign n81501 = pi17 ? n32 : n81500;
  assign n81502 = pi16 ? n32 : n81501;
  assign n81503 = pi18 ? n814 : ~n1477;
  assign n81504 = pi17 ? n32 : n81503;
  assign n81505 = pi16 ? n32 : n81504;
  assign n81506 = pi15 ? n81502 : n81505;
  assign n81507 = pi14 ? n81506 : n81505;
  assign n81508 = pi18 ? n237 : ~n751;
  assign n81509 = pi17 ? n32 : n81508;
  assign n81510 = pi16 ? n32 : n81509;
  assign n81511 = pi15 ? n81510 : n10136;
  assign n81512 = pi14 ? n81511 : n10136;
  assign n81513 = pi13 ? n81507 : n81512;
  assign n81514 = pi12 ? n81499 : n81513;
  assign n81515 = pi11 ? n81474 : n81514;
  assign n81516 = pi18 ? n618 : ~n341;
  assign n81517 = pi17 ? n32 : n81516;
  assign n81518 = pi16 ? n32 : n81517;
  assign n81519 = pi15 ? n10147 : n81518;
  assign n81520 = pi14 ? n10147 : n81519;
  assign n81521 = pi18 ? n618 : ~n2962;
  assign n81522 = pi17 ? n32 : n81521;
  assign n81523 = pi16 ? n32 : n81522;
  assign n81524 = pi18 ? n618 : ~n1965;
  assign n81525 = pi17 ? n32 : n81524;
  assign n81526 = pi16 ? n32 : n81525;
  assign n81527 = pi15 ? n81523 : n81526;
  assign n81528 = pi14 ? n10157 : n81527;
  assign n81529 = pi13 ? n81520 : n81528;
  assign n81530 = pi18 ? n1676 : ~n1965;
  assign n81531 = pi17 ? n32 : n81530;
  assign n81532 = pi16 ? n32 : n81531;
  assign n81533 = pi17 ? n3155 : ~n2733;
  assign n81534 = pi16 ? n32 : n81533;
  assign n81535 = pi14 ? n81532 : n81534;
  assign n81536 = pi17 ? n3155 : ~n2839;
  assign n81537 = pi16 ? n32 : n81536;
  assign n81538 = pi17 ? n32 : ~n2839;
  assign n81539 = pi16 ? n32 : n81538;
  assign n81540 = pi15 ? n81537 : n81539;
  assign n81541 = pi17 ? n3569 : ~n2850;
  assign n81542 = pi16 ? n32 : n81541;
  assign n81543 = pi15 ? n10199 : n81542;
  assign n81544 = pi14 ? n81540 : n81543;
  assign n81545 = pi13 ? n81535 : n81544;
  assign n81546 = pi12 ? n81529 : n81545;
  assign n81547 = pi17 ? n3569 : ~n4245;
  assign n81548 = pi16 ? n32 : n81547;
  assign n81549 = pi14 ? n81548 : n10219;
  assign n81550 = pi15 ? n10226 : n10235;
  assign n81551 = pi14 ? n10223 : n81550;
  assign n81552 = pi13 ? n81549 : n81551;
  assign n81553 = pi17 ? n32 : n48014;
  assign n81554 = pi16 ? n32 : n81553;
  assign n81555 = pi18 ? n1813 : ~n2754;
  assign n81556 = pi17 ? n32 : n81555;
  assign n81557 = pi16 ? n32 : n81556;
  assign n81558 = pi15 ? n81554 : n81557;
  assign n81559 = pi14 ? n81558 : n10250;
  assign n81560 = pi13 ? n10244 : n81559;
  assign n81561 = pi12 ? n81552 : n81560;
  assign n81562 = pi11 ? n81546 : n81561;
  assign n81563 = pi10 ? n81515 : n81562;
  assign n81564 = pi09 ? n81446 : n81563;
  assign n81565 = pi18 ? n590 : ~n936;
  assign n81566 = pi17 ? n32 : n81565;
  assign n81567 = pi16 ? n32 : n81566;
  assign n81568 = pi15 ? n32 : n81567;
  assign n81569 = pi18 ? n2849 : ~n1575;
  assign n81570 = pi17 ? n32 : n81569;
  assign n81571 = pi16 ? n32 : n81570;
  assign n81572 = pi18 ? n697 : ~n1575;
  assign n81573 = pi17 ? n32 : n81572;
  assign n81574 = pi16 ? n32 : n81573;
  assign n81575 = pi15 ? n81571 : n81574;
  assign n81576 = pi14 ? n81568 : n81575;
  assign n81577 = pi13 ? n32 : n81576;
  assign n81578 = pi12 ? n32 : n81577;
  assign n81579 = pi11 ? n32 : n81578;
  assign n81580 = pi10 ? n32 : n81579;
  assign n81581 = pi18 ? n2615 : ~n1575;
  assign n81582 = pi17 ? n32 : n81581;
  assign n81583 = pi16 ? n32 : n81582;
  assign n81584 = pi18 ? n1750 : ~n1575;
  assign n81585 = pi17 ? n32 : n81584;
  assign n81586 = pi16 ? n32 : n81585;
  assign n81587 = pi15 ? n81583 : n81586;
  assign n81588 = pi15 ? n81586 : n81303;
  assign n81589 = pi14 ? n81587 : n81588;
  assign n81590 = pi15 ? n81303 : n81440;
  assign n81591 = pi14 ? n81590 : n81316;
  assign n81592 = pi13 ? n81589 : n81591;
  assign n81593 = pi14 ? n81072 : n81319;
  assign n81594 = pi18 ? n2413 : ~n2142;
  assign n81595 = pi17 ? n32 : n81594;
  assign n81596 = pi16 ? n32 : n81595;
  assign n81597 = pi18 ? n2424 : ~n2142;
  assign n81598 = pi17 ? n32 : n81597;
  assign n81599 = pi16 ? n32 : n81598;
  assign n81600 = pi15 ? n81596 : n81599;
  assign n81601 = pi18 ? n418 : ~n2142;
  assign n81602 = pi17 ? n32 : n81601;
  assign n81603 = pi16 ? n32 : n81602;
  assign n81604 = pi14 ? n81600 : n81603;
  assign n81605 = pi13 ? n81593 : n81604;
  assign n81606 = pi12 ? n81592 : n81605;
  assign n81607 = pi18 ? n418 : ~n863;
  assign n81608 = pi17 ? n32 : n81607;
  assign n81609 = pi16 ? n32 : n81608;
  assign n81610 = pi18 ? n3786 : ~n863;
  assign n81611 = pi17 ? n32 : n81610;
  assign n81612 = pi16 ? n32 : n81611;
  assign n81613 = pi15 ? n81609 : n81612;
  assign n81614 = pi18 ? n532 : ~n1592;
  assign n81615 = pi17 ? n32 : n81614;
  assign n81616 = pi16 ? n32 : n81615;
  assign n81617 = pi15 ? n81612 : n81616;
  assign n81618 = pi14 ? n81613 : n81617;
  assign n81619 = pi18 ? n2298 : ~n1592;
  assign n81620 = pi17 ? n32 : n81619;
  assign n81621 = pi16 ? n32 : n81620;
  assign n81622 = pi15 ? n81616 : n81621;
  assign n81623 = pi18 ? n2298 : ~n1841;
  assign n81624 = pi17 ? n32 : n81623;
  assign n81625 = pi16 ? n32 : n81624;
  assign n81626 = pi15 ? n81621 : n81625;
  assign n81627 = pi14 ? n81622 : n81626;
  assign n81628 = pi13 ? n81618 : n81627;
  assign n81629 = pi18 ? n430 : ~n1841;
  assign n81630 = pi17 ? n32 : n81629;
  assign n81631 = pi16 ? n32 : n81630;
  assign n81632 = pi18 ? n430 : ~n1477;
  assign n81633 = pi17 ? n32 : n81632;
  assign n81634 = pi16 ? n32 : n81633;
  assign n81635 = pi15 ? n81631 : n81634;
  assign n81636 = pi18 ? n2304 : ~n1477;
  assign n81637 = pi17 ? n32 : n81636;
  assign n81638 = pi16 ? n32 : n81637;
  assign n81639 = pi18 ? n3336 : ~n1477;
  assign n81640 = pi17 ? n32 : n81639;
  assign n81641 = pi16 ? n32 : n81640;
  assign n81642 = pi15 ? n81638 : n81641;
  assign n81643 = pi14 ? n81635 : n81642;
  assign n81644 = pi18 ? n350 : ~n751;
  assign n81645 = pi17 ? n32 : n81644;
  assign n81646 = pi16 ? n32 : n81645;
  assign n81647 = pi18 ? n350 : ~n1970;
  assign n81648 = pi17 ? n32 : n81647;
  assign n81649 = pi16 ? n32 : n81648;
  assign n81650 = pi15 ? n81646 : n81649;
  assign n81651 = pi15 ? n81649 : n10385;
  assign n81652 = pi14 ? n81650 : n81651;
  assign n81653 = pi13 ? n81643 : n81652;
  assign n81654 = pi12 ? n81628 : n81653;
  assign n81655 = pi11 ? n81606 : n81654;
  assign n81656 = pi15 ? n10385 : n10393;
  assign n81657 = pi14 ? n10385 : n81656;
  assign n81658 = pi18 ? n814 : ~n2962;
  assign n81659 = pi17 ? n32 : n81658;
  assign n81660 = pi16 ? n32 : n81659;
  assign n81661 = pi15 ? n10393 : n81660;
  assign n81662 = pi15 ? n81660 : n10114;
  assign n81663 = pi14 ? n81661 : n81662;
  assign n81664 = pi13 ? n81657 : n81663;
  assign n81665 = pi18 ? n1942 : ~n1965;
  assign n81666 = pi17 ? n32 : n81665;
  assign n81667 = pi16 ? n32 : n81666;
  assign n81668 = pi15 ? n81667 : n10402;
  assign n81669 = pi18 ? n1676 : ~n684;
  assign n81670 = pi17 ? n32 : n81669;
  assign n81671 = pi16 ? n32 : n81670;
  assign n81672 = pi18 ? n237 : ~n590;
  assign n81673 = pi17 ? n32 : n81672;
  assign n81674 = pi16 ? n32 : n81673;
  assign n81675 = pi15 ? n81671 : n81674;
  assign n81676 = pi14 ? n81668 : n81675;
  assign n81677 = pi18 ? n237 : ~n2849;
  assign n81678 = pi17 ? n32 : n81677;
  assign n81679 = pi16 ? n32 : n81678;
  assign n81680 = pi15 ? n10433 : n81679;
  assign n81681 = pi14 ? n10429 : n81680;
  assign n81682 = pi13 ? n81676 : n81681;
  assign n81683 = pi12 ? n81664 : n81682;
  assign n81684 = pi18 ? n237 : ~n4244;
  assign n81685 = pi17 ? n32 : n81684;
  assign n81686 = pi16 ? n32 : n81685;
  assign n81687 = pi18 ? n237 : ~n2730;
  assign n81688 = pi17 ? n32 : n81687;
  assign n81689 = pi16 ? n32 : n81688;
  assign n81690 = pi15 ? n81686 : n81689;
  assign n81691 = pi14 ? n81690 : n10455;
  assign n81692 = pi15 ? n10466 : n10475;
  assign n81693 = pi14 ? n10463 : n81692;
  assign n81694 = pi13 ? n81691 : n81693;
  assign n81695 = pi18 ? n344 : ~n2754;
  assign n81696 = pi17 ? n32 : n81695;
  assign n81697 = pi16 ? n32 : n81696;
  assign n81698 = pi15 ? n10484 : n39445;
  assign n81699 = pi14 ? n81697 : n81698;
  assign n81700 = pi13 ? n10481 : n81699;
  assign n81701 = pi12 ? n81694 : n81700;
  assign n81702 = pi11 ? n81683 : n81701;
  assign n81703 = pi10 ? n81655 : n81702;
  assign n81704 = pi09 ? n81580 : n81703;
  assign n81705 = pi08 ? n81564 : n81704;
  assign n81706 = pi16 ? n32 : n1042;
  assign n81707 = pi15 ? n32 : n81706;
  assign n81708 = pi18 ? n2830 : ~n1575;
  assign n81709 = pi17 ? n32 : n81708;
  assign n81710 = pi16 ? n32 : n81709;
  assign n81711 = pi18 ? n496 : ~n1575;
  assign n81712 = pi17 ? n32 : n81711;
  assign n81713 = pi16 ? n32 : n81712;
  assign n81714 = pi15 ? n81710 : n81713;
  assign n81715 = pi14 ? n81707 : n81714;
  assign n81716 = pi13 ? n32 : n81715;
  assign n81717 = pi12 ? n32 : n81716;
  assign n81718 = pi11 ? n32 : n81717;
  assign n81719 = pi10 ? n32 : n81718;
  assign n81720 = pi18 ? n4244 : ~n1575;
  assign n81721 = pi17 ? n32 : n81720;
  assign n81722 = pi16 ? n32 : n81721;
  assign n81723 = pi18 ? n962 : ~n1575;
  assign n81724 = pi17 ? n32 : n81723;
  assign n81725 = pi16 ? n32 : n81724;
  assign n81726 = pi15 ? n81722 : n81725;
  assign n81727 = pi15 ? n81725 : n81437;
  assign n81728 = pi14 ? n81726 : n81727;
  assign n81729 = pi15 ? n81437 : n81574;
  assign n81730 = pi14 ? n81729 : n81453;
  assign n81731 = pi13 ? n81728 : n81730;
  assign n81732 = pi15 ? n81181 : n81458;
  assign n81733 = pi14 ? n81452 : n81732;
  assign n81734 = pi18 ? n508 : ~n2142;
  assign n81735 = pi17 ? n32 : n81734;
  assign n81736 = pi16 ? n32 : n81735;
  assign n81737 = pi18 ? n2291 : ~n2142;
  assign n81738 = pi17 ? n32 : n81737;
  assign n81739 = pi16 ? n32 : n81738;
  assign n81740 = pi15 ? n81736 : n81739;
  assign n81741 = pi18 ? n797 : ~n2142;
  assign n81742 = pi17 ? n32 : n81741;
  assign n81743 = pi16 ? n32 : n81742;
  assign n81744 = pi14 ? n81740 : n81743;
  assign n81745 = pi13 ? n81733 : n81744;
  assign n81746 = pi12 ? n81731 : n81745;
  assign n81747 = pi18 ? n797 : ~n863;
  assign n81748 = pi17 ? n32 : n81747;
  assign n81749 = pi16 ? n32 : n81748;
  assign n81750 = pi18 ? n2413 : ~n863;
  assign n81751 = pi17 ? n32 : n81750;
  assign n81752 = pi16 ? n32 : n81751;
  assign n81753 = pi15 ? n81749 : n81752;
  assign n81754 = pi18 ? n2413 : ~n1592;
  assign n81755 = pi17 ? n32 : n81754;
  assign n81756 = pi16 ? n32 : n81755;
  assign n81757 = pi15 ? n81752 : n81756;
  assign n81758 = pi14 ? n81753 : n81757;
  assign n81759 = pi18 ? n605 : ~n1592;
  assign n81760 = pi17 ? n32 : n81759;
  assign n81761 = pi16 ? n32 : n81760;
  assign n81762 = pi18 ? n2424 : ~n1592;
  assign n81763 = pi17 ? n32 : n81762;
  assign n81764 = pi16 ? n32 : n81763;
  assign n81765 = pi15 ? n81761 : n81764;
  assign n81766 = pi18 ? n2424 : ~n1841;
  assign n81767 = pi17 ? n32 : n81766;
  assign n81768 = pi16 ? n32 : n81767;
  assign n81769 = pi15 ? n81764 : n81768;
  assign n81770 = pi14 ? n81765 : n81769;
  assign n81771 = pi13 ? n81758 : n81770;
  assign n81772 = pi18 ? n418 : ~n1841;
  assign n81773 = pi17 ? n32 : n81772;
  assign n81774 = pi16 ? n32 : n81773;
  assign n81775 = pi18 ? n418 : ~n1477;
  assign n81776 = pi17 ? n32 : n81775;
  assign n81777 = pi16 ? n32 : n81776;
  assign n81778 = pi15 ? n81774 : n81777;
  assign n81779 = pi18 ? n3786 : ~n1477;
  assign n81780 = pi17 ? n32 : n81779;
  assign n81781 = pi16 ? n32 : n81780;
  assign n81782 = pi14 ? n81778 : n81781;
  assign n81783 = pi18 ? n532 : ~n751;
  assign n81784 = pi17 ? n32 : n81783;
  assign n81785 = pi16 ? n32 : n81784;
  assign n81786 = pi18 ? n532 : ~n1970;
  assign n81787 = pi17 ? n32 : n81786;
  assign n81788 = pi16 ? n32 : n81787;
  assign n81789 = pi15 ? n81785 : n81788;
  assign n81790 = pi18 ? n532 : ~n245;
  assign n81791 = pi17 ? n32 : n81790;
  assign n81792 = pi16 ? n32 : n81791;
  assign n81793 = pi15 ? n81788 : n81792;
  assign n81794 = pi14 ? n81789 : n81793;
  assign n81795 = pi13 ? n81782 : n81794;
  assign n81796 = pi12 ? n81771 : n81795;
  assign n81797 = pi11 ? n81746 : n81796;
  assign n81798 = pi18 ? n2298 : ~n245;
  assign n81799 = pi17 ? n32 : n81798;
  assign n81800 = pi16 ? n32 : n81799;
  assign n81801 = pi15 ? n81792 : n81800;
  assign n81802 = pi15 ? n10623 : n10631;
  assign n81803 = pi14 ? n81801 : n81802;
  assign n81804 = pi18 ? n1548 : ~n2962;
  assign n81805 = pi17 ? n32 : n81804;
  assign n81806 = pi16 ? n32 : n81805;
  assign n81807 = pi15 ? n10631 : n81806;
  assign n81808 = pi15 ? n81806 : n10640;
  assign n81809 = pi14 ? n81807 : n81808;
  assign n81810 = pi13 ? n81803 : n81809;
  assign n81811 = pi15 ? n10640 : n10626;
  assign n81812 = pi18 ? n3336 : ~n684;
  assign n81813 = pi17 ? n32 : n81812;
  assign n81814 = pi16 ? n32 : n81813;
  assign n81815 = pi15 ? n81814 : n10659;
  assign n81816 = pi14 ? n81811 : n81815;
  assign n81817 = pi15 ? n10669 : n50763;
  assign n81818 = pi14 ? n10659 : n81817;
  assign n81819 = pi13 ? n81816 : n81818;
  assign n81820 = pi12 ? n81810 : n81819;
  assign n81821 = pi14 ? n10683 : n10691;
  assign n81822 = pi15 ? n10695 : n10708;
  assign n81823 = pi14 ? n81822 : n10708;
  assign n81824 = pi13 ? n81821 : n81823;
  assign n81825 = pi18 ? n2298 : ~n508;
  assign n81826 = pi17 ? n32 : n81825;
  assign n81827 = pi16 ? n32 : n81826;
  assign n81828 = pi15 ? n81827 : n10716;
  assign n81829 = pi14 ? n10709 : n81828;
  assign n81830 = pi14 ? n10716 : n10729;
  assign n81831 = pi13 ? n81829 : n81830;
  assign n81832 = pi12 ? n81824 : n81831;
  assign n81833 = pi11 ? n81820 : n81832;
  assign n81834 = pi10 ? n81797 : n81833;
  assign n81835 = pi09 ? n81719 : n81834;
  assign n81836 = pi18 ? n751 : ~n936;
  assign n81837 = pi17 ? n32 : n81836;
  assign n81838 = pi16 ? n32 : n81837;
  assign n81839 = pi15 ? n32 : n81838;
  assign n81840 = pi18 ? n684 : ~n1575;
  assign n81841 = pi17 ? n32 : n81840;
  assign n81842 = pi16 ? n32 : n81841;
  assign n81843 = pi15 ? n81710 : n81842;
  assign n81844 = pi14 ? n81839 : n81843;
  assign n81845 = pi13 ? n32 : n81844;
  assign n81846 = pi12 ? n32 : n81845;
  assign n81847 = pi11 ? n32 : n81846;
  assign n81848 = pi10 ? n32 : n81847;
  assign n81849 = pi18 ? n2835 : ~n1575;
  assign n81850 = pi17 ? n32 : n81849;
  assign n81851 = pi16 ? n32 : n81850;
  assign n81852 = pi18 ? n590 : ~n1575;
  assign n81853 = pi17 ? n32 : n81852;
  assign n81854 = pi16 ? n32 : n81853;
  assign n81855 = pi15 ? n81851 : n81854;
  assign n81856 = pi15 ? n81854 : n81571;
  assign n81857 = pi14 ? n81855 : n81856;
  assign n81858 = pi15 ? n81571 : n81713;
  assign n81859 = pi14 ? n81858 : n81587;
  assign n81860 = pi13 ? n81857 : n81859;
  assign n81861 = pi14 ? n81586 : n81303;
  assign n81862 = pi18 ? n702 : ~n2142;
  assign n81863 = pi17 ? n32 : n81862;
  assign n81864 = pi16 ? n32 : n81863;
  assign n81865 = pi18 ? n4098 : ~n2142;
  assign n81866 = pi17 ? n32 : n81865;
  assign n81867 = pi16 ? n32 : n81866;
  assign n81868 = pi15 ? n81864 : n81867;
  assign n81869 = pi18 ? n595 : ~n2142;
  assign n81870 = pi17 ? n32 : n81869;
  assign n81871 = pi16 ? n32 : n81870;
  assign n81872 = pi14 ? n81868 : n81871;
  assign n81873 = pi13 ? n81861 : n81872;
  assign n81874 = pi12 ? n81860 : n81873;
  assign n81875 = pi18 ? n595 : ~n863;
  assign n81876 = pi17 ? n32 : n81875;
  assign n81877 = pi16 ? n32 : n81876;
  assign n81878 = pi18 ? n2627 : ~n863;
  assign n81879 = pi17 ? n32 : n81878;
  assign n81880 = pi16 ? n32 : n81879;
  assign n81881 = pi15 ? n81877 : n81880;
  assign n81882 = pi18 ? n508 : ~n1592;
  assign n81883 = pi17 ? n32 : n81882;
  assign n81884 = pi16 ? n32 : n81883;
  assign n81885 = pi14 ? n81881 : n81884;
  assign n81886 = pi18 ? n323 : ~n1592;
  assign n81887 = pi17 ? n32 : n81886;
  assign n81888 = pi16 ? n32 : n81887;
  assign n81889 = pi18 ? n2291 : ~n1592;
  assign n81890 = pi17 ? n32 : n81889;
  assign n81891 = pi16 ? n32 : n81890;
  assign n81892 = pi15 ? n81888 : n81891;
  assign n81893 = pi18 ? n2291 : ~n1841;
  assign n81894 = pi17 ? n32 : n81893;
  assign n81895 = pi16 ? n32 : n81894;
  assign n81896 = pi14 ? n81892 : n81895;
  assign n81897 = pi13 ? n81885 : n81896;
  assign n81898 = pi18 ? n797 : ~n1841;
  assign n81899 = pi17 ? n32 : n81898;
  assign n81900 = pi16 ? n32 : n81899;
  assign n81901 = pi18 ? n797 : ~n1477;
  assign n81902 = pi17 ? n32 : n81901;
  assign n81903 = pi16 ? n32 : n81902;
  assign n81904 = pi15 ? n81900 : n81903;
  assign n81905 = pi18 ? n2413 : ~n1477;
  assign n81906 = pi17 ? n32 : n81905;
  assign n81907 = pi16 ? n32 : n81906;
  assign n81908 = pi15 ? n81903 : n81907;
  assign n81909 = pi14 ? n81904 : n81908;
  assign n81910 = pi18 ? n605 : ~n751;
  assign n81911 = pi17 ? n32 : n81910;
  assign n81912 = pi16 ? n32 : n81911;
  assign n81913 = pi18 ? n605 : ~n1970;
  assign n81914 = pi17 ? n32 : n81913;
  assign n81915 = pi16 ? n32 : n81914;
  assign n81916 = pi15 ? n81912 : n81915;
  assign n81917 = pi18 ? n605 : ~n245;
  assign n81918 = pi17 ? n32 : n81917;
  assign n81919 = pi16 ? n32 : n81918;
  assign n81920 = pi15 ? n81915 : n81919;
  assign n81921 = pi14 ? n81916 : n81920;
  assign n81922 = pi13 ? n81909 : n81921;
  assign n81923 = pi12 ? n81897 : n81922;
  assign n81924 = pi11 ? n81874 : n81923;
  assign n81925 = pi15 ? n81919 : n10851;
  assign n81926 = pi18 ? n418 : ~n366;
  assign n81927 = pi17 ? n32 : n81926;
  assign n81928 = pi16 ? n32 : n81927;
  assign n81929 = pi15 ? n10851 : n81928;
  assign n81930 = pi14 ? n81925 : n81929;
  assign n81931 = pi18 ? n418 : ~n2962;
  assign n81932 = pi17 ? n32 : n81931;
  assign n81933 = pi16 ? n32 : n81932;
  assign n81934 = pi15 ? n81928 : n81933;
  assign n81935 = pi18 ? n418 : ~n1965;
  assign n81936 = pi17 ? n32 : n81935;
  assign n81937 = pi16 ? n32 : n81936;
  assign n81938 = pi15 ? n81933 : n81937;
  assign n81939 = pi14 ? n81934 : n81938;
  assign n81940 = pi13 ? n81930 : n81939;
  assign n81941 = pi18 ? n3786 : ~n1965;
  assign n81942 = pi17 ? n32 : n81941;
  assign n81943 = pi16 ? n32 : n81942;
  assign n81944 = pi18 ? n2304 : ~n684;
  assign n81945 = pi17 ? n32 : n81944;
  assign n81946 = pi16 ? n32 : n81945;
  assign n81947 = pi15 ? n81943 : n81946;
  assign n81948 = pi18 ? n2304 : ~n590;
  assign n81949 = pi17 ? n32 : n81948;
  assign n81950 = pi16 ? n32 : n81949;
  assign n81951 = pi14 ? n81947 : n81950;
  assign n81952 = pi18 ? n532 : ~n2849;
  assign n81953 = pi17 ? n32 : n81952;
  assign n81954 = pi16 ? n32 : n81953;
  assign n81955 = pi18 ? n2298 : ~n4244;
  assign n81956 = pi17 ? n32 : n81955;
  assign n81957 = pi16 ? n32 : n81956;
  assign n81958 = pi15 ? n81954 : n81957;
  assign n81959 = pi14 ? n81950 : n81958;
  assign n81960 = pi13 ? n81951 : n81959;
  assign n81961 = pi12 ? n81940 : n81960;
  assign n81962 = pi14 ? n10921 : n36497;
  assign n81963 = pi15 ? n10935 : n10942;
  assign n81964 = pi18 ? n2424 : ~n4098;
  assign n81965 = pi17 ? n32 : n81964;
  assign n81966 = pi16 ? n32 : n81965;
  assign n81967 = pi15 ? n10942 : n81966;
  assign n81968 = pi14 ? n81963 : n81967;
  assign n81969 = pi13 ? n81962 : n81968;
  assign n81970 = pi18 ? n2424 : ~n2627;
  assign n81971 = pi17 ? n32 : n81970;
  assign n81972 = pi16 ? n32 : n81971;
  assign n81973 = pi15 ? n10942 : n81972;
  assign n81974 = pi14 ? n81973 : n10958;
  assign n81975 = pi13 ? n81974 : n10968;
  assign n81976 = pi12 ? n81969 : n81975;
  assign n81977 = pi11 ? n81961 : n81976;
  assign n81978 = pi10 ? n81924 : n81977;
  assign n81979 = pi09 ? n81848 : n81978;
  assign n81980 = pi08 ? n81835 : n81979;
  assign n81981 = pi07 ? n81705 : n81980;
  assign n81982 = pi18 ? n1592 : ~n936;
  assign n81983 = pi17 ? n32 : n81982;
  assign n81984 = pi16 ? n32 : n81983;
  assign n81985 = pi15 ? n32 : n81984;
  assign n81986 = pi18 ? n1970 : ~n1575;
  assign n81987 = pi17 ? n32 : n81986;
  assign n81988 = pi16 ? n32 : n81987;
  assign n81989 = pi18 ? n209 : ~n1575;
  assign n81990 = pi17 ? n32 : n81989;
  assign n81991 = pi16 ? n32 : n81990;
  assign n81992 = pi15 ? n81988 : n81991;
  assign n81993 = pi14 ? n81985 : n81992;
  assign n81994 = pi13 ? n32 : n81993;
  assign n81995 = pi12 ? n32 : n81994;
  assign n81996 = pi11 ? n32 : n81995;
  assign n81997 = pi10 ? n32 : n81996;
  assign n81998 = pi18 ? n245 : ~n1575;
  assign n81999 = pi17 ? n32 : n81998;
  assign n82000 = pi16 ? n32 : n81999;
  assign n82001 = pi18 ? n341 : ~n1575;
  assign n82002 = pi17 ? n32 : n82001;
  assign n82003 = pi16 ? n32 : n82002;
  assign n82004 = pi15 ? n82000 : n82003;
  assign n82005 = pi18 ? n366 : ~n1575;
  assign n82006 = pi17 ? n32 : n82005;
  assign n82007 = pi16 ? n32 : n82006;
  assign n82008 = pi15 ? n82003 : n82007;
  assign n82009 = pi14 ? n82004 : n82008;
  assign n82010 = pi15 ? n82007 : n81842;
  assign n82011 = pi14 ? n82010 : n81726;
  assign n82012 = pi13 ? n82009 : n82011;
  assign n82013 = pi14 ? n81725 : n81437;
  assign n82014 = pi18 ? n697 : ~n2142;
  assign n82015 = pi17 ? n32 : n82014;
  assign n82016 = pi16 ? n32 : n82015;
  assign n82017 = pi18 ? n2615 : ~n2142;
  assign n82018 = pi17 ? n32 : n82017;
  assign n82019 = pi16 ? n32 : n82018;
  assign n82020 = pi15 ? n82016 : n82019;
  assign n82021 = pi18 ? n1750 : ~n2142;
  assign n82022 = pi17 ? n32 : n82021;
  assign n82023 = pi16 ? n32 : n82022;
  assign n82024 = pi14 ? n82020 : n82023;
  assign n82025 = pi13 ? n82013 : n82024;
  assign n82026 = pi12 ? n82012 : n82025;
  assign n82027 = pi18 ? n1750 : ~n863;
  assign n82028 = pi17 ? n32 : n82027;
  assign n82029 = pi16 ? n32 : n82028;
  assign n82030 = pi18 ? n2622 : ~n863;
  assign n82031 = pi17 ? n32 : n82030;
  assign n82032 = pi16 ? n32 : n82031;
  assign n82033 = pi15 ? n82029 : n82032;
  assign n82034 = pi18 ? n2622 : ~n1592;
  assign n82035 = pi17 ? n32 : n82034;
  assign n82036 = pi16 ? n32 : n82035;
  assign n82037 = pi18 ? n702 : ~n1592;
  assign n82038 = pi17 ? n32 : n82037;
  assign n82039 = pi16 ? n32 : n82038;
  assign n82040 = pi15 ? n82036 : n82039;
  assign n82041 = pi14 ? n82033 : n82040;
  assign n82042 = pi18 ? n4098 : ~n1592;
  assign n82043 = pi17 ? n32 : n82042;
  assign n82044 = pi16 ? n32 : n82043;
  assign n82045 = pi15 ? n82039 : n82044;
  assign n82046 = pi18 ? n4098 : ~n1841;
  assign n82047 = pi17 ? n32 : n82046;
  assign n82048 = pi16 ? n32 : n82047;
  assign n82049 = pi14 ? n82045 : n82048;
  assign n82050 = pi13 ? n82041 : n82049;
  assign n82051 = pi18 ? n595 : ~n1477;
  assign n82052 = pi17 ? n32 : n82051;
  assign n82053 = pi16 ? n32 : n82052;
  assign n82054 = pi18 ? n2627 : ~n1477;
  assign n82055 = pi17 ? n32 : n82054;
  assign n82056 = pi16 ? n32 : n82055;
  assign n82057 = pi15 ? n82053 : n82056;
  assign n82058 = pi18 ? n2754 : ~n1477;
  assign n82059 = pi17 ? n32 : n82058;
  assign n82060 = pi16 ? n32 : n82059;
  assign n82061 = pi15 ? n82056 : n82060;
  assign n82062 = pi14 ? n82057 : n82061;
  assign n82063 = pi18 ? n323 : ~n1970;
  assign n82064 = pi17 ? n32 : n82063;
  assign n82065 = pi16 ? n32 : n82064;
  assign n82066 = pi14 ? n82065 : n11081;
  assign n82067 = pi13 ? n82062 : n82066;
  assign n82068 = pi12 ? n82050 : n82067;
  assign n82069 = pi11 ? n82026 : n82068;
  assign n82070 = pi18 ? n797 : ~n366;
  assign n82071 = pi17 ? n32 : n82070;
  assign n82072 = pi16 ? n32 : n82071;
  assign n82073 = pi15 ? n11085 : n82072;
  assign n82074 = pi14 ? n11081 : n82073;
  assign n82075 = pi18 ? n797 : ~n2962;
  assign n82076 = pi17 ? n32 : n82075;
  assign n82077 = pi16 ? n32 : n82076;
  assign n82078 = pi18 ? n797 : ~n1965;
  assign n82079 = pi17 ? n32 : n82078;
  assign n82080 = pi16 ? n32 : n82079;
  assign n82081 = pi15 ? n82077 : n82080;
  assign n82082 = pi14 ? n82077 : n82081;
  assign n82083 = pi13 ? n82074 : n82082;
  assign n82084 = pi18 ? n3786 : ~n590;
  assign n82085 = pi17 ? n32 : n82084;
  assign n82086 = pi16 ? n32 : n82085;
  assign n82087 = pi15 ? n10565 : n82086;
  assign n82088 = pi18 ? n2413 : ~n590;
  assign n82089 = pi17 ? n32 : n82088;
  assign n82090 = pi16 ? n32 : n82089;
  assign n82091 = pi15 ? n82086 : n82090;
  assign n82092 = pi14 ? n82087 : n82091;
  assign n82093 = pi18 ? n2413 : ~n496;
  assign n82094 = pi17 ? n32 : n82093;
  assign n82095 = pi16 ? n32 : n82094;
  assign n82096 = pi15 ? n82090 : n82095;
  assign n82097 = pi18 ? n2413 : ~n2730;
  assign n82098 = pi17 ? n32 : n82097;
  assign n82099 = pi16 ? n32 : n82098;
  assign n82100 = pi15 ? n82099 : n11160;
  assign n82101 = pi14 ? n82096 : n82100;
  assign n82102 = pi13 ? n82092 : n82101;
  assign n82103 = pi12 ? n82083 : n82102;
  assign n82104 = pi15 ? n36508 : n11167;
  assign n82105 = pi14 ? n11160 : n82104;
  assign n82106 = pi13 ? n82105 : n11179;
  assign n82107 = pi18 ? n323 : ~n2627;
  assign n82108 = pi17 ? n32 : n82107;
  assign n82109 = pi16 ? n32 : n82108;
  assign n82110 = pi15 ? n82109 : n11194;
  assign n82111 = pi14 ? n82110 : n11194;
  assign n82112 = pi13 ? n82111 : n11207;
  assign n82113 = pi12 ? n82106 : n82112;
  assign n82114 = pi11 ? n82103 : n82113;
  assign n82115 = pi10 ? n82069 : n82114;
  assign n82116 = pi09 ? n81997 : n82115;
  assign n82117 = pi18 ? n2142 : ~n936;
  assign n82118 = pi17 ? n32 : n82117;
  assign n82119 = pi16 ? n32 : n82118;
  assign n82120 = pi15 ? n32 : n82119;
  assign n82121 = pi18 ? n1841 : ~n1575;
  assign n82122 = pi17 ? n32 : n82121;
  assign n82123 = pi16 ? n32 : n82122;
  assign n82124 = pi18 ? n940 : ~n1575;
  assign n82125 = pi17 ? n32 : n82124;
  assign n82126 = pi16 ? n32 : n82125;
  assign n82127 = pi15 ? n82123 : n82126;
  assign n82128 = pi14 ? n82120 : n82127;
  assign n82129 = pi13 ? n32 : n82128;
  assign n82130 = pi12 ? n32 : n82129;
  assign n82131 = pi11 ? n32 : n82130;
  assign n82132 = pi10 ? n32 : n82131;
  assign n82133 = pi18 ? n1477 : ~n1575;
  assign n82134 = pi17 ? n32 : n82133;
  assign n82135 = pi16 ? n32 : n82134;
  assign n82136 = pi18 ? n751 : ~n1575;
  assign n82137 = pi17 ? n32 : n82136;
  assign n82138 = pi16 ? n32 : n82137;
  assign n82139 = pi15 ? n82135 : n82138;
  assign n82140 = pi15 ? n82138 : n81988;
  assign n82141 = pi14 ? n82139 : n82140;
  assign n82142 = pi15 ? n81988 : n81842;
  assign n82143 = pi14 ? n82142 : n81855;
  assign n82144 = pi13 ? n82141 : n82143;
  assign n82145 = pi14 ? n81854 : n81571;
  assign n82146 = pi18 ? n496 : ~n2142;
  assign n82147 = pi17 ? n32 : n82146;
  assign n82148 = pi16 ? n32 : n82147;
  assign n82149 = pi18 ? n4244 : ~n2142;
  assign n82150 = pi17 ? n32 : n82149;
  assign n82151 = pi16 ? n32 : n82150;
  assign n82152 = pi15 ? n82148 : n82151;
  assign n82153 = pi18 ? n962 : ~n2142;
  assign n82154 = pi17 ? n32 : n82153;
  assign n82155 = pi16 ? n32 : n82154;
  assign n82156 = pi14 ? n82152 : n82155;
  assign n82157 = pi13 ? n82145 : n82156;
  assign n82158 = pi12 ? n82144 : n82157;
  assign n82159 = pi18 ? n962 : ~n863;
  assign n82160 = pi17 ? n32 : n82159;
  assign n82161 = pi16 ? n32 : n82160;
  assign n82162 = pi18 ? n2730 : ~n863;
  assign n82163 = pi17 ? n32 : n82162;
  assign n82164 = pi16 ? n32 : n82163;
  assign n82165 = pi15 ? n82161 : n82164;
  assign n82166 = pi18 ? n2730 : ~n1592;
  assign n82167 = pi17 ? n32 : n82166;
  assign n82168 = pi16 ? n32 : n82167;
  assign n82169 = pi18 ? n697 : ~n1592;
  assign n82170 = pi17 ? n32 : n82169;
  assign n82171 = pi16 ? n32 : n82170;
  assign n82172 = pi15 ? n82168 : n82171;
  assign n82173 = pi14 ? n82165 : n82172;
  assign n82174 = pi18 ? n2615 : ~n1592;
  assign n82175 = pi17 ? n32 : n82174;
  assign n82176 = pi16 ? n32 : n82175;
  assign n82177 = pi15 ? n82171 : n82176;
  assign n82178 = pi18 ? n2615 : ~n1841;
  assign n82179 = pi17 ? n32 : n82178;
  assign n82180 = pi16 ? n32 : n82179;
  assign n82181 = pi14 ? n82177 : n82180;
  assign n82182 = pi13 ? n82173 : n82181;
  assign n82183 = pi18 ? n1750 : ~n1477;
  assign n82184 = pi17 ? n32 : n82183;
  assign n82185 = pi16 ? n32 : n82184;
  assign n82186 = pi18 ? n2622 : ~n1477;
  assign n82187 = pi17 ? n32 : n82186;
  assign n82188 = pi16 ? n32 : n82187;
  assign n82189 = pi14 ? n82185 : n82188;
  assign n82190 = pi18 ? n702 : ~n1970;
  assign n82191 = pi17 ? n32 : n82190;
  assign n82192 = pi16 ? n32 : n82191;
  assign n82193 = pi14 ? n82192 : n11308;
  assign n82194 = pi13 ? n82189 : n82193;
  assign n82195 = pi12 ? n82182 : n82194;
  assign n82196 = pi11 ? n82158 : n82195;
  assign n82197 = pi18 ? n520 : ~n366;
  assign n82198 = pi17 ? n32 : n82197;
  assign n82199 = pi16 ? n32 : n82198;
  assign n82200 = pi15 ? n11320 : n82199;
  assign n82201 = pi14 ? n11316 : n82200;
  assign n82202 = pi18 ? n520 : ~n2962;
  assign n82203 = pi17 ? n32 : n82202;
  assign n82204 = pi16 ? n32 : n82203;
  assign n82205 = pi18 ? n520 : ~n1965;
  assign n82206 = pi17 ? n32 : n82205;
  assign n82207 = pi16 ? n32 : n82206;
  assign n82208 = pi15 ? n82204 : n82207;
  assign n82209 = pi14 ? n82204 : n82208;
  assign n82210 = pi13 ? n82201 : n82209;
  assign n82211 = pi18 ? n520 : ~n684;
  assign n82212 = pi17 ? n32 : n82211;
  assign n82213 = pi16 ? n32 : n82212;
  assign n82214 = pi18 ? n2754 : ~n590;
  assign n82215 = pi17 ? n32 : n82214;
  assign n82216 = pi16 ? n32 : n82215;
  assign n82217 = pi15 ? n82213 : n82216;
  assign n82218 = pi14 ? n82217 : n82216;
  assign n82219 = pi18 ? n2754 : ~n496;
  assign n82220 = pi17 ? n32 : n82219;
  assign n82221 = pi16 ? n32 : n82220;
  assign n82222 = pi15 ? n82216 : n82221;
  assign n82223 = pi18 ? n2754 : ~n2730;
  assign n82224 = pi17 ? n32 : n82223;
  assign n82225 = pi16 ? n32 : n82224;
  assign n82226 = pi15 ? n82225 : n11385;
  assign n82227 = pi14 ? n82222 : n82226;
  assign n82228 = pi13 ? n82218 : n82227;
  assign n82229 = pi12 ? n82210 : n82228;
  assign n82230 = pi18 ? n323 : ~n2615;
  assign n82231 = pi17 ? n32 : n82230;
  assign n82232 = pi16 ? n32 : n82231;
  assign n82233 = pi15 ? n82232 : n11401;
  assign n82234 = pi14 ? n11385 : n82233;
  assign n82235 = pi13 ? n82234 : n11401;
  assign n82236 = pi15 ? n11414 : n11198;
  assign n82237 = pi15 ? n11198 : n11418;
  assign n82238 = pi14 ? n82236 : n82237;
  assign n82239 = pi15 ? n11418 : n11423;
  assign n82240 = pi14 ? n82239 : n11430;
  assign n82241 = pi13 ? n82238 : n82240;
  assign n82242 = pi12 ? n82235 : n82241;
  assign n82243 = pi11 ? n82229 : n82242;
  assign n82244 = pi10 ? n82196 : n82243;
  assign n82245 = pi09 ? n82132 : n82244;
  assign n82246 = pi08 ? n82116 : n82245;
  assign n82247 = pi19 ? n1105 : ~n594;
  assign n82248 = pi18 ? n32 : n82247;
  assign n82249 = pi17 ? n32 : n82248;
  assign n82250 = pi16 ? n32 : n82249;
  assign n82251 = pi15 ? n32 : n82250;
  assign n82252 = pi18 ? n2142 : ~n1575;
  assign n82253 = pi17 ? n32 : n82252;
  assign n82254 = pi16 ? n32 : n82253;
  assign n82255 = pi18 ? n863 : ~n1575;
  assign n82256 = pi17 ? n32 : n82255;
  assign n82257 = pi16 ? n32 : n82256;
  assign n82258 = pi15 ? n82254 : n82257;
  assign n82259 = pi14 ? n82251 : n82258;
  assign n82260 = pi13 ? n32 : n82259;
  assign n82261 = pi12 ? n32 : n82260;
  assign n82262 = pi11 ? n32 : n82261;
  assign n82263 = pi10 ? n32 : n82262;
  assign n82264 = pi18 ? n1592 : ~n1575;
  assign n82265 = pi17 ? n32 : n82264;
  assign n82266 = pi16 ? n32 : n82265;
  assign n82267 = pi15 ? n82257 : n82266;
  assign n82268 = pi15 ? n82266 : n82123;
  assign n82269 = pi14 ? n82267 : n82268;
  assign n82270 = pi15 ? n82123 : n81991;
  assign n82271 = pi14 ? n82270 : n82004;
  assign n82272 = pi13 ? n82269 : n82271;
  assign n82273 = pi14 ? n82003 : n82007;
  assign n82274 = pi18 ? n684 : ~n2142;
  assign n82275 = pi17 ? n32 : n82274;
  assign n82276 = pi16 ? n32 : n82275;
  assign n82277 = pi18 ? n2835 : ~n2142;
  assign n82278 = pi17 ? n32 : n82277;
  assign n82279 = pi16 ? n32 : n82278;
  assign n82280 = pi15 ? n82276 : n82279;
  assign n82281 = pi18 ? n590 : ~n2142;
  assign n82282 = pi17 ? n32 : n82281;
  assign n82283 = pi16 ? n32 : n82282;
  assign n82284 = pi14 ? n82280 : n82283;
  assign n82285 = pi13 ? n82273 : n82284;
  assign n82286 = pi12 ? n82272 : n82285;
  assign n82287 = pi18 ? n590 : ~n863;
  assign n82288 = pi17 ? n32 : n82287;
  assign n82289 = pi16 ? n32 : n82288;
  assign n82290 = pi18 ? n2849 : ~n863;
  assign n82291 = pi17 ? n32 : n82290;
  assign n82292 = pi16 ? n32 : n82291;
  assign n82293 = pi15 ? n82289 : n82292;
  assign n82294 = pi18 ? n2849 : ~n1592;
  assign n82295 = pi17 ? n32 : n82294;
  assign n82296 = pi16 ? n32 : n82295;
  assign n82297 = pi18 ? n496 : ~n1592;
  assign n82298 = pi17 ? n32 : n82297;
  assign n82299 = pi16 ? n32 : n82298;
  assign n82300 = pi15 ? n82296 : n82299;
  assign n82301 = pi14 ? n82293 : n82300;
  assign n82302 = pi18 ? n4244 : ~n1592;
  assign n82303 = pi17 ? n32 : n82302;
  assign n82304 = pi16 ? n32 : n82303;
  assign n82305 = pi15 ? n82299 : n82304;
  assign n82306 = pi18 ? n4244 : ~n1841;
  assign n82307 = pi17 ? n32 : n82306;
  assign n82308 = pi16 ? n32 : n82307;
  assign n82309 = pi14 ? n82305 : n82308;
  assign n82310 = pi13 ? n82301 : n82309;
  assign n82311 = pi18 ? n962 : ~n1477;
  assign n82312 = pi17 ? n32 : n82311;
  assign n82313 = pi16 ? n32 : n82312;
  assign n82314 = pi18 ? n2730 : ~n1477;
  assign n82315 = pi17 ? n32 : n82314;
  assign n82316 = pi16 ? n32 : n82315;
  assign n82317 = pi14 ? n82313 : n82316;
  assign n82318 = pi18 ? n697 : ~n1970;
  assign n82319 = pi17 ? n32 : n82318;
  assign n82320 = pi16 ? n32 : n82319;
  assign n82321 = pi14 ? n82320 : n11530;
  assign n82322 = pi13 ? n82317 : n82321;
  assign n82323 = pi12 ? n82310 : n82322;
  assign n82324 = pi11 ? n82286 : n82323;
  assign n82325 = pi18 ? n2615 : ~n245;
  assign n82326 = pi17 ? n32 : n82325;
  assign n82327 = pi16 ? n32 : n82326;
  assign n82328 = pi15 ? n11530 : n82327;
  assign n82329 = pi14 ? n82328 : n11558;
  assign n82330 = pi18 ? n595 : ~n2830;
  assign n82331 = pi17 ? n32 : n82330;
  assign n82332 = pi16 ? n32 : n82331;
  assign n82333 = pi15 ? n11557 : n82332;
  assign n82334 = pi14 ? n11557 : n82333;
  assign n82335 = pi13 ? n82329 : n82334;
  assign n82336 = pi18 ? n2622 : ~n590;
  assign n82337 = pi17 ? n32 : n82336;
  assign n82338 = pi16 ? n32 : n82337;
  assign n82339 = pi18 ? n2627 : ~n590;
  assign n82340 = pi17 ? n32 : n82339;
  assign n82341 = pi16 ? n32 : n82340;
  assign n82342 = pi15 ? n82338 : n82341;
  assign n82343 = pi14 ? n82342 : n82341;
  assign n82344 = pi15 ? n82341 : n11609;
  assign n82345 = pi18 ? n508 : ~n2730;
  assign n82346 = pi17 ? n32 : n82345;
  assign n82347 = pi16 ? n32 : n82346;
  assign n82348 = pi15 ? n11613 : n82347;
  assign n82349 = pi14 ? n82344 : n82348;
  assign n82350 = pi13 ? n82343 : n82349;
  assign n82351 = pi12 ? n82335 : n82350;
  assign n82352 = pi14 ? n82347 : n11632;
  assign n82353 = pi13 ? n82352 : n11631;
  assign n82354 = pi12 ? n82353 : n11660;
  assign n82355 = pi11 ? n82351 : n82354;
  assign n82356 = pi10 ? n82324 : n82355;
  assign n82357 = pi09 ? n82263 : n82356;
  assign n82358 = pi19 ? n1941 : ~n594;
  assign n82359 = pi18 ? n32 : n82358;
  assign n82360 = pi17 ? n32 : n82359;
  assign n82361 = pi16 ? n32 : n82360;
  assign n82362 = pi15 ? n32 : n82361;
  assign n82363 = pi19 ? n1105 : ~n1574;
  assign n82364 = pi18 ? n32 : n82363;
  assign n82365 = pi17 ? n32 : n82364;
  assign n82366 = pi16 ? n32 : n82365;
  assign n82367 = pi18 ? n32 : ~n1575;
  assign n82368 = pi17 ? n32 : n82367;
  assign n82369 = pi16 ? n32 : n82368;
  assign n82370 = pi15 ? n82366 : n82369;
  assign n82371 = pi14 ? n82362 : n82370;
  assign n82372 = pi13 ? n32 : n82371;
  assign n82373 = pi12 ? n32 : n82372;
  assign n82374 = pi11 ? n32 : n82373;
  assign n82375 = pi10 ? n32 : n82374;
  assign n82376 = pi18 ? n1575 : ~n1575;
  assign n82377 = pi17 ? n32 : n82376;
  assign n82378 = pi16 ? n32 : n82377;
  assign n82379 = pi15 ? n82369 : n82378;
  assign n82380 = pi15 ? n82378 : n82254;
  assign n82381 = pi14 ? n82379 : n82380;
  assign n82382 = pi15 ? n82257 : n82126;
  assign n82383 = pi14 ? n82382 : n82139;
  assign n82384 = pi13 ? n82381 : n82383;
  assign n82385 = pi14 ? n82138 : n81988;
  assign n82386 = pi18 ? n209 : ~n2142;
  assign n82387 = pi17 ? n32 : n82386;
  assign n82388 = pi16 ? n32 : n82387;
  assign n82389 = pi18 ? n245 : ~n2142;
  assign n82390 = pi17 ? n32 : n82389;
  assign n82391 = pi16 ? n32 : n82390;
  assign n82392 = pi15 ? n82388 : n82391;
  assign n82393 = pi18 ? n341 : ~n2142;
  assign n82394 = pi17 ? n32 : n82393;
  assign n82395 = pi16 ? n32 : n82394;
  assign n82396 = pi14 ? n82392 : n82395;
  assign n82397 = pi13 ? n82385 : n82396;
  assign n82398 = pi12 ? n82384 : n82397;
  assign n82399 = pi16 ? n32 : n1039;
  assign n82400 = pi16 ? n32 : n1239;
  assign n82401 = pi15 ? n82399 : n82400;
  assign n82402 = pi16 ? n32 : n1875;
  assign n82403 = pi18 ? n684 : ~n1592;
  assign n82404 = pi17 ? n32 : n82403;
  assign n82405 = pi16 ? n32 : n82404;
  assign n82406 = pi15 ? n82402 : n82405;
  assign n82407 = pi14 ? n82401 : n82406;
  assign n82408 = pi18 ? n2835 : ~n1592;
  assign n82409 = pi17 ? n32 : n82408;
  assign n82410 = pi16 ? n32 : n82409;
  assign n82411 = pi15 ? n82405 : n82410;
  assign n82412 = pi18 ? n2835 : ~n1841;
  assign n82413 = pi17 ? n32 : n82412;
  assign n82414 = pi16 ? n32 : n82413;
  assign n82415 = pi14 ? n82411 : n82414;
  assign n82416 = pi13 ? n82407 : n82415;
  assign n82417 = pi18 ? n590 : ~n1477;
  assign n82418 = pi17 ? n32 : n82417;
  assign n82419 = pi16 ? n32 : n82418;
  assign n82420 = pi18 ? n2849 : ~n1477;
  assign n82421 = pi17 ? n32 : n82420;
  assign n82422 = pi16 ? n32 : n82421;
  assign n82423 = pi14 ? n82419 : n82422;
  assign n82424 = pi14 ? n11746 : n11750;
  assign n82425 = pi13 ? n82423 : n82424;
  assign n82426 = pi12 ? n82416 : n82425;
  assign n82427 = pi11 ? n82398 : n82426;
  assign n82428 = pi18 ? n4244 : ~n245;
  assign n82429 = pi17 ? n32 : n82428;
  assign n82430 = pi16 ? n32 : n82429;
  assign n82431 = pi15 ? n11750 : n82430;
  assign n82432 = pi18 ? n4244 : ~n366;
  assign n82433 = pi17 ? n32 : n82432;
  assign n82434 = pi16 ? n32 : n82433;
  assign n82435 = pi15 ? n82434 : n11775;
  assign n82436 = pi14 ? n82431 : n82435;
  assign n82437 = pi18 ? n962 : ~n2830;
  assign n82438 = pi17 ? n32 : n82437;
  assign n82439 = pi16 ? n32 : n82438;
  assign n82440 = pi15 ? n11775 : n82439;
  assign n82441 = pi14 ? n11775 : n82440;
  assign n82442 = pi13 ? n82436 : n82441;
  assign n82443 = pi15 ? n12033 : n82338;
  assign n82444 = pi14 ? n82443 : n82338;
  assign n82445 = pi18 ? n2730 : ~n2849;
  assign n82446 = pi17 ? n32 : n82445;
  assign n82447 = pi16 ? n32 : n82446;
  assign n82448 = pi15 ? n82447 : n11815;
  assign n82449 = pi14 ? n82448 : n11820;
  assign n82450 = pi13 ? n82444 : n82449;
  assign n82451 = pi12 ? n82442 : n82450;
  assign n82452 = pi14 ? n11819 : n11835;
  assign n82453 = pi18 ? n496 : ~n4098;
  assign n82454 = pi17 ? n32 : n82453;
  assign n82455 = pi16 ? n32 : n82454;
  assign n82456 = pi15 ? n82455 : n11839;
  assign n82457 = pi14 ? n11834 : n82456;
  assign n82458 = pi13 ? n82452 : n82457;
  assign n82459 = pi12 ? n82458 : n11866;
  assign n82460 = pi11 ? n82451 : n82459;
  assign n82461 = pi10 ? n82427 : n82460;
  assign n82462 = pi09 ? n82375 : n82461;
  assign n82463 = pi08 ? n82357 : n82462;
  assign n82464 = pi07 ? n82246 : n82463;
  assign n82465 = pi06 ? n81981 : n82464;
  assign n82466 = pi19 ? n1941 : ~n1574;
  assign n82467 = pi18 ? n32 : n82466;
  assign n82468 = pi17 ? n32 : n82467;
  assign n82469 = pi16 ? n32 : n82468;
  assign n82470 = pi19 ? n236 : ~n1574;
  assign n82471 = pi18 ? n32 : n82470;
  assign n82472 = pi17 ? n32 : n82471;
  assign n82473 = pi16 ? n32 : n82472;
  assign n82474 = pi15 ? n82469 : n82473;
  assign n82475 = pi14 ? n82362 : n82474;
  assign n82476 = pi13 ? n32 : n82475;
  assign n82477 = pi12 ? n32 : n82476;
  assign n82478 = pi11 ? n32 : n82477;
  assign n82479 = pi10 ? n32 : n82478;
  assign n82480 = pi19 ? n2614 : ~n1574;
  assign n82481 = pi18 ? n32 : n82480;
  assign n82482 = pi17 ? n32 : n82481;
  assign n82483 = pi16 ? n32 : n82482;
  assign n82484 = pi15 ? n82473 : n82483;
  assign n82485 = pi19 ? n617 : ~n1574;
  assign n82486 = pi18 ? n32 : n82485;
  assign n82487 = pi17 ? n32 : n82486;
  assign n82488 = pi16 ? n32 : n82487;
  assign n82489 = pi15 ? n82488 : n82369;
  assign n82490 = pi14 ? n82484 : n82489;
  assign n82491 = pi15 ? n82369 : n82257;
  assign n82492 = pi18 ? n1321 : ~n1575;
  assign n82493 = pi17 ? n32 : n82492;
  assign n82494 = pi16 ? n32 : n82493;
  assign n82495 = pi14 ? n82491 : n82494;
  assign n82496 = pi13 ? n82490 : n82495;
  assign n82497 = pi14 ? n82266 : n82123;
  assign n82498 = pi18 ? n940 : ~n2142;
  assign n82499 = pi17 ? n32 : n82498;
  assign n82500 = pi16 ? n32 : n82499;
  assign n82501 = pi18 ? n1477 : ~n2142;
  assign n82502 = pi17 ? n32 : n82501;
  assign n82503 = pi16 ? n32 : n82502;
  assign n82504 = pi15 ? n82500 : n82503;
  assign n82505 = pi18 ? n751 : ~n2142;
  assign n82506 = pi17 ? n32 : n82505;
  assign n82507 = pi16 ? n32 : n82506;
  assign n82508 = pi14 ? n82504 : n82507;
  assign n82509 = pi13 ? n82497 : n82508;
  assign n82510 = pi12 ? n82496 : n82509;
  assign n82511 = pi18 ? n751 : ~n863;
  assign n82512 = pi17 ? n32 : n82511;
  assign n82513 = pi16 ? n32 : n82512;
  assign n82514 = pi18 ? n1970 : ~n863;
  assign n82515 = pi17 ? n32 : n82514;
  assign n82516 = pi16 ? n32 : n82515;
  assign n82517 = pi15 ? n82513 : n82516;
  assign n82518 = pi18 ? n1970 : ~n1592;
  assign n82519 = pi17 ? n32 : n82518;
  assign n82520 = pi16 ? n32 : n82519;
  assign n82521 = pi18 ? n209 : ~n1592;
  assign n82522 = pi17 ? n32 : n82521;
  assign n82523 = pi16 ? n32 : n82522;
  assign n82524 = pi15 ? n82520 : n82523;
  assign n82525 = pi14 ? n82517 : n82524;
  assign n82526 = pi18 ? n245 : ~n1592;
  assign n82527 = pi17 ? n32 : n82526;
  assign n82528 = pi16 ? n32 : n82527;
  assign n82529 = pi15 ? n82523 : n82528;
  assign n82530 = pi18 ? n245 : ~n1841;
  assign n82531 = pi17 ? n32 : n82530;
  assign n82532 = pi16 ? n32 : n82531;
  assign n82533 = pi14 ? n82529 : n82532;
  assign n82534 = pi13 ? n82525 : n82533;
  assign n82535 = pi18 ? n341 : ~n1477;
  assign n82536 = pi17 ? n32 : n82535;
  assign n82537 = pi16 ? n32 : n82536;
  assign n82538 = pi18 ? n2830 : ~n1477;
  assign n82539 = pi17 ? n32 : n82538;
  assign n82540 = pi16 ? n32 : n82539;
  assign n82541 = pi14 ? n82537 : n82540;
  assign n82542 = pi18 ? n684 : ~n245;
  assign n82543 = pi17 ? n32 : n82542;
  assign n82544 = pi16 ? n32 : n82543;
  assign n82545 = pi14 ? n11984 : n82544;
  assign n82546 = pi13 ? n82541 : n82545;
  assign n82547 = pi12 ? n82534 : n82546;
  assign n82548 = pi11 ? n82510 : n82547;
  assign n82549 = pi18 ? n2835 : ~n245;
  assign n82550 = pi17 ? n32 : n82549;
  assign n82551 = pi16 ? n32 : n82550;
  assign n82552 = pi15 ? n82544 : n82551;
  assign n82553 = pi15 ? n12007 : n12017;
  assign n82554 = pi14 ? n82552 : n82553;
  assign n82555 = pi15 ? n12017 : n12027;
  assign n82556 = pi14 ? n12017 : n82555;
  assign n82557 = pi13 ? n82554 : n82556;
  assign n82558 = pi14 ? n12037 : n12036;
  assign n82559 = pi18 ? n2849 : ~n2849;
  assign n82560 = pi17 ? n32 : n82559;
  assign n82561 = pi16 ? n32 : n82560;
  assign n82562 = pi15 ? n82561 : n12040;
  assign n82563 = pi14 ? n82562 : n12050;
  assign n82564 = pi13 ? n82558 : n82563;
  assign n82565 = pi12 ? n82557 : n82564;
  assign n82566 = pi15 ? n12059 : n12070;
  assign n82567 = pi14 ? n12059 : n82566;
  assign n82568 = pi13 ? n12061 : n82567;
  assign n82569 = pi17 ? n32 : n46312;
  assign n82570 = pi16 ? n32 : n82569;
  assign n82571 = pi15 ? n82570 : n12079;
  assign n82572 = pi14 ? n82571 : n12084;
  assign n82573 = pi13 ? n82572 : n12100;
  assign n82574 = pi12 ? n82568 : n82573;
  assign n82575 = pi11 ? n82565 : n82574;
  assign n82576 = pi10 ? n82548 : n82575;
  assign n82577 = pi09 ? n82479 : n82576;
  assign n82578 = pi19 ? n2848 : ~n594;
  assign n82579 = pi18 ? n32 : n82578;
  assign n82580 = pi17 ? n32 : n82579;
  assign n82581 = pi16 ? n32 : n82580;
  assign n82582 = pi15 ? n32 : n82581;
  assign n82583 = pi19 ? n2848 : ~n1574;
  assign n82584 = pi18 ? n32 : n82583;
  assign n82585 = pi17 ? n32 : n82584;
  assign n82586 = pi16 ? n32 : n82585;
  assign n82587 = pi19 ? n349 : ~n1574;
  assign n82588 = pi18 ? n32 : n82587;
  assign n82589 = pi17 ? n32 : n82588;
  assign n82590 = pi16 ? n32 : n82589;
  assign n82591 = pi15 ? n82586 : n82590;
  assign n82592 = pi14 ? n82582 : n82591;
  assign n82593 = pi13 ? n32 : n82592;
  assign n82594 = pi12 ? n32 : n82593;
  assign n82595 = pi11 ? n32 : n82594;
  assign n82596 = pi10 ? n32 : n82595;
  assign n82597 = pi19 ? n813 : ~n1574;
  assign n82598 = pi18 ? n32 : n82597;
  assign n82599 = pi17 ? n32 : n82598;
  assign n82600 = pi16 ? n32 : n82599;
  assign n82601 = pi15 ? n82590 : n82600;
  assign n82602 = pi14 ? n82601 : n82474;
  assign n82603 = pi15 ? n82473 : n82369;
  assign n82604 = pi14 ? n82603 : n82378;
  assign n82605 = pi13 ? n82602 : n82604;
  assign n82606 = pi14 ? n82378 : n82258;
  assign n82607 = pi18 ? n863 : ~n2142;
  assign n82608 = pi17 ? n32 : n82607;
  assign n82609 = pi16 ? n32 : n82608;
  assign n82610 = pi18 ? n1321 : ~n2142;
  assign n82611 = pi17 ? n32 : n82610;
  assign n82612 = pi16 ? n32 : n82611;
  assign n82613 = pi15 ? n82609 : n82612;
  assign n82614 = pi18 ? n1592 : ~n2142;
  assign n82615 = pi17 ? n32 : n82614;
  assign n82616 = pi16 ? n32 : n82615;
  assign n82617 = pi15 ? n82612 : n82616;
  assign n82618 = pi14 ? n82613 : n82617;
  assign n82619 = pi13 ? n82606 : n82618;
  assign n82620 = pi12 ? n82605 : n82619;
  assign n82621 = pi18 ? n1592 : ~n863;
  assign n82622 = pi17 ? n32 : n82621;
  assign n82623 = pi16 ? n32 : n82622;
  assign n82624 = pi18 ? n1841 : ~n863;
  assign n82625 = pi17 ? n32 : n82624;
  assign n82626 = pi16 ? n32 : n82625;
  assign n82627 = pi15 ? n82623 : n82626;
  assign n82628 = pi18 ? n1841 : ~n1592;
  assign n82629 = pi17 ? n32 : n82628;
  assign n82630 = pi16 ? n32 : n82629;
  assign n82631 = pi18 ? n940 : ~n1592;
  assign n82632 = pi17 ? n32 : n82631;
  assign n82633 = pi16 ? n32 : n82632;
  assign n82634 = pi15 ? n82630 : n82633;
  assign n82635 = pi14 ? n82627 : n82634;
  assign n82636 = pi18 ? n1477 : ~n1592;
  assign n82637 = pi17 ? n32 : n82636;
  assign n82638 = pi16 ? n32 : n82637;
  assign n82639 = pi15 ? n82633 : n82638;
  assign n82640 = pi18 ? n1477 : ~n1841;
  assign n82641 = pi17 ? n32 : n82640;
  assign n82642 = pi16 ? n32 : n82641;
  assign n82643 = pi14 ? n82639 : n82642;
  assign n82644 = pi13 ? n82635 : n82643;
  assign n82645 = pi18 ? n751 : ~n1477;
  assign n82646 = pi17 ? n32 : n82645;
  assign n82647 = pi16 ? n32 : n82646;
  assign n82648 = pi18 ? n1970 : ~n1477;
  assign n82649 = pi17 ? n32 : n82648;
  assign n82650 = pi16 ? n32 : n82649;
  assign n82651 = pi14 ? n82647 : n82650;
  assign n82652 = pi18 ? n209 : ~n1970;
  assign n82653 = pi17 ? n32 : n82652;
  assign n82654 = pi16 ? n32 : n82653;
  assign n82655 = pi15 ? n82654 : n12203;
  assign n82656 = pi14 ? n82655 : n12203;
  assign n82657 = pi13 ? n82651 : n82656;
  assign n82658 = pi12 ? n82644 : n82657;
  assign n82659 = pi11 ? n82620 : n82658;
  assign n82660 = pi18 ? n2962 : ~n341;
  assign n82661 = pi17 ? n32 : n82660;
  assign n82662 = pi16 ? n32 : n82661;
  assign n82663 = pi15 ? n12203 : n82662;
  assign n82664 = pi15 ? n12219 : n12227;
  assign n82665 = pi14 ? n82663 : n82664;
  assign n82666 = pi15 ? n12230 : n12237;
  assign n82667 = pi14 ? n12227 : n82666;
  assign n82668 = pi13 ? n82665 : n82667;
  assign n82669 = pi15 ? n12257 : n51144;
  assign n82670 = pi14 ? n12258 : n82669;
  assign n82671 = pi13 ? n12243 : n82670;
  assign n82672 = pi12 ? n82668 : n82671;
  assign n82673 = pi15 ? n51144 : n12261;
  assign n82674 = pi14 ? n82673 : n12272;
  assign n82675 = pi15 ? n12271 : n12283;
  assign n82676 = pi14 ? n12271 : n82675;
  assign n82677 = pi13 ? n82674 : n82676;
  assign n82678 = pi15 ? n32885 : n12083;
  assign n82679 = pi14 ? n82678 : n12293;
  assign n82680 = pi13 ? n82679 : n12309;
  assign n82681 = pi12 ? n82677 : n82680;
  assign n82682 = pi11 ? n82672 : n82681;
  assign n82683 = pi10 ? n82659 : n82682;
  assign n82684 = pi09 ? n82596 : n82683;
  assign n82685 = pi08 ? n82577 : n82684;
  assign n82686 = pi19 ? n2303 : ~n594;
  assign n82687 = pi18 ? n32 : n82686;
  assign n82688 = pi17 ? n32 : n82687;
  assign n82689 = pi16 ? n32 : n82688;
  assign n82690 = pi15 ? n32 : n82689;
  assign n82691 = pi19 ? n2303 : ~n1574;
  assign n82692 = pi18 ? n32 : n82691;
  assign n82693 = pi17 ? n32 : n82692;
  assign n82694 = pi16 ? n32 : n82693;
  assign n82695 = pi19 ? n2317 : ~n1574;
  assign n82696 = pi18 ? n32 : n82695;
  assign n82697 = pi17 ? n32 : n82696;
  assign n82698 = pi16 ? n32 : n82697;
  assign n82699 = pi15 ? n82694 : n82698;
  assign n82700 = pi14 ? n82690 : n82699;
  assign n82701 = pi13 ? n32 : n82700;
  assign n82702 = pi12 ? n32 : n82701;
  assign n82703 = pi11 ? n32 : n82702;
  assign n82704 = pi10 ? n32 : n82703;
  assign n82705 = pi15 ? n82698 : n82586;
  assign n82706 = pi14 ? n82705 : n82590;
  assign n82707 = pi14 ? n82473 : n82483;
  assign n82708 = pi13 ? n82706 : n82707;
  assign n82709 = pi15 ? n82483 : n82488;
  assign n82710 = pi14 ? n82709 : n82369;
  assign n82711 = pi18 ? n32 : ~n2142;
  assign n82712 = pi17 ? n32 : n82711;
  assign n82713 = pi16 ? n32 : n82712;
  assign n82714 = pi18 ? n1575 : ~n2142;
  assign n82715 = pi17 ? n32 : n82714;
  assign n82716 = pi16 ? n32 : n82715;
  assign n82717 = pi15 ? n82713 : n82716;
  assign n82718 = pi14 ? n82717 : n82716;
  assign n82719 = pi13 ? n82710 : n82718;
  assign n82720 = pi12 ? n82708 : n82719;
  assign n82721 = pi18 ? n1575 : ~n863;
  assign n82722 = pi17 ? n32 : n82721;
  assign n82723 = pi16 ? n32 : n82722;
  assign n82724 = pi18 ? n2142 : ~n863;
  assign n82725 = pi17 ? n32 : n82724;
  assign n82726 = pi16 ? n32 : n82725;
  assign n82727 = pi15 ? n82723 : n82726;
  assign n82728 = pi18 ? n863 : ~n1592;
  assign n82729 = pi17 ? n32 : n82728;
  assign n82730 = pi16 ? n32 : n82729;
  assign n82731 = pi14 ? n82727 : n82730;
  assign n82732 = pi18 ? n1321 : ~n1841;
  assign n82733 = pi17 ? n32 : n82732;
  assign n82734 = pi16 ? n32 : n82733;
  assign n82735 = pi14 ? n82730 : n82734;
  assign n82736 = pi13 ? n82731 : n82735;
  assign n82737 = pi18 ? n1592 : ~n1477;
  assign n82738 = pi17 ? n32 : n82737;
  assign n82739 = pi16 ? n32 : n82738;
  assign n82740 = pi18 ? n1841 : ~n1477;
  assign n82741 = pi17 ? n32 : n82740;
  assign n82742 = pi16 ? n32 : n82741;
  assign n82743 = pi14 ? n82739 : n82742;
  assign n82744 = pi18 ? n940 : ~n1970;
  assign n82745 = pi17 ? n32 : n82744;
  assign n82746 = pi16 ? n32 : n82745;
  assign n82747 = pi15 ? n82746 : n12454;
  assign n82748 = pi14 ? n82747 : n12454;
  assign n82749 = pi13 ? n82743 : n82748;
  assign n82750 = pi12 ? n82736 : n82749;
  assign n82751 = pi11 ? n82720 : n82750;
  assign n82752 = pi18 ? n1477 : ~n2962;
  assign n82753 = pi17 ? n32 : n82752;
  assign n82754 = pi16 ? n32 : n82753;
  assign n82755 = pi18 ? n751 : ~n2962;
  assign n82756 = pi17 ? n32 : n82755;
  assign n82757 = pi16 ? n32 : n82756;
  assign n82758 = pi15 ? n82754 : n82757;
  assign n82759 = pi14 ? n12458 : n82758;
  assign n82760 = pi18 ? n751 : ~n590;
  assign n82761 = pi17 ? n32 : n82760;
  assign n82762 = pi16 ? n32 : n82761;
  assign n82763 = pi15 ? n12472 : n82762;
  assign n82764 = pi14 ? n82757 : n82763;
  assign n82765 = pi13 ? n82759 : n82764;
  assign n82766 = pi18 ? n366 : ~n2730;
  assign n82767 = pi17 ? n32 : n82766;
  assign n82768 = pi16 ? n32 : n82767;
  assign n82769 = pi15 ? n12486 : n82768;
  assign n82770 = pi15 ? n12491 : n82768;
  assign n82771 = pi14 ? n82769 : n82770;
  assign n82772 = pi13 ? n12481 : n82771;
  assign n82773 = pi12 ? n82765 : n82772;
  assign n82774 = pi18 ? n863 : ~n2298;
  assign n82775 = pi17 ? n32 : n82774;
  assign n82776 = pi16 ? n32 : n82775;
  assign n82777 = pi15 ? n12542 : n82776;
  assign n82778 = pi14 ? n12539 : n82777;
  assign n82779 = pi13 ? n12532 : n82778;
  assign n82780 = pi12 ? n12521 : n82779;
  assign n82781 = pi11 ? n82773 : n82780;
  assign n82782 = pi10 ? n82751 : n82781;
  assign n82783 = pi09 ? n82704 : n82782;
  assign n82784 = pi19 ? n429 : ~n594;
  assign n82785 = pi18 ? n32 : n82784;
  assign n82786 = pi17 ? n32 : n82785;
  assign n82787 = pi16 ? n32 : n82786;
  assign n82788 = pi15 ? n32 : n82787;
  assign n82789 = pi19 ? n429 : ~n1574;
  assign n82790 = pi18 ? n32 : n82789;
  assign n82791 = pi17 ? n32 : n82790;
  assign n82792 = pi16 ? n32 : n82791;
  assign n82793 = pi14 ? n82788 : n82792;
  assign n82794 = pi13 ? n32 : n82793;
  assign n82795 = pi12 ? n32 : n82794;
  assign n82796 = pi11 ? n32 : n82795;
  assign n82797 = pi10 ? n32 : n82796;
  assign n82798 = pi19 ? n343 : ~n1574;
  assign n82799 = pi18 ? n32 : n82798;
  assign n82800 = pi17 ? n32 : n82799;
  assign n82801 = pi16 ? n32 : n82800;
  assign n82802 = pi15 ? n82792 : n82801;
  assign n82803 = pi14 ? n82802 : n82801;
  assign n82804 = pi19 ? n1812 : ~n1574;
  assign n82805 = pi18 ? n32 : n82804;
  assign n82806 = pi17 ? n32 : n82805;
  assign n82807 = pi16 ? n32 : n82806;
  assign n82808 = pi14 ? n82590 : n82807;
  assign n82809 = pi13 ? n82803 : n82808;
  assign n82810 = pi15 ? n82600 : n82469;
  assign n82811 = pi14 ? n82810 : n82473;
  assign n82812 = pi19 ? n236 : ~n2141;
  assign n82813 = pi18 ? n32 : n82812;
  assign n82814 = pi17 ? n32 : n82813;
  assign n82815 = pi16 ? n32 : n82814;
  assign n82816 = pi19 ? n2614 : ~n2141;
  assign n82817 = pi18 ? n32 : n82816;
  assign n82818 = pi17 ? n32 : n82817;
  assign n82819 = pi16 ? n32 : n82818;
  assign n82820 = pi15 ? n82815 : n82819;
  assign n82821 = pi14 ? n82820 : n82819;
  assign n82822 = pi13 ? n82811 : n82821;
  assign n82823 = pi12 ? n82809 : n82822;
  assign n82824 = pi19 ? n617 : ~n507;
  assign n82825 = pi18 ? n32 : n82824;
  assign n82826 = pi17 ? n32 : n82825;
  assign n82827 = pi16 ? n32 : n82826;
  assign n82828 = pi15 ? n82827 : n12638;
  assign n82829 = pi18 ? n32 : ~n1592;
  assign n82830 = pi17 ? n32 : n82829;
  assign n82831 = pi16 ? n32 : n82830;
  assign n82832 = pi14 ? n82828 : n82831;
  assign n82833 = pi18 ? n32 : ~n1841;
  assign n82834 = pi17 ? n32 : n82833;
  assign n82835 = pi16 ? n32 : n82834;
  assign n82836 = pi14 ? n82831 : n82835;
  assign n82837 = pi13 ? n82832 : n82836;
  assign n82838 = pi18 ? n936 : ~n1477;
  assign n82839 = pi17 ? n32 : n82838;
  assign n82840 = pi16 ? n32 : n82839;
  assign n82841 = pi15 ? n82840 : n12665;
  assign n82842 = pi14 ? n82841 : n12665;
  assign n82843 = pi18 ? n2142 : ~n1970;
  assign n82844 = pi17 ? n32 : n82843;
  assign n82845 = pi16 ? n32 : n82844;
  assign n82846 = pi15 ? n82845 : n12687;
  assign n82847 = pi14 ? n82846 : n12687;
  assign n82848 = pi13 ? n82842 : n82847;
  assign n82849 = pi12 ? n82837 : n82848;
  assign n82850 = pi11 ? n82823 : n82849;
  assign n82851 = pi18 ? n1321 : ~n2962;
  assign n82852 = pi17 ? n32 : n82851;
  assign n82853 = pi16 ? n32 : n82852;
  assign n82854 = pi18 ? n1592 : ~n2962;
  assign n82855 = pi17 ? n32 : n82854;
  assign n82856 = pi16 ? n32 : n82855;
  assign n82857 = pi15 ? n82853 : n82856;
  assign n82858 = pi14 ? n12696 : n82857;
  assign n82859 = pi18 ? n1592 : ~n590;
  assign n82860 = pi17 ? n32 : n82859;
  assign n82861 = pi16 ? n32 : n82860;
  assign n82862 = pi15 ? n12715 : n82861;
  assign n82863 = pi14 ? n82856 : n82862;
  assign n82864 = pi13 ? n82858 : n82863;
  assign n82865 = pi18 ? n1970 : ~n590;
  assign n82866 = pi17 ? n32 : n82865;
  assign n82867 = pi16 ? n32 : n82866;
  assign n82868 = pi18 ? n1841 : ~n590;
  assign n82869 = pi17 ? n32 : n82868;
  assign n82870 = pi16 ? n32 : n82869;
  assign n82871 = pi15 ? n82870 : n12727;
  assign n82872 = pi14 ? n82867 : n82871;
  assign n82873 = pi15 ? n12732 : n12739;
  assign n82874 = pi14 ? n82873 : n12743;
  assign n82875 = pi13 ? n82872 : n82874;
  assign n82876 = pi12 ? n82864 : n82875;
  assign n82877 = pi11 ? n82876 : n12795;
  assign n82878 = pi10 ? n82850 : n82877;
  assign n82879 = pi09 ? n82797 : n82878;
  assign n82880 = pi08 ? n82783 : n82879;
  assign n82881 = pi07 ? n82685 : n82880;
  assign n82882 = pi19 ? n531 : ~n594;
  assign n82883 = pi18 ? n32 : n82882;
  assign n82884 = pi17 ? n32 : n82883;
  assign n82885 = pi16 ? n32 : n82884;
  assign n82886 = pi15 ? n32 : n82885;
  assign n82887 = pi19 ? n531 : ~n1574;
  assign n82888 = pi18 ? n32 : n82887;
  assign n82889 = pi17 ? n32 : n82888;
  assign n82890 = pi16 ? n32 : n82889;
  assign n82891 = pi14 ? n82886 : n82890;
  assign n82892 = pi13 ? n32 : n82891;
  assign n82893 = pi12 ? n32 : n82892;
  assign n82894 = pi11 ? n32 : n82893;
  assign n82895 = pi10 ? n32 : n82894;
  assign n82896 = pi19 ? n2297 : ~n1574;
  assign n82897 = pi18 ? n32 : n82896;
  assign n82898 = pi17 ? n32 : n82897;
  assign n82899 = pi16 ? n32 : n82898;
  assign n82900 = pi15 ? n82890 : n82899;
  assign n82901 = pi14 ? n82900 : n82899;
  assign n82902 = pi19 ? n589 : ~n1574;
  assign n82903 = pi18 ? n32 : n82902;
  assign n82904 = pi17 ? n32 : n82903;
  assign n82905 = pi16 ? n32 : n82904;
  assign n82906 = pi14 ? n82801 : n82905;
  assign n82907 = pi13 ? n82901 : n82906;
  assign n82908 = pi14 ? n82591 : n82590;
  assign n82909 = pi18 ? n32 : n18492;
  assign n82910 = pi17 ? n32 : n82909;
  assign n82911 = pi16 ? n32 : n82910;
  assign n82912 = pi19 ? n1812 : ~n2141;
  assign n82913 = pi18 ? n32 : n82912;
  assign n82914 = pi17 ? n32 : n82913;
  assign n82915 = pi16 ? n32 : n82914;
  assign n82916 = pi15 ? n82911 : n82915;
  assign n82917 = pi19 ? n813 : ~n2141;
  assign n82918 = pi18 ? n32 : n82917;
  assign n82919 = pi17 ? n32 : n82918;
  assign n82920 = pi16 ? n32 : n82919;
  assign n82921 = pi15 ? n82915 : n82920;
  assign n82922 = pi14 ? n82916 : n82921;
  assign n82923 = pi13 ? n82908 : n82922;
  assign n82924 = pi12 ? n82907 : n82923;
  assign n82925 = pi19 ? n1941 : ~n507;
  assign n82926 = pi18 ? n32 : n82925;
  assign n82927 = pi17 ? n32 : n82926;
  assign n82928 = pi16 ? n32 : n82927;
  assign n82929 = pi15 ? n82928 : n12893;
  assign n82930 = pi19 ? n236 : ~n519;
  assign n82931 = pi18 ? n32 : n82930;
  assign n82932 = pi17 ? n32 : n82931;
  assign n82933 = pi16 ? n32 : n82932;
  assign n82934 = pi14 ? n82929 : n82933;
  assign n82935 = pi19 ? n2614 : ~n1476;
  assign n82936 = pi18 ? n32 : n82935;
  assign n82937 = pi17 ? n32 : n82936;
  assign n82938 = pi16 ? n32 : n82937;
  assign n82939 = pi15 ? n12918 : n82938;
  assign n82940 = pi14 ? n82933 : n82939;
  assign n82941 = pi13 ? n82934 : n82940;
  assign n82942 = pi19 ? n1105 : ~n1476;
  assign n82943 = pi18 ? n32 : n82942;
  assign n82944 = pi17 ? n32 : n82943;
  assign n82945 = pi16 ? n32 : n82944;
  assign n82946 = pi19 ? n1105 : ~n750;
  assign n82947 = pi18 ? n32 : n82946;
  assign n82948 = pi17 ? n32 : n82947;
  assign n82949 = pi16 ? n32 : n82948;
  assign n82950 = pi15 ? n82945 : n82949;
  assign n82951 = pi14 ? n82945 : n82950;
  assign n82952 = pi19 ? n1105 : ~n244;
  assign n82953 = pi18 ? n32 : n82952;
  assign n82954 = pi17 ? n32 : n82953;
  assign n82955 = pi16 ? n32 : n82954;
  assign n82956 = pi18 ? n32 : ~n245;
  assign n82957 = pi17 ? n32 : n82956;
  assign n82958 = pi16 ? n32 : n82957;
  assign n82959 = pi15 ? n82955 : n82958;
  assign n82960 = pi14 ? n82955 : n82959;
  assign n82961 = pi13 ? n82951 : n82960;
  assign n82962 = pi12 ? n82941 : n82961;
  assign n82963 = pi11 ? n82924 : n82962;
  assign n82964 = pi18 ? n1575 : ~n2962;
  assign n82965 = pi17 ? n32 : n82964;
  assign n82966 = pi16 ? n32 : n82965;
  assign n82967 = pi15 ? n12969 : n82966;
  assign n82968 = pi14 ? n82967 : n82966;
  assign n82969 = pi18 ? n936 : ~n590;
  assign n82970 = pi17 ? n32 : n82969;
  assign n82971 = pi16 ? n32 : n82970;
  assign n82972 = pi15 ? n12991 : n82971;
  assign n82973 = pi14 ? n12981 : n82972;
  assign n82974 = pi13 ? n82968 : n82973;
  assign n82975 = pi15 ? n13000 : n13006;
  assign n82976 = pi14 ? n13000 : n82975;
  assign n82977 = pi13 ? n82976 : n13020;
  assign n82978 = pi12 ? n82974 : n82977;
  assign n82979 = pi11 ? n82978 : n13093;
  assign n82980 = pi10 ? n82963 : n82979;
  assign n82981 = pi09 ? n82895 : n82980;
  assign n82982 = pi19 ? n340 : ~n594;
  assign n82983 = pi18 ? n32 : n82982;
  assign n82984 = pi17 ? n32 : n82983;
  assign n82985 = pi16 ? n32 : n82984;
  assign n82986 = pi15 ? n32 : n82985;
  assign n82987 = pi19 ? n340 : ~n1574;
  assign n82988 = pi18 ? n32 : n82987;
  assign n82989 = pi17 ? n32 : n82988;
  assign n82990 = pi16 ? n32 : n82989;
  assign n82991 = pi14 ? n82986 : n82990;
  assign n82992 = pi13 ? n32 : n82991;
  assign n82993 = pi12 ? n32 : n82992;
  assign n82994 = pi11 ? n32 : n82993;
  assign n82995 = pi10 ? n32 : n82994;
  assign n82996 = pi19 ? n365 : ~n1574;
  assign n82997 = pi18 ? n32 : n82996;
  assign n82998 = pi17 ? n32 : n82997;
  assign n82999 = pi16 ? n32 : n82998;
  assign n83000 = pi15 ? n82999 : n82890;
  assign n83001 = pi14 ? n83000 : n82890;
  assign n83002 = pi13 ? n83001 : n82694;
  assign n83003 = pi19 ? n343 : ~n2141;
  assign n83004 = pi18 ? n32 : n83003;
  assign n83005 = pi17 ? n32 : n83004;
  assign n83006 = pi16 ? n32 : n83005;
  assign n83007 = pi19 ? n589 : ~n2141;
  assign n83008 = pi18 ? n32 : n83007;
  assign n83009 = pi17 ? n32 : n83008;
  assign n83010 = pi16 ? n32 : n83009;
  assign n83011 = pi15 ? n83006 : n83010;
  assign n83012 = pi19 ? n2848 : ~n2141;
  assign n83013 = pi18 ? n32 : n83012;
  assign n83014 = pi17 ? n32 : n83013;
  assign n83015 = pi16 ? n32 : n83014;
  assign n83016 = pi15 ? n83010 : n83015;
  assign n83017 = pi14 ? n83011 : n83016;
  assign n83018 = pi13 ? n82801 : n83017;
  assign n83019 = pi12 ? n83002 : n83018;
  assign n83020 = pi18 ? n32 : n31093;
  assign n83021 = pi17 ? n32 : n83020;
  assign n83022 = pi16 ? n32 : n83021;
  assign n83023 = pi19 ? n349 : ~n519;
  assign n83024 = pi18 ? n32 : n83023;
  assign n83025 = pi17 ? n32 : n83024;
  assign n83026 = pi16 ? n32 : n83025;
  assign n83027 = pi14 ? n83022 : n83026;
  assign n83028 = pi19 ? n813 : ~n1476;
  assign n83029 = pi18 ? n32 : n83028;
  assign n83030 = pi17 ? n32 : n83029;
  assign n83031 = pi16 ? n32 : n83030;
  assign n83032 = pi15 ? n13200 : n83031;
  assign n83033 = pi14 ? n83026 : n83032;
  assign n83034 = pi13 ? n83027 : n83033;
  assign n83035 = pi19 ? n1941 : ~n1476;
  assign n83036 = pi18 ? n32 : n83035;
  assign n83037 = pi17 ? n32 : n83036;
  assign n83038 = pi16 ? n32 : n83037;
  assign n83039 = pi15 ? n83038 : n13220;
  assign n83040 = pi14 ? n83038 : n83039;
  assign n83041 = pi19 ? n1941 : ~n244;
  assign n83042 = pi18 ? n32 : n83041;
  assign n83043 = pi17 ? n32 : n83042;
  assign n83044 = pi16 ? n32 : n83043;
  assign n83045 = pi19 ? n236 : ~n244;
  assign n83046 = pi18 ? n32 : n83045;
  assign n83047 = pi17 ? n32 : n83046;
  assign n83048 = pi16 ? n32 : n83047;
  assign n83049 = pi19 ? n2614 : ~n244;
  assign n83050 = pi18 ? n32 : n83049;
  assign n83051 = pi17 ? n32 : n83050;
  assign n83052 = pi16 ? n32 : n83051;
  assign n83053 = pi15 ? n83048 : n83052;
  assign n83054 = pi14 ? n83044 : n83053;
  assign n83055 = pi13 ? n83040 : n83054;
  assign n83056 = pi12 ? n83034 : n83055;
  assign n83057 = pi11 ? n83019 : n83056;
  assign n83058 = pi19 ? n2614 : ~n2297;
  assign n83059 = pi18 ? n32 : n83058;
  assign n83060 = pi17 ? n32 : n83059;
  assign n83061 = pi16 ? n32 : n83060;
  assign n83062 = pi15 ? n13244 : n83061;
  assign n83063 = pi14 ? n83062 : n83061;
  assign n83064 = pi15 ? n83061 : n13255;
  assign n83065 = pi19 ? n617 : ~n2317;
  assign n83066 = pi18 ? n32 : n83065;
  assign n83067 = pi17 ? n32 : n83066;
  assign n83068 = pi16 ? n32 : n83067;
  assign n83069 = pi15 ? n83068 : n13285;
  assign n83070 = pi14 ? n83064 : n83069;
  assign n83071 = pi13 ? n83063 : n83070;
  assign n83072 = pi15 ? n13285 : n13293;
  assign n83073 = pi14 ? n13285 : n83072;
  assign n83074 = pi19 ? n2614 : ~n1941;
  assign n83075 = pi18 ? n32 : n83074;
  assign n83076 = pi17 ? n32 : n83075;
  assign n83077 = pi16 ? n32 : n83076;
  assign n83078 = pi15 ? n13299 : n83077;
  assign n83079 = pi15 ? n13309 : n83077;
  assign n83080 = pi14 ? n83078 : n83079;
  assign n83081 = pi13 ? n83073 : n83080;
  assign n83082 = pi12 ? n83071 : n83081;
  assign n83083 = pi14 ? n13338 : n13350;
  assign n83084 = pi13 ? n13329 : n83083;
  assign n83085 = pi12 ? n83084 : n13395;
  assign n83086 = pi11 ? n83082 : n83085;
  assign n83087 = pi10 ? n83057 : n83086;
  assign n83088 = pi09 ? n82995 : n83087;
  assign n83089 = pi08 ? n82981 : n83088;
  assign n83090 = pi19 ? n1969 : ~n594;
  assign n83091 = pi18 ? n32 : n83090;
  assign n83092 = pi17 ? n32 : n83091;
  assign n83093 = pi16 ? n32 : n83092;
  assign n83094 = pi15 ? n32 : n83093;
  assign n83095 = pi19 ? n1969 : ~n1574;
  assign n83096 = pi18 ? n32 : n83095;
  assign n83097 = pi17 ? n32 : n83096;
  assign n83098 = pi16 ? n32 : n83097;
  assign n83099 = pi14 ? n83094 : n83098;
  assign n83100 = pi13 ? n32 : n83099;
  assign n83101 = pi12 ? n32 : n83100;
  assign n83102 = pi11 ? n32 : n83101;
  assign n83103 = pi10 ? n32 : n83102;
  assign n83104 = pi19 ? n208 : ~n1574;
  assign n83105 = pi18 ? n32 : n83104;
  assign n83106 = pi17 ? n32 : n83105;
  assign n83107 = pi16 ? n32 : n83106;
  assign n83108 = pi19 ? n244 : ~n1574;
  assign n83109 = pi18 ? n32 : n83108;
  assign n83110 = pi17 ? n32 : n83109;
  assign n83111 = pi16 ? n32 : n83110;
  assign n83112 = pi15 ? n83107 : n83111;
  assign n83113 = pi14 ? n83112 : n82990;
  assign n83114 = pi13 ? n83113 : n82899;
  assign n83115 = pi15 ? n82899 : n82792;
  assign n83116 = pi14 ? n82899 : n83115;
  assign n83117 = pi19 ? n2303 : ~n2141;
  assign n83118 = pi18 ? n32 : n83117;
  assign n83119 = pi17 ? n32 : n83118;
  assign n83120 = pi16 ? n32 : n83119;
  assign n83121 = pi13 ? n83116 : n83120;
  assign n83122 = pi12 ? n83114 : n83121;
  assign n83123 = pi18 ? n32 : n56298;
  assign n83124 = pi17 ? n32 : n83123;
  assign n83125 = pi16 ? n32 : n83124;
  assign n83126 = pi18 ? n32 : n28423;
  assign n83127 = pi17 ? n32 : n83126;
  assign n83128 = pi16 ? n32 : n83127;
  assign n83129 = pi14 ? n83125 : n83128;
  assign n83130 = pi19 ? n2317 : ~n519;
  assign n83131 = pi18 ? n32 : n83130;
  assign n83132 = pi17 ? n32 : n83131;
  assign n83133 = pi16 ? n32 : n83132;
  assign n83134 = pi15 ? n83128 : n83133;
  assign n83135 = pi19 ? n2317 : ~n1840;
  assign n83136 = pi18 ? n32 : n83135;
  assign n83137 = pi17 ? n32 : n83136;
  assign n83138 = pi16 ? n32 : n83137;
  assign n83139 = pi19 ? n589 : ~n1476;
  assign n83140 = pi18 ? n32 : n83139;
  assign n83141 = pi17 ? n32 : n83140;
  assign n83142 = pi16 ? n32 : n83141;
  assign n83143 = pi15 ? n83138 : n83142;
  assign n83144 = pi14 ? n83134 : n83143;
  assign n83145 = pi13 ? n83129 : n83144;
  assign n83146 = pi19 ? n2848 : ~n1476;
  assign n83147 = pi18 ? n32 : n83146;
  assign n83148 = pi17 ? n32 : n83147;
  assign n83149 = pi16 ? n32 : n83148;
  assign n83150 = pi19 ? n2848 : ~n750;
  assign n83151 = pi18 ? n32 : n83150;
  assign n83152 = pi17 ? n32 : n83151;
  assign n83153 = pi16 ? n32 : n83152;
  assign n83154 = pi15 ? n83149 : n83153;
  assign n83155 = pi14 ? n83149 : n83154;
  assign n83156 = pi19 ? n2848 : ~n244;
  assign n83157 = pi18 ? n32 : n83156;
  assign n83158 = pi17 ? n32 : n83157;
  assign n83159 = pi16 ? n32 : n83158;
  assign n83160 = pi19 ? n349 : ~n244;
  assign n83161 = pi18 ? n32 : n83160;
  assign n83162 = pi17 ? n32 : n83161;
  assign n83163 = pi16 ? n32 : n83162;
  assign n83164 = pi19 ? n1812 : ~n244;
  assign n83165 = pi18 ? n32 : n83164;
  assign n83166 = pi17 ? n32 : n83165;
  assign n83167 = pi16 ? n32 : n83166;
  assign n83168 = pi15 ? n83163 : n83167;
  assign n83169 = pi14 ? n83159 : n83168;
  assign n83170 = pi13 ? n83155 : n83169;
  assign n83171 = pi12 ? n83145 : n83170;
  assign n83172 = pi11 ? n83122 : n83171;
  assign n83173 = pi19 ? n1812 : ~n340;
  assign n83174 = pi18 ? n32 : n83173;
  assign n83175 = pi17 ? n32 : n83174;
  assign n83176 = pi16 ? n32 : n83175;
  assign n83177 = pi15 ? n83176 : n13556;
  assign n83178 = pi14 ? n83177 : n13556;
  assign n83179 = pi19 ? n813 : ~n2317;
  assign n83180 = pi18 ? n32 : n83179;
  assign n83181 = pi17 ? n32 : n83180;
  assign n83182 = pi16 ? n32 : n83181;
  assign n83183 = pi15 ? n83182 : n13575;
  assign n83184 = pi14 ? n13561 : n83183;
  assign n83185 = pi13 ? n83178 : n83184;
  assign n83186 = pi19 ? n1941 : ~n1812;
  assign n83187 = pi18 ? n32 : n83186;
  assign n83188 = pi17 ? n32 : n83187;
  assign n83189 = pi16 ? n32 : n83188;
  assign n83190 = pi15 ? n83189 : n13595;
  assign n83191 = pi14 ? n13575 : n83190;
  assign n83192 = pi13 ? n83191 : n13611;
  assign n83193 = pi12 ? n83185 : n83192;
  assign n83194 = pi11 ? n83193 : n13688;
  assign n83195 = pi10 ? n83172 : n83194;
  assign n83196 = pi09 ? n83103 : n83195;
  assign n83197 = pi19 ? n1476 : ~n594;
  assign n83198 = pi18 ? n32 : n83197;
  assign n83199 = pi17 ? n32 : n83198;
  assign n83200 = pi16 ? n32 : n83199;
  assign n83201 = pi15 ? n32 : n83200;
  assign n83202 = pi19 ? n1476 : ~n1574;
  assign n83203 = pi18 ? n32 : n83202;
  assign n83204 = pi17 ? n32 : n83203;
  assign n83205 = pi16 ? n32 : n83204;
  assign n83206 = pi14 ? n83201 : n83205;
  assign n83207 = pi13 ? n32 : n83206;
  assign n83208 = pi12 ? n32 : n83207;
  assign n83209 = pi11 ? n32 : n83208;
  assign n83210 = pi10 ? n32 : n83209;
  assign n83211 = pi19 ? n750 : ~n1574;
  assign n83212 = pi18 ? n32 : n83211;
  assign n83213 = pi17 ? n32 : n83212;
  assign n83214 = pi16 ? n32 : n83213;
  assign n83215 = pi15 ? n83214 : n83098;
  assign n83216 = pi15 ? n83098 : n82990;
  assign n83217 = pi14 ? n83215 : n83216;
  assign n83218 = pi13 ? n83217 : n82999;
  assign n83219 = pi19 ? n2297 : ~n2141;
  assign n83220 = pi18 ? n32 : n83219;
  assign n83221 = pi17 ? n32 : n83220;
  assign n83222 = pi16 ? n32 : n83221;
  assign n83223 = pi13 ? n82890 : n83222;
  assign n83224 = pi12 ? n83218 : n83223;
  assign n83225 = pi19 ? n2297 : ~n507;
  assign n83226 = pi18 ? n32 : n83225;
  assign n83227 = pi17 ? n32 : n83226;
  assign n83228 = pi16 ? n32 : n83227;
  assign n83229 = pi19 ? n2297 : ~n519;
  assign n83230 = pi18 ? n32 : n83229;
  assign n83231 = pi17 ? n32 : n83230;
  assign n83232 = pi16 ? n32 : n83231;
  assign n83233 = pi15 ? n83228 : n83232;
  assign n83234 = pi19 ? n429 : ~n519;
  assign n83235 = pi18 ? n32 : n83234;
  assign n83236 = pi17 ? n32 : n83235;
  assign n83237 = pi16 ? n32 : n83236;
  assign n83238 = pi15 ? n83232 : n83237;
  assign n83239 = pi14 ? n83233 : n83238;
  assign n83240 = pi19 ? n429 : ~n1840;
  assign n83241 = pi18 ? n32 : n83240;
  assign n83242 = pi17 ? n32 : n83241;
  assign n83243 = pi16 ? n32 : n83242;
  assign n83244 = pi15 ? n83237 : n83243;
  assign n83245 = pi19 ? n429 : ~n1476;
  assign n83246 = pi18 ? n32 : n83245;
  assign n83247 = pi17 ? n32 : n83246;
  assign n83248 = pi16 ? n32 : n83247;
  assign n83249 = pi14 ? n83244 : n83248;
  assign n83250 = pi13 ? n83239 : n83249;
  assign n83251 = pi19 ? n2303 : ~n1476;
  assign n83252 = pi18 ? n32 : n83251;
  assign n83253 = pi17 ? n32 : n83252;
  assign n83254 = pi16 ? n32 : n83253;
  assign n83255 = pi19 ? n2303 : ~n750;
  assign n83256 = pi18 ? n32 : n83255;
  assign n83257 = pi17 ? n32 : n83256;
  assign n83258 = pi16 ? n32 : n83257;
  assign n83259 = pi19 ? n2303 : ~n244;
  assign n83260 = pi18 ? n32 : n83259;
  assign n83261 = pi17 ? n32 : n83260;
  assign n83262 = pi16 ? n32 : n83261;
  assign n83263 = pi15 ? n83258 : n83262;
  assign n83264 = pi14 ? n83254 : n83263;
  assign n83265 = pi19 ? n343 : ~n244;
  assign n83266 = pi18 ? n32 : n83265;
  assign n83267 = pi17 ? n32 : n83266;
  assign n83268 = pi16 ? n32 : n83267;
  assign n83269 = pi15 ? n83262 : n83268;
  assign n83270 = pi19 ? n2317 : ~n244;
  assign n83271 = pi18 ? n32 : n83270;
  assign n83272 = pi17 ? n32 : n83271;
  assign n83273 = pi16 ? n32 : n83272;
  assign n83274 = pi15 ? n83268 : n83273;
  assign n83275 = pi14 ? n83269 : n83274;
  assign n83276 = pi13 ? n83264 : n83275;
  assign n83277 = pi12 ? n83250 : n83276;
  assign n83278 = pi11 ? n83224 : n83277;
  assign n83279 = pi15 ? n13830 : n13839;
  assign n83280 = pi14 ? n83279 : n13839;
  assign n83281 = pi19 ? n589 : ~n2317;
  assign n83282 = pi18 ? n32 : n83281;
  assign n83283 = pi17 ? n32 : n83282;
  assign n83284 = pi16 ? n32 : n83283;
  assign n83285 = pi15 ? n83284 : n13869;
  assign n83286 = pi14 ? n13850 : n83285;
  assign n83287 = pi13 ? n83280 : n83286;
  assign n83288 = pi14 ? n13869 : n13879;
  assign n83289 = pi13 ? n83288 : n13894;
  assign n83290 = pi12 ? n83287 : n83289;
  assign n83291 = pi11 ? n83290 : n13956;
  assign n83292 = pi10 ? n83278 : n83291;
  assign n83293 = pi09 ? n83210 : n83292;
  assign n83294 = pi08 ? n83196 : n83293;
  assign n83295 = pi07 ? n83089 : n83294;
  assign n83296 = pi06 ? n82881 : n83295;
  assign n83297 = pi05 ? n82465 : n83296;
  assign n83298 = pi04 ? n81430 : n83297;
  assign n83299 = pi19 ? n1840 : ~n594;
  assign n83300 = pi18 ? n32 : n83299;
  assign n83301 = pi17 ? n32 : n83300;
  assign n83302 = pi16 ? n32 : n83301;
  assign n83303 = pi15 ? n32 : n83302;
  assign n83304 = pi19 ? n1840 : ~n1574;
  assign n83305 = pi18 ? n32 : n83304;
  assign n83306 = pi17 ? n32 : n83305;
  assign n83307 = pi16 ? n32 : n83306;
  assign n83308 = pi14 ? n83303 : n83307;
  assign n83309 = pi13 ? n32 : n83308;
  assign n83310 = pi12 ? n32 : n83309;
  assign n83311 = pi11 ? n32 : n83310;
  assign n83312 = pi10 ? n32 : n83311;
  assign n83313 = pi19 ? n322 : ~n1574;
  assign n83314 = pi18 ? n32 : n83313;
  assign n83315 = pi17 ? n32 : n83314;
  assign n83316 = pi16 ? n32 : n83315;
  assign n83317 = pi15 ? n83316 : n83205;
  assign n83318 = pi15 ? n83205 : n83098;
  assign n83319 = pi14 ? n83317 : n83318;
  assign n83320 = pi13 ? n83319 : n83107;
  assign n83321 = pi14 ? n83111 : n82990;
  assign n83322 = pi19 ? n365 : ~n2141;
  assign n83323 = pi18 ? n32 : n83322;
  assign n83324 = pi17 ? n32 : n83323;
  assign n83325 = pi16 ? n32 : n83324;
  assign n83326 = pi13 ? n83321 : n83325;
  assign n83327 = pi12 ? n83320 : n83326;
  assign n83328 = pi19 ? n531 : ~n507;
  assign n83329 = pi18 ? n32 : n83328;
  assign n83330 = pi17 ? n32 : n83329;
  assign n83331 = pi16 ? n32 : n83330;
  assign n83332 = pi19 ? n531 : ~n519;
  assign n83333 = pi18 ? n32 : n83332;
  assign n83334 = pi17 ? n32 : n83333;
  assign n83335 = pi16 ? n32 : n83334;
  assign n83336 = pi15 ? n83331 : n83335;
  assign n83337 = pi14 ? n83336 : n83335;
  assign n83338 = pi19 ? n531 : ~n1840;
  assign n83339 = pi18 ? n32 : n83338;
  assign n83340 = pi17 ? n32 : n83339;
  assign n83341 = pi16 ? n32 : n83340;
  assign n83342 = pi15 ? n83335 : n83341;
  assign n83343 = pi19 ? n531 : ~n1476;
  assign n83344 = pi18 ? n32 : n83343;
  assign n83345 = pi17 ? n32 : n83344;
  assign n83346 = pi16 ? n32 : n83345;
  assign n83347 = pi14 ? n83342 : n83346;
  assign n83348 = pi13 ? n83337 : n83347;
  assign n83349 = pi19 ? n531 : ~n750;
  assign n83350 = pi18 ? n32 : n83349;
  assign n83351 = pi17 ? n32 : n83350;
  assign n83352 = pi16 ? n32 : n83351;
  assign n83353 = pi19 ? n2297 : ~n244;
  assign n83354 = pi18 ? n32 : n83353;
  assign n83355 = pi17 ? n32 : n83354;
  assign n83356 = pi16 ? n32 : n83355;
  assign n83357 = pi15 ? n83352 : n83356;
  assign n83358 = pi14 ? n83346 : n83357;
  assign n83359 = pi15 ? n83356 : n14064;
  assign n83360 = pi14 ? n83356 : n83359;
  assign n83361 = pi13 ? n83358 : n83360;
  assign n83362 = pi12 ? n83348 : n83361;
  assign n83363 = pi11 ? n83327 : n83362;
  assign n83364 = pi15 ? n13733 : n14096;
  assign n83365 = pi15 ? n14096 : n14105;
  assign n83366 = pi14 ? n83364 : n83365;
  assign n83367 = pi13 ? n14087 : n83366;
  assign n83368 = pi19 ? n2303 : ~n1941;
  assign n83369 = pi18 ? n32 : n83368;
  assign n83370 = pi17 ? n32 : n83369;
  assign n83371 = pi16 ? n32 : n83370;
  assign n83372 = pi15 ? n14116 : n83371;
  assign n83373 = pi14 ? n14112 : n83372;
  assign n83374 = pi13 ? n83373 : n14133;
  assign n83375 = pi12 ? n83367 : n83374;
  assign n83376 = pi14 ? n14157 : n14164;
  assign n83377 = pi13 ? n14149 : n83376;
  assign n83378 = pi12 ? n83377 : n32;
  assign n83379 = pi11 ? n83375 : n83378;
  assign n83380 = pi10 ? n83363 : n83379;
  assign n83381 = pi09 ? n83312 : n83380;
  assign n83382 = pi19 ? n519 : ~n594;
  assign n83383 = pi18 ? n32 : n83382;
  assign n83384 = pi17 ? n32 : n83383;
  assign n83385 = pi16 ? n32 : n83384;
  assign n83386 = pi15 ? n32 : n83385;
  assign n83387 = pi19 ? n519 : ~n1574;
  assign n83388 = pi18 ? n32 : n83387;
  assign n83389 = pi17 ? n32 : n83388;
  assign n83390 = pi16 ? n32 : n83389;
  assign n83391 = pi14 ? n83386 : n83390;
  assign n83392 = pi13 ? n32 : n83391;
  assign n83393 = pi12 ? n32 : n83392;
  assign n83394 = pi11 ? n32 : n83393;
  assign n83395 = pi10 ? n32 : n83394;
  assign n83396 = pi15 ? n83390 : n83307;
  assign n83397 = pi15 ? n83307 : n83205;
  assign n83398 = pi14 ? n83396 : n83397;
  assign n83399 = pi13 ? n83398 : n83214;
  assign n83400 = pi18 ? n32 : n18856;
  assign n83401 = pi17 ? n32 : n83400;
  assign n83402 = pi16 ? n32 : n83401;
  assign n83403 = pi13 ? n83098 : n83402;
  assign n83404 = pi12 ? n83399 : n83403;
  assign n83405 = pi19 ? n244 : ~n507;
  assign n83406 = pi18 ? n32 : n83405;
  assign n83407 = pi17 ? n32 : n83406;
  assign n83408 = pi16 ? n32 : n83407;
  assign n83409 = pi19 ? n244 : ~n519;
  assign n83410 = pi18 ? n32 : n83409;
  assign n83411 = pi17 ? n32 : n83410;
  assign n83412 = pi16 ? n32 : n83411;
  assign n83413 = pi15 ? n83408 : n83412;
  assign n83414 = pi19 ? n340 : ~n519;
  assign n83415 = pi18 ? n32 : n83414;
  assign n83416 = pi17 ? n32 : n83415;
  assign n83417 = pi16 ? n32 : n83416;
  assign n83418 = pi14 ? n83413 : n83417;
  assign n83419 = pi19 ? n340 : ~n1840;
  assign n83420 = pi18 ? n32 : n83419;
  assign n83421 = pi17 ? n32 : n83420;
  assign n83422 = pi16 ? n32 : n83421;
  assign n83423 = pi15 ? n83417 : n83422;
  assign n83424 = pi19 ? n340 : ~n1476;
  assign n83425 = pi18 ? n32 : n83424;
  assign n83426 = pi17 ? n32 : n83425;
  assign n83427 = pi16 ? n32 : n83426;
  assign n83428 = pi14 ? n83423 : n83427;
  assign n83429 = pi13 ? n83418 : n83428;
  assign n83430 = pi19 ? n365 : ~n1476;
  assign n83431 = pi18 ? n32 : n83430;
  assign n83432 = pi17 ? n32 : n83431;
  assign n83433 = pi16 ? n32 : n83432;
  assign n83434 = pi19 ? n365 : ~n750;
  assign n83435 = pi18 ? n32 : n83434;
  assign n83436 = pi17 ? n32 : n83435;
  assign n83437 = pi16 ? n32 : n83436;
  assign n83438 = pi19 ? n365 : ~n244;
  assign n83439 = pi18 ? n32 : n83438;
  assign n83440 = pi17 ? n32 : n83439;
  assign n83441 = pi16 ? n32 : n83440;
  assign n83442 = pi15 ? n83437 : n83441;
  assign n83443 = pi14 ? n83433 : n83442;
  assign n83444 = pi19 ? n340 : ~n340;
  assign n83445 = pi18 ? n32 : n83444;
  assign n83446 = pi17 ? n32 : n83445;
  assign n83447 = pi16 ? n32 : n83446;
  assign n83448 = pi15 ? n83441 : n83447;
  assign n83449 = pi14 ? n83441 : n83448;
  assign n83450 = pi13 ? n83443 : n83449;
  assign n83451 = pi12 ? n83429 : n83450;
  assign n83452 = pi11 ? n83404 : n83451;
  assign n83453 = pi15 ? n14315 : n14306;
  assign n83454 = pi15 ? n14306 : n14315;
  assign n83455 = pi14 ? n83453 : n83454;
  assign n83456 = pi15 ? n14005 : n14327;
  assign n83457 = pi14 ? n83456 : n14333;
  assign n83458 = pi13 ? n83455 : n83457;
  assign n83459 = pi19 ? n365 : ~n1812;
  assign n83460 = pi18 ? n32 : n83459;
  assign n83461 = pi17 ? n32 : n83460;
  assign n83462 = pi16 ? n32 : n83461;
  assign n83463 = pi15 ? n14339 : n83462;
  assign n83464 = pi14 ? n83463 : n14349;
  assign n83465 = pi14 ? n14359 : n40239;
  assign n83466 = pi13 ? n83464 : n83465;
  assign n83467 = pi12 ? n83458 : n83466;
  assign n83468 = pi11 ? n83467 : n14408;
  assign n83469 = pi10 ? n83452 : n83468;
  assign n83470 = pi09 ? n83395 : n83469;
  assign n83471 = pi08 ? n83381 : n83470;
  assign n83472 = pi19 ? n507 : ~n594;
  assign n83473 = pi18 ? n32 : n83472;
  assign n83474 = pi17 ? n32 : n83473;
  assign n83475 = pi16 ? n32 : n83474;
  assign n83476 = pi15 ? n32 : n83475;
  assign n83477 = pi18 ? n32 : n18997;
  assign n83478 = pi17 ? n32 : n83477;
  assign n83479 = pi16 ? n32 : n83478;
  assign n83480 = pi14 ? n83476 : n83479;
  assign n83481 = pi13 ? n32 : n83480;
  assign n83482 = pi12 ? n32 : n83481;
  assign n83483 = pi11 ? n32 : n83482;
  assign n83484 = pi10 ? n32 : n83483;
  assign n83485 = pi19 ? n1320 : ~n1574;
  assign n83486 = pi18 ? n32 : n83485;
  assign n83487 = pi17 ? n32 : n83486;
  assign n83488 = pi16 ? n32 : n83487;
  assign n83489 = pi15 ? n83488 : n83390;
  assign n83490 = pi14 ? n83489 : n83396;
  assign n83491 = pi13 ? n83490 : n83316;
  assign n83492 = pi19 ? n750 : ~n2141;
  assign n83493 = pi18 ? n32 : n83492;
  assign n83494 = pi17 ? n32 : n83493;
  assign n83495 = pi16 ? n32 : n83494;
  assign n83496 = pi13 ? n83205 : n83495;
  assign n83497 = pi12 ? n83491 : n83496;
  assign n83498 = pi19 ? n1969 : ~n507;
  assign n83499 = pi18 ? n32 : n83498;
  assign n83500 = pi17 ? n32 : n83499;
  assign n83501 = pi16 ? n32 : n83500;
  assign n83502 = pi19 ? n1969 : ~n519;
  assign n83503 = pi18 ? n32 : n83502;
  assign n83504 = pi17 ? n32 : n83503;
  assign n83505 = pi16 ? n32 : n83504;
  assign n83506 = pi15 ? n83501 : n83505;
  assign n83507 = pi14 ? n83506 : n83505;
  assign n83508 = pi19 ? n1969 : ~n1840;
  assign n83509 = pi18 ? n32 : n83508;
  assign n83510 = pi17 ? n32 : n83509;
  assign n83511 = pi16 ? n32 : n83510;
  assign n83512 = pi15 ? n83505 : n83511;
  assign n83513 = pi19 ? n1969 : ~n1476;
  assign n83514 = pi18 ? n32 : n83513;
  assign n83515 = pi17 ? n32 : n83514;
  assign n83516 = pi16 ? n32 : n83515;
  assign n83517 = pi14 ? n83512 : n83516;
  assign n83518 = pi13 ? n83507 : n83517;
  assign n83519 = pi19 ? n208 : ~n1476;
  assign n83520 = pi18 ? n32 : n83519;
  assign n83521 = pi17 ? n32 : n83520;
  assign n83522 = pi16 ? n32 : n83521;
  assign n83523 = pi19 ? n244 : ~n750;
  assign n83524 = pi18 ? n32 : n83523;
  assign n83525 = pi17 ? n32 : n83524;
  assign n83526 = pi16 ? n32 : n83525;
  assign n83527 = pi19 ? n244 : ~n244;
  assign n83528 = pi18 ? n32 : n83527;
  assign n83529 = pi17 ? n32 : n83528;
  assign n83530 = pi16 ? n32 : n83529;
  assign n83531 = pi15 ? n83526 : n83530;
  assign n83532 = pi14 ? n83522 : n83531;
  assign n83533 = pi15 ? n83530 : n13423;
  assign n83534 = pi14 ? n83530 : n83533;
  assign n83535 = pi13 ? n83532 : n83534;
  assign n83536 = pi12 ? n83518 : n83535;
  assign n83537 = pi11 ? n83497 : n83536;
  assign n83538 = pi19 ? n244 : ~n2297;
  assign n83539 = pi18 ? n32 : n83538;
  assign n83540 = pi17 ? n32 : n83539;
  assign n83541 = pi16 ? n32 : n83540;
  assign n83542 = pi15 ? n83541 : n14219;
  assign n83543 = pi14 ? n83541 : n83542;
  assign n83544 = pi15 ? n14207 : n14488;
  assign n83545 = pi19 ? n340 : ~n589;
  assign n83546 = pi18 ? n32 : n83545;
  assign n83547 = pi17 ? n32 : n83546;
  assign n83548 = pi16 ? n32 : n83547;
  assign n83549 = pi19 ? n340 : ~n1812;
  assign n83550 = pi18 ? n32 : n83549;
  assign n83551 = pi17 ? n32 : n83550;
  assign n83552 = pi16 ? n32 : n83551;
  assign n83553 = pi15 ? n83548 : n83552;
  assign n83554 = pi14 ? n83544 : n83553;
  assign n83555 = pi13 ? n83543 : n83554;
  assign n83556 = pi15 ? n14566 : n24443;
  assign n83557 = pi14 ? n83556 : n14576;
  assign n83558 = pi13 ? n83557 : n14586;
  assign n83559 = pi12 ? n83555 : n83558;
  assign n83560 = pi11 ? n83559 : n14616;
  assign n83561 = pi10 ? n83537 : n83560;
  assign n83562 = pi09 ? n83484 : n83561;
  assign n83563 = pi19 ? n594 : ~n594;
  assign n83564 = pi18 ? n32 : n83563;
  assign n83565 = pi17 ? n32 : n83564;
  assign n83566 = pi16 ? n32 : n83565;
  assign n83567 = pi15 ? n32 : n83566;
  assign n83568 = pi19 ? n594 : ~n1574;
  assign n83569 = pi18 ? n32 : n83568;
  assign n83570 = pi17 ? n32 : n83569;
  assign n83571 = pi16 ? n32 : n83570;
  assign n83572 = pi14 ? n83567 : n83571;
  assign n83573 = pi13 ? n32 : n83572;
  assign n83574 = pi12 ? n32 : n83573;
  assign n83575 = pi11 ? n32 : n83574;
  assign n83576 = pi10 ? n32 : n83575;
  assign n83577 = pi19 ? n2141 : ~n1574;
  assign n83578 = pi18 ? n32 : n83577;
  assign n83579 = pi17 ? n32 : n83578;
  assign n83580 = pi16 ? n32 : n83579;
  assign n83581 = pi15 ? n83580 : n83479;
  assign n83582 = pi15 ? n83479 : n83390;
  assign n83583 = pi14 ? n83581 : n83582;
  assign n83584 = pi13 ? n83583 : n83307;
  assign n83585 = pi19 ? n322 : ~n2141;
  assign n83586 = pi18 ? n32 : n83585;
  assign n83587 = pi17 ? n32 : n83586;
  assign n83588 = pi16 ? n32 : n83587;
  assign n83589 = pi13 ? n83307 : n83588;
  assign n83590 = pi12 ? n83584 : n83589;
  assign n83591 = pi19 ? n1476 : ~n507;
  assign n83592 = pi18 ? n32 : n83591;
  assign n83593 = pi17 ? n32 : n83592;
  assign n83594 = pi16 ? n32 : n83593;
  assign n83595 = pi19 ? n1476 : ~n519;
  assign n83596 = pi18 ? n32 : n83595;
  assign n83597 = pi17 ? n32 : n83596;
  assign n83598 = pi16 ? n32 : n83597;
  assign n83599 = pi15 ? n83594 : n83598;
  assign n83600 = pi14 ? n83599 : n83598;
  assign n83601 = pi19 ? n1476 : ~n1840;
  assign n83602 = pi18 ? n32 : n83601;
  assign n83603 = pi17 ? n32 : n83602;
  assign n83604 = pi16 ? n32 : n83603;
  assign n83605 = pi15 ? n83598 : n83604;
  assign n83606 = pi19 ? n1476 : ~n1476;
  assign n83607 = pi18 ? n32 : n83606;
  assign n83608 = pi17 ? n32 : n83607;
  assign n83609 = pi16 ? n32 : n83608;
  assign n83610 = pi14 ? n83605 : n83609;
  assign n83611 = pi13 ? n83600 : n83610;
  assign n83612 = pi19 ? n750 : ~n1476;
  assign n83613 = pi18 ? n32 : n83612;
  assign n83614 = pi17 ? n32 : n83613;
  assign n83615 = pi16 ? n32 : n83614;
  assign n83616 = pi19 ? n750 : ~n750;
  assign n83617 = pi18 ? n32 : n83616;
  assign n83618 = pi17 ? n32 : n83617;
  assign n83619 = pi16 ? n32 : n83618;
  assign n83620 = pi19 ? n750 : ~n244;
  assign n83621 = pi18 ? n32 : n83620;
  assign n83622 = pi17 ? n32 : n83621;
  assign n83623 = pi16 ? n32 : n83622;
  assign n83624 = pi15 ? n83619 : n83623;
  assign n83625 = pi14 ? n83615 : n83624;
  assign n83626 = pi19 ? n1969 : ~n244;
  assign n83627 = pi18 ? n32 : n83626;
  assign n83628 = pi17 ? n32 : n83627;
  assign n83629 = pi16 ? n32 : n83628;
  assign n83630 = pi15 ? n83629 : n13710;
  assign n83631 = pi14 ? n83623 : n83630;
  assign n83632 = pi13 ? n83625 : n83631;
  assign n83633 = pi12 ? n83611 : n83632;
  assign n83634 = pi11 ? n83590 : n83633;
  assign n83635 = pi19 ? n1969 : ~n2297;
  assign n83636 = pi18 ? n32 : n83635;
  assign n83637 = pi17 ? n32 : n83636;
  assign n83638 = pi16 ? n32 : n83637;
  assign n83639 = pi19 ? n750 : ~n2297;
  assign n83640 = pi18 ? n32 : n83639;
  assign n83641 = pi17 ? n32 : n83640;
  assign n83642 = pi16 ? n32 : n83641;
  assign n83643 = pi15 ? n83638 : n83642;
  assign n83644 = pi15 ? n83638 : n13404;
  assign n83645 = pi14 ? n83643 : n83644;
  assign n83646 = pi15 ? n13404 : n14744;
  assign n83647 = pi15 ? n55212 : n14758;
  assign n83648 = pi14 ? n83646 : n83647;
  assign n83649 = pi13 ? n83645 : n83648;
  assign n83650 = pi19 ? n1969 : ~n1812;
  assign n83651 = pi18 ? n32 : n83650;
  assign n83652 = pi17 ? n32 : n83651;
  assign n83653 = pi16 ? n32 : n83652;
  assign n83654 = pi15 ? n83653 : n14758;
  assign n83655 = pi19 ? n1476 : ~n2614;
  assign n83656 = pi18 ? n32 : n83655;
  assign n83657 = pi17 ? n32 : n83656;
  assign n83658 = pi16 ? n32 : n83657;
  assign n83659 = pi15 ? n14765 : n83658;
  assign n83660 = pi14 ? n83654 : n83659;
  assign n83661 = pi13 ? n83660 : n14777;
  assign n83662 = pi12 ? n83649 : n83661;
  assign n83663 = pi11 ? n83662 : n14802;
  assign n83664 = pi10 ? n83634 : n83663;
  assign n83665 = pi09 ? n83576 : n83664;
  assign n83666 = pi08 ? n83562 : n83665;
  assign n83667 = pi07 ? n83471 : n83666;
  assign n83668 = pi15 ? n83571 : n83580;
  assign n83669 = pi14 ? n83668 : n83479;
  assign n83670 = pi13 ? n83669 : n83488;
  assign n83671 = pi19 ? n1840 : ~n2141;
  assign n83672 = pi18 ? n32 : n83671;
  assign n83673 = pi17 ? n32 : n83672;
  assign n83674 = pi16 ? n32 : n83673;
  assign n83675 = pi13 ? n83390 : n83674;
  assign n83676 = pi12 ? n83670 : n83675;
  assign n83677 = pi19 ? n1840 : ~n507;
  assign n83678 = pi18 ? n32 : n83677;
  assign n83679 = pi17 ? n32 : n83678;
  assign n83680 = pi16 ? n32 : n83679;
  assign n83681 = pi19 ? n1840 : ~n519;
  assign n83682 = pi18 ? n32 : n83681;
  assign n83683 = pi17 ? n32 : n83682;
  assign n83684 = pi16 ? n32 : n83683;
  assign n83685 = pi15 ? n83680 : n83684;
  assign n83686 = pi14 ? n83685 : n83684;
  assign n83687 = pi19 ? n1840 : ~n1840;
  assign n83688 = pi18 ? n32 : n83687;
  assign n83689 = pi17 ? n32 : n83688;
  assign n83690 = pi16 ? n32 : n83689;
  assign n83691 = pi15 ? n83684 : n83690;
  assign n83692 = pi19 ? n1840 : ~n1476;
  assign n83693 = pi18 ? n32 : n83692;
  assign n83694 = pi17 ? n32 : n83693;
  assign n83695 = pi16 ? n32 : n83694;
  assign n83696 = pi14 ? n83691 : n83695;
  assign n83697 = pi13 ? n83686 : n83696;
  assign n83698 = pi19 ? n322 : ~n1476;
  assign n83699 = pi18 ? n32 : n83698;
  assign n83700 = pi17 ? n32 : n83699;
  assign n83701 = pi16 ? n32 : n83700;
  assign n83702 = pi19 ? n322 : ~n750;
  assign n83703 = pi18 ? n32 : n83702;
  assign n83704 = pi17 ? n32 : n83703;
  assign n83705 = pi16 ? n32 : n83704;
  assign n83706 = pi15 ? n83705 : n14900;
  assign n83707 = pi14 ? n83701 : n83706;
  assign n83708 = pi15 ? n14900 : n13978;
  assign n83709 = pi14 ? n14900 : n83708;
  assign n83710 = pi13 ? n83707 : n83709;
  assign n83711 = pi12 ? n83697 : n83710;
  assign n83712 = pi11 ? n83676 : n83711;
  assign n83713 = pi15 ? n14895 : n14651;
  assign n83714 = pi14 ? n14909 : n83713;
  assign n83715 = pi17 ? n32 : n67116;
  assign n83716 = pi16 ? n32 : n83715;
  assign n83717 = pi15 ? n14651 : n83716;
  assign n83718 = pi14 ? n83717 : n14933;
  assign n83719 = pi13 ? n83714 : n83718;
  assign n83720 = pi19 ? n1840 : ~n2614;
  assign n83721 = pi18 ? n32 : n83720;
  assign n83722 = pi17 ? n32 : n83721;
  assign n83723 = pi16 ? n32 : n83722;
  assign n83724 = pi15 ? n25466 : n83723;
  assign n83725 = pi14 ? n14932 : n83724;
  assign n83726 = pi14 ? n14952 : n14958;
  assign n83727 = pi13 ? n83725 : n83726;
  assign n83728 = pi12 ? n83719 : n83727;
  assign n83729 = pi11 ? n83728 : n14978;
  assign n83730 = pi10 ? n83712 : n83729;
  assign n83731 = pi09 ? n83576 : n83730;
  assign n83732 = pi18 ? n32 : n29542;
  assign n83733 = pi17 ? n32 : n83732;
  assign n83734 = pi16 ? n32 : n83733;
  assign n83735 = pi15 ? n32 : n83734;
  assign n83736 = pi18 ? n32 : n29807;
  assign n83737 = pi17 ? n32 : n83736;
  assign n83738 = pi16 ? n32 : n83737;
  assign n83739 = pi14 ? n83735 : n83738;
  assign n83740 = pi13 ? n32 : n83739;
  assign n83741 = pi12 ? n32 : n83740;
  assign n83742 = pi11 ? n32 : n83741;
  assign n83743 = pi10 ? n32 : n83742;
  assign n83744 = pi19 ? n1574 : ~n1574;
  assign n83745 = pi18 ? n32 : n83744;
  assign n83746 = pi17 ? n32 : n83745;
  assign n83747 = pi16 ? n32 : n83746;
  assign n83748 = pi15 ? n83747 : n83571;
  assign n83749 = pi14 ? n83748 : n83580;
  assign n83750 = pi13 ? n83749 : n83580;
  assign n83751 = pi19 ? n1320 : ~n2141;
  assign n83752 = pi18 ? n32 : n83751;
  assign n83753 = pi17 ? n32 : n83752;
  assign n83754 = pi16 ? n32 : n83753;
  assign n83755 = pi13 ? n83479 : n83754;
  assign n83756 = pi12 ? n83750 : n83755;
  assign n83757 = pi19 ? n519 : ~n507;
  assign n83758 = pi18 ? n32 : n83757;
  assign n83759 = pi17 ? n32 : n83758;
  assign n83760 = pi16 ? n32 : n83759;
  assign n83761 = pi19 ? n519 : ~n519;
  assign n83762 = pi18 ? n32 : n83761;
  assign n83763 = pi17 ? n32 : n83762;
  assign n83764 = pi16 ? n32 : n83763;
  assign n83765 = pi15 ? n83760 : n83764;
  assign n83766 = pi14 ? n83765 : n83764;
  assign n83767 = pi19 ? n519 : ~n1840;
  assign n83768 = pi18 ? n32 : n83767;
  assign n83769 = pi17 ? n32 : n83768;
  assign n83770 = pi16 ? n32 : n83769;
  assign n83771 = pi15 ? n83764 : n83770;
  assign n83772 = pi14 ? n83771 : n72982;
  assign n83773 = pi13 ? n83766 : n83772;
  assign n83774 = pi19 ? n1840 : ~n244;
  assign n83775 = pi18 ? n32 : n83774;
  assign n83776 = pi17 ? n32 : n83775;
  assign n83777 = pi16 ? n32 : n83776;
  assign n83778 = pi15 ? n15046 : n83777;
  assign n83779 = pi14 ? n72982 : n83778;
  assign n83780 = pi19 ? n519 : ~n244;
  assign n83781 = pi18 ? n32 : n83780;
  assign n83782 = pi17 ? n32 : n83781;
  assign n83783 = pi16 ? n32 : n83782;
  assign n83784 = pi14 ? n83783 : n14179;
  assign n83785 = pi13 ? n83779 : n83784;
  assign n83786 = pi12 ? n83773 : n83785;
  assign n83787 = pi11 ? n83756 : n83786;
  assign n83788 = pi19 ? n519 : ~n2297;
  assign n83789 = pi18 ? n32 : n83788;
  assign n83790 = pi17 ? n32 : n83789;
  assign n83791 = pi16 ? n32 : n83790;
  assign n83792 = pi15 ? n83791 : n15066;
  assign n83793 = pi14 ? n83792 : n15075;
  assign n83794 = pi15 ? n15075 : n36095;
  assign n83795 = pi14 ? n83794 : n15091;
  assign n83796 = pi13 ? n83793 : n83795;
  assign n83797 = pi15 ? n73131 : n15090;
  assign n83798 = pi14 ? n83797 : n15110;
  assign n83799 = pi13 ? n83798 : n15124;
  assign n83800 = pi12 ? n83796 : n83799;
  assign n83801 = pi11 ? n83800 : n15130;
  assign n83802 = pi10 ? n83787 : n83801;
  assign n83803 = pi09 ? n83743 : n83802;
  assign n83804 = pi08 ? n83731 : n83803;
  assign n83805 = pi20 ? n339 : ~n428;
  assign n83806 = pi19 ? n32 : n83805;
  assign n83807 = pi18 ? n32 : n83806;
  assign n83808 = pi17 ? n32 : n83807;
  assign n83809 = pi16 ? n32 : n83808;
  assign n83810 = pi15 ? n32 : n83809;
  assign n83811 = pi20 ? n339 : ~n101;
  assign n83812 = pi19 ? n32 : n83811;
  assign n83813 = pi18 ? n32 : n83812;
  assign n83814 = pi17 ? n32 : n83813;
  assign n83815 = pi16 ? n32 : n83814;
  assign n83816 = pi14 ? n83810 : n83815;
  assign n83817 = pi13 ? n32 : n83816;
  assign n83818 = pi12 ? n32 : n83817;
  assign n83819 = pi11 ? n32 : n83818;
  assign n83820 = pi10 ? n32 : n83819;
  assign n83821 = pi20 ? n141 : ~n101;
  assign n83822 = pi19 ? n32 : n83821;
  assign n83823 = pi18 ? n32 : n83822;
  assign n83824 = pi17 ? n32 : n83823;
  assign n83825 = pi16 ? n32 : n83824;
  assign n83826 = pi15 ? n83825 : n83738;
  assign n83827 = pi14 ? n83826 : n83571;
  assign n83828 = pi13 ? n83827 : n83580;
  assign n83829 = pi19 ? n2141 : ~n2141;
  assign n83830 = pi18 ? n32 : n83829;
  assign n83831 = pi17 ? n32 : n83830;
  assign n83832 = pi16 ? n32 : n83831;
  assign n83833 = pi13 ? n83580 : n83832;
  assign n83834 = pi12 ? n83828 : n83833;
  assign n83835 = pi19 ? n507 : ~n507;
  assign n83836 = pi18 ? n32 : n83835;
  assign n83837 = pi17 ? n32 : n83836;
  assign n83838 = pi16 ? n32 : n83837;
  assign n83839 = pi15 ? n83838 : n15182;
  assign n83840 = pi14 ? n83839 : n15182;
  assign n83841 = pi14 ? n15187 : n15191;
  assign n83842 = pi13 ? n83840 : n83841;
  assign n83843 = pi19 ? n1320 : ~n208;
  assign n83844 = pi18 ? n32 : n83843;
  assign n83845 = pi17 ? n32 : n83844;
  assign n83846 = pi16 ? n32 : n83845;
  assign n83847 = pi15 ? n83846 : n15206;
  assign n83848 = pi14 ? n15198 : n83847;
  assign n83849 = pi14 ? n15206 : n14426;
  assign n83850 = pi13 ? n83848 : n83849;
  assign n83851 = pi12 ? n83842 : n83850;
  assign n83852 = pi11 ? n83834 : n83851;
  assign n83853 = pi15 ? n15221 : n37998;
  assign n83854 = pi14 ? n83853 : n15230;
  assign n83855 = pi13 ? n83854 : n15250;
  assign n83856 = pi12 ? n83855 : n15265;
  assign n83857 = pi11 ? n83856 : n15270;
  assign n83858 = pi10 ? n83852 : n83857;
  assign n83859 = pi09 ? n83820 : n83858;
  assign n83860 = pi14 ? n83815 : n83738;
  assign n83861 = pi13 ? n83860 : n83747;
  assign n83862 = pi13 ? n83571 : n83832;
  assign n83863 = pi12 ? n83861 : n83862;
  assign n83864 = pi15 ? n15296 : n15307;
  assign n83865 = pi14 ? n83864 : n15307;
  assign n83866 = pi14 ? n15312 : n15316;
  assign n83867 = pi13 ? n83865 : n83866;
  assign n83868 = pi19 ? n2141 : ~n208;
  assign n83869 = pi18 ? n32 : n83868;
  assign n83870 = pi17 ? n32 : n83869;
  assign n83871 = pi16 ? n32 : n83870;
  assign n83872 = pi15 ? n83871 : n15331;
  assign n83873 = pi14 ? n15323 : n83872;
  assign n83874 = pi14 ? n15338 : n14633;
  assign n83875 = pi13 ? n83873 : n83874;
  assign n83876 = pi12 ? n83867 : n83875;
  assign n83877 = pi11 ? n83863 : n83876;
  assign n83878 = pi19 ? n2141 : ~n429;
  assign n83879 = pi18 ? n32 : n83878;
  assign n83880 = pi17 ? n32 : n83879;
  assign n83881 = pi16 ? n32 : n83880;
  assign n83882 = pi15 ? n15347 : n83881;
  assign n83883 = pi14 ? n83882 : n15235;
  assign n83884 = pi13 ? n83883 : n15368;
  assign n83885 = pi12 ? n83884 : n15392;
  assign n83886 = pi11 ? n83885 : n32;
  assign n83887 = pi10 ? n83877 : n83886;
  assign n83888 = pi09 ? n83820 : n83887;
  assign n83889 = pi08 ? n83859 : n83888;
  assign n83890 = pi07 ? n83804 : n83889;
  assign n83891 = pi06 ? n83667 : n83890;
  assign n83892 = pi19 ? n32 : n13323;
  assign n83893 = pi18 ? n32 : n83892;
  assign n83894 = pi17 ? n32 : n83893;
  assign n83895 = pi16 ? n32 : n83894;
  assign n83896 = pi15 ? n32 : n83895;
  assign n83897 = pi19 ? n32 : n25089;
  assign n83898 = pi18 ? n32 : n83897;
  assign n83899 = pi17 ? n32 : n83898;
  assign n83900 = pi16 ? n32 : n83899;
  assign n83901 = pi20 ? n243 : ~n101;
  assign n83902 = pi19 ? n32 : n83901;
  assign n83903 = pi18 ? n32 : n83902;
  assign n83904 = pi17 ? n32 : n83903;
  assign n83905 = pi16 ? n32 : n83904;
  assign n83906 = pi15 ? n83900 : n83905;
  assign n83907 = pi14 ? n83896 : n83906;
  assign n83908 = pi13 ? n32 : n83907;
  assign n83909 = pi12 ? n32 : n83908;
  assign n83910 = pi11 ? n32 : n83909;
  assign n83911 = pi10 ? n32 : n83910;
  assign n83912 = pi15 ? n83905 : n83815;
  assign n83913 = pi14 ? n83912 : n83815;
  assign n83914 = pi13 ? n83913 : n83825;
  assign n83915 = pi19 ? n1574 : ~n2141;
  assign n83916 = pi18 ? n32 : n83915;
  assign n83917 = pi17 ? n32 : n83916;
  assign n83918 = pi16 ? n32 : n83917;
  assign n83919 = pi13 ? n83738 : n83918;
  assign n83920 = pi12 ? n83914 : n83919;
  assign n83921 = pi15 ? n15444 : n15459;
  assign n83922 = pi14 ? n83921 : n15459;
  assign n83923 = pi15 ? n15459 : n15316;
  assign n83924 = pi14 ? n83923 : n15316;
  assign n83925 = pi13 ? n83922 : n83924;
  assign n83926 = pi19 ? n594 : ~n244;
  assign n83927 = pi18 ? n32 : n83926;
  assign n83928 = pi17 ? n32 : n83927;
  assign n83929 = pi16 ? n32 : n83928;
  assign n83930 = pi15 ? n15476 : n83929;
  assign n83931 = pi14 ? n15477 : n83930;
  assign n83932 = pi13 ? n83931 : n15490;
  assign n83933 = pi12 ? n83925 : n83932;
  assign n83934 = pi11 ? n83920 : n83933;
  assign n83935 = pi10 ? n83934 : n15524;
  assign n83936 = pi09 ? n83911 : n83935;
  assign n83937 = pi19 ? n32 : n6323;
  assign n83938 = pi18 ? n32 : n83937;
  assign n83939 = pi17 ? n32 : n83938;
  assign n83940 = pi16 ? n32 : n83939;
  assign n83941 = pi15 ? n32 : n83940;
  assign n83942 = pi19 ? n32 : n66184;
  assign n83943 = pi18 ? n32 : n83942;
  assign n83944 = pi17 ? n32 : n83943;
  assign n83945 = pi16 ? n32 : n83944;
  assign n83946 = pi14 ? n83941 : n83945;
  assign n83947 = pi13 ? n32 : n83946;
  assign n83948 = pi12 ? n32 : n83947;
  assign n83949 = pi11 ? n32 : n83948;
  assign n83950 = pi10 ? n32 : n83949;
  assign n83951 = pi15 ? n83945 : n83815;
  assign n83952 = pi14 ? n83951 : n83815;
  assign n83953 = pi13 ? n83952 : n83825;
  assign n83954 = pi15 ? n83825 : n83815;
  assign n83955 = pi14 ? n83825 : n83954;
  assign n83956 = pi20 ? n141 : ~n2140;
  assign n83957 = pi19 ? n32 : n83956;
  assign n83958 = pi18 ? n32 : n83957;
  assign n83959 = pi17 ? n32 : n83958;
  assign n83960 = pi16 ? n32 : n83959;
  assign n83961 = pi13 ? n83955 : n83960;
  assign n83962 = pi12 ? n83953 : n83961;
  assign n83963 = pi15 ? n15573 : n15588;
  assign n83964 = pi14 ? n83963 : n15588;
  assign n83965 = pi15 ? n15588 : n71673;
  assign n83966 = pi14 ? n83965 : n71673;
  assign n83967 = pi13 ? n83964 : n83966;
  assign n83968 = pi19 ? n1574 : ~n244;
  assign n83969 = pi18 ? n32 : n83968;
  assign n83970 = pi17 ? n32 : n83969;
  assign n83971 = pi16 ? n32 : n83970;
  assign n83972 = pi15 ? n15608 : n83971;
  assign n83973 = pi14 ? n15609 : n83972;
  assign n83974 = pi15 ? n15620 : n14995;
  assign n83975 = pi14 ? n83974 : n14995;
  assign n83976 = pi13 ? n83973 : n83975;
  assign n83977 = pi12 ? n83967 : n83976;
  assign n83978 = pi11 ? n83962 : n83977;
  assign n83979 = pi15 ? n27528 : n24700;
  assign n83980 = pi15 ? n24700 : n15643;
  assign n83981 = pi14 ? n83979 : n83980;
  assign n83982 = pi13 ? n83981 : n15657;
  assign n83983 = pi12 ? n83982 : n15668;
  assign n83984 = pi11 ? n83983 : n32;
  assign n83985 = pi10 ? n83978 : n83984;
  assign n83986 = pi09 ? n83950 : n83985;
  assign n83987 = pi08 ? n83936 : n83986;
  assign n83988 = pi20 ? n1475 : ~n428;
  assign n83989 = pi19 ? n32 : n83988;
  assign n83990 = pi18 ? n32 : n83989;
  assign n83991 = pi17 ? n32 : n83990;
  assign n83992 = pi16 ? n32 : n83991;
  assign n83993 = pi15 ? n32 : n83992;
  assign n83994 = pi14 ? n83993 : n83945;
  assign n83995 = pi13 ? n32 : n83994;
  assign n83996 = pi12 ? n32 : n83995;
  assign n83997 = pi11 ? n32 : n83996;
  assign n83998 = pi10 ? n32 : n83997;
  assign n83999 = pi20 ? n1940 : ~n101;
  assign n84000 = pi19 ? n32 : n83999;
  assign n84001 = pi18 ? n32 : n84000;
  assign n84002 = pi17 ? n32 : n84001;
  assign n84003 = pi16 ? n32 : n84002;
  assign n84004 = pi15 ? n83945 : n84003;
  assign n84005 = pi14 ? n84004 : n84003;
  assign n84006 = pi14 ? n83906 : n83912;
  assign n84007 = pi13 ? n84005 : n84006;
  assign n84008 = pi13 ? n83815 : n83960;
  assign n84009 = pi12 ? n84007 : n84008;
  assign n84010 = pi20 ? n141 : ~n342;
  assign n84011 = pi19 ? n32 : n84010;
  assign n84012 = pi18 ? n32 : n84011;
  assign n84013 = pi17 ? n32 : n84012;
  assign n84014 = pi16 ? n32 : n84013;
  assign n84015 = pi20 ? n141 : ~n518;
  assign n84016 = pi19 ? n32 : n84015;
  assign n84017 = pi18 ? n32 : n84016;
  assign n84018 = pi17 ? n32 : n84017;
  assign n84019 = pi16 ? n32 : n84018;
  assign n84020 = pi15 ? n84014 : n84019;
  assign n84021 = pi14 ? n84020 : n84019;
  assign n84022 = pi15 ? n15755 : n73452;
  assign n84023 = pi14 ? n84022 : n73452;
  assign n84024 = pi13 ? n84021 : n84023;
  assign n84025 = pi20 ? n141 : ~n243;
  assign n84026 = pi19 ? n32 : n84025;
  assign n84027 = pi18 ? n32 : n84026;
  assign n84028 = pi17 ? n32 : n84027;
  assign n84029 = pi16 ? n32 : n84028;
  assign n84030 = pi15 ? n15779 : n84029;
  assign n84031 = pi14 ? n15780 : n84030;
  assign n84032 = pi20 ? n141 : ~n339;
  assign n84033 = pi19 ? n32 : n84032;
  assign n84034 = pi18 ? n32 : n84033;
  assign n84035 = pi17 ? n32 : n84034;
  assign n84036 = pi16 ? n32 : n84035;
  assign n84037 = pi15 ? n84036 : n15150;
  assign n84038 = pi14 ? n84037 : n15150;
  assign n84039 = pi13 ? n84031 : n84038;
  assign n84040 = pi12 ? n84024 : n84039;
  assign n84041 = pi11 ? n84009 : n84040;
  assign n84042 = pi15 ? n15810 : n15643;
  assign n84043 = pi14 ? n84042 : n15643;
  assign n84044 = pi13 ? n84043 : n15838;
  assign n84045 = pi12 ? n84044 : n32;
  assign n84046 = pi11 ? n84045 : n32;
  assign n84047 = pi10 ? n84041 : n84046;
  assign n84048 = pi09 ? n83998 : n84047;
  assign n84049 = pi18 ? n32 : n61714;
  assign n84050 = pi17 ? n32 : n84049;
  assign n84051 = pi16 ? n32 : n84050;
  assign n84052 = pi15 ? n32 : n84051;
  assign n84053 = pi19 ? n32 : n35513;
  assign n84054 = pi18 ? n32 : n84053;
  assign n84055 = pi17 ? n32 : n84054;
  assign n84056 = pi16 ? n32 : n84055;
  assign n84057 = pi14 ? n84052 : n84056;
  assign n84058 = pi13 ? n32 : n84057;
  assign n84059 = pi12 ? n32 : n84058;
  assign n84060 = pi11 ? n32 : n84059;
  assign n84061 = pi10 ? n32 : n84060;
  assign n84062 = pi15 ? n84056 : n84003;
  assign n84063 = pi15 ? n84003 : n83900;
  assign n84064 = pi14 ? n84062 : n84063;
  assign n84065 = pi15 ? n83900 : n84003;
  assign n84066 = pi14 ? n84065 : n84003;
  assign n84067 = pi13 ? n84064 : n84066;
  assign n84068 = pi19 ? n32 : n22751;
  assign n84069 = pi18 ? n32 : n84068;
  assign n84070 = pi17 ? n32 : n84069;
  assign n84071 = pi16 ? n32 : n84070;
  assign n84072 = pi20 ? n243 : ~n2140;
  assign n84073 = pi19 ? n32 : n84072;
  assign n84074 = pi18 ? n32 : n84073;
  assign n84075 = pi17 ? n32 : n84074;
  assign n84076 = pi16 ? n32 : n84075;
  assign n84077 = pi15 ? n84071 : n84076;
  assign n84078 = pi19 ? n32 : n61029;
  assign n84079 = pi18 ? n32 : n84078;
  assign n84080 = pi17 ? n32 : n84079;
  assign n84081 = pi16 ? n32 : n84080;
  assign n84082 = pi15 ? n84076 : n84081;
  assign n84083 = pi14 ? n84077 : n84082;
  assign n84084 = pi13 ? n84003 : n84083;
  assign n84085 = pi12 ? n84067 : n84084;
  assign n84086 = pi15 ? n73452 : n15766;
  assign n84087 = pi14 ? n73452 : n84086;
  assign n84088 = pi13 ? n15755 : n84087;
  assign n84089 = pi15 ? n15916 : n73544;
  assign n84090 = pi14 ? n15916 : n84089;
  assign n84091 = pi14 ? n15707 : n16086;
  assign n84092 = pi13 ? n84090 : n84091;
  assign n84093 = pi12 ? n84088 : n84092;
  assign n84094 = pi11 ? n84085 : n84093;
  assign n84095 = pi15 ? n73574 : n15966;
  assign n84096 = pi14 ? n15947 : n84095;
  assign n84097 = pi13 ? n84096 : n15969;
  assign n84098 = pi12 ? n84097 : n32;
  assign n84099 = pi11 ? n84098 : n32;
  assign n84100 = pi10 ? n84094 : n84099;
  assign n84101 = pi09 ? n84061 : n84100;
  assign n84102 = pi08 ? n84048 : n84101;
  assign n84103 = pi07 ? n83987 : n84102;
  assign n84104 = pi20 ? n1839 : ~n428;
  assign n84105 = pi19 ? n32 : n84104;
  assign n84106 = pi18 ? n32 : n84105;
  assign n84107 = pi17 ? n32 : n84106;
  assign n84108 = pi16 ? n32 : n84107;
  assign n84109 = pi15 ? n32 : n84108;
  assign n84110 = pi20 ? n1839 : ~n101;
  assign n84111 = pi19 ? n32 : n84110;
  assign n84112 = pi18 ? n32 : n84111;
  assign n84113 = pi17 ? n32 : n84112;
  assign n84114 = pi16 ? n32 : n84113;
  assign n84115 = pi14 ? n84109 : n84114;
  assign n84116 = pi13 ? n32 : n84115;
  assign n84117 = pi12 ? n32 : n84116;
  assign n84118 = pi11 ? n32 : n84117;
  assign n84119 = pi10 ? n32 : n84118;
  assign n84120 = pi20 ? n1475 : ~n101;
  assign n84121 = pi19 ? n32 : n84120;
  assign n84122 = pi18 ? n32 : n84121;
  assign n84123 = pi17 ? n32 : n84122;
  assign n84124 = pi16 ? n32 : n84123;
  assign n84125 = pi15 ? n84114 : n84124;
  assign n84126 = pi14 ? n84125 : n83945;
  assign n84127 = pi14 ? n83945 : n84003;
  assign n84128 = pi13 ? n84126 : n84127;
  assign n84129 = pi13 ? n84003 : n84071;
  assign n84130 = pi12 ? n84128 : n84129;
  assign n84131 = pi20 ? n1940 : ~n518;
  assign n84132 = pi19 ? n32 : n84131;
  assign n84133 = pi18 ? n32 : n84132;
  assign n84134 = pi17 ? n32 : n84133;
  assign n84135 = pi16 ? n32 : n84134;
  assign n84136 = pi19 ? n32 : n8907;
  assign n84137 = pi18 ? n32 : n84136;
  assign n84138 = pi17 ? n32 : n84137;
  assign n84139 = pi16 ? n32 : n84138;
  assign n84140 = pi15 ? n84139 : n84135;
  assign n84141 = pi14 ? n84135 : n84140;
  assign n84142 = pi19 ? n32 : n23553;
  assign n84143 = pi18 ? n32 : n84142;
  assign n84144 = pi17 ? n32 : n84143;
  assign n84145 = pi16 ? n32 : n84144;
  assign n84146 = pi20 ? n1940 : ~n1475;
  assign n84147 = pi19 ? n32 : n84146;
  assign n84148 = pi18 ? n32 : n84147;
  assign n84149 = pi17 ? n32 : n84148;
  assign n84150 = pi16 ? n32 : n84149;
  assign n84151 = pi15 ? n84145 : n84150;
  assign n84152 = pi19 ? n32 : n13057;
  assign n84153 = pi18 ? n32 : n84152;
  assign n84154 = pi17 ? n32 : n84153;
  assign n84155 = pi16 ? n32 : n84154;
  assign n84156 = pi15 ? n84145 : n84155;
  assign n84157 = pi14 ? n84151 : n84156;
  assign n84158 = pi13 ? n84141 : n84157;
  assign n84159 = pi20 ? n243 : ~n207;
  assign n84160 = pi19 ? n32 : n84159;
  assign n84161 = pi18 ? n32 : n84160;
  assign n84162 = pi17 ? n32 : n84161;
  assign n84163 = pi16 ? n32 : n84162;
  assign n84164 = pi15 ? n84163 : n16070;
  assign n84165 = pi14 ? n84163 : n84164;
  assign n84166 = pi13 ? n84165 : n84091;
  assign n84167 = pi12 ? n84158 : n84166;
  assign n84168 = pi11 ? n84130 : n84167;
  assign n84169 = pi15 ? n15947 : n16101;
  assign n84170 = pi15 ? n16215 : n16105;
  assign n84171 = pi14 ? n84169 : n84170;
  assign n84172 = pi13 ? n84171 : n16111;
  assign n84173 = pi12 ? n84172 : n32;
  assign n84174 = pi11 ? n84173 : n32;
  assign n84175 = pi10 ? n84168 : n84174;
  assign n84176 = pi09 ? n84119 : n84175;
  assign n84177 = pi15 ? n84114 : n84056;
  assign n84178 = pi14 ? n84177 : n84124;
  assign n84179 = pi13 ? n84178 : n84124;
  assign n84180 = pi15 ? n84124 : n83945;
  assign n84181 = pi14 ? n84124 : n84180;
  assign n84182 = pi20 ? n749 : ~n2140;
  assign n84183 = pi19 ? n32 : n84182;
  assign n84184 = pi18 ? n32 : n84183;
  assign n84185 = pi17 ? n32 : n84184;
  assign n84186 = pi16 ? n32 : n84185;
  assign n84187 = pi20 ? n1940 : ~n2140;
  assign n84188 = pi19 ? n32 : n84187;
  assign n84189 = pi18 ? n32 : n84188;
  assign n84190 = pi17 ? n32 : n84189;
  assign n84191 = pi16 ? n32 : n84190;
  assign n84192 = pi15 ? n84186 : n84191;
  assign n84193 = pi14 ? n84186 : n84192;
  assign n84194 = pi13 ? n84181 : n84193;
  assign n84195 = pi12 ? n84179 : n84194;
  assign n84196 = pi20 ? n1940 : ~n1839;
  assign n84197 = pi19 ? n32 : n84196;
  assign n84198 = pi18 ? n32 : n84197;
  assign n84199 = pi17 ? n32 : n84198;
  assign n84200 = pi16 ? n32 : n84199;
  assign n84201 = pi15 ? n84135 : n84200;
  assign n84202 = pi14 ? n84135 : n84201;
  assign n84203 = pi15 ? n84150 : n73628;
  assign n84204 = pi14 ? n84150 : n84203;
  assign n84205 = pi13 ? n84202 : n84204;
  assign n84206 = pi20 ? n16195 : ~n207;
  assign n84207 = pi19 ? n32 : n84206;
  assign n84208 = pi18 ? n32 : n84207;
  assign n84209 = pi17 ? n32 : n84208;
  assign n84210 = pi16 ? n32 : n84209;
  assign n84211 = pi20 ? n1940 : ~n339;
  assign n84212 = pi19 ? n32 : n84211;
  assign n84213 = pi18 ? n32 : n84212;
  assign n84214 = pi17 ? n32 : n84213;
  assign n84215 = pi16 ? n32 : n84214;
  assign n84216 = pi15 ? n84210 : n84215;
  assign n84217 = pi14 ? n16286 : n84216;
  assign n84218 = pi14 ? n15403 : n16205;
  assign n84219 = pi13 ? n84217 : n84218;
  assign n84220 = pi12 ? n84205 : n84219;
  assign n84221 = pi11 ? n84195 : n84220;
  assign n84222 = pi10 ? n84221 : n16222;
  assign n84223 = pi09 ? n84119 : n84222;
  assign n84224 = pi08 ? n84176 : n84223;
  assign n84225 = pi20 ? n518 : ~n428;
  assign n84226 = pi19 ? n32 : n84225;
  assign n84227 = pi18 ? n32 : n84226;
  assign n84228 = pi17 ? n32 : n84227;
  assign n84229 = pi16 ? n32 : n84228;
  assign n84230 = pi15 ? n32 : n84229;
  assign n84231 = pi20 ? n518 : ~n101;
  assign n84232 = pi19 ? n32 : n84231;
  assign n84233 = pi18 ? n32 : n84232;
  assign n84234 = pi17 ? n32 : n84233;
  assign n84235 = pi16 ? n32 : n84234;
  assign n84236 = pi14 ? n84230 : n84235;
  assign n84237 = pi13 ? n32 : n84236;
  assign n84238 = pi12 ? n32 : n84237;
  assign n84239 = pi11 ? n32 : n84238;
  assign n84240 = pi10 ? n32 : n84239;
  assign n84241 = pi15 ? n84056 : n84124;
  assign n84242 = pi14 ? n84177 : n84241;
  assign n84243 = pi14 ? n84124 : n84056;
  assign n84244 = pi13 ? n84242 : n84243;
  assign n84245 = pi14 ? n84056 : n84241;
  assign n84246 = pi15 ? n16246 : n84186;
  assign n84247 = pi14 ? n16246 : n84246;
  assign n84248 = pi13 ? n84245 : n84247;
  assign n84249 = pi12 ? n84244 : n84248;
  assign n84250 = pi20 ? n1475 : ~n518;
  assign n84251 = pi19 ? n32 : n84250;
  assign n84252 = pi18 ? n32 : n84251;
  assign n84253 = pi17 ? n32 : n84252;
  assign n84254 = pi16 ? n32 : n84253;
  assign n84255 = pi20 ? n1475 : ~n1839;
  assign n84256 = pi19 ? n32 : n84255;
  assign n84257 = pi18 ? n32 : n84256;
  assign n84258 = pi17 ? n32 : n84257;
  assign n84259 = pi16 ? n32 : n84258;
  assign n84260 = pi15 ? n84254 : n84259;
  assign n84261 = pi14 ? n84254 : n84260;
  assign n84262 = pi15 ? n73741 : n16278;
  assign n84263 = pi14 ? n73741 : n84262;
  assign n84264 = pi13 ? n84261 : n84263;
  assign n84265 = pi14 ? n16286 : n16287;
  assign n84266 = pi20 ? n26667 : n32;
  assign n84267 = pi19 ? n32 : n84266;
  assign n84268 = pi18 ? n32 : n84267;
  assign n84269 = pi17 ? n32 : n84268;
  assign n84270 = pi16 ? n32 : n84269;
  assign n84271 = pi15 ? n84270 : n16298;
  assign n84272 = pi14 ? n15531 : n84271;
  assign n84273 = pi13 ? n84265 : n84272;
  assign n84274 = pi12 ? n84264 : n84273;
  assign n84275 = pi11 ? n84249 : n84274;
  assign n84276 = pi15 ? n16298 : n16314;
  assign n84277 = pi14 ? n84276 : n27740;
  assign n84278 = pi13 ? n84277 : n16322;
  assign n84279 = pi12 ? n84278 : n32;
  assign n84280 = pi11 ? n84279 : n32;
  assign n84281 = pi10 ? n84275 : n84280;
  assign n84282 = pi09 ? n84240 : n84281;
  assign n84283 = pi15 ? n84235 : n84114;
  assign n84284 = pi14 ? n84283 : n84177;
  assign n84285 = pi13 ? n84284 : n84056;
  assign n84286 = pi13 ? n84056 : n16246;
  assign n84287 = pi12 ? n84285 : n84286;
  assign n84288 = pi15 ? n84254 : n68552;
  assign n84289 = pi15 ? n68552 : n73734;
  assign n84290 = pi14 ? n84288 : n84289;
  assign n84291 = pi14 ? n73774 : n73775;
  assign n84292 = pi13 ? n84290 : n84291;
  assign n84293 = pi14 ? n73782 : n16356;
  assign n84294 = pi15 ? n84270 : n16293;
  assign n84295 = pi14 ? n16232 : n84294;
  assign n84296 = pi13 ? n84293 : n84295;
  assign n84297 = pi12 ? n84292 : n84296;
  assign n84298 = pi11 ? n84287 : n84297;
  assign n84299 = pi10 ? n84298 : n27763;
  assign n84300 = pi09 ? n84240 : n84299;
  assign n84301 = pi08 ? n84282 : n84300;
  assign n84302 = pi07 ? n84224 : n84301;
  assign n84303 = pi06 ? n84103 : n84302;
  assign n84304 = pi05 ? n83891 : n84303;
  assign n84305 = pi20 ? n1319 : ~n428;
  assign n84306 = pi19 ? n32 : n84305;
  assign n84307 = pi18 ? n32 : n84306;
  assign n84308 = pi17 ? n32 : n84307;
  assign n84309 = pi16 ? n32 : n84308;
  assign n84310 = pi15 ? n32 : n84309;
  assign n84311 = pi20 ? n1319 : ~n101;
  assign n84312 = pi19 ? n32 : n84311;
  assign n84313 = pi18 ? n32 : n84312;
  assign n84314 = pi17 ? n32 : n84313;
  assign n84315 = pi16 ? n32 : n84314;
  assign n84316 = pi14 ? n84310 : n84315;
  assign n84317 = pi13 ? n32 : n84316;
  assign n84318 = pi12 ? n32 : n84317;
  assign n84319 = pi11 ? n32 : n84318;
  assign n84320 = pi10 ? n32 : n84319;
  assign n84321 = pi15 ? n72946 : n69136;
  assign n84322 = pi14 ? n72946 : n84321;
  assign n84323 = pi13 ? n84114 : n84322;
  assign n84324 = pi12 ? n84114 : n84323;
  assign n84325 = pi14 ? n68552 : n84289;
  assign n84326 = pi15 ? n67879 : n16352;
  assign n84327 = pi14 ? n67879 : n84326;
  assign n84328 = pi13 ? n84325 : n84327;
  assign n84329 = pi14 ? n16334 : n26447;
  assign n84330 = pi13 ? n16448 : n84329;
  assign n84331 = pi12 ? n84328 : n84330;
  assign n84332 = pi11 ? n84324 : n84331;
  assign n84333 = pi10 ? n84332 : n16461;
  assign n84334 = pi09 ? n84320 : n84333;
  assign n84335 = pi14 ? n84235 : n84283;
  assign n84336 = pi13 ? n84335 : n84114;
  assign n84337 = pi20 ? n1839 : ~n2140;
  assign n84338 = pi19 ? n32 : n84337;
  assign n84339 = pi18 ? n32 : n84338;
  assign n84340 = pi17 ? n32 : n84339;
  assign n84341 = pi16 ? n32 : n84340;
  assign n84342 = pi15 ? n72946 : n16559;
  assign n84343 = pi14 ? n84341 : n84342;
  assign n84344 = pi13 ? n84114 : n84343;
  assign n84345 = pi12 ? n84336 : n84344;
  assign n84346 = pi20 ? n1839 : ~n518;
  assign n84347 = pi19 ? n32 : n84346;
  assign n84348 = pi18 ? n32 : n84347;
  assign n84349 = pi17 ? n32 : n84348;
  assign n84350 = pi16 ? n32 : n84349;
  assign n84351 = pi20 ? n1839 : ~n1839;
  assign n84352 = pi19 ? n32 : n84351;
  assign n84353 = pi18 ? n32 : n84352;
  assign n84354 = pi17 ? n32 : n84353;
  assign n84355 = pi16 ? n32 : n84354;
  assign n84356 = pi15 ? n84350 : n84355;
  assign n84357 = pi14 ? n84350 : n84356;
  assign n84358 = pi15 ? n16582 : n16413;
  assign n84359 = pi14 ? n16582 : n84358;
  assign n84360 = pi13 ? n84357 : n84359;
  assign n84361 = pi14 ? n16413 : n16554;
  assign n84362 = pi14 ? n73888 : n16527;
  assign n84363 = pi13 ? n84361 : n84362;
  assign n84364 = pi12 ? n84360 : n84363;
  assign n84365 = pi11 ? n84345 : n84364;
  assign n84366 = pi10 ? n84365 : n32;
  assign n84367 = pi09 ? n84320 : n84366;
  assign n84368 = pi08 ? n84334 : n84367;
  assign n84369 = pi18 ? n32 : n19001;
  assign n84370 = pi17 ? n32 : n84369;
  assign n84371 = pi16 ? n32 : n84370;
  assign n84372 = pi15 ? n32 : n84371;
  assign n84373 = pi19 ? n32 : n24750;
  assign n84374 = pi18 ? n32 : n84373;
  assign n84375 = pi17 ? n32 : n84374;
  assign n84376 = pi16 ? n32 : n84375;
  assign n84377 = pi14 ? n84372 : n84376;
  assign n84378 = pi13 ? n32 : n84377;
  assign n84379 = pi12 ? n32 : n84378;
  assign n84380 = pi11 ? n32 : n84379;
  assign n84381 = pi10 ? n32 : n84380;
  assign n84382 = pi15 ? n84315 : n84235;
  assign n84383 = pi14 ? n84315 : n84382;
  assign n84384 = pi13 ? n84383 : n84235;
  assign n84385 = pi15 ? n84341 : n16559;
  assign n84386 = pi14 ? n84341 : n84385;
  assign n84387 = pi13 ? n84235 : n84386;
  assign n84388 = pi12 ? n84384 : n84387;
  assign n84389 = pi15 ? n16582 : n16595;
  assign n84390 = pi14 ? n16582 : n84389;
  assign n84391 = pi13 ? n84357 : n84390;
  assign n84392 = pi15 ? n16629 : n16546;
  assign n84393 = pi14 ? n16595 : n84392;
  assign n84394 = pi13 ? n84393 : n16608;
  assign n84395 = pi12 ? n84391 : n84394;
  assign n84396 = pi11 ? n84388 : n84395;
  assign n84397 = pi10 ? n84396 : n32;
  assign n84398 = pi09 ? n84381 : n84397;
  assign n84399 = pi15 ? n84235 : n84315;
  assign n84400 = pi14 ? n84235 : n84399;
  assign n84401 = pi20 ? n518 : ~n2140;
  assign n84402 = pi19 ? n32 : n84401;
  assign n84403 = pi18 ? n32 : n84402;
  assign n84404 = pi17 ? n32 : n84403;
  assign n84405 = pi16 ? n32 : n84404;
  assign n84406 = pi20 ? n518 : ~n342;
  assign n84407 = pi19 ? n32 : n84406;
  assign n84408 = pi18 ? n32 : n84407;
  assign n84409 = pi17 ? n32 : n84408;
  assign n84410 = pi16 ? n32 : n84409;
  assign n84411 = pi15 ? n84405 : n84410;
  assign n84412 = pi14 ? n84405 : n84411;
  assign n84413 = pi13 ? n84400 : n84412;
  assign n84414 = pi12 ? n84384 : n84413;
  assign n84415 = pi20 ? n518 : ~n1839;
  assign n84416 = pi19 ? n32 : n84415;
  assign n84417 = pi18 ? n32 : n84416;
  assign n84418 = pi17 ? n32 : n84417;
  assign n84419 = pi16 ? n32 : n84418;
  assign n84420 = pi15 ? n16634 : n84419;
  assign n84421 = pi14 ? n16634 : n84420;
  assign n84422 = pi15 ? n16645 : n16595;
  assign n84423 = pi14 ? n16645 : n84422;
  assign n84424 = pi13 ? n84421 : n84423;
  assign n84425 = pi13 ? n84393 : n16657;
  assign n84426 = pi12 ? n84424 : n84425;
  assign n84427 = pi11 ? n84414 : n84426;
  assign n84428 = pi10 ? n84427 : n32;
  assign n84429 = pi09 ? n84381 : n84428;
  assign n84430 = pi08 ? n84398 : n84429;
  assign n84431 = pi07 ? n84368 : n84430;
  assign n84432 = pi20 ? n2140 : ~n428;
  assign n84433 = pi19 ? n32 : n84432;
  assign n84434 = pi18 ? n32 : n84433;
  assign n84435 = pi17 ? n32 : n84434;
  assign n84436 = pi16 ? n32 : n84435;
  assign n84437 = pi15 ? n32 : n84436;
  assign n84438 = pi19 ? n32 : n13126;
  assign n84439 = pi18 ? n32 : n84438;
  assign n84440 = pi17 ? n32 : n84439;
  assign n84441 = pi16 ? n32 : n84440;
  assign n84442 = pi14 ? n84437 : n84441;
  assign n84443 = pi13 ? n32 : n84442;
  assign n84444 = pi12 ? n32 : n84443;
  assign n84445 = pi11 ? n32 : n84444;
  assign n84446 = pi10 ? n32 : n84445;
  assign n84447 = pi15 ? n84376 : n84315;
  assign n84448 = pi14 ? n84376 : n84447;
  assign n84449 = pi13 ? n84448 : n84315;
  assign n84450 = pi13 ? n84315 : n84412;
  assign n84451 = pi12 ? n84449 : n84450;
  assign n84452 = pi15 ? n16634 : n16645;
  assign n84453 = pi14 ? n16634 : n84452;
  assign n84454 = pi15 ? n16645 : n16706;
  assign n84455 = pi14 ? n84454 : n16711;
  assign n84456 = pi13 ? n84453 : n84455;
  assign n84457 = pi15 ? n16711 : n16724;
  assign n84458 = pi14 ? n84457 : n16725;
  assign n84459 = pi13 ? n84458 : n16727;
  assign n84460 = pi12 ? n84456 : n84459;
  assign n84461 = pi11 ? n84451 : n84460;
  assign n84462 = pi10 ? n84461 : n32;
  assign n84463 = pi09 ? n84446 : n84462;
  assign n84464 = pi20 ? n428 : ~n428;
  assign n84465 = pi19 ? n32 : n84464;
  assign n84466 = pi18 ? n32 : n84465;
  assign n84467 = pi17 ? n32 : n84466;
  assign n84468 = pi16 ? n32 : n84467;
  assign n84469 = pi15 ? n32 : n84468;
  assign n84470 = pi20 ? n428 : ~n101;
  assign n84471 = pi19 ? n32 : n84470;
  assign n84472 = pi18 ? n32 : n84471;
  assign n84473 = pi17 ? n32 : n84472;
  assign n84474 = pi16 ? n32 : n84473;
  assign n84475 = pi15 ? n84474 : n84441;
  assign n84476 = pi14 ? n84469 : n84475;
  assign n84477 = pi13 ? n32 : n84476;
  assign n84478 = pi12 ? n32 : n84477;
  assign n84479 = pi11 ? n32 : n84478;
  assign n84480 = pi10 ? n32 : n84479;
  assign n84481 = pi14 ? n84315 : n84376;
  assign n84482 = pi20 ? n1319 : ~n342;
  assign n84483 = pi19 ? n32 : n84482;
  assign n84484 = pi18 ? n32 : n84483;
  assign n84485 = pi17 ? n32 : n84484;
  assign n84486 = pi16 ? n32 : n84485;
  assign n84487 = pi15 ? n16812 : n84486;
  assign n84488 = pi14 ? n16812 : n84487;
  assign n84489 = pi13 ? n84481 : n84488;
  assign n84490 = pi12 ? n84449 : n84489;
  assign n84491 = pi20 ? n1319 : ~n518;
  assign n84492 = pi19 ? n32 : n84491;
  assign n84493 = pi18 ? n32 : n84492;
  assign n84494 = pi17 ? n32 : n84493;
  assign n84495 = pi16 ? n32 : n84494;
  assign n84496 = pi15 ? n84495 : n16706;
  assign n84497 = pi14 ? n84495 : n84496;
  assign n84498 = pi14 ? n16706 : n16711;
  assign n84499 = pi13 ? n84497 : n84498;
  assign n84500 = pi13 ? n84458 : n16787;
  assign n84501 = pi12 ? n84499 : n84500;
  assign n84502 = pi11 ? n84490 : n84501;
  assign n84503 = pi10 ? n84502 : n32;
  assign n84504 = pi09 ? n84480 : n84503;
  assign n84505 = pi08 ? n84463 : n84504;
  assign n84506 = pi14 ? n84469 : n84474;
  assign n84507 = pi13 ? n32 : n84506;
  assign n84508 = pi12 ? n32 : n84507;
  assign n84509 = pi11 ? n32 : n84508;
  assign n84510 = pi10 ? n32 : n84509;
  assign n84511 = pi15 ? n84441 : n84376;
  assign n84512 = pi14 ? n84441 : n84511;
  assign n84513 = pi13 ? n84512 : n84376;
  assign n84514 = pi13 ? n84376 : n84488;
  assign n84515 = pi12 ? n84513 : n84514;
  assign n84516 = pi14 ? n16824 : n16804;
  assign n84517 = pi13 ? n84497 : n84516;
  assign n84518 = pi12 ? n84517 : n16842;
  assign n84519 = pi11 ? n84515 : n84518;
  assign n84520 = pi10 ? n84519 : n32;
  assign n84521 = pi09 ? n84510 : n84520;
  assign n84522 = pi20 ? n101 : ~n428;
  assign n84523 = pi19 ? n32 : n84522;
  assign n84524 = pi18 ? n32 : n84523;
  assign n84525 = pi17 ? n32 : n84524;
  assign n84526 = pi16 ? n32 : n84525;
  assign n84527 = pi15 ? n32 : n84526;
  assign n84528 = pi20 ? n101 : ~n101;
  assign n84529 = pi19 ? n32 : n84528;
  assign n84530 = pi18 ? n32 : n84529;
  assign n84531 = pi17 ? n32 : n84530;
  assign n84532 = pi16 ? n32 : n84531;
  assign n84533 = pi15 ? n84532 : n84474;
  assign n84534 = pi14 ? n84527 : n84533;
  assign n84535 = pi13 ? n32 : n84534;
  assign n84536 = pi12 ? n32 : n84535;
  assign n84537 = pi11 ? n32 : n84536;
  assign n84538 = pi10 ? n32 : n84537;
  assign n84539 = pi14 ? n84511 : n84441;
  assign n84540 = pi13 ? n84512 : n84539;
  assign n84541 = pi15 ? n16869 : n53963;
  assign n84542 = pi14 ? n16869 : n84541;
  assign n84543 = pi13 ? n84441 : n84542;
  assign n84544 = pi12 ? n84540 : n84543;
  assign n84545 = pi14 ? n53963 : n16824;
  assign n84546 = pi15 ? n16824 : n16804;
  assign n84547 = pi14 ? n84546 : n16804;
  assign n84548 = pi13 ? n84545 : n84547;
  assign n84549 = pi12 ? n84548 : n16902;
  assign n84550 = pi11 ? n84544 : n84549;
  assign n84551 = pi10 ? n84550 : n32;
  assign n84552 = pi09 ? n84538 : n84551;
  assign n84553 = pi08 ? n84521 : n84552;
  assign n84554 = pi07 ? n84505 : n84553;
  assign n84555 = pi06 ? n84431 : n84554;
  assign n84556 = pi14 ? n84527 : n84532;
  assign n84557 = pi13 ? n32 : n84556;
  assign n84558 = pi12 ? n32 : n84557;
  assign n84559 = pi11 ? n32 : n84558;
  assign n84560 = pi10 ? n32 : n84559;
  assign n84561 = pi14 ? n84474 : n84475;
  assign n84562 = pi13 ? n84561 : n84441;
  assign n84563 = pi12 ? n84562 : n84543;
  assign n84564 = pi20 ? n2140 : ~n518;
  assign n84565 = pi19 ? n32 : n84564;
  assign n84566 = pi18 ? n32 : n84565;
  assign n84567 = pi17 ? n32 : n84566;
  assign n84568 = pi16 ? n32 : n84567;
  assign n84569 = pi14 ? n84568 : n16959;
  assign n84570 = pi15 ? n16959 : n16862;
  assign n84571 = pi14 ? n84570 : n16862;
  assign n84572 = pi13 ? n84569 : n84571;
  assign n84573 = pi12 ? n84572 : n16976;
  assign n84574 = pi11 ? n84563 : n84573;
  assign n84575 = pi10 ? n84574 : n32;
  assign n84576 = pi09 ? n84560 : n84575;
  assign n84577 = pi18 ? n32 : n17919;
  assign n84578 = pi17 ? n32 : n84577;
  assign n84579 = pi16 ? n32 : n84578;
  assign n84580 = pi15 ? n32 : n84579;
  assign n84581 = pi14 ? n84580 : n84532;
  assign n84582 = pi13 ? n32 : n84581;
  assign n84583 = pi12 ? n32 : n84582;
  assign n84584 = pi11 ? n32 : n84583;
  assign n84585 = pi10 ? n32 : n84584;
  assign n84586 = pi20 ? n2140 : ~n2140;
  assign n84587 = pi19 ? n32 : n84586;
  assign n84588 = pi18 ? n32 : n84587;
  assign n84589 = pi17 ? n32 : n84588;
  assign n84590 = pi16 ? n32 : n84589;
  assign n84591 = pi15 ? n84590 : n84568;
  assign n84592 = pi14 ? n84590 : n84591;
  assign n84593 = pi13 ? n84474 : n84592;
  assign n84594 = pi12 ? n84474 : n84593;
  assign n84595 = pi14 ? n84570 : n17014;
  assign n84596 = pi13 ? n84569 : n84595;
  assign n84597 = pi12 ? n84596 : n17019;
  assign n84598 = pi11 ? n84594 : n84597;
  assign n84599 = pi10 ? n84598 : n32;
  assign n84600 = pi09 ? n84585 : n84599;
  assign n84601 = pi08 ? n84576 : n84600;
  assign n84602 = pi18 ? n32 : n18023;
  assign n84603 = pi17 ? n32 : n84602;
  assign n84604 = pi16 ? n32 : n84603;
  assign n84605 = pi14 ? n84580 : n84604;
  assign n84606 = pi13 ? n32 : n84605;
  assign n84607 = pi12 ? n32 : n84606;
  assign n84608 = pi11 ? n32 : n84607;
  assign n84609 = pi10 ? n32 : n84608;
  assign n84610 = pi14 ? n84533 : n84474;
  assign n84611 = pi13 ? n84532 : n84610;
  assign n84612 = pi20 ? n428 : ~n2140;
  assign n84613 = pi19 ? n32 : n84612;
  assign n84614 = pi18 ? n32 : n84613;
  assign n84615 = pi17 ? n32 : n84614;
  assign n84616 = pi16 ? n32 : n84615;
  assign n84617 = pi15 ? n84616 : n53119;
  assign n84618 = pi14 ? n84616 : n84617;
  assign n84619 = pi13 ? n84474 : n84618;
  assign n84620 = pi12 ? n84611 : n84619;
  assign n84621 = pi15 ? n17056 : n16959;
  assign n84622 = pi14 ? n53119 : n84621;
  assign n84623 = pi14 ? n74153 : n17067;
  assign n84624 = pi13 ? n84622 : n84623;
  assign n84625 = pi12 ? n84624 : n17072;
  assign n84626 = pi11 ? n84620 : n84625;
  assign n84627 = pi10 ? n84626 : n32;
  assign n84628 = pi09 ? n84609 : n84627;
  assign n84629 = pi16 ? n32 : n66825;
  assign n84630 = pi15 ? n32 : n84629;
  assign n84631 = pi14 ? n84630 : n84604;
  assign n84632 = pi13 ? n32 : n84631;
  assign n84633 = pi12 ? n32 : n84632;
  assign n84634 = pi11 ? n32 : n84633;
  assign n84635 = pi10 ? n32 : n84634;
  assign n84636 = pi14 ? n84532 : n84604;
  assign n84637 = pi15 ? n84604 : n84532;
  assign n84638 = pi14 ? n84637 : n84533;
  assign n84639 = pi13 ? n84636 : n84638;
  assign n84640 = pi15 ? n74140 : n53119;
  assign n84641 = pi14 ? n74140 : n84640;
  assign n84642 = pi13 ? n84532 : n84641;
  assign n84643 = pi12 ? n84639 : n84642;
  assign n84644 = pi14 ? n53119 : n17056;
  assign n84645 = pi13 ? n84644 : n74169;
  assign n84646 = pi12 ? n84645 : n17102;
  assign n84647 = pi11 ? n84643 : n84646;
  assign n84648 = pi10 ? n84647 : n32;
  assign n84649 = pi09 ? n84635 : n84648;
  assign n84650 = pi08 ? n84628 : n84649;
  assign n84651 = pi07 ? n84601 : n84650;
  assign n84652 = pi21 ? n140 : ~n100;
  assign n84653 = pi20 ? n32 : n84652;
  assign n84654 = pi19 ? n32 : n84653;
  assign n84655 = pi18 ? n32 : n84654;
  assign n84656 = pi17 ? n32 : n84655;
  assign n84657 = pi16 ? n32 : n84656;
  assign n84658 = pi14 ? n84630 : n84657;
  assign n84659 = pi13 ? n32 : n84658;
  assign n84660 = pi12 ? n32 : n84659;
  assign n84661 = pi11 ? n32 : n84660;
  assign n84662 = pi10 ? n32 : n84661;
  assign n84663 = pi14 ? n84604 : n84532;
  assign n84664 = pi13 ? n84604 : n84663;
  assign n84665 = pi15 ? n17193 : n17251;
  assign n84666 = pi14 ? n74140 : n84665;
  assign n84667 = pi13 ? n84532 : n84666;
  assign n84668 = pi12 ? n84664 : n84667;
  assign n84669 = pi15 ? n17251 : n53119;
  assign n84670 = pi14 ? n84669 : n17056;
  assign n84671 = pi14 ? n74185 : n26121;
  assign n84672 = pi13 ? n84670 : n84671;
  assign n84673 = pi12 ? n84672 : n32;
  assign n84674 = pi11 ? n84668 : n84673;
  assign n84675 = pi10 ? n84674 : n32;
  assign n84676 = pi09 ? n84662 : n84675;
  assign n84677 = pi15 ? n84604 : n84657;
  assign n84678 = pi14 ? n84604 : n84677;
  assign n84679 = pi14 ? n84677 : n84532;
  assign n84680 = pi13 ? n84678 : n84679;
  assign n84681 = pi15 ? n84532 : n84604;
  assign n84682 = pi14 ? n84681 : n84604;
  assign n84683 = pi15 ? n17193 : n17286;
  assign n84684 = pi14 ? n17193 : n84683;
  assign n84685 = pi13 ? n84682 : n84684;
  assign n84686 = pi12 ? n84680 : n84685;
  assign n84687 = pi13 ? n17256 : n74186;
  assign n84688 = pi12 ? n84687 : n32;
  assign n84689 = pi11 ? n84686 : n84688;
  assign n84690 = pi10 ? n84689 : n32;
  assign n84691 = pi09 ? n84662 : n84690;
  assign n84692 = pi08 ? n84676 : n84691;
  assign n84693 = pi14 ? n17608 : n84657;
  assign n84694 = pi13 ? n32 : n84693;
  assign n84695 = pi12 ? n32 : n84694;
  assign n84696 = pi11 ? n32 : n84695;
  assign n84697 = pi10 ? n32 : n84696;
  assign n84698 = pi14 ? n84657 : n84604;
  assign n84699 = pi13 ? n84657 : n84698;
  assign n84700 = pi15 ? n17193 : n17205;
  assign n84701 = pi14 ? n17193 : n84700;
  assign n84702 = pi13 ? n84604 : n84701;
  assign n84703 = pi12 ? n84699 : n84702;
  assign n84704 = pi11 ? n84703 : n17265;
  assign n84705 = pi10 ? n84704 : n32;
  assign n84706 = pi09 ? n84697 : n84705;
  assign n84707 = pi15 ? n84657 : n84604;
  assign n84708 = pi14 ? n84657 : n84707;
  assign n84709 = pi13 ? n84657 : n84708;
  assign n84710 = pi14 ? n84707 : n84604;
  assign n84711 = pi15 ? n17278 : n17193;
  assign n84712 = pi14 ? n84711 : n17494;
  assign n84713 = pi13 ? n84710 : n84712;
  assign n84714 = pi12 ? n84709 : n84713;
  assign n84715 = pi15 ? n17255 : n17261;
  assign n84716 = pi14 ? n39553 : n84715;
  assign n84717 = pi13 ? n84716 : n17301;
  assign n84718 = pi12 ? n84717 : n32;
  assign n84719 = pi11 ? n84714 : n84718;
  assign n84720 = pi10 ? n84719 : n32;
  assign n84721 = pi09 ? n84697 : n84720;
  assign n84722 = pi08 ? n84706 : n84721;
  assign n84723 = pi07 ? n84692 : n84722;
  assign n84724 = pi06 ? n84651 : n84723;
  assign n84725 = pi05 ? n84555 : n84724;
  assign n84726 = pi04 ? n84304 : n84725;
  assign n84727 = pi03 ? n83298 : n84726;
  assign n84728 = pi13 ? n84708 : n27844;
  assign n84729 = pi12 ? n84657 : n84728;
  assign n84730 = pi15 ? n17205 : n16850;
  assign n84731 = pi14 ? n84730 : n74233;
  assign n84732 = pi13 ? n84731 : n17301;
  assign n84733 = pi12 ? n84732 : n32;
  assign n84734 = pi11 ? n84729 : n84733;
  assign n84735 = pi10 ? n84734 : n32;
  assign n84736 = pi09 ? n84697 : n84735;
  assign n84737 = pi13 ? n84657 : n27844;
  assign n84738 = pi12 ? n84657 : n84737;
  assign n84739 = pi11 ? n84738 : n74236;
  assign n84740 = pi10 ? n84739 : n32;
  assign n84741 = pi09 ? n84697 : n84740;
  assign n84742 = pi08 ? n84736 : n84741;
  assign n84743 = pi13 ? n84657 : n27929;
  assign n84744 = pi12 ? n84657 : n84743;
  assign n84745 = pi13 ? n27948 : n27935;
  assign n84746 = pi12 ? n84745 : n32;
  assign n84747 = pi11 ? n84744 : n84746;
  assign n84748 = pi10 ? n84747 : n32;
  assign n84749 = pi09 ? n84697 : n84748;
  assign n84750 = pi07 ? n84742 : n84749;
  assign n84751 = pi11 ? n84744 : n27950;
  assign n84752 = pi10 ? n84751 : n32;
  assign n84753 = pi09 ? n84697 : n84752;
  assign n84754 = pi08 ? n84749 : n84753;
  assign n84755 = pi11 ? n84744 : n27943;
  assign n84756 = pi10 ? n84755 : n32;
  assign n84757 = pi09 ? n84697 : n84756;
  assign n84758 = pi08 ? n84753 : n84757;
  assign n84759 = pi07 ? n84754 : n84758;
  assign n84760 = pi06 ? n84750 : n84759;
  assign n84761 = pi11 ? n84744 : n17458;
  assign n84762 = pi10 ? n84761 : n32;
  assign n84763 = pi09 ? n84697 : n84762;
  assign n84764 = pi11 ? n84744 : n17473;
  assign n84765 = pi10 ? n84764 : n32;
  assign n84766 = pi09 ? n84697 : n84765;
  assign n84767 = pi11 ? n84744 : n17480;
  assign n84768 = pi10 ? n84767 : n32;
  assign n84769 = pi09 ? n84697 : n84768;
  assign n84770 = pi08 ? n84766 : n84769;
  assign n84771 = pi07 ? n84763 : n84770;
  assign n84772 = pi15 ? n84657 : n17278;
  assign n84773 = pi14 ? n84772 : n17494;
  assign n84774 = pi13 ? n84657 : n84773;
  assign n84775 = pi12 ? n84657 : n84774;
  assign n84776 = pi11 ? n84775 : n17480;
  assign n84777 = pi10 ? n84776 : n32;
  assign n84778 = pi09 ? n84697 : n84777;
  assign n84779 = pi11 ? n84775 : n17504;
  assign n84780 = pi10 ? n84779 : n32;
  assign n84781 = pi09 ? n84697 : n84780;
  assign n84782 = pi08 ? n84778 : n84781;
  assign n84783 = pi14 ? n84772 : n27978;
  assign n84784 = pi13 ? n84657 : n84783;
  assign n84785 = pi12 ? n84657 : n84784;
  assign n84786 = pi11 ? n84785 : n17521;
  assign n84787 = pi10 ? n84786 : n32;
  assign n84788 = pi09 ? n84697 : n84787;
  assign n84789 = pi07 ? n84782 : n84788;
  assign n84790 = pi06 ? n84771 : n84789;
  assign n84791 = pi05 ? n84760 : n84790;
  assign n84792 = pi14 ? n84772 : n27988;
  assign n84793 = pi13 ? n84657 : n84792;
  assign n84794 = pi12 ? n84657 : n84793;
  assign n84795 = pi11 ? n84794 : n32;
  assign n84796 = pi10 ? n84795 : n32;
  assign n84797 = pi09 ? n84697 : n84796;
  assign n84798 = pi14 ? n84772 : n17357;
  assign n84799 = pi13 ? n84657 : n84798;
  assign n84800 = pi12 ? n84657 : n84799;
  assign n84801 = pi11 ? n84800 : n32;
  assign n84802 = pi10 ? n84801 : n32;
  assign n84803 = pi09 ? n84697 : n84802;
  assign n84804 = pi08 ? n84797 : n84803;
  assign n84805 = pi07 ? n84797 : n84804;
  assign n84806 = pi14 ? n84772 : n32;
  assign n84807 = pi13 ? n84657 : n84806;
  assign n84808 = pi12 ? n84657 : n84807;
  assign n84809 = pi11 ? n84808 : n32;
  assign n84810 = pi10 ? n84809 : n32;
  assign n84811 = pi09 ? n84697 : n84810;
  assign n84812 = pi07 ? n84803 : n84811;
  assign n84813 = pi06 ? n84805 : n84812;
  assign n84814 = pi15 ? n84657 : n32;
  assign n84815 = pi14 ? n84814 : n32;
  assign n84816 = pi13 ? n84657 : n84815;
  assign n84817 = pi12 ? n84657 : n84816;
  assign n84818 = pi11 ? n84817 : n32;
  assign n84819 = pi10 ? n84818 : n32;
  assign n84820 = pi09 ? n84697 : n84819;
  assign n84821 = pi08 ? n84811 : n84820;
  assign n84822 = pi07 ? n84821 : n84820;
  assign n84823 = pi06 ? n84822 : n84820;
  assign n84824 = pi05 ? n84813 : n84823;
  assign n84825 = pi04 ? n84791 : n84824;
  assign n84826 = pi03 ? n84825 : n84820;
  assign n84827 = pi02 ? n84727 : n84826;
  assign n84828 = pi14 ? n84657 : n32;
  assign n84829 = pi13 ? n84657 : n84828;
  assign n84830 = pi12 ? n84657 : n84829;
  assign n84831 = pi11 ? n84830 : n32;
  assign n84832 = pi10 ? n84831 : n32;
  assign n84833 = pi09 ? n84697 : n84832;
  assign n84834 = pi07 ? n84820 : n84833;
  assign n84835 = pi06 ? n84834 : n84833;
  assign n84836 = pi05 ? n84820 : n84835;
  assign n84837 = pi04 ? n84836 : n84833;
  assign n84838 = pi14 ? n17619 : n84657;
  assign n84839 = pi13 ? n32 : n84838;
  assign n84840 = pi12 ? n32 : n84839;
  assign n84841 = pi11 ? n32 : n84840;
  assign n84842 = pi10 ? n32 : n84841;
  assign n84843 = pi09 ? n84842 : n84832;
  assign n84844 = pi08 ? n84833 : n84843;
  assign n84845 = pi14 ? n32 : n84657;
  assign n84846 = pi13 ? n32 : n84845;
  assign n84847 = pi12 ? n32 : n84846;
  assign n84848 = pi11 ? n32 : n84847;
  assign n84849 = pi10 ? n32 : n84848;
  assign n84850 = pi09 ? n84849 : n84832;
  assign n84851 = pi08 ? n84850 : n32;
  assign n84852 = pi07 ? n84844 : n84851;
  assign n84853 = pi06 ? n84833 : n84852;
  assign n84854 = pi05 ? n84853 : n32;
  assign n84855 = pi04 ? n84833 : n84854;
  assign n84856 = pi03 ? n84837 : n84855;
  assign n84857 = pi02 ? n84856 : n32;
  assign n84858 = pi01 ? n84827 : n84857;
  assign n84859 = pi00 ? n79456 : n84858;
  assign po0 = ~n17634;
  assign po1 = ~n28012;
  assign po2 = ~n40904;
  assign po3 = ~n56011;
  assign po4 = ~n74331;
  assign po5 = ~n84859;
endmodule


