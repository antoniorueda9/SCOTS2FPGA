// Benchmark "DD" written by ABC on Wed Jun 26 12:38:34 2019

module DD ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    po0  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23;
  output po0;
  wire n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
    n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
    n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
    n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
    n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
    n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
    n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
    n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
    n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
    n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
    n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
    n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
    n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361;
  assign n26 = 1'b1;
  assign n27 = pi23 ? n26 : ~n26;
  assign n28 = pi22 ? n27 : n26;
  assign n29 = pi21 ? n28 : n26;
  assign n30 = pi20 ? n26 : n29;
  assign n31 = pi19 ? n26 : n30;
  assign n32 = pi18 ? n26 : n31;
  assign n33 = pi17 ? n26 : n32;
  assign n34 = pi16 ? n33 : n32;
  assign n35 = pi15 ? n34 : n32;
  assign n36 = pi14 ? n26 : n35;
  assign n37 = pi22 ? n26 : n27;
  assign n38 = pi21 ? n26 : n37;
  assign n39 = pi20 ? n26 : n38;
  assign n40 = pi19 ? n39 : n26;
  assign n41 = pi18 ? n40 : n26;
  assign n42 = pi17 ? n26 : n41;
  assign n43 = pi16 ? n26 : n42;
  assign n44 = pi21 ? n26 : n28;
  assign n45 = pi20 ? n26 : n44;
  assign n46 = pi19 ? n45 : n26;
  assign n47 = pi18 ? n46 : n26;
  assign n48 = pi16 ? n41 : n47;
  assign n49 = pi15 ? n43 : n48;
  assign n50 = pi21 ? n37 : n26;
  assign n51 = pi20 ? n26 : n50;
  assign n52 = pi19 ? n51 : n26;
  assign n53 = pi18 ? n52 : n26;
  assign n54 = pi22 ? n26 : ~n27;
  assign n55 = pi21 ? n54 : n26;
  assign n56 = pi20 ? n26 : n55;
  assign n57 = pi19 ? n56 : n26;
  assign n58 = pi18 ? n57 : n26;
  assign n59 = pi19 ? n30 : n26;
  assign n60 = pi18 ? n59 : n26;
  assign n61 = pi17 ? n58 : n60;
  assign n62 = pi16 ? n53 : n61;
  assign n63 = pi20 ? n29 : n26;
  assign n64 = pi19 ? n26 : n63;
  assign n65 = pi18 ? n64 : n26;
  assign n66 = pi16 ? n60 : n65;
  assign n67 = pi15 ? n62 : n66;
  assign n68 = pi14 ? n49 : n67;
  assign n69 = pi13 ? n36 : n68;
  assign n70 = pi12 ? n26 : n69;
  assign n71 = pi11 ? n26 : n70;
  assign n72 = pi17 ? n32 : n41;
  assign n73 = pi16 ? n32 : n72;
  assign n74 = pi15 ? n73 : n48;
  assign n75 = pi14 ? n74 : n67;
  assign n76 = pi13 ? n36 : n75;
  assign n77 = pi12 ? n26 : n76;
  assign n78 = pi10 ? n71 : n77;
  assign n79 = pi09 ? n26 : n78;
  assign n80 = pi08 ? n26 : n79;
  assign n81 = pi16 ? n26 : n32;
  assign n82 = pi15 ? n81 : n32;
  assign n83 = pi14 ? n26 : n82;
  assign n84 = pi13 ? n83 : n75;
  assign n85 = pi12 ? n26 : n84;
  assign n86 = pi11 ? n77 : n85;
  assign n87 = pi16 ? n26 : n33;
  assign n88 = pi15 ? n87 : n32;
  assign n89 = pi14 ? n26 : n88;
  assign n90 = pi13 ? n89 : n75;
  assign n91 = pi12 ? n26 : n90;
  assign n92 = pi11 ? n85 : n91;
  assign n93 = pi10 ? n86 : n92;
  assign n94 = pi20 ? n38 : n26;
  assign n95 = pi19 ? n26 : n94;
  assign n96 = pi18 ? n95 : n26;
  assign n97 = pi17 ? n32 : n96;
  assign n98 = pi16 ? n32 : n97;
  assign n99 = pi15 ? n98 : n48;
  assign n100 = pi16 ? n53 : n58;
  assign n101 = pi15 ? n100 : n66;
  assign n102 = pi14 ? n99 : n101;
  assign n103 = pi13 ? n89 : n102;
  assign n104 = pi12 ? n26 : n103;
  assign n105 = pi15 ? n26 : n32;
  assign n106 = pi14 ? n26 : n105;
  assign n107 = pi18 ? n26 : n64;
  assign n108 = pi16 ? n32 : n107;
  assign n109 = pi15 ? n108 : n48;
  assign n110 = pi14 ? n109 : n101;
  assign n111 = pi13 ? n106 : n110;
  assign n112 = pi12 ? n26 : n111;
  assign n113 = pi11 ? n104 : n112;
  assign n114 = pi16 ? n107 : n32;
  assign n115 = pi15 ? n26 : n114;
  assign n116 = pi14 ? n26 : n115;
  assign n117 = pi15 ? n32 : n96;
  assign n118 = pi21 ? n26 : n54;
  assign n119 = pi20 ? n26 : n118;
  assign n120 = pi19 ? n119 : n26;
  assign n121 = pi18 ? n120 : n26;
  assign n122 = pi16 ? n41 : n121;
  assign n123 = pi16 ? n53 : n60;
  assign n124 = pi15 ? n122 : n123;
  assign n125 = pi14 ? n117 : n124;
  assign n126 = pi13 ? n116 : n125;
  assign n127 = pi12 ? n26 : n126;
  assign n128 = pi17 ? n26 : n107;
  assign n129 = pi16 ? n128 : n32;
  assign n130 = pi15 ? n26 : n129;
  assign n131 = pi14 ? n26 : n130;
  assign n132 = pi17 ? n96 : n41;
  assign n133 = pi16 ? n96 : n132;
  assign n134 = pi15 ? n32 : n133;
  assign n135 = pi17 ? n53 : n60;
  assign n136 = pi16 ? n53 : n135;
  assign n137 = pi15 ? n122 : n136;
  assign n138 = pi14 ? n134 : n137;
  assign n139 = pi13 ? n131 : n138;
  assign n140 = pi12 ? n26 : n139;
  assign n141 = pi11 ? n127 : n140;
  assign n142 = pi10 ? n113 : n141;
  assign n143 = pi09 ? n93 : n142;
  assign n144 = pi15 ? n26 : n81;
  assign n145 = pi14 ? n26 : n144;
  assign n146 = pi17 ? n121 : n41;
  assign n147 = pi16 ? n41 : n146;
  assign n148 = pi17 ? n41 : n121;
  assign n149 = pi16 ? n148 : n26;
  assign n150 = pi15 ? n147 : n149;
  assign n151 = pi14 ? n32 : n150;
  assign n152 = pi13 ? n145 : n151;
  assign n153 = pi12 ? n26 : n152;
  assign n154 = pi19 ? n26 : n119;
  assign n155 = pi18 ? n26 : n154;
  assign n156 = pi17 ? n155 : n32;
  assign n157 = pi16 ? n156 : n32;
  assign n158 = pi15 ? n157 : n32;
  assign n159 = pi14 ? n158 : n26;
  assign n160 = pi13 ? n26 : n159;
  assign n161 = pi12 ? n26 : n160;
  assign n162 = pi11 ? n153 : n161;
  assign n163 = pi10 ? n162 : n26;
  assign n164 = pi13 ? n83 : n68;
  assign n165 = pi12 ? n26 : n164;
  assign n166 = pi11 ? n26 : n165;
  assign n167 = pi10 ? n166 : n92;
  assign n168 = pi09 ? n163 : n167;
  assign n169 = pi08 ? n143 : n168;
  assign n170 = pi07 ? n80 : n169;
  assign n171 = pi09 ? n142 : n163;
  assign n172 = pi09 ? n167 : n142;
  assign n173 = pi08 ? n171 : n172;
  assign n174 = pi19 ? n26 : n51;
  assign n175 = pi18 ? n26 : n174;
  assign n176 = pi17 ? n26 : n175;
  assign n177 = pi16 ? n176 : n155;
  assign n178 = pi16 ? n175 : n32;
  assign n179 = pi15 ? n177 : n178;
  assign n180 = pi14 ? n26 : n179;
  assign n181 = pi15 ? n43 : n41;
  assign n182 = pi14 ? n181 : n124;
  assign n183 = pi13 ? n180 : n182;
  assign n184 = pi12 ? n26 : n183;
  assign n185 = pi11 ? n26 : n184;
  assign n186 = pi17 ? n175 : n32;
  assign n187 = pi16 ? n175 : n186;
  assign n188 = pi15 ? n177 : n187;
  assign n189 = pi14 ? n26 : n188;
  assign n190 = pi15 ? n73 : n41;
  assign n191 = pi14 ? n190 : n124;
  assign n192 = pi13 ? n189 : n191;
  assign n193 = pi12 ? n26 : n192;
  assign n194 = pi17 ? n175 : n155;
  assign n195 = pi16 ? n175 : n194;
  assign n196 = pi15 ? n177 : n195;
  assign n197 = pi14 ? n26 : n196;
  assign n198 = pi15 ? n98 : n41;
  assign n199 = pi14 ? n198 : n124;
  assign n200 = pi13 ? n197 : n199;
  assign n201 = pi12 ? n26 : n200;
  assign n202 = pi11 ? n193 : n201;
  assign n203 = pi10 ? n185 : n202;
  assign n204 = pi09 ? n163 : n203;
  assign n205 = pi15 ? n32 : n41;
  assign n206 = pi14 ? n205 : n124;
  assign n207 = pi13 ? n180 : n206;
  assign n208 = pi12 ? n26 : n207;
  assign n209 = pi16 ? n33 : n155;
  assign n210 = pi15 ? n209 : n178;
  assign n211 = pi14 ? n26 : n210;
  assign n212 = pi17 ? n32 : n175;
  assign n213 = pi16 ? n212 : n32;
  assign n214 = pi15 ? n213 : n41;
  assign n215 = pi14 ? n214 : n124;
  assign n216 = pi13 ? n211 : n215;
  assign n217 = pi12 ? n26 : n216;
  assign n218 = pi11 ? n208 : n217;
  assign n219 = pi15 ? n213 : n133;
  assign n220 = pi14 ? n219 : n124;
  assign n221 = pi13 ? n211 : n220;
  assign n222 = pi12 ? n26 : n221;
  assign n223 = pi19 ? n26 : n39;
  assign n224 = pi18 ? n26 : n223;
  assign n225 = pi17 ? n26 : n224;
  assign n226 = pi16 ? n225 : n155;
  assign n227 = pi15 ? n226 : n178;
  assign n228 = pi14 ? n26 : n227;
  assign n229 = pi16 ? n96 : n41;
  assign n230 = pi15 ? n213 : n229;
  assign n231 = pi16 ? n148 : n121;
  assign n232 = pi15 ? n231 : n123;
  assign n233 = pi14 ? n230 : n232;
  assign n234 = pi13 ? n228 : n233;
  assign n235 = pi12 ? n26 : n234;
  assign n236 = pi11 ? n222 : n235;
  assign n237 = pi10 ? n218 : n236;
  assign n238 = pi17 ? n224 : n175;
  assign n239 = pi16 ? n238 : n32;
  assign n240 = pi15 ? n226 : n239;
  assign n241 = pi14 ? n26 : n240;
  assign n242 = pi15 ? n213 : n32;
  assign n243 = pi14 ? n242 : n124;
  assign n244 = pi13 ? n241 : n243;
  assign n245 = pi12 ? n26 : n244;
  assign n246 = pi17 ? n26 : n60;
  assign n247 = pi16 ? n246 : n26;
  assign n248 = pi16 ? n225 : n26;
  assign n249 = pi15 ? n247 : n248;
  assign n250 = pi16 ? n225 : n224;
  assign n251 = pi17 ? n224 : n107;
  assign n252 = pi16 ? n251 : n186;
  assign n253 = pi15 ? n250 : n252;
  assign n254 = pi14 ? n249 : n253;
  assign n255 = pi17 ? n224 : n32;
  assign n256 = pi16 ? n212 : n255;
  assign n257 = pi15 ? n256 : n32;
  assign n258 = pi16 ? n41 : n148;
  assign n259 = pi17 ? n121 : n26;
  assign n260 = pi16 ? n53 : n259;
  assign n261 = pi15 ? n258 : n260;
  assign n262 = pi14 ? n257 : n261;
  assign n263 = pi13 ? n254 : n262;
  assign n264 = pi12 ? n26 : n263;
  assign n265 = pi11 ? n245 : n264;
  assign n266 = pi17 ? n53 : n121;
  assign n267 = pi16 ? n26 : n266;
  assign n268 = pi15 ? n26 : n267;
  assign n269 = pi14 ? n26 : n268;
  assign n270 = pi13 ? n26 : n269;
  assign n271 = pi17 ? n60 : n26;
  assign n272 = pi16 ? n271 : n26;
  assign n273 = pi15 ? n123 : n272;
  assign n274 = pi17 ? n224 : n26;
  assign n275 = pi16 ? n26 : n274;
  assign n276 = pi17 ? n32 : n155;
  assign n277 = pi16 ? n225 : n276;
  assign n278 = pi15 ? n275 : n277;
  assign n279 = pi14 ? n273 : n278;
  assign n280 = pi16 ? n175 : n255;
  assign n281 = pi15 ? n280 : n32;
  assign n282 = pi15 ? n43 : n26;
  assign n283 = pi14 ? n281 : n282;
  assign n284 = pi13 ? n279 : n283;
  assign n285 = pi12 ? n270 : n284;
  assign n286 = pi16 ? n42 : n121;
  assign n287 = pi15 ? n26 : n286;
  assign n288 = pi14 ? n26 : n287;
  assign n289 = pi13 ? n26 : n288;
  assign n290 = pi17 ? n60 : n65;
  assign n291 = pi16 ? n290 : n26;
  assign n292 = pi15 ? n100 : n291;
  assign n293 = pi16 ? n26 : n155;
  assign n294 = pi15 ? n26 : n293;
  assign n295 = pi14 ? n292 : n294;
  assign n296 = pi19 ? n26 : n56;
  assign n297 = pi18 ? n26 : n296;
  assign n298 = pi17 ? n297 : n224;
  assign n299 = pi16 ? n175 : n298;
  assign n300 = pi17 ? n297 : n26;
  assign n301 = pi16 ? n32 : n300;
  assign n302 = pi15 ? n299 : n301;
  assign n303 = pi14 ? n302 : n26;
  assign n304 = pi13 ? n295 : n303;
  assign n305 = pi12 ? n289 : n304;
  assign n306 = pi11 ? n285 : n305;
  assign n307 = pi10 ? n265 : n306;
  assign n308 = pi09 ? n237 : n307;
  assign n309 = pi08 ? n204 : n308;
  assign n310 = pi07 ? n173 : n309;
  assign n311 = pi06 ? n170 : n310;
  assign n312 = pi05 ? n26 : n311;
  assign n313 = pi14 ? n26 : n32;
  assign n314 = pi16 ? n121 : n47;
  assign n315 = pi15 ? n41 : n314;
  assign n316 = pi15 ? n123 : n66;
  assign n317 = pi14 ? n315 : n316;
  assign n318 = pi13 ? n313 : n317;
  assign n319 = pi12 ? n26 : n318;
  assign n320 = pi11 ? n26 : n319;
  assign n321 = pi16 ? n121 : n58;
  assign n322 = pi15 ? n41 : n321;
  assign n323 = pi15 ? n60 : n66;
  assign n324 = pi14 ? n322 : n323;
  assign n325 = pi13 ? n313 : n324;
  assign n326 = pi12 ? n26 : n325;
  assign n327 = pi13 ? n36 : n324;
  assign n328 = pi12 ? n26 : n327;
  assign n329 = pi11 ? n326 : n328;
  assign n330 = pi10 ? n320 : n329;
  assign n331 = pi09 ? n26 : n330;
  assign n332 = pi08 ? n26 : n331;
  assign n333 = pi16 ? n107 : n96;
  assign n334 = pi15 ? n34 : n333;
  assign n335 = pi14 ? n26 : n334;
  assign n336 = pi13 ? n335 : n324;
  assign n337 = pi12 ? n26 : n336;
  assign n338 = pi15 ? n81 : n333;
  assign n339 = pi14 ? n26 : n338;
  assign n340 = pi13 ? n339 : n324;
  assign n341 = pi12 ? n26 : n340;
  assign n342 = pi11 ? n337 : n341;
  assign n343 = pi17 ? n32 : n107;
  assign n344 = pi16 ? n26 : n343;
  assign n345 = pi15 ? n344 : n333;
  assign n346 = pi14 ? n26 : n345;
  assign n347 = pi16 ? n290 : n65;
  assign n348 = pi15 ? n60 : n347;
  assign n349 = pi14 ? n315 : n348;
  assign n350 = pi13 ? n346 : n349;
  assign n351 = pi12 ? n26 : n350;
  assign n352 = pi16 ? n26 : n128;
  assign n353 = pi15 ? n352 : n333;
  assign n354 = pi14 ? n26 : n353;
  assign n355 = pi18 ? n26 : n95;
  assign n356 = pi17 ? n65 : n355;
  assign n357 = pi16 ? n290 : n356;
  assign n358 = pi15 ? n123 : n357;
  assign n359 = pi14 ? n315 : n358;
  assign n360 = pi13 ? n354 : n359;
  assign n361 = pi12 ? n26 : n360;
  assign n362 = pi11 ? n351 : n361;
  assign n363 = pi10 ? n342 : n362;
  assign n364 = pi16 ? n148 : n47;
  assign n365 = pi15 ? n41 : n364;
  assign n366 = pi14 ? n365 : n358;
  assign n367 = pi13 ? n354 : n366;
  assign n368 = pi12 ? n26 : n367;
  assign n369 = pi15 ? n26 : n333;
  assign n370 = pi14 ? n26 : n369;
  assign n371 = pi15 ? n100 : n357;
  assign n372 = pi14 ? n365 : n371;
  assign n373 = pi13 ? n370 : n372;
  assign n374 = pi12 ? n26 : n373;
  assign n375 = pi11 ? n368 : n374;
  assign n376 = pi15 ? n41 : n48;
  assign n377 = pi16 ? n60 : n356;
  assign n378 = pi15 ? n100 : n377;
  assign n379 = pi14 ? n376 : n378;
  assign n380 = pi13 ? n370 : n379;
  assign n381 = pi12 ? n26 : n380;
  assign n382 = pi16 ? n176 : n32;
  assign n383 = pi15 ? n26 : n382;
  assign n384 = pi14 ? n26 : n383;
  assign n385 = pi16 ? n41 : n96;
  assign n386 = pi15 ? n41 : n385;
  assign n387 = pi15 ? n122 : n100;
  assign n388 = pi14 ? n386 : n387;
  assign n389 = pi13 ? n384 : n388;
  assign n390 = pi12 ? n26 : n389;
  assign n391 = pi11 ? n381 : n390;
  assign n392 = pi10 ? n375 : n391;
  assign n393 = pi09 ? n363 : n392;
  assign n394 = pi16 ? n26 : n186;
  assign n395 = pi15 ? n26 : n394;
  assign n396 = pi14 ? n26 : n395;
  assign n397 = pi16 ? n32 : n343;
  assign n398 = pi15 ? n397 : n333;
  assign n399 = pi16 ? n121 : n259;
  assign n400 = pi15 ? n41 : n399;
  assign n401 = pi14 ? n398 : n400;
  assign n402 = pi13 ? n396 : n401;
  assign n403 = pi12 ? n26 : n402;
  assign n404 = pi17 ? n26 : n155;
  assign n405 = pi16 ? n26 : n404;
  assign n406 = pi15 ? n26 : n405;
  assign n407 = pi14 ? n26 : n406;
  assign n408 = pi15 ? n157 : n114;
  assign n409 = pi15 ? n73 : n26;
  assign n410 = pi14 ? n408 : n409;
  assign n411 = pi13 ? n407 : n410;
  assign n412 = pi12 ? n26 : n411;
  assign n413 = pi11 ? n403 : n412;
  assign n414 = pi10 ? n413 : n26;
  assign n415 = pi13 ? n83 : n317;
  assign n416 = pi12 ? n26 : n415;
  assign n417 = pi11 ? n26 : n416;
  assign n418 = pi10 ? n417 : n362;
  assign n419 = pi09 ? n414 : n418;
  assign n420 = pi08 ? n393 : n419;
  assign n421 = pi07 ? n332 : n420;
  assign n422 = pi09 ? n392 : n414;
  assign n423 = pi09 ? n418 : n392;
  assign n424 = pi08 ? n422 : n423;
  assign n425 = pi15 ? n178 : n32;
  assign n426 = pi14 ? n26 : n425;
  assign n427 = pi15 ? n122 : n66;
  assign n428 = pi14 ? n41 : n427;
  assign n429 = pi13 ? n426 : n428;
  assign n430 = pi12 ? n26 : n429;
  assign n431 = pi11 ? n26 : n430;
  assign n432 = pi16 ? n41 : n58;
  assign n433 = pi15 ? n432 : n60;
  assign n434 = pi14 ? n190 : n433;
  assign n435 = pi13 ? n313 : n434;
  assign n436 = pi12 ? n26 : n435;
  assign n437 = pi17 ? n297 : n41;
  assign n438 = pi16 ? n32 : n437;
  assign n439 = pi15 ? n438 : n41;
  assign n440 = pi14 ? n439 : n433;
  assign n441 = pi13 ? n313 : n440;
  assign n442 = pi12 ? n26 : n441;
  assign n443 = pi11 ? n436 : n442;
  assign n444 = pi10 ? n431 : n443;
  assign n445 = pi09 ? n414 : n444;
  assign n446 = pi17 ? n297 : n96;
  assign n447 = pi16 ? n32 : n446;
  assign n448 = pi15 ? n447 : n41;
  assign n449 = pi14 ? n448 : n433;
  assign n450 = pi13 ? n313 : n449;
  assign n451 = pi12 ? n26 : n450;
  assign n452 = pi17 ? n297 : n32;
  assign n453 = pi16 ? n156 : n452;
  assign n454 = pi15 ? n453 : n32;
  assign n455 = pi14 ? n406 : n454;
  assign n456 = pi16 ? n32 : n452;
  assign n457 = pi15 ? n456 : n229;
  assign n458 = pi14 ? n457 : n124;
  assign n459 = pi13 ? n455 : n458;
  assign n460 = pi12 ? n26 : n459;
  assign n461 = pi17 ? n155 : n224;
  assign n462 = pi16 ? n26 : n461;
  assign n463 = pi15 ? n26 : n462;
  assign n464 = pi16 ? n224 : n461;
  assign n465 = pi15 ? n464 : n32;
  assign n466 = pi14 ? n463 : n465;
  assign n467 = pi16 ? n32 : n298;
  assign n468 = pi15 ? n467 : n133;
  assign n469 = pi14 ? n468 : n124;
  assign n470 = pi13 ? n466 : n469;
  assign n471 = pi12 ? n26 : n470;
  assign n472 = pi11 ? n460 : n471;
  assign n473 = pi10 ? n451 : n472;
  assign n474 = pi15 ? n26 : n250;
  assign n475 = pi16 ? n224 : n155;
  assign n476 = pi17 ? n107 : n32;
  assign n477 = pi16 ? n476 : n32;
  assign n478 = pi15 ? n475 : n477;
  assign n479 = pi14 ? n474 : n478;
  assign n480 = pi16 ? n32 : n96;
  assign n481 = pi15 ? n467 : n480;
  assign n482 = pi17 ? n47 : n60;
  assign n483 = pi16 ? n482 : n60;
  assign n484 = pi15 ? n231 : n483;
  assign n485 = pi14 ? n481 : n484;
  assign n486 = pi13 ? n479 : n485;
  assign n487 = pi12 ? n26 : n486;
  assign n488 = pi17 ? n26 : n58;
  assign n489 = pi16 ? n26 : n488;
  assign n490 = pi15 ? n26 : n489;
  assign n491 = pi14 ? n26 : n490;
  assign n492 = pi13 ? n26 : n491;
  assign n493 = pi16 ? n60 : n224;
  assign n494 = pi15 ? n493 : n224;
  assign n495 = pi15 ? n224 : n187;
  assign n496 = pi14 ? n494 : n495;
  assign n497 = pi15 ? n467 : n32;
  assign n498 = pi22 ? n27 : ~n26;
  assign n499 = pi21 ? n26 : ~n498;
  assign n500 = pi20 ? n26 : n499;
  assign n501 = pi19 ? n500 : n26;
  assign n502 = pi18 ? n501 : n26;
  assign n503 = pi16 ? n502 : n135;
  assign n504 = pi15 ? n122 : n503;
  assign n505 = pi14 ? n497 : n504;
  assign n506 = pi13 ? n496 : n505;
  assign n507 = pi12 ? n492 : n506;
  assign n508 = pi11 ? n487 : n507;
  assign n509 = pi16 ? n65 : n224;
  assign n510 = pi15 ? n509 : n475;
  assign n511 = pi14 ? n101 : n510;
  assign n512 = pi16 ? n156 : n298;
  assign n513 = pi15 ? n512 : n32;
  assign n514 = pi15 ? n438 : n149;
  assign n515 = pi14 ? n513 : n514;
  assign n516 = pi13 ? n511 : n515;
  assign n517 = pi12 ? n289 : n516;
  assign n518 = pi17 ? n26 : n96;
  assign n519 = pi16 ? n518 : n41;
  assign n520 = pi15 ? n26 : n519;
  assign n521 = pi14 ? n26 : n520;
  assign n522 = pi13 ? n26 : n521;
  assign n523 = pi15 ? n100 : n347;
  assign n524 = pi16 ? n65 : n26;
  assign n525 = pi15 ? n524 : n226;
  assign n526 = pi14 ? n523 : n525;
  assign n527 = pi16 ? n175 : n461;
  assign n528 = pi17 ? n297 : n155;
  assign n529 = pi16 ? n32 : n528;
  assign n530 = pi15 ? n527 : n529;
  assign n531 = pi14 ? n530 : n26;
  assign n532 = pi13 ? n526 : n531;
  assign n533 = pi12 ? n522 : n532;
  assign n534 = pi11 ? n517 : n533;
  assign n535 = pi10 ? n508 : n534;
  assign n536 = pi09 ? n473 : n535;
  assign n537 = pi08 ? n445 : n536;
  assign n538 = pi07 ? n424 : n537;
  assign n539 = pi06 ? n421 : n538;
  assign n540 = pi14 ? n26 : n134;
  assign n541 = pi17 ? n47 : n502;
  assign n542 = pi16 ? n541 : n58;
  assign n543 = pi15 ? n122 : n542;
  assign n544 = pi16 ? n60 : n61;
  assign n545 = pi17 ? n355 : n224;
  assign n546 = pi16 ? n545 : n224;
  assign n547 = pi15 ? n544 : n546;
  assign n548 = pi14 ? n543 : n547;
  assign n549 = pi13 ? n540 : n548;
  assign n550 = pi12 ? n26 : n549;
  assign n551 = pi11 ? n26 : n550;
  assign n552 = pi16 ? n26 : n518;
  assign n553 = pi15 ? n26 : n552;
  assign n554 = pi16 ? n96 : n32;
  assign n555 = pi16 ? n32 : n132;
  assign n556 = pi15 ? n554 : n555;
  assign n557 = pi14 ? n553 : n556;
  assign n558 = pi16 ? n545 : n65;
  assign n559 = pi15 ? n493 : n558;
  assign n560 = pi14 ? n543 : n559;
  assign n561 = pi13 ? n557 : n560;
  assign n562 = pi12 ? n26 : n561;
  assign n563 = pi17 ? n96 : n32;
  assign n564 = pi16 ? n563 : n32;
  assign n565 = pi15 ? n564 : n555;
  assign n566 = pi14 ? n26 : n565;
  assign n567 = pi13 ? n566 : n560;
  assign n568 = pi12 ? n26 : n567;
  assign n569 = pi11 ? n562 : n568;
  assign n570 = pi10 ? n551 : n569;
  assign n571 = pi09 ? n26 : n570;
  assign n572 = pi08 ? n26 : n571;
  assign n573 = pi16 ? n41 : n32;
  assign n574 = pi16 ? n107 : n41;
  assign n575 = pi15 ? n573 : n574;
  assign n576 = pi14 ? n26 : n575;
  assign n577 = pi13 ? n576 : n560;
  assign n578 = pi12 ? n26 : n577;
  assign n579 = pi16 ? n518 : n32;
  assign n580 = pi15 ? n579 : n574;
  assign n581 = pi14 ? n26 : n580;
  assign n582 = pi13 ? n581 : n560;
  assign n583 = pi12 ? n26 : n582;
  assign n584 = pi11 ? n578 : n583;
  assign n585 = pi15 ? n519 : n229;
  assign n586 = pi14 ? n26 : n585;
  assign n587 = pi15 ? n493 : n546;
  assign n588 = pi14 ? n543 : n587;
  assign n589 = pi13 ? n586 : n588;
  assign n590 = pi12 ? n26 : n589;
  assign n591 = pi16 ? n26 : n41;
  assign n592 = pi15 ? n591 : n229;
  assign n593 = pi14 ? n26 : n592;
  assign n594 = pi13 ? n593 : n588;
  assign n595 = pi12 ? n26 : n594;
  assign n596 = pi11 ? n590 : n595;
  assign n597 = pi10 ? n584 : n596;
  assign n598 = pi16 ? n26 : n132;
  assign n599 = pi15 ? n598 : n229;
  assign n600 = pi14 ? n26 : n599;
  assign n601 = pi13 ? n600 : n588;
  assign n602 = pi12 ? n26 : n601;
  assign n603 = pi15 ? n43 : n229;
  assign n604 = pi14 ? n26 : n603;
  assign n605 = pi13 ? n604 : n588;
  assign n606 = pi12 ? n26 : n605;
  assign n607 = pi11 ? n602 : n606;
  assign n608 = pi15 ? n26 : n96;
  assign n609 = pi14 ? n26 : n608;
  assign n610 = pi16 ? n60 : n355;
  assign n611 = pi15 ? n100 : n610;
  assign n612 = pi14 ? n376 : n611;
  assign n613 = pi13 ? n609 : n612;
  assign n614 = pi12 ? n26 : n613;
  assign n615 = pi15 ? n26 : n187;
  assign n616 = pi14 ? n26 : n615;
  assign n617 = pi14 ? n386 : n232;
  assign n618 = pi13 ? n616 : n617;
  assign n619 = pi12 ? n26 : n618;
  assign n620 = pi11 ? n614 : n619;
  assign n621 = pi10 ? n607 : n620;
  assign n622 = pi09 ? n597 : n621;
  assign n623 = pi16 ? n176 : n186;
  assign n624 = pi15 ? n26 : n623;
  assign n625 = pi14 ? n26 : n624;
  assign n626 = pi17 ? n121 : n60;
  assign n627 = pi16 ? n121 : n626;
  assign n628 = pi15 ? n41 : n627;
  assign n629 = pi14 ? n398 : n628;
  assign n630 = pi13 ? n625 : n629;
  assign n631 = pi12 ? n26 : n630;
  assign n632 = pi14 ? n26 : n294;
  assign n633 = pi14 ? n408 : n514;
  assign n634 = pi13 ? n632 : n633;
  assign n635 = pi12 ? n26 : n634;
  assign n636 = pi11 ? n631 : n635;
  assign n637 = pi10 ? n636 : n26;
  assign n638 = pi15 ? n34 : n133;
  assign n639 = pi14 ? n26 : n638;
  assign n640 = pi13 ? n639 : n548;
  assign n641 = pi12 ? n26 : n640;
  assign n642 = pi11 ? n26 : n641;
  assign n643 = pi16 ? n42 : n41;
  assign n644 = pi15 ? n643 : n229;
  assign n645 = pi14 ? n26 : n644;
  assign n646 = pi13 ? n645 : n588;
  assign n647 = pi12 ? n26 : n646;
  assign n648 = pi11 ? n647 : n595;
  assign n649 = pi10 ? n642 : n648;
  assign n650 = pi09 ? n637 : n649;
  assign n651 = pi08 ? n622 : n650;
  assign n652 = pi07 ? n572 : n651;
  assign n653 = pi09 ? n621 : n637;
  assign n654 = pi09 ? n649 : n621;
  assign n655 = pi08 ? n653 : n654;
  assign n656 = pi15 ? n26 : n87;
  assign n657 = pi14 ? n656 : n32;
  assign n658 = pi15 ? n432 : n66;
  assign n659 = pi14 ? n41 : n658;
  assign n660 = pi13 ? n657 : n659;
  assign n661 = pi12 ? n26 : n660;
  assign n662 = pi11 ? n26 : n661;
  assign n663 = pi13 ? n657 : n434;
  assign n664 = pi12 ? n26 : n663;
  assign n665 = pi14 ? n205 : n433;
  assign n666 = pi13 ? n657 : n665;
  assign n667 = pi12 ? n26 : n666;
  assign n668 = pi11 ? n664 : n667;
  assign n669 = pi10 ? n662 : n668;
  assign n670 = pi09 ? n637 : n669;
  assign n671 = pi14 ? n553 : n32;
  assign n672 = pi13 ? n671 : n665;
  assign n673 = pi12 ? n26 : n672;
  assign n674 = pi16 ? n26 : n276;
  assign n675 = pi15 ? n26 : n674;
  assign n676 = pi19 ? n26 : n500;
  assign n677 = pi18 ? n26 : n676;
  assign n678 = pi16 ? n677 : n32;
  assign n679 = pi15 ? n678 : n32;
  assign n680 = pi14 ? n675 : n679;
  assign n681 = pi13 ? n680 : n665;
  assign n682 = pi12 ? n26 : n681;
  assign n683 = pi11 ? n673 : n682;
  assign n684 = pi14 ? n294 : n425;
  assign n685 = pi15 ? n32 : n229;
  assign n686 = pi14 ? n685 : n658;
  assign n687 = pi13 ? n684 : n686;
  assign n688 = pi12 ? n26 : n687;
  assign n689 = pi16 ? n225 : n461;
  assign n690 = pi15 ? n26 : n689;
  assign n691 = pi16 ? n238 : n461;
  assign n692 = pi15 ? n691 : n32;
  assign n693 = pi14 ? n690 : n692;
  assign n694 = pi16 ? n41 : n626;
  assign n695 = pi15 ? n694 : n377;
  assign n696 = pi14 ? n134 : n695;
  assign n697 = pi13 ? n693 : n696;
  assign n698 = pi12 ? n26 : n697;
  assign n699 = pi11 ? n688 : n698;
  assign n700 = pi10 ? n683 : n699;
  assign n701 = pi16 ? n26 : n224;
  assign n702 = pi15 ? n701 : n224;
  assign n703 = pi15 ? n475 : n32;
  assign n704 = pi14 ? n702 : n703;
  assign n705 = pi16 ? n32 : n41;
  assign n706 = pi15 ? n32 : n705;
  assign n707 = pi17 ? n121 : n58;
  assign n708 = pi16 ? n41 : n707;
  assign n709 = pi15 ? n708 : n377;
  assign n710 = pi14 ? n706 : n709;
  assign n711 = pi13 ? n704 : n710;
  assign n712 = pi12 ? n26 : n711;
  assign n713 = pi16 ? n26 : n58;
  assign n714 = pi15 ? n26 : n713;
  assign n715 = pi14 ? n26 : n714;
  assign n716 = pi13 ? n26 : n715;
  assign n717 = pi16 ? n60 : n135;
  assign n718 = pi16 ? n461 : n224;
  assign n719 = pi15 ? n717 : n718;
  assign n720 = pi15 ? n475 : n678;
  assign n721 = pi14 ? n719 : n720;
  assign n722 = pi16 ? n502 : n58;
  assign n723 = pi15 ? n122 : n722;
  assign n724 = pi14 ? n32 : n723;
  assign n725 = pi13 ? n721 : n724;
  assign n726 = pi12 ? n716 : n725;
  assign n727 = pi11 ? n712 : n726;
  assign n728 = pi15 ? n722 : n66;
  assign n729 = pi14 ? n728 : n510;
  assign n730 = pi16 ? n148 : n259;
  assign n731 = pi15 ? n147 : n730;
  assign n732 = pi14 ? n425 : n731;
  assign n733 = pi13 ? n729 : n732;
  assign n734 = pi12 ? n289 : n733;
  assign n735 = pi16 ? n128 : n132;
  assign n736 = pi15 ? n26 : n735;
  assign n737 = pi14 ? n26 : n736;
  assign n738 = pi13 ? n26 : n737;
  assign n739 = pi16 ? n65 : n60;
  assign n740 = pi17 ? n60 : n224;
  assign n741 = pi16 ? n740 : n461;
  assign n742 = pi15 ? n739 : n741;
  assign n743 = pi14 ? n658 : n742;
  assign n744 = pi16 ? n238 : n155;
  assign n745 = pi15 ? n744 : n32;
  assign n746 = pi17 ? n32 : n26;
  assign n747 = pi16 ? n32 : n746;
  assign n748 = pi15 ? n747 : n26;
  assign n749 = pi14 ? n745 : n748;
  assign n750 = pi13 ? n743 : n749;
  assign n751 = pi12 ? n738 : n750;
  assign n752 = pi11 ? n734 : n751;
  assign n753 = pi10 ? n727 : n752;
  assign n754 = pi09 ? n700 : n753;
  assign n755 = pi08 ? n670 : n754;
  assign n756 = pi07 ? n655 : n755;
  assign n757 = pi06 ? n652 : n756;
  assign n758 = pi05 ? n539 : n757;
  assign n759 = pi04 ? n312 : n758;
  assign n760 = pi03 ? n26 : n759;
  assign n761 = pi02 ? n26 : n760;
  assign n762 = pi14 ? n656 : n117;
  assign n763 = pi16 ? n60 : n58;
  assign n764 = pi15 ? n122 : n763;
  assign n765 = pi14 ? n764 : n547;
  assign n766 = pi13 ? n762 : n765;
  assign n767 = pi12 ? n26 : n766;
  assign n768 = pi11 ? n26 : n767;
  assign n769 = pi14 ? n553 : n117;
  assign n770 = pi15 ? n122 : n60;
  assign n771 = pi16 ? n740 : n224;
  assign n772 = pi15 ? n771 : n224;
  assign n773 = pi14 ? n770 : n772;
  assign n774 = pi13 ? n769 : n773;
  assign n775 = pi12 ? n26 : n774;
  assign n776 = pi14 ? n770 : n224;
  assign n777 = pi13 ? n769 : n776;
  assign n778 = pi12 ? n26 : n777;
  assign n779 = pi11 ? n775 : n778;
  assign n780 = pi10 ? n768 : n779;
  assign n781 = pi09 ? n26 : n780;
  assign n782 = pi08 ? n26 : n781;
  assign n783 = pi15 ? n573 : n41;
  assign n784 = pi14 ? n553 : n783;
  assign n785 = pi14 ? n433 : n224;
  assign n786 = pi13 ? n784 : n785;
  assign n787 = pi12 ? n26 : n786;
  assign n788 = pi17 ? n47 : n96;
  assign n789 = pi16 ? n788 : n41;
  assign n790 = pi15 ? n789 : n41;
  assign n791 = pi14 ? n26 : n790;
  assign n792 = pi13 ? n791 : n785;
  assign n793 = pi12 ? n26 : n792;
  assign n794 = pi11 ? n787 : n793;
  assign n795 = pi15 ? n643 : n258;
  assign n796 = pi14 ? n26 : n795;
  assign n797 = pi14 ? n378 : n224;
  assign n798 = pi13 ? n796 : n797;
  assign n799 = pi12 ? n26 : n798;
  assign n800 = pi15 ? n591 : n258;
  assign n801 = pi14 ? n26 : n800;
  assign n802 = pi15 ? n100 : n493;
  assign n803 = pi14 ? n802 : n224;
  assign n804 = pi13 ? n801 : n803;
  assign n805 = pi12 ? n26 : n804;
  assign n806 = pi11 ? n799 : n805;
  assign n807 = pi10 ? n794 : n806;
  assign n808 = pi16 ? n32 : n186;
  assign n809 = pi15 ? n405 : n808;
  assign n810 = pi14 ? n26 : n809;
  assign n811 = pi15 ? n385 : n229;
  assign n812 = pi14 ? n811 : n124;
  assign n813 = pi13 ? n810 : n812;
  assign n814 = pi12 ? n26 : n813;
  assign n815 = pi11 ? n26 : n814;
  assign n816 = pi10 ? n26 : n815;
  assign n817 = pi09 ? n807 : n816;
  assign n818 = pi15 ? n405 : n187;
  assign n819 = pi14 ? n26 : n818;
  assign n820 = pi15 ? n231 : n136;
  assign n821 = pi14 ? n398 : n820;
  assign n822 = pi13 ? n819 : n821;
  assign n823 = pi12 ? n26 : n822;
  assign n824 = pi15 ? n26 : n226;
  assign n825 = pi14 ? n26 : n824;
  assign n826 = pi15 ? n438 : n730;
  assign n827 = pi14 ? n408 : n826;
  assign n828 = pi13 ? n825 : n827;
  assign n829 = pi12 ? n26 : n828;
  assign n830 = pi11 ? n823 : n829;
  assign n831 = pi10 ? n830 : n26;
  assign n832 = pi15 ? n34 : n96;
  assign n833 = pi14 ? n26 : n832;
  assign n834 = pi14 ? n770 : n547;
  assign n835 = pi13 ? n833 : n834;
  assign n836 = pi12 ? n26 : n835;
  assign n837 = pi11 ? n26 : n836;
  assign n838 = pi15 ? n519 : n258;
  assign n839 = pi14 ? n26 : n838;
  assign n840 = pi15 ? n546 : n224;
  assign n841 = pi14 ? n378 : n840;
  assign n842 = pi13 ? n839 : n841;
  assign n843 = pi12 ? n26 : n842;
  assign n844 = pi11 ? n843 : n805;
  assign n845 = pi10 ? n837 : n844;
  assign n846 = pi09 ? n831 : n845;
  assign n847 = pi08 ? n817 : n846;
  assign n848 = pi07 ? n782 : n847;
  assign n849 = pi09 ? n816 : n831;
  assign n850 = pi09 ? n845 : n816;
  assign n851 = pi08 ? n849 : n850;
  assign n852 = pi14 ? n144 : n32;
  assign n853 = pi17 ? n65 : n58;
  assign n854 = pi16 ? n53 : n853;
  assign n855 = pi15 ? n854 : n493;
  assign n856 = pi14 ? n365 : n855;
  assign n857 = pi13 ? n852 : n856;
  assign n858 = pi12 ? n26 : n857;
  assign n859 = pi11 ? n26 : n858;
  assign n860 = pi15 ? n147 : n364;
  assign n861 = pi14 ? n860 : n855;
  assign n862 = pi13 ? n852 : n861;
  assign n863 = pi12 ? n26 : n862;
  assign n864 = pi10 ? n859 : n863;
  assign n865 = pi09 ? n831 : n864;
  assign n866 = pi16 ? n128 : n276;
  assign n867 = pi15 ? n26 : n866;
  assign n868 = pi14 ? n867 : n32;
  assign n869 = pi13 ? n868 : n861;
  assign n870 = pi12 ? n26 : n869;
  assign n871 = pi11 ? n863 : n870;
  assign n872 = pi14 ? n824 : n425;
  assign n873 = pi15 ? n854 : n66;
  assign n874 = pi14 ? n860 : n873;
  assign n875 = pi13 ? n872 : n874;
  assign n876 = pi12 ? n26 : n875;
  assign n877 = pi15 ? n405 : n475;
  assign n878 = pi14 ? n877 : n454;
  assign n879 = pi13 ? n878 : n861;
  assign n880 = pi12 ? n26 : n879;
  assign n881 = pi11 ? n876 : n880;
  assign n882 = pi10 ? n871 : n881;
  assign n883 = pi15 ? n250 : n475;
  assign n884 = pi14 ? n883 : n679;
  assign n885 = pi14 ? n860 : n611;
  assign n886 = pi13 ? n884 : n885;
  assign n887 = pi12 ? n26 : n886;
  assign n888 = pi14 ? n26 : n474;
  assign n889 = pi13 ? n26 : n888;
  assign n890 = pi15 ? n224 : n475;
  assign n891 = pi14 ? n890 : n679;
  assign n892 = pi16 ? n41 : n224;
  assign n893 = pi16 ? n224 : n47;
  assign n894 = pi15 ? n892 : n893;
  assign n895 = pi14 ? n894 : n611;
  assign n896 = pi13 ? n891 : n895;
  assign n897 = pi12 ? n889 : n896;
  assign n898 = pi11 ? n887 : n897;
  assign n899 = pi15 ? n60 : n224;
  assign n900 = pi14 ? n723 : n899;
  assign n901 = pi15 ? n224 : n678;
  assign n902 = pi15 ? n32 : n224;
  assign n903 = pi14 ? n901 : n902;
  assign n904 = pi13 ? n900 : n903;
  assign n905 = pi12 ? n889 : n904;
  assign n906 = pi16 ? n518 : n132;
  assign n907 = pi15 ? n26 : n906;
  assign n908 = pi14 ? n26 : n907;
  assign n909 = pi13 ? n26 : n908;
  assign n910 = pi15 ? n60 : n771;
  assign n911 = pi14 ? n723 : n910;
  assign n912 = pi15 ? n32 : n26;
  assign n913 = pi14 ? n901 : n912;
  assign n914 = pi13 ? n911 : n913;
  assign n915 = pi12 ? n909 : n914;
  assign n916 = pi11 ? n905 : n915;
  assign n917 = pi10 ? n898 : n916;
  assign n918 = pi09 ? n882 : n917;
  assign n919 = pi08 ? n865 : n918;
  assign n920 = pi07 ? n851 : n919;
  assign n921 = pi06 ? n848 : n920;
  assign n922 = pi14 ? n144 : n685;
  assign n923 = pi16 ? n502 : n60;
  assign n924 = pi15 ? n122 : n923;
  assign n925 = pi16 ? n545 : n461;
  assign n926 = pi15 ? n60 : n925;
  assign n927 = pi14 ? n924 : n926;
  assign n928 = pi13 ? n922 : n927;
  assign n929 = pi12 ? n26 : n928;
  assign n930 = pi11 ? n26 : n929;
  assign n931 = pi14 ? n770 : n840;
  assign n932 = pi13 ? n922 : n931;
  assign n933 = pi12 ? n26 : n932;
  assign n934 = pi16 ? n26 : n96;
  assign n935 = pi15 ? n26 : n934;
  assign n936 = pi16 ? n96 : n148;
  assign n937 = pi15 ? n32 : n936;
  assign n938 = pi14 ? n935 : n937;
  assign n939 = pi15 ? n464 : n546;
  assign n940 = pi14 ? n770 : n939;
  assign n941 = pi13 ? n938 : n940;
  assign n942 = pi12 ? n26 : n941;
  assign n943 = pi11 ? n933 : n942;
  assign n944 = pi10 ? n930 : n943;
  assign n945 = pi09 ? n26 : n944;
  assign n946 = pi08 ? n26 : n945;
  assign n947 = pi16 ? n41 : n97;
  assign n948 = pi15 ? n947 : n258;
  assign n949 = pi14 ? n935 : n948;
  assign n950 = pi14 ? n378 : n939;
  assign n951 = pi13 ? n949 : n950;
  assign n952 = pi12 ? n26 : n951;
  assign n953 = pi14 ? n553 : n41;
  assign n954 = pi14 ? n802 : n939;
  assign n955 = pi13 ? n953 : n954;
  assign n956 = pi12 ? n26 : n955;
  assign n957 = pi11 ? n952 : n956;
  assign n958 = pi15 ? n41 : n122;
  assign n959 = pi14 ? n26 : n958;
  assign n960 = pi15 ? n100 : n771;
  assign n961 = pi16 ? n255 : n461;
  assign n962 = pi17 ? n224 : n155;
  assign n963 = pi16 ? n545 : n962;
  assign n964 = pi15 ? n961 : n963;
  assign n965 = pi14 ? n960 : n964;
  assign n966 = pi13 ? n959 : n965;
  assign n967 = pi12 ? n26 : n966;
  assign n968 = pi17 ? n96 : n121;
  assign n969 = pi16 ? n518 : n968;
  assign n970 = pi15 ? n969 : n542;
  assign n971 = pi14 ? n26 : n970;
  assign n972 = pi16 ? n677 : n300;
  assign n973 = pi15 ? n961 : n972;
  assign n974 = pi14 ? n494 : n973;
  assign n975 = pi13 ? n971 : n974;
  assign n976 = pi12 ? n26 : n975;
  assign n977 = pi11 ? n967 : n976;
  assign n978 = pi10 ? n957 : n977;
  assign n979 = pi16 ? n53 : n626;
  assign n980 = pi15 ? n979 : n66;
  assign n981 = pi14 ? n811 : n980;
  assign n982 = pi13 ? n36 : n981;
  assign n983 = pi12 ? n26 : n982;
  assign n984 = pi11 ? n26 : n983;
  assign n985 = pi10 ? n26 : n984;
  assign n986 = pi09 ? n978 : n985;
  assign n987 = pi15 ? n293 : n114;
  assign n988 = pi14 ? n26 : n987;
  assign n989 = pi16 ? n107 : n132;
  assign n990 = pi15 ? n397 : n989;
  assign n991 = pi17 ? n53 : n65;
  assign n992 = pi16 ? n991 : n60;
  assign n993 = pi15 ? n231 : n992;
  assign n994 = pi14 ? n990 : n993;
  assign n995 = pi13 ? n988 : n994;
  assign n996 = pi12 ? n26 : n995;
  assign n997 = pi16 ? n186 : n32;
  assign n998 = pi15 ? n293 : n997;
  assign n999 = pi14 ? n26 : n998;
  assign n1000 = pi16 ? n107 : n72;
  assign n1001 = pi15 ? n32 : n1000;
  assign n1002 = pi14 ? n1001 : n232;
  assign n1003 = pi13 ? n999 : n1002;
  assign n1004 = pi12 ? n26 : n1003;
  assign n1005 = pi11 ? n996 : n1004;
  assign n1006 = pi10 ? n1005 : n26;
  assign n1007 = pi16 ? n33 : n107;
  assign n1008 = pi15 ? n1007 : n229;
  assign n1009 = pi14 ? n26 : n1008;
  assign n1010 = pi14 ? n101 : n926;
  assign n1011 = pi13 ? n1009 : n1010;
  assign n1012 = pi12 ? n26 : n1011;
  assign n1013 = pi11 ? n26 : n1012;
  assign n1014 = pi16 ? n224 : n962;
  assign n1015 = pi15 ? n546 : n1014;
  assign n1016 = pi14 ? n371 : n1015;
  assign n1017 = pi13 ? n959 : n1016;
  assign n1018 = pi12 ? n26 : n1017;
  assign n1019 = pi16 ? n42 : n968;
  assign n1020 = pi15 ? n1019 : n542;
  assign n1021 = pi14 ? n26 : n1020;
  assign n1022 = pi15 ? n464 : n972;
  assign n1023 = pi14 ? n494 : n1022;
  assign n1024 = pi13 ? n1021 : n1023;
  assign n1025 = pi12 ? n26 : n1024;
  assign n1026 = pi11 ? n1018 : n1025;
  assign n1027 = pi10 ? n1013 : n1026;
  assign n1028 = pi09 ? n1006 : n1027;
  assign n1029 = pi08 ? n986 : n1028;
  assign n1030 = pi07 ? n946 : n1029;
  assign n1031 = pi09 ? n985 : n1006;
  assign n1032 = pi09 ? n1027 : n985;
  assign n1033 = pi08 ? n1031 : n1032;
  assign n1034 = pi15 ? n32 : n554;
  assign n1035 = pi14 ? n130 : n1034;
  assign n1036 = pi14 ? n723 : n547;
  assign n1037 = pi13 ? n1035 : n1036;
  assign n1038 = pi12 ? n26 : n1037;
  assign n1039 = pi11 ? n26 : n1038;
  assign n1040 = pi15 ? n32 : n555;
  assign n1041 = pi14 ? n130 : n1040;
  assign n1042 = pi13 ? n1041 : n1036;
  assign n1043 = pi12 ? n26 : n1042;
  assign n1044 = pi15 ? n26 : n579;
  assign n1045 = pi14 ? n1044 : n1040;
  assign n1046 = pi13 ? n1045 : n1036;
  assign n1047 = pi12 ? n26 : n1046;
  assign n1048 = pi11 ? n1043 : n1047;
  assign n1049 = pi10 ? n1039 : n1048;
  assign n1050 = pi09 ? n1006 : n1049;
  assign n1051 = pi17 ? n107 : n175;
  assign n1052 = pi16 ? n1051 : n186;
  assign n1053 = pi15 ? n26 : n1052;
  assign n1054 = pi14 ? n1053 : n1040;
  assign n1055 = pi13 ? n1054 : n1036;
  assign n1056 = pi12 ? n26 : n1055;
  assign n1057 = pi11 ? n1043 : n1056;
  assign n1058 = pi14 ? n615 : n1040;
  assign n1059 = pi13 ? n1058 : n1036;
  assign n1060 = pi12 ? n26 : n1059;
  assign n1061 = pi15 ? n462 : n187;
  assign n1062 = pi15 ? n456 : n555;
  assign n1063 = pi14 ? n1061 : n1062;
  assign n1064 = pi16 ? n355 : n224;
  assign n1065 = pi15 ? n544 : n1064;
  assign n1066 = pi14 ? n723 : n1065;
  assign n1067 = pi13 ? n1063 : n1066;
  assign n1068 = pi12 ? n26 : n1067;
  assign n1069 = pi11 ? n1060 : n1068;
  assign n1070 = pi10 ? n1057 : n1069;
  assign n1071 = pi19 ? n26 : n45;
  assign n1072 = pi18 ? n26 : n1071;
  assign n1073 = pi16 ? n1072 : n32;
  assign n1074 = pi15 ? n250 : n1073;
  assign n1075 = pi14 ? n1074 : n1040;
  assign n1076 = pi15 ? n544 : n493;
  assign n1077 = pi14 ? n723 : n1076;
  assign n1078 = pi13 ? n1075 : n1077;
  assign n1079 = pi12 ? n26 : n1078;
  assign n1080 = pi15 ? n224 : n1073;
  assign n1081 = pi16 ? n32 : n224;
  assign n1082 = pi15 ? n32 : n1081;
  assign n1083 = pi14 ? n1080 : n1082;
  assign n1084 = pi14 ? n723 : n493;
  assign n1085 = pi13 ? n1083 : n1084;
  assign n1086 = pi12 ? n889 : n1085;
  assign n1087 = pi11 ? n1079 : n1086;
  assign n1088 = pi16 ? n225 : n32;
  assign n1089 = pi15 ? n26 : n1088;
  assign n1090 = pi14 ? n26 : n1089;
  assign n1091 = pi13 ? n26 : n1090;
  assign n1092 = pi15 ? n892 : n122;
  assign n1093 = pi15 ? n722 : n224;
  assign n1094 = pi14 ? n1092 : n1093;
  assign n1095 = pi15 ? n178 : n224;
  assign n1096 = pi14 ? n890 : n1095;
  assign n1097 = pi13 ? n1094 : n1096;
  assign n1098 = pi12 ? n1091 : n1097;
  assign n1099 = pi15 ? n26 : n34;
  assign n1100 = pi14 ? n26 : n1099;
  assign n1101 = pi13 ? n26 : n1100;
  assign n1102 = pi15 ? n147 : n122;
  assign n1103 = pi15 ? n722 : n771;
  assign n1104 = pi14 ? n1102 : n1103;
  assign n1105 = pi15 ? n178 : n26;
  assign n1106 = pi14 ? n890 : n1105;
  assign n1107 = pi13 ? n1104 : n1106;
  assign n1108 = pi12 ? n1101 : n1107;
  assign n1109 = pi11 ? n1098 : n1108;
  assign n1110 = pi10 ? n1087 : n1109;
  assign n1111 = pi09 ? n1070 : n1110;
  assign n1112 = pi08 ? n1050 : n1111;
  assign n1113 = pi07 ? n1033 : n1112;
  assign n1114 = pi06 ? n1030 : n1113;
  assign n1115 = pi05 ? n921 : n1114;
  assign n1116 = pi14 ? n130 : n937;
  assign n1117 = pi16 ? n545 : n155;
  assign n1118 = pi15 ? n544 : n1117;
  assign n1119 = pi14 ? n924 : n1118;
  assign n1120 = pi13 ? n1116 : n1119;
  assign n1121 = pi12 ? n26 : n1120;
  assign n1122 = pi11 ? n26 : n1121;
  assign n1123 = pi15 ? n573 : n122;
  assign n1124 = pi14 ? n130 : n1123;
  assign n1125 = pi15 ? n100 : n60;
  assign n1126 = pi15 ? n493 : n961;
  assign n1127 = pi14 ? n1125 : n1126;
  assign n1128 = pi13 ? n1124 : n1127;
  assign n1129 = pi12 ? n26 : n1128;
  assign n1130 = pi16 ? n518 : n96;
  assign n1131 = pi15 ? n26 : n1130;
  assign n1132 = pi14 ? n1131 : n958;
  assign n1133 = pi13 ? n1132 : n950;
  assign n1134 = pi12 ? n26 : n1133;
  assign n1135 = pi11 ? n1129 : n1134;
  assign n1136 = pi10 ? n1122 : n1135;
  assign n1137 = pi09 ? n26 : n1136;
  assign n1138 = pi08 ? n26 : n1137;
  assign n1139 = pi15 ? n475 : n224;
  assign n1140 = pi14 ? n802 : n1139;
  assign n1141 = pi13 ? n1132 : n1140;
  assign n1142 = pi12 ? n26 : n1141;
  assign n1143 = pi17 ? n41 : n96;
  assign n1144 = pi16 ? n42 : n1143;
  assign n1145 = pi15 ? n26 : n1144;
  assign n1146 = pi14 ? n1145 : n958;
  assign n1147 = pi14 ? n960 : n1139;
  assign n1148 = pi13 ? n1146 : n1147;
  assign n1149 = pi12 ? n26 : n1148;
  assign n1150 = pi11 ? n1142 : n1149;
  assign n1151 = pi17 ? n53 : n96;
  assign n1152 = pi16 ? n26 : n1151;
  assign n1153 = pi15 ? n26 : n1152;
  assign n1154 = pi14 ? n1153 : n958;
  assign n1155 = pi15 ? n123 : n224;
  assign n1156 = pi16 ? n224 : n274;
  assign n1157 = pi15 ? n475 : n1156;
  assign n1158 = pi14 ? n1155 : n1157;
  assign n1159 = pi13 ? n1154 : n1158;
  assign n1160 = pi12 ? n26 : n1159;
  assign n1161 = pi17 ? n47 : n41;
  assign n1162 = pi16 ? n1161 : n121;
  assign n1163 = pi15 ? n1162 : n542;
  assign n1164 = pi14 ? n490 : n1163;
  assign n1165 = pi15 ? n493 : n464;
  assign n1166 = pi16 ? n255 : n155;
  assign n1167 = pi17 ? n155 : n677;
  assign n1168 = pi16 ? n1167 : n26;
  assign n1169 = pi15 ? n1166 : n1168;
  assign n1170 = pi14 ? n1165 : n1169;
  assign n1171 = pi13 ? n1164 : n1170;
  assign n1172 = pi12 ? n26 : n1171;
  assign n1173 = pi11 ? n1160 : n1172;
  assign n1174 = pi10 ? n1150 : n1173;
  assign n1175 = pi15 ? n997 : n32;
  assign n1176 = pi14 ? n26 : n1175;
  assign n1177 = pi15 ? n62 : n610;
  assign n1178 = pi14 ? n376 : n1177;
  assign n1179 = pi13 ? n1176 : n1178;
  assign n1180 = pi12 ? n26 : n1179;
  assign n1181 = pi11 ? n26 : n1180;
  assign n1182 = pi10 ? n26 : n1181;
  assign n1183 = pi09 ? n1174 : n1182;
  assign n1184 = pi15 ? n997 : n114;
  assign n1185 = pi14 ? n26 : n1184;
  assign n1186 = pi15 ? n438 : n48;
  assign n1187 = pi14 ? n1186 : n67;
  assign n1188 = pi13 ? n1185 : n1187;
  assign n1189 = pi12 ? n26 : n1188;
  assign n1190 = pi13 ? n1185 : n75;
  assign n1191 = pi12 ? n26 : n1190;
  assign n1192 = pi11 ? n1189 : n1191;
  assign n1193 = pi15 ? n438 : n364;
  assign n1194 = pi14 ? n1193 : n67;
  assign n1195 = pi13 ? n1185 : n1194;
  assign n1196 = pi12 ? n26 : n1195;
  assign n1197 = pi10 ? n1192 : n1196;
  assign n1198 = pi17 ? n175 : n41;
  assign n1199 = pi16 ? n476 : n1198;
  assign n1200 = pi15 ? n32 : n1199;
  assign n1201 = pi14 ? n26 : n1200;
  assign n1202 = pi15 ? n60 : n65;
  assign n1203 = pi14 ? n232 : n1202;
  assign n1204 = pi13 ? n1201 : n1203;
  assign n1205 = pi12 ? n26 : n1204;
  assign n1206 = pi15 ? n73 : n122;
  assign n1207 = pi14 ? n26 : n1206;
  assign n1208 = pi16 ? n290 : n60;
  assign n1209 = pi15 ? n100 : n1208;
  assign n1210 = pi15 ? n60 : n1117;
  assign n1211 = pi14 ? n1209 : n1210;
  assign n1212 = pi13 ? n1207 : n1211;
  assign n1213 = pi12 ? n26 : n1212;
  assign n1214 = pi11 ? n1205 : n1213;
  assign n1215 = pi17 ? n155 : n26;
  assign n1216 = pi16 ? n255 : n1215;
  assign n1217 = pi15 ? n546 : n1216;
  assign n1218 = pi14 ? n358 : n1217;
  assign n1219 = pi13 ? n959 : n1218;
  assign n1220 = pi12 ? n26 : n1219;
  assign n1221 = pi16 ? n175 : n26;
  assign n1222 = pi15 ? n464 : n1221;
  assign n1223 = pi14 ? n494 : n1222;
  assign n1224 = pi13 ? n971 : n1223;
  assign n1225 = pi12 ? n26 : n1224;
  assign n1226 = pi11 ? n1220 : n1225;
  assign n1227 = pi10 ? n1214 : n1226;
  assign n1228 = pi09 ? n1197 : n1227;
  assign n1229 = pi08 ? n1183 : n1228;
  assign n1230 = pi07 ? n1138 : n1229;
  assign n1231 = pi09 ? n1182 : n1197;
  assign n1232 = pi14 ? n365 : n1177;
  assign n1233 = pi13 ? n1176 : n1232;
  assign n1234 = pi12 ? n26 : n1233;
  assign n1235 = pi11 ? n26 : n1234;
  assign n1236 = pi10 ? n26 : n1235;
  assign n1237 = pi09 ? n1227 : n1236;
  assign n1238 = pi08 ? n1231 : n1237;
  assign n1239 = pi14 ? n26 : n408;
  assign n1240 = pi13 ? n1239 : n1194;
  assign n1241 = pi12 ? n26 : n1240;
  assign n1242 = pi11 ? n1196 : n1241;
  assign n1243 = pi14 ? n406 : n408;
  assign n1244 = pi13 ? n1243 : n1194;
  assign n1245 = pi12 ? n26 : n1244;
  assign n1246 = pi14 ? n294 : n408;
  assign n1247 = pi13 ? n1246 : n1194;
  assign n1248 = pi12 ? n26 : n1247;
  assign n1249 = pi11 ? n1245 : n1248;
  assign n1250 = pi10 ? n1242 : n1249;
  assign n1251 = pi15 ? n26 : n177;
  assign n1252 = pi15 ? n32 : n73;
  assign n1253 = pi14 ? n1251 : n1252;
  assign n1254 = pi14 ? n723 : n323;
  assign n1255 = pi13 ? n1253 : n1254;
  assign n1256 = pi12 ? n26 : n1255;
  assign n1257 = pi16 ? n1051 : n155;
  assign n1258 = pi15 ? n26 : n1257;
  assign n1259 = pi16 ? n476 : n96;
  assign n1260 = pi15 ? n32 : n1259;
  assign n1261 = pi14 ? n1258 : n1260;
  assign n1262 = pi16 ? n482 : n58;
  assign n1263 = pi15 ? n122 : n1262;
  assign n1264 = pi15 ? n60 : n546;
  assign n1265 = pi14 ? n1263 : n1264;
  assign n1266 = pi13 ? n1261 : n1265;
  assign n1267 = pi12 ? n26 : n1266;
  assign n1268 = pi11 ? n1256 : n1267;
  assign n1269 = pi15 ? n26 : n477;
  assign n1270 = pi14 ? n1269 : n205;
  assign n1271 = pi13 ? n1270 : n773;
  assign n1272 = pi12 ? n26 : n1271;
  assign n1273 = pi16 ? n1051 : n32;
  assign n1274 = pi15 ? n26 : n1273;
  assign n1275 = pi14 ? n1274 : n205;
  assign n1276 = pi13 ? n1275 : n776;
  assign n1277 = pi12 ? n26 : n1276;
  assign n1278 = pi11 ? n1272 : n1277;
  assign n1279 = pi10 ? n1268 : n1278;
  assign n1280 = pi09 ? n1250 : n1279;
  assign n1281 = pi16 ? n1051 : n962;
  assign n1282 = pi15 ? n26 : n1281;
  assign n1283 = pi14 ? n1282 : n205;
  assign n1284 = pi13 ? n1283 : n776;
  assign n1285 = pi12 ? n26 : n1284;
  assign n1286 = pi16 ? n175 : n962;
  assign n1287 = pi15 ? n26 : n1286;
  assign n1288 = pi14 ? n1287 : n205;
  assign n1289 = pi13 ? n1288 : n776;
  assign n1290 = pi12 ? n26 : n1289;
  assign n1291 = pi11 ? n1285 : n1290;
  assign n1292 = pi16 ? n156 : n175;
  assign n1293 = pi15 ? n405 : n1292;
  assign n1294 = pi14 ? n1293 : n205;
  assign n1295 = pi13 ? n1294 : n776;
  assign n1296 = pi12 ? n26 : n1295;
  assign n1297 = pi15 ? n293 : n157;
  assign n1298 = pi14 ? n1297 : n205;
  assign n1299 = pi13 ? n1298 : n776;
  assign n1300 = pi12 ? n26 : n1299;
  assign n1301 = pi11 ? n1296 : n1300;
  assign n1302 = pi10 ? n1291 : n1301;
  assign n1303 = pi15 ? n177 : n32;
  assign n1304 = pi14 ? n1303 : n205;
  assign n1305 = pi14 ? n658 : n224;
  assign n1306 = pi13 ? n1304 : n1305;
  assign n1307 = pi12 ? n26 : n1306;
  assign n1308 = pi13 ? n26 : n632;
  assign n1309 = pi15 ? n678 : n480;
  assign n1310 = pi14 ? n1309 : n1102;
  assign n1311 = pi14 ? n101 : n890;
  assign n1312 = pi13 ? n1310 : n1311;
  assign n1313 = pi12 ? n1308 : n1312;
  assign n1314 = pi11 ? n1307 : n1313;
  assign n1315 = pi13 ? n26 : n384;
  assign n1316 = pi14 ? n685 : n723;
  assign n1317 = pi15 ? n544 : n771;
  assign n1318 = pi15 ? n224 : n972;
  assign n1319 = pi14 ? n1317 : n1318;
  assign n1320 = pi13 ? n1316 : n1319;
  assign n1321 = pi12 ? n1315 : n1320;
  assign n1322 = pi17 ? n107 : n41;
  assign n1323 = pi16 ? n1322 : n41;
  assign n1324 = pi15 ? n1323 : n229;
  assign n1325 = pi15 ? n542 : n493;
  assign n1326 = pi14 ? n1324 : n1325;
  assign n1327 = pi16 ? n238 : n528;
  assign n1328 = pi15 ? n1327 : n26;
  assign n1329 = pi14 ? n840 : n1328;
  assign n1330 = pi13 ? n1326 : n1329;
  assign n1331 = pi12 ? n1101 : n1330;
  assign n1332 = pi11 ? n1321 : n1331;
  assign n1333 = pi10 ? n1314 : n1332;
  assign n1334 = pi09 ? n1302 : n1333;
  assign n1335 = pi08 ? n1280 : n1334;
  assign n1336 = pi07 ? n1238 : n1335;
  assign n1337 = pi06 ? n1230 : n1336;
  assign n1338 = pi14 ? n1269 : n1206;
  assign n1339 = pi16 ? n53 : n121;
  assign n1340 = pi15 ? n1339 : n123;
  assign n1341 = pi14 ? n1340 : n1210;
  assign n1342 = pi13 ? n1338 : n1341;
  assign n1343 = pi12 ? n26 : n1342;
  assign n1344 = pi11 ? n26 : n1343;
  assign n1345 = pi16 ? n41 : n72;
  assign n1346 = pi15 ? n1345 : n122;
  assign n1347 = pi14 ? n115 : n1346;
  assign n1348 = pi15 ? n546 : n1166;
  assign n1349 = pi14 ? n378 : n1348;
  assign n1350 = pi13 ? n1347 : n1349;
  assign n1351 = pi12 ? n26 : n1350;
  assign n1352 = pi14 ? n115 : n958;
  assign n1353 = pi15 ? n224 : n1166;
  assign n1354 = pi14 ? n802 : n1353;
  assign n1355 = pi13 ? n1352 : n1354;
  assign n1356 = pi12 ? n26 : n1355;
  assign n1357 = pi11 ? n1351 : n1356;
  assign n1358 = pi10 ? n1344 : n1357;
  assign n1359 = pi09 ? n26 : n1358;
  assign n1360 = pi08 ? n26 : n1359;
  assign n1361 = pi15 ? n26 : n554;
  assign n1362 = pi14 ? n1361 : n958;
  assign n1363 = pi13 ? n1362 : n1147;
  assign n1364 = pi12 ? n26 : n1363;
  assign n1365 = pi14 ? n608 : n958;
  assign n1366 = pi17 ? n224 : n355;
  assign n1367 = pi16 ? n461 : n1366;
  assign n1368 = pi15 ? n475 : n1367;
  assign n1369 = pi14 ? n1155 : n1368;
  assign n1370 = pi13 ? n1365 : n1369;
  assign n1371 = pi12 ? n26 : n1370;
  assign n1372 = pi11 ? n1364 : n1371;
  assign n1373 = pi15 ? n489 : n385;
  assign n1374 = pi15 ? n41 : n432;
  assign n1375 = pi14 ? n1373 : n1374;
  assign n1376 = pi16 ? n461 : n274;
  assign n1377 = pi15 ? n475 : n1376;
  assign n1378 = pi14 ? n899 : n1377;
  assign n1379 = pi13 ? n1375 : n1378;
  assign n1380 = pi12 ? n26 : n1379;
  assign n1381 = pi16 ? n1161 : n1151;
  assign n1382 = pi15 ? n489 : n1381;
  assign n1383 = pi14 ? n1382 : n543;
  assign n1384 = pi16 ? n1215 : n26;
  assign n1385 = pi15 ? n475 : n1384;
  assign n1386 = pi14 ? n494 : n1385;
  assign n1387 = pi13 ? n1383 : n1386;
  assign n1388 = pi12 ? n26 : n1387;
  assign n1389 = pi11 ? n1380 : n1388;
  assign n1390 = pi10 ? n1372 : n1389;
  assign n1391 = pi15 ? n73 : n133;
  assign n1392 = pi14 ? n656 : n1391;
  assign n1393 = pi15 ? n123 : n771;
  assign n1394 = pi14 ? n315 : n1393;
  assign n1395 = pi13 ? n1392 : n1394;
  assign n1396 = pi12 ? n26 : n1395;
  assign n1397 = pi11 ? n26 : n1396;
  assign n1398 = pi10 ? n26 : n1397;
  assign n1399 = pi09 ? n1390 : n1398;
  assign n1400 = pi15 ? n73 : n333;
  assign n1401 = pi14 ? n656 : n1400;
  assign n1402 = pi16 ? n740 : n355;
  assign n1403 = pi15 ? n123 : n1402;
  assign n1404 = pi14 ? n365 : n1403;
  assign n1405 = pi13 ? n1401 : n1404;
  assign n1406 = pi12 ? n26 : n1405;
  assign n1407 = pi14 ? n656 : n398;
  assign n1408 = pi13 ? n1407 : n359;
  assign n1409 = pi12 ? n26 : n1408;
  assign n1410 = pi11 ? n1406 : n1409;
  assign n1411 = pi15 ? n41 : n979;
  assign n1412 = pi15 ? n60 : n357;
  assign n1413 = pi14 ? n1411 : n1412;
  assign n1414 = pi13 ? n1407 : n1413;
  assign n1415 = pi12 ? n26 : n1414;
  assign n1416 = pi14 ? n137 : n1412;
  assign n1417 = pi13 ? n1407 : n1416;
  assign n1418 = pi12 ? n26 : n1417;
  assign n1419 = pi11 ? n1415 : n1418;
  assign n1420 = pi10 ? n1410 : n1419;
  assign n1421 = pi14 ? n656 : n990;
  assign n1422 = pi14 ? n993 : n1412;
  assign n1423 = pi13 ? n1421 : n1422;
  assign n1424 = pi12 ? n26 : n1423;
  assign n1425 = pi14 ? n553 : n1206;
  assign n1426 = pi15 ? n62 : n1208;
  assign n1427 = pi16 ? n355 : n1366;
  assign n1428 = pi15 ? n60 : n1427;
  assign n1429 = pi14 ? n1426 : n1428;
  assign n1430 = pi13 ? n1425 : n1429;
  assign n1431 = pi12 ? n26 : n1430;
  assign n1432 = pi11 ? n1424 : n1431;
  assign n1433 = pi14 ? n553 : n1374;
  assign n1434 = pi16 ? n740 : n356;
  assign n1435 = pi15 ? n60 : n1434;
  assign n1436 = pi15 ? n1064 : n1156;
  assign n1437 = pi14 ? n1435 : n1436;
  assign n1438 = pi13 ? n1433 : n1437;
  assign n1439 = pi12 ? n26 : n1438;
  assign n1440 = pi14 ? n26 : n543;
  assign n1441 = pi15 ? n1064 : n1384;
  assign n1442 = pi14 ? n494 : n1441;
  assign n1443 = pi13 ? n1440 : n1442;
  assign n1444 = pi12 ? n26 : n1443;
  assign n1445 = pi11 ? n1439 : n1444;
  assign n1446 = pi10 ? n1432 : n1445;
  assign n1447 = pi09 ? n1420 : n1446;
  assign n1448 = pi08 ? n1399 : n1447;
  assign n1449 = pi07 ? n1360 : n1448;
  assign n1450 = pi09 ? n1398 : n1420;
  assign n1451 = pi15 ? n258 : n722;
  assign n1452 = pi14 ? n1451 : n910;
  assign n1453 = pi13 ? n1392 : n1452;
  assign n1454 = pi12 ? n26 : n1453;
  assign n1455 = pi11 ? n26 : n1454;
  assign n1456 = pi10 ? n26 : n1455;
  assign n1457 = pi09 ? n1446 : n1456;
  assign n1458 = pi08 ? n1450 : n1457;
  assign n1459 = pi15 ? n60 : n1402;
  assign n1460 = pi14 ? n1451 : n1459;
  assign n1461 = pi13 ? n1401 : n1460;
  assign n1462 = pi12 ? n26 : n1461;
  assign n1463 = pi14 ? n144 : n398;
  assign n1464 = pi14 ? n1451 : n1412;
  assign n1465 = pi13 ? n1463 : n1464;
  assign n1466 = pi12 ? n26 : n1465;
  assign n1467 = pi11 ? n1462 : n1466;
  assign n1468 = pi14 ? n395 : n398;
  assign n1469 = pi13 ? n1468 : n1464;
  assign n1470 = pi12 ? n26 : n1469;
  assign n1471 = pi14 ? n383 : n398;
  assign n1472 = pi14 ? n723 : n1412;
  assign n1473 = pi13 ? n1471 : n1472;
  assign n1474 = pi12 ? n26 : n1473;
  assign n1475 = pi11 ? n1470 : n1474;
  assign n1476 = pi10 ? n1467 : n1475;
  assign n1477 = pi14 ? n615 : n990;
  assign n1478 = pi13 ? n1477 : n1472;
  assign n1479 = pi12 ? n26 : n1478;
  assign n1480 = pi15 ? n26 : n178;
  assign n1481 = pi15 ? n73 : n989;
  assign n1482 = pi14 ? n1480 : n1481;
  assign n1483 = pi14 ? n723 : n926;
  assign n1484 = pi13 ? n1482 : n1483;
  assign n1485 = pi12 ? n26 : n1484;
  assign n1486 = pi11 ? n1479 : n1485;
  assign n1487 = pi14 ? n105 : n190;
  assign n1488 = pi14 ? n770 : n494;
  assign n1489 = pi13 ? n1487 : n1488;
  assign n1490 = pi12 ? n26 : n1489;
  assign n1491 = pi15 ? n43 : n178;
  assign n1492 = pi14 ? n1491 : n190;
  assign n1493 = pi16 ? n60 : n461;
  assign n1494 = pi15 ? n1493 : n546;
  assign n1495 = pi14 ? n770 : n1494;
  assign n1496 = pi13 ? n1492 : n1495;
  assign n1497 = pi12 ? n26 : n1496;
  assign n1498 = pi11 ? n1490 : n1497;
  assign n1499 = pi10 ? n1486 : n1498;
  assign n1500 = pi09 ? n1476 : n1499;
  assign n1501 = pi17 ? n175 : n1072;
  assign n1502 = pi16 ? n1501 : n32;
  assign n1503 = pi15 ? n43 : n1502;
  assign n1504 = pi14 ? n1503 : n190;
  assign n1505 = pi13 ? n1504 : n1495;
  assign n1506 = pi12 ? n26 : n1505;
  assign n1507 = pi16 ? n26 : n563;
  assign n1508 = pi15 ? n1507 : n1073;
  assign n1509 = pi14 ? n1508 : n190;
  assign n1510 = pi17 ? n65 : n224;
  assign n1511 = pi16 ? n1510 : n461;
  assign n1512 = pi15 ? n1511 : n546;
  assign n1513 = pi14 ? n770 : n1512;
  assign n1514 = pi13 ? n1509 : n1513;
  assign n1515 = pi12 ? n26 : n1514;
  assign n1516 = pi11 ? n1506 : n1515;
  assign n1517 = pi17 ? n96 : n155;
  assign n1518 = pi16 ? n26 : n1517;
  assign n1519 = pi17 ? n32 : n1072;
  assign n1520 = pi16 ? n1519 : n32;
  assign n1521 = pi15 ? n1518 : n1520;
  assign n1522 = pi14 ? n1521 : n190;
  assign n1523 = pi13 ? n1522 : n940;
  assign n1524 = pi12 ? n26 : n1523;
  assign n1525 = pi16 ? n33 : n461;
  assign n1526 = pi15 ? n1525 : n808;
  assign n1527 = pi14 ? n1526 : n190;
  assign n1528 = pi13 ? n1527 : n940;
  assign n1529 = pi12 ? n26 : n1528;
  assign n1530 = pi11 ? n1524 : n1529;
  assign n1531 = pi10 ? n1516 : n1530;
  assign n1532 = pi15 ? n382 : n32;
  assign n1533 = pi15 ? n1345 : n41;
  assign n1534 = pi14 ? n1532 : n1533;
  assign n1535 = pi15 ? n961 : n546;
  assign n1536 = pi14 ? n658 : n1535;
  assign n1537 = pi13 ? n1534 : n1536;
  assign n1538 = pi12 ? n26 : n1537;
  assign n1539 = pi13 ? n26 : n407;
  assign n1540 = pi14 ? n454 : n1102;
  assign n1541 = pi16 ? n545 : n1215;
  assign n1542 = pi15 ? n961 : n1541;
  assign n1543 = pi14 ? n873 : n1542;
  assign n1544 = pi13 ? n1540 : n1543;
  assign n1545 = pi12 ? n1539 : n1544;
  assign n1546 = pi11 ? n1538 : n1545;
  assign n1547 = pi13 ? n26 : n396;
  assign n1548 = pi15 ? n573 : n133;
  assign n1549 = pi16 ? n41 : n968;
  assign n1550 = pi15 ? n1549 : n722;
  assign n1551 = pi14 ? n1548 : n1550;
  assign n1552 = pi15 ? n961 : n1221;
  assign n1553 = pi14 ? n1317 : n1552;
  assign n1554 = pi13 ? n1551 : n1553;
  assign n1555 = pi12 ? n1547 : n1554;
  assign n1556 = pi16 ? n33 : n186;
  assign n1557 = pi15 ? n26 : n1556;
  assign n1558 = pi14 ? n26 : n1557;
  assign n1559 = pi13 ? n26 : n1558;
  assign n1560 = pi16 ? n1322 : n146;
  assign n1561 = pi15 ? n1560 : n133;
  assign n1562 = pi15 ? n122 : n377;
  assign n1563 = pi14 ? n1561 : n1562;
  assign n1564 = pi16 ? n255 : n224;
  assign n1565 = pi15 ? n1564 : n26;
  assign n1566 = pi14 ? n494 : n1565;
  assign n1567 = pi13 ? n1563 : n1566;
  assign n1568 = pi12 ? n1559 : n1567;
  assign n1569 = pi11 ? n1555 : n1568;
  assign n1570 = pi10 ? n1546 : n1569;
  assign n1571 = pi09 ? n1531 : n1570;
  assign n1572 = pi08 ? n1500 : n1571;
  assign n1573 = pi07 ? n1458 : n1572;
  assign n1574 = pi06 ? n1449 : n1573;
  assign n1575 = pi05 ? n1337 : n1574;
  assign n1576 = pi04 ? n1115 : n1575;
  assign n1577 = pi14 ? n105 : n1206;
  assign n1578 = pi14 ? n101 : n1210;
  assign n1579 = pi13 ? n1577 : n1578;
  assign n1580 = pi12 ? n26 : n1579;
  assign n1581 = pi11 ? n26 : n1580;
  assign n1582 = pi14 ? n105 : n1346;
  assign n1583 = pi15 ? n493 : n475;
  assign n1584 = pi14 ? n101 : n1583;
  assign n1585 = pi13 ? n1582 : n1584;
  assign n1586 = pi12 ? n26 : n1585;
  assign n1587 = pi15 ? n552 : n32;
  assign n1588 = pi14 ? n1587 : n958;
  assign n1589 = pi17 ? n355 : n32;
  assign n1590 = pi16 ? n1589 : n155;
  assign n1591 = pi15 ? n464 : n1590;
  assign n1592 = pi14 ? n523 : n1591;
  assign n1593 = pi13 ? n1588 : n1592;
  assign n1594 = pi12 ? n26 : n1593;
  assign n1595 = pi11 ? n1586 : n1594;
  assign n1596 = pi10 ? n1581 : n1595;
  assign n1597 = pi09 ? n26 : n1596;
  assign n1598 = pi08 ? n26 : n1597;
  assign n1599 = pi15 ? n552 : n554;
  assign n1600 = pi14 ? n1599 : n1374;
  assign n1601 = pi15 ? n224 : n961;
  assign n1602 = pi14 ? n910 : n1601;
  assign n1603 = pi13 ? n1600 : n1602;
  assign n1604 = pi12 ? n26 : n1603;
  assign n1605 = pi15 ? n598 : n96;
  assign n1606 = pi16 ? n1161 : n58;
  assign n1607 = pi15 ? n41 : n1606;
  assign n1608 = pi14 ? n1605 : n1607;
  assign n1609 = pi16 ? n212 : n274;
  assign n1610 = pi15 ? n224 : n1609;
  assign n1611 = pi14 ? n899 : n1610;
  assign n1612 = pi13 ? n1608 : n1611;
  assign n1613 = pi12 ? n26 : n1612;
  assign n1614 = pi11 ? n1604 : n1613;
  assign n1615 = pi15 ? n598 : n385;
  assign n1616 = pi15 ? n122 : n432;
  assign n1617 = pi14 ? n1615 : n1616;
  assign n1618 = pi15 ? n475 : n1221;
  assign n1619 = pi14 ? n899 : n1618;
  assign n1620 = pi13 ? n1617 : n1619;
  assign n1621 = pi12 ? n26 : n1620;
  assign n1622 = pi16 ? n41 : n1143;
  assign n1623 = pi15 ? n906 : n1622;
  assign n1624 = pi14 ? n1623 : n543;
  assign n1625 = pi15 ? n1166 : n1384;
  assign n1626 = pi14 ? n494 : n1625;
  assign n1627 = pi13 ? n1624 : n1626;
  assign n1628 = pi12 ? n26 : n1627;
  assign n1629 = pi11 ? n1621 : n1628;
  assign n1630 = pi10 ? n1614 : n1629;
  assign n1631 = pi15 ? n43 : n96;
  assign n1632 = pi14 ? n144 : n1631;
  assign n1633 = pi16 ? n60 : n26;
  assign n1634 = pi15 ? n1633 : n250;
  assign n1635 = pi14 ? n387 : n1634;
  assign n1636 = pi13 ? n1632 : n1635;
  assign n1637 = pi12 ? n26 : n1636;
  assign n1638 = pi11 ? n26 : n1637;
  assign n1639 = pi10 ? n26 : n1638;
  assign n1640 = pi09 ? n1630 : n1639;
  assign n1641 = pi15 ? n41 : n96;
  assign n1642 = pi14 ? n144 : n1641;
  assign n1643 = pi14 ? n137 : n494;
  assign n1644 = pi13 ? n1642 : n1643;
  assign n1645 = pi12 ? n26 : n1644;
  assign n1646 = pi14 ? n387 : n494;
  assign n1647 = pi13 ? n1642 : n1646;
  assign n1648 = pi12 ? n26 : n1647;
  assign n1649 = pi11 ? n1645 : n1648;
  assign n1650 = pi14 ? n124 : n494;
  assign n1651 = pi13 ? n1642 : n1650;
  assign n1652 = pi12 ? n26 : n1651;
  assign n1653 = pi15 ? n41 : n229;
  assign n1654 = pi14 ? n144 : n1653;
  assign n1655 = pi14 ? n232 : n494;
  assign n1656 = pi13 ? n1654 : n1655;
  assign n1657 = pi12 ? n26 : n1656;
  assign n1658 = pi11 ? n1652 : n1657;
  assign n1659 = pi10 ? n1649 : n1658;
  assign n1660 = pi14 ? n144 : n41;
  assign n1661 = pi16 ? n53 : n65;
  assign n1662 = pi15 ? n1661 : n66;
  assign n1663 = pi14 ? n1662 : n494;
  assign n1664 = pi13 ? n1660 : n1663;
  assign n1665 = pi12 ? n26 : n1664;
  assign n1666 = pi15 ? n26 : n1507;
  assign n1667 = pi14 ? n1666 : n958;
  assign n1668 = pi15 ? n493 : n1156;
  assign n1669 = pi14 ? n67 : n1668;
  assign n1670 = pi13 ? n1667 : n1669;
  assign n1671 = pi12 ? n26 : n1670;
  assign n1672 = pi11 ? n1665 : n1671;
  assign n1673 = pi15 ? n26 : n598;
  assign n1674 = pi14 ? n1673 : n1374;
  assign n1675 = pi16 ? n224 : n26;
  assign n1676 = pi15 ? n224 : n1675;
  assign n1677 = pi14 ? n910 : n1676;
  assign n1678 = pi13 ? n1674 : n1677;
  assign n1679 = pi12 ? n26 : n1678;
  assign n1680 = pi14 ? n553 : n543;
  assign n1681 = pi15 ? n224 : n1384;
  assign n1682 = pi14 ? n1634 : n1681;
  assign n1683 = pi13 ? n1680 : n1682;
  assign n1684 = pi12 ? n26 : n1683;
  assign n1685 = pi11 ? n1679 : n1684;
  assign n1686 = pi10 ? n1672 : n1685;
  assign n1687 = pi09 ? n1659 : n1686;
  assign n1688 = pi08 ? n1640 : n1687;
  assign n1689 = pi07 ? n1598 : n1688;
  assign n1690 = pi09 ? n1639 : n1659;
  assign n1691 = pi14 ? n723 : n1634;
  assign n1692 = pi13 ? n1632 : n1691;
  assign n1693 = pi12 ? n26 : n1692;
  assign n1694 = pi11 ? n26 : n1693;
  assign n1695 = pi10 ? n26 : n1694;
  assign n1696 = pi09 ? n1686 : n1695;
  assign n1697 = pi08 ? n1690 : n1696;
  assign n1698 = pi14 ? n723 : n494;
  assign n1699 = pi13 ? n1642 : n1698;
  assign n1700 = pi12 ? n26 : n1699;
  assign n1701 = pi14 ? n130 : n1641;
  assign n1702 = pi13 ? n1701 : n1698;
  assign n1703 = pi12 ? n26 : n1702;
  assign n1704 = pi11 ? n1700 : n1703;
  assign n1705 = pi14 ? n383 : n1641;
  assign n1706 = pi13 ? n1705 : n1698;
  assign n1707 = pi12 ? n26 : n1706;
  assign n1708 = pi16 ? n1501 : n186;
  assign n1709 = pi15 ? n26 : n1708;
  assign n1710 = pi14 ? n1709 : n1653;
  assign n1711 = pi13 ? n1710 : n1698;
  assign n1712 = pi12 ? n26 : n1711;
  assign n1713 = pi11 ? n1707 : n1712;
  assign n1714 = pi10 ? n1704 : n1713;
  assign n1715 = pi15 ? n26 : n1520;
  assign n1716 = pi14 ? n1715 : n41;
  assign n1717 = pi13 ? n1716 : n1698;
  assign n1718 = pi12 ? n26 : n1717;
  assign n1719 = pi15 ? n87 : n808;
  assign n1720 = pi14 ? n1719 : n41;
  assign n1721 = pi14 ? n723 : n1583;
  assign n1722 = pi13 ? n1720 : n1721;
  assign n1723 = pi12 ? n26 : n1722;
  assign n1724 = pi11 ? n1718 : n1723;
  assign n1725 = pi14 ? n88 : n1653;
  assign n1726 = pi15 ? n493 : n1166;
  assign n1727 = pi14 ? n723 : n1726;
  assign n1728 = pi13 ? n1725 : n1727;
  assign n1729 = pi12 ? n26 : n1728;
  assign n1730 = pi13 ? n1725 : n1698;
  assign n1731 = pi12 ? n26 : n1730;
  assign n1732 = pi11 ? n1729 : n1731;
  assign n1733 = pi10 ? n1724 : n1732;
  assign n1734 = pi09 ? n1714 : n1733;
  assign n1735 = pi16 ? n1510 : n155;
  assign n1736 = pi15 ? n1735 : n224;
  assign n1737 = pi14 ? n924 : n1736;
  assign n1738 = pi13 ? n1725 : n1737;
  assign n1739 = pi12 ? n26 : n1738;
  assign n1740 = pi15 ? n87 : n1073;
  assign n1741 = pi14 ? n1740 : n1653;
  assign n1742 = pi14 ? n924 : n1139;
  assign n1743 = pi13 ? n1741 : n1742;
  assign n1744 = pi12 ? n26 : n1743;
  assign n1745 = pi11 ? n1739 : n1744;
  assign n1746 = pi15 ? n81 : n1073;
  assign n1747 = pi14 ? n1746 : n1653;
  assign n1748 = pi14 ? n770 : n1139;
  assign n1749 = pi13 ? n1747 : n1748;
  assign n1750 = pi12 ? n26 : n1749;
  assign n1751 = pi14 ? n35 : n1653;
  assign n1752 = pi14 ? n1562 : n1139;
  assign n1753 = pi13 ? n1751 : n1752;
  assign n1754 = pi12 ? n26 : n1753;
  assign n1755 = pi11 ? n1750 : n1754;
  assign n1756 = pi10 ? n1745 : n1755;
  assign n1757 = pi14 ? n1532 : n41;
  assign n1758 = pi16 ? n224 : n1366;
  assign n1759 = pi15 ? n475 : n1758;
  assign n1760 = pi14 ? n802 : n1759;
  assign n1761 = pi13 ? n1757 : n1760;
  assign n1762 = pi12 ? n26 : n1761;
  assign n1763 = pi15 ? n477 : n32;
  assign n1764 = pi14 ? n1763 : n958;
  assign n1765 = pi15 ? n854 : n771;
  assign n1766 = pi14 ? n1765 : n1157;
  assign n1767 = pi13 ? n1764 : n1766;
  assign n1768 = pi12 ? n26 : n1767;
  assign n1769 = pi11 ? n1762 : n1768;
  assign n1770 = pi13 ? n26 : n145;
  assign n1771 = pi14 ? n134 : n1550;
  assign n1772 = pi14 ? n910 : n1385;
  assign n1773 = pi13 ? n1771 : n1772;
  assign n1774 = pi12 ? n1770 : n1773;
  assign n1775 = pi16 ? n128 : n186;
  assign n1776 = pi15 ? n26 : n1775;
  assign n1777 = pi14 ? n26 : n1776;
  assign n1778 = pi13 ? n26 : n1777;
  assign n1779 = pi15 ? n122 : n483;
  assign n1780 = pi14 ? n1631 : n1779;
  assign n1781 = pi15 ? n1633 : n689;
  assign n1782 = pi15 ? n475 : n26;
  assign n1783 = pi14 ? n1781 : n1782;
  assign n1784 = pi13 ? n1780 : n1783;
  assign n1785 = pi12 ? n1778 : n1784;
  assign n1786 = pi11 ? n1774 : n1785;
  assign n1787 = pi10 ? n1769 : n1786;
  assign n1788 = pi09 ? n1756 : n1787;
  assign n1789 = pi08 ? n1734 : n1788;
  assign n1790 = pi07 ? n1697 : n1789;
  assign n1791 = pi06 ? n1689 : n1790;
  assign n1792 = pi15 ? n438 : n122;
  assign n1793 = pi14 ? n88 : n1792;
  assign n1794 = pi13 ? n1793 : n1578;
  assign n1795 = pi12 ? n26 : n1794;
  assign n1796 = pi11 ? n26 : n1795;
  assign n1797 = pi14 ? n88 : n958;
  assign n1798 = pi14 ? n101 : n1726;
  assign n1799 = pi13 ? n1797 : n1798;
  assign n1800 = pi12 ? n26 : n1799;
  assign n1801 = pi15 ? n598 : n32;
  assign n1802 = pi14 ? n1801 : n958;
  assign n1803 = pi16 ? n290 : n224;
  assign n1804 = pi15 ? n100 : n1803;
  assign n1805 = pi14 ? n1804 : n890;
  assign n1806 = pi13 ? n1802 : n1805;
  assign n1807 = pi12 ? n26 : n1806;
  assign n1808 = pi11 ? n1800 : n1807;
  assign n1809 = pi10 ? n1796 : n1808;
  assign n1810 = pi09 ? n26 : n1809;
  assign n1811 = pi08 ? n26 : n1810;
  assign n1812 = pi14 ? n1801 : n1374;
  assign n1813 = pi17 ? n155 : n355;
  assign n1814 = pi16 ? n255 : n1813;
  assign n1815 = pi15 ? n475 : n1814;
  assign n1816 = pi14 ? n910 : n1815;
  assign n1817 = pi13 ? n1812 : n1816;
  assign n1818 = pi12 ? n26 : n1817;
  assign n1819 = pi15 ? n519 : n554;
  assign n1820 = pi15 ? n41 : n542;
  assign n1821 = pi14 ? n1819 : n1820;
  assign n1822 = pi16 ? n1051 : n274;
  assign n1823 = pi15 ? n475 : n1822;
  assign n1824 = pi14 ? n899 : n1823;
  assign n1825 = pi13 ? n1821 : n1824;
  assign n1826 = pi12 ? n26 : n1825;
  assign n1827 = pi11 ? n1818 : n1826;
  assign n1828 = pi15 ? n1130 : n41;
  assign n1829 = pi14 ? n1828 : n1616;
  assign n1830 = pi17 ? n175 : n224;
  assign n1831 = pi16 ? n1830 : n26;
  assign n1832 = pi15 ? n475 : n1831;
  assign n1833 = pi14 ? n899 : n1832;
  assign n1834 = pi13 ? n1829 : n1833;
  assign n1835 = pi12 ? n26 : n1834;
  assign n1836 = pi16 ? n41 : n132;
  assign n1837 = pi15 ? n96 : n1836;
  assign n1838 = pi14 ? n1837 : n543;
  assign n1839 = pi13 ? n1838 : n1386;
  assign n1840 = pi12 ? n26 : n1839;
  assign n1841 = pi11 ? n1835 : n1840;
  assign n1842 = pi10 ? n1827 : n1841;
  assign n1843 = pi09 ? n1842 : n26;
  assign n1844 = pi08 ? n1843 : n26;
  assign n1845 = pi07 ? n1811 : n1844;
  assign n1846 = pi06 ? n1845 : n26;
  assign n1847 = pi05 ? n1791 : n1846;
  assign n1848 = pi14 ? n101 : n1264;
  assign n1849 = pi13 ? n1793 : n1848;
  assign n1850 = pi12 ? n26 : n1849;
  assign n1851 = pi11 ? n26 : n1850;
  assign n1852 = pi15 ? n546 : n475;
  assign n1853 = pi14 ? n101 : n1852;
  assign n1854 = pi13 ? n1797 : n1853;
  assign n1855 = pi12 ? n26 : n1854;
  assign n1856 = pi14 ? n82 : n958;
  assign n1857 = pi13 ? n1856 : n1354;
  assign n1858 = pi12 ? n26 : n1857;
  assign n1859 = pi11 ? n1855 : n1858;
  assign n1860 = pi10 ? n1851 : n1859;
  assign n1861 = pi09 ? n26 : n1860;
  assign n1862 = pi08 ? n26 : n1861;
  assign n1863 = pi14 ? n82 : n1374;
  assign n1864 = pi15 ? n224 : n1814;
  assign n1865 = pi14 ? n910 : n1864;
  assign n1866 = pi13 ? n1863 : n1865;
  assign n1867 = pi12 ? n26 : n1866;
  assign n1868 = pi15 ? n579 : n480;
  assign n1869 = pi14 ? n1868 : n1820;
  assign n1870 = pi16 ? n175 : n274;
  assign n1871 = pi15 ? n224 : n1870;
  assign n1872 = pi14 ? n899 : n1871;
  assign n1873 = pi13 ? n1869 : n1872;
  assign n1874 = pi12 ? n26 : n1873;
  assign n1875 = pi11 ? n1867 : n1874;
  assign n1876 = pi14 ? n790 : n1616;
  assign n1877 = pi13 ? n1876 : n1833;
  assign n1878 = pi12 ? n26 : n1877;
  assign n1879 = pi14 ? n26 : n553;
  assign n1880 = pi13 ? n26 : n1879;
  assign n1881 = pi14 ? n41 : n543;
  assign n1882 = pi13 ? n1881 : n1386;
  assign n1883 = pi12 ? n1880 : n1882;
  assign n1884 = pi11 ? n1878 : n1883;
  assign n1885 = pi10 ? n1875 : n1884;
  assign n1886 = pi09 ? n1885 : n26;
  assign n1887 = pi08 ? n1886 : n26;
  assign n1888 = pi07 ? n1862 : n1887;
  assign n1889 = pi06 ? n1888 : n26;
  assign n1890 = pi14 ? n82 : n1792;
  assign n1891 = pi13 ? n1890 : n1578;
  assign n1892 = pi12 ? n26 : n1891;
  assign n1893 = pi11 ? n26 : n1892;
  assign n1894 = pi13 ? n1856 : n1584;
  assign n1895 = pi12 ? n26 : n1894;
  assign n1896 = pi15 ? n579 : n32;
  assign n1897 = pi14 ? n1896 : n958;
  assign n1898 = pi15 ? n224 : n1117;
  assign n1899 = pi14 ? n960 : n1898;
  assign n1900 = pi13 ? n1897 : n1899;
  assign n1901 = pi12 ? n26 : n1900;
  assign n1902 = pi11 ? n1895 : n1901;
  assign n1903 = pi10 ? n1893 : n1902;
  assign n1904 = pi09 ? n26 : n1903;
  assign n1905 = pi08 ? n26 : n1904;
  assign n1906 = pi14 ? n1896 : n1374;
  assign n1907 = pi13 ? n1906 : n1865;
  assign n1908 = pi12 ? n26 : n1907;
  assign n1909 = pi15 ? n554 : n480;
  assign n1910 = pi14 ? n1909 : n1820;
  assign n1911 = pi16 ? n238 : n274;
  assign n1912 = pi15 ? n224 : n1911;
  assign n1913 = pi14 ? n899 : n1912;
  assign n1914 = pi13 ? n1910 : n1913;
  assign n1915 = pi12 ? n26 : n1914;
  assign n1916 = pi11 ? n1908 : n1915;
  assign n1917 = pi14 ? n783 : n1616;
  assign n1918 = pi13 ? n1917 : n1833;
  assign n1919 = pi12 ? n1880 : n1918;
  assign n1920 = pi14 ? n26 : n935;
  assign n1921 = pi13 ? n26 : n1920;
  assign n1922 = pi12 ? n1921 : n1882;
  assign n1923 = pi11 ? n1919 : n1922;
  assign n1924 = pi10 ? n1916 : n1923;
  assign n1925 = pi14 ? n26 : n1131;
  assign n1926 = pi13 ? n26 : n1925;
  assign n1927 = pi15 ? n41 : n258;
  assign n1928 = pi15 ? n722 : n493;
  assign n1929 = pi14 ? n1927 : n1928;
  assign n1930 = pi17 ? n1072 : n32;
  assign n1931 = pi16 ? n1930 : n300;
  assign n1932 = pi15 ? n1931 : n26;
  assign n1933 = pi14 ? n840 : n1932;
  assign n1934 = pi13 ? n1929 : n1933;
  assign n1935 = pi12 ? n1926 : n1934;
  assign n1936 = pi14 ? n543 : n494;
  assign n1937 = pi16 ? n1167 : n32;
  assign n1938 = pi15 ? n464 : n1937;
  assign n1939 = pi14 ? n1938 : n26;
  assign n1940 = pi13 ? n1936 : n1939;
  assign n1941 = pi12 ? n1926 : n1940;
  assign n1942 = pi11 ? n1935 : n1941;
  assign n1943 = pi16 ? n1051 : n300;
  assign n1944 = pi15 ? n475 : n1943;
  assign n1945 = pi14 ? n1944 : n26;
  assign n1946 = pi13 ? n1936 : n1945;
  assign n1947 = pi12 ? n1926 : n1946;
  assign n1948 = pi14 ? n1618 : n26;
  assign n1949 = pi13 ? n1936 : n1948;
  assign n1950 = pi12 ? n1926 : n1949;
  assign n1951 = pi11 ? n1947 : n1950;
  assign n1952 = pi10 ? n1942 : n1951;
  assign n1953 = pi09 ? n1924 : n1952;
  assign n1954 = pi14 ? n1681 : n26;
  assign n1955 = pi13 ? n1936 : n1954;
  assign n1956 = pi12 ? n1926 : n1955;
  assign n1957 = pi08 ? n1953 : n1956;
  assign n1958 = pi07 ? n1905 : n1957;
  assign n1959 = pi12 ? n522 : n1955;
  assign n1960 = pi14 ? n543 : n1634;
  assign n1961 = pi13 ? n1960 : n1954;
  assign n1962 = pi12 ? n522 : n1961;
  assign n1963 = pi11 ? n1959 : n1962;
  assign n1964 = pi10 ? n1956 : n1963;
  assign n1965 = pi09 ? n1956 : n1964;
  assign n1966 = pi08 ? n1956 : n1965;
  assign n1967 = pi07 ? n1956 : n1966;
  assign n1968 = pi06 ? n1958 : n1967;
  assign n1969 = pi05 ? n1889 : n1968;
  assign n1970 = pi04 ? n1847 : n1969;
  assign n1971 = pi03 ? n1576 : n1970;
  assign n1972 = pi15 ? n62 : n771;
  assign n1973 = pi14 ? n1972 : n890;
  assign n1974 = pi13 ? n1897 : n1973;
  assign n1975 = pi12 ? n26 : n1974;
  assign n1976 = pi11 ? n1895 : n1975;
  assign n1977 = pi10 ? n1893 : n1976;
  assign n1978 = pi09 ? n26 : n1977;
  assign n1979 = pi08 ? n26 : n1978;
  assign n1980 = pi16 ? n42 : n32;
  assign n1981 = pi15 ? n1980 : n32;
  assign n1982 = pi14 ? n1981 : n1374;
  assign n1983 = pi16 ? n224 : n1813;
  assign n1984 = pi15 ? n224 : n1983;
  assign n1985 = pi14 ? n910 : n1984;
  assign n1986 = pi13 ? n1982 : n1985;
  assign n1987 = pi12 ? n26 : n1986;
  assign n1988 = pi17 ? n41 : n32;
  assign n1989 = pi16 ? n1988 : n32;
  assign n1990 = pi15 ? n1989 : n480;
  assign n1991 = pi14 ? n1990 : n1820;
  assign n1992 = pi15 ? n224 : n1156;
  assign n1993 = pi14 ? n899 : n1992;
  assign n1994 = pi13 ? n1991 : n1993;
  assign n1995 = pi12 ? n26 : n1994;
  assign n1996 = pi11 ? n1987 : n1995;
  assign n1997 = pi15 ? n573 : n989;
  assign n1998 = pi14 ? n1997 : n1616;
  assign n1999 = pi15 ? n475 : n1675;
  assign n2000 = pi14 ? n899 : n1999;
  assign n2001 = pi13 ? n1998 : n2000;
  assign n2002 = pi12 ? n1880 : n2001;
  assign n2003 = pi15 ? n385 : n41;
  assign n2004 = pi14 ? n2003 : n543;
  assign n2005 = pi13 ? n2004 : n1386;
  assign n2006 = pi12 ? n1921 : n2005;
  assign n2007 = pi11 ? n2002 : n2006;
  assign n2008 = pi10 ? n1996 : n2007;
  assign n2009 = pi15 ? n722 : n377;
  assign n2010 = pi14 ? n958 : n2009;
  assign n2011 = pi16 ? n175 : n746;
  assign n2012 = pi15 ? n2011 : n26;
  assign n2013 = pi14 ? n890 : n2012;
  assign n2014 = pi13 ? n2010 : n2013;
  assign n2015 = pi12 ? n1926 : n2014;
  assign n2016 = pi14 ? n958 : n1103;
  assign n2017 = pi15 ? n1221 : n26;
  assign n2018 = pi14 ? n890 : n2017;
  assign n2019 = pi13 ? n2016 : n2018;
  assign n2020 = pi12 ? n1926 : n2019;
  assign n2021 = pi11 ? n2015 : n2020;
  assign n2022 = pi14 ? n958 : n1393;
  assign n2023 = pi16 ? n251 : n155;
  assign n2024 = pi15 ? n224 : n2023;
  assign n2025 = pi14 ? n2024 : n26;
  assign n2026 = pi13 ? n2022 : n2025;
  assign n2027 = pi12 ? n1926 : n2026;
  assign n2028 = pi14 ? n1374 : n1393;
  assign n2029 = pi16 ? n224 : n300;
  assign n2030 = pi15 ? n224 : n2029;
  assign n2031 = pi14 ? n2030 : n26;
  assign n2032 = pi13 ? n2028 : n2031;
  assign n2033 = pi12 ? n1926 : n2032;
  assign n2034 = pi11 ? n2027 : n2033;
  assign n2035 = pi10 ? n2021 : n2034;
  assign n2036 = pi09 ? n2008 : n2035;
  assign n2037 = pi14 ? n1374 : n899;
  assign n2038 = pi14 ? n1992 : n26;
  assign n2039 = pi13 ? n2037 : n2038;
  assign n2040 = pi12 ? n1926 : n2039;
  assign n2041 = pi14 ? n1676 : n26;
  assign n2042 = pi13 ? n2037 : n2041;
  assign n2043 = pi12 ? n1926 : n2042;
  assign n2044 = pi11 ? n2040 : n2043;
  assign n2045 = pi15 ? n41 : n121;
  assign n2046 = pi14 ? n2045 : n899;
  assign n2047 = pi13 ? n2046 : n2041;
  assign n2048 = pi12 ? n1926 : n2047;
  assign n2049 = pi10 ? n2044 : n2048;
  assign n2050 = pi09 ? n2049 : n2048;
  assign n2051 = pi08 ? n2036 : n2050;
  assign n2052 = pi07 ? n1979 : n2051;
  assign n2053 = pi14 ? n2045 : n910;
  assign n2054 = pi13 ? n2053 : n2041;
  assign n2055 = pi12 ? n1926 : n2054;
  assign n2056 = pi11 ? n2048 : n2055;
  assign n2057 = pi10 ? n2048 : n2056;
  assign n2058 = pi09 ? n2048 : n2057;
  assign n2059 = pi08 ? n2048 : n2058;
  assign n2060 = pi07 ? n2048 : n2059;
  assign n2061 = pi06 ? n2052 : n2060;
  assign n2062 = pi14 ? n35 : n1792;
  assign n2063 = pi13 ? n2062 : n1848;
  assign n2064 = pi12 ? n26 : n2063;
  assign n2065 = pi11 ? n26 : n2064;
  assign n2066 = pi14 ? n35 : n958;
  assign n2067 = pi13 ? n2066 : n1584;
  assign n2068 = pi12 ? n26 : n2067;
  assign n2069 = pi15 ? n1989 : n32;
  assign n2070 = pi14 ? n2069 : n958;
  assign n2071 = pi13 ? n2070 : n1973;
  assign n2072 = pi12 ? n26 : n2071;
  assign n2073 = pi11 ? n2068 : n2072;
  assign n2074 = pi10 ? n2065 : n2073;
  assign n2075 = pi09 ? n26 : n2074;
  assign n2076 = pi08 ? n26 : n2075;
  assign n2077 = pi14 ? n32 : n1374;
  assign n2078 = pi15 ? n224 : n1758;
  assign n2079 = pi14 ? n910 : n2078;
  assign n2080 = pi13 ? n2077 : n2079;
  assign n2081 = pi12 ? n26 : n2080;
  assign n2082 = pi15 ? n32 : n480;
  assign n2083 = pi14 ? n2082 : n1820;
  assign n2084 = pi13 ? n2083 : n1993;
  assign n2085 = pi12 ? n1880 : n2084;
  assign n2086 = pi11 ? n2081 : n2085;
  assign n2087 = pi14 ? n26 : n656;
  assign n2088 = pi13 ? n26 : n2087;
  assign n2089 = pi16 ? n343 : n132;
  assign n2090 = pi15 ? n41 : n2089;
  assign n2091 = pi14 ? n2090 : n1616;
  assign n2092 = pi16 ? n461 : n26;
  assign n2093 = pi15 ? n475 : n2092;
  assign n2094 = pi14 ? n899 : n2093;
  assign n2095 = pi13 ? n2091 : n2094;
  assign n2096 = pi12 ? n2088 : n2095;
  assign n2097 = pi11 ? n2096 : n1922;
  assign n2098 = pi10 ? n2086 : n2097;
  assign n2099 = pi13 ? n26 : n131;
  assign n2100 = pi15 ? n1323 : n122;
  assign n2101 = pi15 ? n722 : n60;
  assign n2102 = pi14 ? n2100 : n2101;
  assign n2103 = pi16 ? n175 : n224;
  assign n2104 = pi15 ? n2103 : n26;
  assign n2105 = pi14 ? n1583 : n2104;
  assign n2106 = pi13 ? n2102 : n2105;
  assign n2107 = pi12 ? n2099 : n2106;
  assign n2108 = pi14 ? n958 : n728;
  assign n2109 = pi14 ? n1583 : n2017;
  assign n2110 = pi13 ? n2108 : n2109;
  assign n2111 = pi12 ? n1101 : n2110;
  assign n2112 = pi11 ? n2107 : n2111;
  assign n2113 = pi14 ? n2100 : n523;
  assign n2114 = pi16 ? n224 : n276;
  assign n2115 = pi15 ? n1064 : n2114;
  assign n2116 = pi17 ? n1072 : n26;
  assign n2117 = pi16 ? n2116 : n26;
  assign n2118 = pi15 ? n2117 : n26;
  assign n2119 = pi14 ? n2115 : n2118;
  assign n2120 = pi13 ? n2113 : n2119;
  assign n2121 = pi12 ? n1101 : n2120;
  assign n2122 = pi15 ? n136 : n347;
  assign n2123 = pi14 ? n958 : n2122;
  assign n2124 = pi14 ? n2115 : n26;
  assign n2125 = pi13 ? n2123 : n2124;
  assign n2126 = pi12 ? n1101 : n2125;
  assign n2127 = pi11 ? n2121 : n2126;
  assign n2128 = pi10 ? n2112 : n2127;
  assign n2129 = pi09 ? n2098 : n2128;
  assign n2130 = pi15 ? n136 : n66;
  assign n2131 = pi14 ? n958 : n2130;
  assign n2132 = pi15 ? n1064 : n1758;
  assign n2133 = pi14 ? n2132 : n26;
  assign n2134 = pi13 ? n2131 : n2133;
  assign n2135 = pi12 ? n1101 : n2134;
  assign n2136 = pi15 ? n123 : n347;
  assign n2137 = pi14 ? n958 : n2136;
  assign n2138 = pi16 ? n224 : n1215;
  assign n2139 = pi15 ? n1064 : n2138;
  assign n2140 = pi14 ? n2139 : n26;
  assign n2141 = pi13 ? n2137 : n2140;
  assign n2142 = pi12 ? n1101 : n2141;
  assign n2143 = pi11 ? n2135 : n2142;
  assign n2144 = pi14 ? n2045 : n348;
  assign n2145 = pi14 ? n1436 : n26;
  assign n2146 = pi13 ? n2144 : n2145;
  assign n2147 = pi12 ? n1101 : n2146;
  assign n2148 = pi10 ? n2143 : n2147;
  assign n2149 = pi09 ? n2148 : n2147;
  assign n2150 = pi08 ? n2129 : n2149;
  assign n2151 = pi07 ? n2076 : n2150;
  assign n2152 = pi14 ? n26 : n1044;
  assign n2153 = pi13 ? n26 : n2152;
  assign n2154 = pi12 ? n2153 : n2146;
  assign n2155 = pi13 ? n2144 : n2038;
  assign n2156 = pi12 ? n2153 : n2155;
  assign n2157 = pi11 ? n2154 : n2156;
  assign n2158 = pi13 ? n2053 : n2038;
  assign n2159 = pi12 ? n2153 : n2158;
  assign n2160 = pi10 ? n2157 : n2159;
  assign n2161 = pi09 ? n2147 : n2160;
  assign n2162 = pi08 ? n2147 : n2161;
  assign n2163 = pi07 ? n2147 : n2162;
  assign n2164 = pi06 ? n2151 : n2163;
  assign n2165 = pi05 ? n2061 : n2164;
  assign n2166 = pi15 ? n43 : n122;
  assign n2167 = pi14 ? n35 : n2166;
  assign n2168 = pi14 ? n101 : n1634;
  assign n2169 = pi13 ? n2167 : n2168;
  assign n2170 = pi12 ? n26 : n2169;
  assign n2171 = pi11 ? n26 : n2170;
  assign n2172 = pi14 ? n1532 : n958;
  assign n2173 = pi13 ? n2172 : n1973;
  assign n2174 = pi12 ? n26 : n2173;
  assign n2175 = pi11 ? n2068 : n2174;
  assign n2176 = pi10 ? n2171 : n2175;
  assign n2177 = pi09 ? n26 : n2176;
  assign n2178 = pi08 ? n26 : n2177;
  assign n2179 = pi13 ? n2077 : n1985;
  assign n2180 = pi12 ? n26 : n2179;
  assign n2181 = pi14 ? n910 : n1992;
  assign n2182 = pi13 ? n2083 : n2181;
  assign n2183 = pi12 ? n26 : n2182;
  assign n2184 = pi11 ? n2180 : n2183;
  assign n2185 = pi15 ? n32 : n2089;
  assign n2186 = pi14 ? n2185 : n1616;
  assign n2187 = pi13 ? n2186 : n1677;
  assign n2188 = pi12 ? n2088 : n2187;
  assign n2189 = pi14 ? n205 : n543;
  assign n2190 = pi14 ? n910 : n1681;
  assign n2191 = pi13 ? n2189 : n2190;
  assign n2192 = pi12 ? n1770 : n2191;
  assign n2193 = pi11 ? n2188 : n2192;
  assign n2194 = pi10 ? n2184 : n2193;
  assign n2195 = pi14 ? n205 : n770;
  assign n2196 = pi16 ? n740 : n155;
  assign n2197 = pi15 ? n60 : n2196;
  assign n2198 = pi15 ? n224 : n26;
  assign n2199 = pi14 ? n2197 : n2198;
  assign n2200 = pi13 ? n2195 : n2199;
  assign n2201 = pi12 ? n2099 : n2200;
  assign n2202 = pi14 ? n205 : n427;
  assign n2203 = pi15 ? n60 : n1735;
  assign n2204 = pi15 ? n1156 : n26;
  assign n2205 = pi14 ? n2203 : n2204;
  assign n2206 = pi13 ? n2202 : n2205;
  assign n2207 = pi12 ? n1101 : n2206;
  assign n2208 = pi11 ? n2201 : n2207;
  assign n2209 = pi14 ? n190 : n728;
  assign n2210 = pi17 ? n155 : n175;
  assign n2211 = pi16 ? n740 : n2210;
  assign n2212 = pi15 ? n60 : n2211;
  assign n2213 = pi14 ? n2212 : n2118;
  assign n2214 = pi13 ? n2209 : n2213;
  assign n2215 = pi12 ? n1101 : n2214;
  assign n2216 = pi16 ? n1510 : n238;
  assign n2217 = pi15 ? n60 : n2216;
  assign n2218 = pi14 ? n2217 : n2118;
  assign n2219 = pi13 ? n2209 : n2218;
  assign n2220 = pi12 ? n1101 : n2219;
  assign n2221 = pi11 ? n2215 : n2220;
  assign n2222 = pi10 ? n2208 : n2221;
  assign n2223 = pi09 ? n2194 : n2222;
  assign n2224 = pi14 ? n1206 : n728;
  assign n2225 = pi17 ? n355 : n26;
  assign n2226 = pi16 ? n2225 : n26;
  assign n2227 = pi15 ? n2226 : n26;
  assign n2228 = pi14 ? n2203 : n2227;
  assign n2229 = pi13 ? n2224 : n2228;
  assign n2230 = pi12 ? n1101 : n2229;
  assign n2231 = pi14 ? n2203 : n26;
  assign n2232 = pi13 ? n2224 : n2231;
  assign n2233 = pi12 ? n1101 : n2232;
  assign n2234 = pi11 ? n2230 : n2233;
  assign n2235 = pi16 ? n1510 : n1366;
  assign n2236 = pi15 ? n60 : n2235;
  assign n2237 = pi14 ? n2236 : n26;
  assign n2238 = pi13 ? n2224 : n2237;
  assign n2239 = pi12 ? n1101 : n2238;
  assign n2240 = pi10 ? n2234 : n2239;
  assign n2241 = pi09 ? n2240 : n2239;
  assign n2242 = pi08 ? n2223 : n2241;
  assign n2243 = pi07 ? n2178 : n2242;
  assign n2244 = pi14 ? n1206 : n2101;
  assign n2245 = pi16 ? n740 : n1366;
  assign n2246 = pi15 ? n60 : n2245;
  assign n2247 = pi14 ? n2246 : n26;
  assign n2248 = pi13 ? n2244 : n2247;
  assign n2249 = pi12 ? n1101 : n2248;
  assign n2250 = pi15 ? n1560 : n122;
  assign n2251 = pi14 ? n2250 : n2101;
  assign n2252 = pi16 ? n224 : n355;
  assign n2253 = pi15 ? n493 : n2252;
  assign n2254 = pi14 ? n2253 : n26;
  assign n2255 = pi13 ? n2251 : n2254;
  assign n2256 = pi12 ? n2153 : n2255;
  assign n2257 = pi11 ? n2249 : n2256;
  assign n2258 = pi14 ? n2250 : n728;
  assign n2259 = pi15 ? n224 : n2252;
  assign n2260 = pi14 ? n2259 : n26;
  assign n2261 = pi13 ? n2258 : n2260;
  assign n2262 = pi12 ? n1101 : n2261;
  assign n2263 = pi14 ? n2078 : n26;
  assign n2264 = pi13 ? n2258 : n2263;
  assign n2265 = pi12 ? n1101 : n2264;
  assign n2266 = pi11 ? n2262 : n2265;
  assign n2267 = pi10 ? n2257 : n2266;
  assign n2268 = pi09 ? n2239 : n2267;
  assign n2269 = pi08 ? n2239 : n2268;
  assign n2270 = pi07 ? n2239 : n2269;
  assign n2271 = pi06 ? n2243 : n2270;
  assign n2272 = pi16 ? n32 : n1198;
  assign n2273 = pi15 ? n32 : n2272;
  assign n2274 = pi17 ? n47 : n53;
  assign n2275 = pi16 ? n2274 : n60;
  assign n2276 = pi15 ? n122 : n2275;
  assign n2277 = pi14 ? n2273 : n2276;
  assign n2278 = pi17 ? n65 : n26;
  assign n2279 = pi16 ? n2278 : n26;
  assign n2280 = pi15 ? n2279 : n26;
  assign n2281 = pi14 ? n323 : n2280;
  assign n2282 = pi13 ? n2277 : n2281;
  assign n2283 = pi12 ? n1101 : n2282;
  assign n2284 = pi11 ? n26 : n2283;
  assign n2285 = pi10 ? n26 : n2284;
  assign n2286 = pi14 ? n2185 : n2276;
  assign n2287 = pi14 ? n1202 : n2227;
  assign n2288 = pi13 ? n2286 : n2287;
  assign n2289 = pi12 ? n1101 : n2288;
  assign n2290 = pi15 ? n694 : n739;
  assign n2291 = pi14 ? n205 : n2290;
  assign n2292 = pi16 ? n224 : n65;
  assign n2293 = pi15 ? n60 : n2292;
  assign n2294 = pi14 ? n2293 : n2227;
  assign n2295 = pi13 ? n2291 : n2294;
  assign n2296 = pi12 ? n1101 : n2295;
  assign n2297 = pi11 ? n2289 : n2296;
  assign n2298 = pi15 ? n32 : n122;
  assign n2299 = pi16 ? n502 : n626;
  assign n2300 = pi15 ? n2299 : n66;
  assign n2301 = pi14 ? n2298 : n2300;
  assign n2302 = pi14 ? n224 : n2227;
  assign n2303 = pi13 ? n2301 : n2302;
  assign n2304 = pi12 ? n1101 : n2303;
  assign n2305 = pi13 ? n2258 : n2302;
  assign n2306 = pi12 ? n1101 : n2305;
  assign n2307 = pi11 ? n2304 : n2306;
  assign n2308 = pi10 ? n2297 : n2307;
  assign n2309 = pi09 ? n2285 : n2308;
  assign n2310 = pi08 ? n26 : n2309;
  assign n2311 = pi07 ? n26 : n2310;
  assign n2312 = pi06 ? n26 : n2311;
  assign n2313 = pi05 ? n2271 : n2312;
  assign n2314 = pi04 ? n2165 : n2313;
  assign n2315 = pi16 ? n186 : n452;
  assign n2316 = pi15 ? n2315 : n32;
  assign n2317 = pi15 ? n438 : n231;
  assign n2318 = pi14 ? n2316 : n2317;
  assign n2319 = pi16 ? n60 : n2278;
  assign n2320 = pi15 ? n2319 : n26;
  assign n2321 = pi14 ? n1662 : n2320;
  assign n2322 = pi13 ? n2318 : n2321;
  assign n2323 = pi12 ? n1308 : n2322;
  assign n2324 = pi11 ? n26 : n2323;
  assign n2325 = pi10 ? n26 : n2324;
  assign n2326 = pi16 ? n476 : n452;
  assign n2327 = pi15 ? n2326 : n32;
  assign n2328 = pi15 ? n231 : n503;
  assign n2329 = pi14 ? n2327 : n2328;
  assign n2330 = pi15 ? n1633 : n26;
  assign n2331 = pi14 ? n323 : n2330;
  assign n2332 = pi13 ? n2329 : n2331;
  assign n2333 = pi12 ? n1315 : n2332;
  assign n2334 = pi15 ? n2326 : n555;
  assign n2335 = pi15 ? n231 : n923;
  assign n2336 = pi14 ? n2334 : n2335;
  assign n2337 = pi14 ? n899 : n2330;
  assign n2338 = pi13 ? n2336 : n2337;
  assign n2339 = pi12 ? n1101 : n2338;
  assign n2340 = pi11 ? n2333 : n2339;
  assign n2341 = pi15 ? n32 : n989;
  assign n2342 = pi17 ? n121 : n53;
  assign n2343 = pi16 ? n2342 : n60;
  assign n2344 = pi15 ? n122 : n2343;
  assign n2345 = pi14 ? n2341 : n2344;
  assign n2346 = pi16 ? n274 : n26;
  assign n2347 = pi15 ? n2346 : n26;
  assign n2348 = pi14 ? n494 : n2347;
  assign n2349 = pi13 ? n2345 : n2348;
  assign n2350 = pi12 ? n1101 : n2349;
  assign n2351 = pi15 ? n1323 : n41;
  assign n2352 = pi14 ? n2351 : n2276;
  assign n2353 = pi13 ? n2352 : n2348;
  assign n2354 = pi12 ? n1559 : n2353;
  assign n2355 = pi11 ? n2350 : n2354;
  assign n2356 = pi10 ? n2340 : n2355;
  assign n2357 = pi09 ? n2325 : n2356;
  assign n2358 = pi08 ? n26 : n2357;
  assign n2359 = pi07 ? n26 : n2358;
  assign n2360 = pi06 ? n26 : n2359;
  assign n2361 = pi14 ? n49 : n101;
  assign n2362 = pi13 ? n426 : n2361;
  assign n2363 = pi12 ? n26 : n2362;
  assign n2364 = pi11 ? n26 : n2363;
  assign n2365 = pi14 ? n74 : n101;
  assign n2366 = pi13 ? n426 : n2365;
  assign n2367 = pi12 ? n26 : n2366;
  assign n2368 = pi10 ? n2364 : n2367;
  assign n2369 = pi09 ? n26 : n2368;
  assign n2370 = pi08 ? n26 : n2369;
  assign n2371 = pi13 ? n1176 : n2365;
  assign n2372 = pi12 ? n26 : n2371;
  assign n2373 = pi11 ? n2367 : n2372;
  assign n2374 = pi10 ? n2367 : n2373;
  assign n2375 = pi11 ? n2372 : n2367;
  assign n2376 = pi10 ? n2375 : n2367;
  assign n2377 = pi09 ? n2374 : n2376;
  assign n2378 = pi08 ? n2367 : n2377;
  assign n2379 = pi07 ? n2370 : n2378;
  assign n2380 = pi16 ? n175 : n452;
  assign n2381 = pi15 ? n2380 : n32;
  assign n2382 = pi14 ? n406 : n2381;
  assign n2383 = pi15 ? n100 : n2319;
  assign n2384 = pi14 ? n74 : n2383;
  assign n2385 = pi13 ? n2382 : n2384;
  assign n2386 = pi12 ? n26 : n2385;
  assign n2387 = pi11 ? n2367 : n2386;
  assign n2388 = pi10 ? n2367 : n2387;
  assign n2389 = pi09 ? n2367 : n2388;
  assign n2390 = pi17 ? n355 : n175;
  assign n2391 = pi16 ? n2390 : n452;
  assign n2392 = pi15 ? n2391 : n32;
  assign n2393 = pi14 ? n294 : n2392;
  assign n2394 = pi15 ? n73 : n364;
  assign n2395 = pi14 ? n2394 : n292;
  assign n2396 = pi13 ? n2393 : n2395;
  assign n2397 = pi12 ? n26 : n2396;
  assign n2398 = pi14 ? n824 : n454;
  assign n2399 = pi15 ? n62 : n2279;
  assign n2400 = pi14 ? n1193 : n2399;
  assign n2401 = pi13 ? n2398 : n2400;
  assign n2402 = pi12 ? n26 : n2401;
  assign n2403 = pi11 ? n2397 : n2402;
  assign n2404 = pi16 ? n1072 : n186;
  assign n2405 = pi15 ? n250 : n2404;
  assign n2406 = pi14 ? n2405 : n1200;
  assign n2407 = pi15 ? n66 : n26;
  assign n2408 = pi14 ? n232 : n2407;
  assign n2409 = pi13 ? n2406 : n2408;
  assign n2410 = pi12 ? n26 : n2409;
  assign n2411 = pi15 ? n178 : n808;
  assign n2412 = pi14 ? n2411 : n2317;
  assign n2413 = pi14 ? n1426 : n2407;
  assign n2414 = pi13 ? n2412 : n2413;
  assign n2415 = pi12 ? n1539 : n2414;
  assign n2416 = pi11 ? n2410 : n2415;
  assign n2417 = pi10 ? n2403 : n2416;
  assign n2418 = pi16 ? n2274 : n626;
  assign n2419 = pi15 ? n258 : n2418;
  assign n2420 = pi14 ? n242 : n2419;
  assign n2421 = pi14 ? n323 : n2320;
  assign n2422 = pi13 ? n2420 : n2421;
  assign n2423 = pi12 ? n1770 : n2422;
  assign n2424 = pi15 ? n231 : n321;
  assign n2425 = pi14 ? n2327 : n2424;
  assign n2426 = pi16 ? n224 : n2278;
  assign n2427 = pi15 ? n2426 : n26;
  assign n2428 = pi14 ? n2293 : n2427;
  assign n2429 = pi13 ? n2425 : n2428;
  assign n2430 = pi12 ? n1315 : n2429;
  assign n2431 = pi11 ? n2423 : n2430;
  assign n2432 = pi16 ? n176 : n1830;
  assign n2433 = pi15 ? n26 : n2432;
  assign n2434 = pi14 ? n26 : n2433;
  assign n2435 = pi13 ? n26 : n2434;
  assign n2436 = pi14 ? n1548 : n2335;
  assign n2437 = pi15 ? n1675 : n26;
  assign n2438 = pi14 ? n494 : n2437;
  assign n2439 = pi13 ? n2436 : n2438;
  assign n2440 = pi12 ? n2435 : n2439;
  assign n2441 = pi13 ? n26 : n625;
  assign n2442 = pi14 ? n1561 : n924;
  assign n2443 = pi13 ? n2442 : n2438;
  assign n2444 = pi12 ? n2441 : n2443;
  assign n2445 = pi11 ? n2440 : n2444;
  assign n2446 = pi10 ? n2431 : n2445;
  assign n2447 = pi09 ? n2417 : n2446;
  assign n2448 = pi08 ? n2389 : n2447;
  assign n2449 = pi07 ? n2367 : n2448;
  assign n2450 = pi06 ? n2379 : n2449;
  assign n2451 = pi05 ? n2360 : n2450;
  assign n2452 = pi14 ? n376 : n316;
  assign n2453 = pi13 ? n657 : n2452;
  assign n2454 = pi12 ? n26 : n2453;
  assign n2455 = pi11 ? n26 : n2454;
  assign n2456 = pi15 ? n32 : n114;
  assign n2457 = pi14 ? n656 : n2456;
  assign n2458 = pi13 ? n2457 : n2452;
  assign n2459 = pi12 ? n26 : n2458;
  assign n2460 = pi10 ? n2455 : n2459;
  assign n2461 = pi09 ? n26 : n2460;
  assign n2462 = pi08 ? n26 : n2461;
  assign n2463 = pi15 ? n213 : n114;
  assign n2464 = pi14 ? n656 : n2463;
  assign n2465 = pi13 ? n2464 : n2452;
  assign n2466 = pi12 ? n26 : n2465;
  assign n2467 = pi11 ? n2466 : n2459;
  assign n2468 = pi10 ? n2459 : n2467;
  assign n2469 = pi09 ? n2468 : n2459;
  assign n2470 = pi08 ? n2459 : n2469;
  assign n2471 = pi07 ? n2462 : n2470;
  assign n2472 = pi14 ? n406 : n2456;
  assign n2473 = pi13 ? n2472 : n2452;
  assign n2474 = pi12 ? n26 : n2473;
  assign n2475 = pi11 ? n2459 : n2474;
  assign n2476 = pi14 ? n144 : n2456;
  assign n2477 = pi13 ? n2476 : n2452;
  assign n2478 = pi12 ? n26 : n2477;
  assign n2479 = pi14 ? n294 : n2456;
  assign n2480 = pi15 ? n123 : n2319;
  assign n2481 = pi14 ? n365 : n2480;
  assign n2482 = pi13 ? n2479 : n2481;
  assign n2483 = pi12 ? n26 : n2482;
  assign n2484 = pi11 ? n2478 : n2483;
  assign n2485 = pi10 ? n2475 : n2484;
  assign n2486 = pi09 ? n2459 : n2485;
  assign n2487 = pi17 ? n175 : n355;
  assign n2488 = pi16 ? n176 : n2487;
  assign n2489 = pi15 ? n26 : n2488;
  assign n2490 = pi14 ? n2489 : n2456;
  assign n2491 = pi16 ? n53 : n47;
  assign n2492 = pi15 ? n41 : n2491;
  assign n2493 = pi15 ? n123 : n291;
  assign n2494 = pi14 ? n2492 : n2493;
  assign n2495 = pi13 ? n2490 : n2494;
  assign n2496 = pi12 ? n26 : n2495;
  assign n2497 = pi15 ? n405 : n1073;
  assign n2498 = pi14 ? n2497 : n2456;
  assign n2499 = pi15 ? n60 : n2279;
  assign n2500 = pi14 ? n820 : n2499;
  assign n2501 = pi13 ? n2498 : n2500;
  assign n2502 = pi12 ? n26 : n2501;
  assign n2503 = pi11 ? n2496 : n2502;
  assign n2504 = pi15 ? n701 : n1073;
  assign n2505 = pi14 ? n2504 : n2341;
  assign n2506 = pi15 ? n65 : n26;
  assign n2507 = pi14 ? n124 : n2506;
  assign n2508 = pi13 ? n2505 : n2507;
  assign n2509 = pi12 ? n26 : n2508;
  assign n2510 = pi14 ? n425 : n1206;
  assign n2511 = pi15 ? n62 : n739;
  assign n2512 = pi14 ? n2511 : n2506;
  assign n2513 = pi13 ? n2510 : n2512;
  assign n2514 = pi12 ? n26 : n2513;
  assign n2515 = pi11 ? n2509 : n2514;
  assign n2516 = pi10 ? n2503 : n2515;
  assign n2517 = pi14 ? n242 : n958;
  assign n2518 = pi16 ? n355 : n274;
  assign n2519 = pi15 ? n2518 : n26;
  assign n2520 = pi14 ? n1202 : n2519;
  assign n2521 = pi13 ? n2517 : n2520;
  assign n2522 = pi12 ? n1770 : n2521;
  assign n2523 = pi16 ? n128 : n1830;
  assign n2524 = pi15 ? n26 : n2523;
  assign n2525 = pi14 ? n26 : n2524;
  assign n2526 = pi13 ? n26 : n2525;
  assign n2527 = pi16 ? n41 : n53;
  assign n2528 = pi15 ? n41 : n2527;
  assign n2529 = pi14 ? n1763 : n2528;
  assign n2530 = pi13 ? n2529 : n2520;
  assign n2531 = pi12 ? n2526 : n2530;
  assign n2532 = pi11 ? n2522 : n2531;
  assign n2533 = pi15 ? n231 : n722;
  assign n2534 = pi14 ? n134 : n2533;
  assign n2535 = pi14 ? n899 : n2437;
  assign n2536 = pi13 ? n2534 : n2535;
  assign n2537 = pi12 ? n2435 : n2536;
  assign n2538 = pi14 ? n1653 : n2533;
  assign n2539 = pi13 ? n2538 : n2438;
  assign n2540 = pi12 ? n2441 : n2539;
  assign n2541 = pi11 ? n2537 : n2540;
  assign n2542 = pi10 ? n2532 : n2541;
  assign n2543 = pi09 ? n2516 : n2542;
  assign n2544 = pi08 ? n2486 : n2543;
  assign n2545 = pi07 ? n2459 : n2544;
  assign n2546 = pi06 ? n2471 : n2545;
  assign n2547 = pi15 ? n73 : n96;
  assign n2548 = pi14 ? n144 : n2547;
  assign n2549 = pi15 ? n123 : n546;
  assign n2550 = pi14 ? n315 : n2549;
  assign n2551 = pi13 ? n2548 : n2550;
  assign n2552 = pi12 ? n26 : n2551;
  assign n2553 = pi11 ? n26 : n2552;
  assign n2554 = pi14 ? n144 : n1400;
  assign n2555 = pi13 ? n2554 : n2550;
  assign n2556 = pi12 ? n26 : n2555;
  assign n2557 = pi10 ? n2553 : n2556;
  assign n2558 = pi09 ? n26 : n2557;
  assign n2559 = pi08 ? n26 : n2558;
  assign n2560 = pi15 ? n438 : n333;
  assign n2561 = pi14 ? n144 : n2560;
  assign n2562 = pi13 ? n2561 : n1394;
  assign n2563 = pi12 ? n26 : n2562;
  assign n2564 = pi11 ? n2556 : n2563;
  assign n2565 = pi10 ? n2556 : n2564;
  assign n2566 = pi15 ? n32 : n333;
  assign n2567 = pi14 ? n144 : n2566;
  assign n2568 = pi13 ? n2567 : n1394;
  assign n2569 = pi12 ? n26 : n2568;
  assign n2570 = pi16 ? n107 : n563;
  assign n2571 = pi15 ? n32 : n2570;
  assign n2572 = pi14 ? n144 : n2571;
  assign n2573 = pi13 ? n2572 : n1394;
  assign n2574 = pi12 ? n26 : n2573;
  assign n2575 = pi11 ? n2569 : n2574;
  assign n2576 = pi15 ? n123 : n558;
  assign n2577 = pi14 ? n315 : n2576;
  assign n2578 = pi13 ? n2567 : n2577;
  assign n2579 = pi12 ? n26 : n2578;
  assign n2580 = pi13 ? n2554 : n2577;
  assign n2581 = pi12 ? n26 : n2580;
  assign n2582 = pi11 ? n2579 : n2581;
  assign n2583 = pi10 ? n2575 : n2582;
  assign n2584 = pi09 ? n2565 : n2583;
  assign n2585 = pi08 ? n2556 : n2584;
  assign n2586 = pi07 ? n2559 : n2585;
  assign n2587 = pi14 ? n395 : n1400;
  assign n2588 = pi14 ? n365 : n2549;
  assign n2589 = pi13 ? n2587 : n2588;
  assign n2590 = pi12 ? n26 : n2589;
  assign n2591 = pi11 ? n2556 : n2590;
  assign n2592 = pi14 ? n1776 : n1400;
  assign n2593 = pi16 ? n545 : n355;
  assign n2594 = pi15 ? n60 : n2593;
  assign n2595 = pi14 ? n315 : n2594;
  assign n2596 = pi13 ? n2592 : n2595;
  assign n2597 = pi12 ? n26 : n2596;
  assign n2598 = pi16 ? n176 : n255;
  assign n2599 = pi15 ? n26 : n2598;
  assign n2600 = pi14 ? n2599 : n1400;
  assign n2601 = pi16 ? n545 : n274;
  assign n2602 = pi15 ? n60 : n2601;
  assign n2603 = pi14 ? n628 : n2602;
  assign n2604 = pi13 ? n2600 : n2603;
  assign n2605 = pi12 ? n26 : n2604;
  assign n2606 = pi11 ? n2597 : n2605;
  assign n2607 = pi10 ? n2591 : n2606;
  assign n2608 = pi09 ? n2556 : n2607;
  assign n2609 = pi16 ? n1072 : n255;
  assign n2610 = pi15 ? n26 : n2609;
  assign n2611 = pi14 ? n2610 : n1400;
  assign n2612 = pi16 ? n545 : n26;
  assign n2613 = pi15 ? n60 : n2612;
  assign n2614 = pi14 ? n124 : n2613;
  assign n2615 = pi13 ? n2611 : n2614;
  assign n2616 = pi12 ? n26 : n2615;
  assign n2617 = pi15 ? n405 : n2609;
  assign n2618 = pi14 ? n2617 : n1481;
  assign n2619 = pi17 ? n355 : n65;
  assign n2620 = pi16 ? n2619 : n26;
  assign n2621 = pi15 ? n60 : n2620;
  assign n2622 = pi14 ? n124 : n2621;
  assign n2623 = pi13 ? n2618 : n2622;
  assign n2624 = pi12 ? n26 : n2623;
  assign n2625 = pi11 ? n2616 : n2624;
  assign n2626 = pi16 ? n33 : n298;
  assign n2627 = pi16 ? n32 : n194;
  assign n2628 = pi15 ? n2626 : n2627;
  assign n2629 = pi14 ? n2628 : n190;
  assign n2630 = pi15 ? n65 : n2346;
  assign n2631 = pi14 ? n1340 : n2630;
  assign n2632 = pi13 ? n2629 : n2631;
  assign n2633 = pi12 ? n26 : n2632;
  assign n2634 = pi14 ? n425 : n1792;
  assign n2635 = pi15 ? n65 : n2279;
  assign n2636 = pi14 ? n1125 : n2635;
  assign n2637 = pi13 ? n2634 : n2636;
  assign n2638 = pi12 ? n26 : n2637;
  assign n2639 = pi11 ? n2633 : n2638;
  assign n2640 = pi10 ? n2625 : n2639;
  assign n2641 = pi15 ? n41 : n231;
  assign n2642 = pi14 ? n32 : n2641;
  assign n2643 = pi15 ? n123 : n65;
  assign n2644 = pi15 ? n1064 : n26;
  assign n2645 = pi14 ? n2643 : n2644;
  assign n2646 = pi13 ? n2642 : n2645;
  assign n2647 = pi12 ? n1539 : n2646;
  assign n2648 = pi16 ? n26 : n1830;
  assign n2649 = pi15 ? n26 : n2648;
  assign n2650 = pi14 ? n26 : n2649;
  assign n2651 = pi13 ? n26 : n2650;
  assign n2652 = pi16 ? n476 : n437;
  assign n2653 = pi15 ? n2652 : n32;
  assign n2654 = pi14 ? n2653 : n958;
  assign n2655 = pi16 ? n740 : n65;
  assign n2656 = pi15 ? n123 : n2655;
  assign n2657 = pi14 ? n2656 : n2644;
  assign n2658 = pi13 ? n2654 : n2657;
  assign n2659 = pi12 ? n2651 : n2658;
  assign n2660 = pi11 ? n2647 : n2659;
  assign n2661 = pi14 ? n1548 : n723;
  assign n2662 = pi14 ? n910 : n2204;
  assign n2663 = pi13 ? n2661 : n2662;
  assign n2664 = pi12 ? n2435 : n2663;
  assign n2665 = pi15 ? n1323 : n96;
  assign n2666 = pi14 ? n2665 : n723;
  assign n2667 = pi14 ? n494 : n2204;
  assign n2668 = pi13 ? n2666 : n2667;
  assign n2669 = pi12 ? n2441 : n2668;
  assign n2670 = pi11 ? n2664 : n2669;
  assign n2671 = pi10 ? n2660 : n2670;
  assign n2672 = pi09 ? n2640 : n2671;
  assign n2673 = pi08 ? n2608 : n2672;
  assign n2674 = pi07 ? n2556 : n2673;
  assign n2675 = pi06 ? n2586 : n2674;
  assign n2676 = pi05 ? n2546 : n2675;
  assign n2677 = pi04 ? n2451 : n2676;
  assign n2678 = pi03 ? n2314 : n2677;
  assign n2679 = pi02 ? n1971 : n2678;
  assign n2680 = pi01 ? n761 : n2679;
  assign n2681 = pi14 ? n130 : n1631;
  assign n2682 = pi13 ? n2681 : n1691;
  assign n2683 = pi12 ? n26 : n2682;
  assign n2684 = pi11 ? n26 : n2683;
  assign n2685 = pi10 ? n2684 : n1703;
  assign n2686 = pi09 ? n26 : n2685;
  assign n2687 = pi08 ? n26 : n2686;
  assign n2688 = pi14 ? n1776 : n1641;
  assign n2689 = pi13 ? n2688 : n1698;
  assign n2690 = pi12 ? n26 : n2689;
  assign n2691 = pi11 ? n2690 : n1703;
  assign n2692 = pi10 ? n1703 : n2691;
  assign n2693 = pi14 ? n130 : n117;
  assign n2694 = pi14 ? n723 : n1264;
  assign n2695 = pi13 ? n2693 : n2694;
  assign n2696 = pi12 ? n26 : n2695;
  assign n2697 = pi15 ? n573 : n96;
  assign n2698 = pi14 ? n1044 : n2697;
  assign n2699 = pi15 ? n60 : n1064;
  assign n2700 = pi14 ? n723 : n2699;
  assign n2701 = pi13 ? n2698 : n2700;
  assign n2702 = pi12 ? n26 : n2701;
  assign n2703 = pi11 ? n2702 : n1703;
  assign n2704 = pi10 ? n2696 : n2703;
  assign n2705 = pi09 ? n2692 : n2704;
  assign n2706 = pi08 ? n1703 : n2705;
  assign n2707 = pi07 ? n2687 : n2706;
  assign n2708 = pi13 ? n1701 : n1646;
  assign n2709 = pi12 ? n26 : n2708;
  assign n2710 = pi13 ? n1705 : n1643;
  assign n2711 = pi12 ? n26 : n2710;
  assign n2712 = pi11 ? n2709 : n2711;
  assign n2713 = pi14 ? n1053 : n1653;
  assign n2714 = pi14 ? n723 : n2253;
  assign n2715 = pi13 ? n2713 : n2714;
  assign n2716 = pi12 ? n26 : n2715;
  assign n2717 = pi14 ? n723 : n1668;
  assign n2718 = pi13 ? n1710 : n2717;
  assign n2719 = pi12 ? n26 : n2718;
  assign n2720 = pi11 ? n2716 : n2719;
  assign n2721 = pi10 ? n2712 : n2720;
  assign n2722 = pi09 ? n1703 : n2721;
  assign n2723 = pi15 ? n26 : n2404;
  assign n2724 = pi14 ? n2723 : n1653;
  assign n2725 = pi15 ? n493 : n1675;
  assign n2726 = pi14 ? n924 : n2725;
  assign n2727 = pi13 ? n2724 : n2726;
  assign n2728 = pi12 ? n26 : n2727;
  assign n2729 = pi15 ? n462 : n2404;
  assign n2730 = pi15 ? n41 : n133;
  assign n2731 = pi14 ? n2729 : n2730;
  assign n2732 = pi15 ? n493 : n2346;
  assign n2733 = pi14 ? n924 : n2732;
  assign n2734 = pi13 ? n2731 : n2733;
  assign n2735 = pi12 ? n26 : n2734;
  assign n2736 = pi11 ? n2728 : n2735;
  assign n2737 = pi16 ? n33 : n452;
  assign n2738 = pi15 ? n2737 : n808;
  assign n2739 = pi14 ? n2738 : n41;
  assign n2740 = pi14 ? n1125 : n2732;
  assign n2741 = pi13 ? n2739 : n2740;
  assign n2742 = pi12 ? n26 : n2741;
  assign n2743 = pi14 ? n425 : n958;
  assign n2744 = pi14 ? n378 : n2198;
  assign n2745 = pi13 ? n2743 : n2744;
  assign n2746 = pi12 ? n26 : n2745;
  assign n2747 = pi11 ? n2742 : n2746;
  assign n2748 = pi10 ? n2736 : n2747;
  assign n2749 = pi15 ? n123 : n493;
  assign n2750 = pi14 ? n2749 : n2198;
  assign n2751 = pi13 ? n2517 : n2750;
  assign n2752 = pi12 ? n2088 : n2751;
  assign n2753 = pi14 ? n32 : n958;
  assign n2754 = pi14 ? n1393 : n2198;
  assign n2755 = pi13 ? n2753 : n2754;
  assign n2756 = pi12 ? n1770 : n2755;
  assign n2757 = pi11 ? n2752 : n2756;
  assign n2758 = pi14 ? n117 : n723;
  assign n2759 = pi13 ? n2758 : n2662;
  assign n2760 = pi12 ? n2526 : n2759;
  assign n2761 = pi14 ? n1631 : n723;
  assign n2762 = pi14 ? n1634 : n2204;
  assign n2763 = pi13 ? n2761 : n2762;
  assign n2764 = pi12 ? n1315 : n2763;
  assign n2765 = pi11 ? n2760 : n2764;
  assign n2766 = pi10 ? n2757 : n2765;
  assign n2767 = pi09 ? n2748 : n2766;
  assign n2768 = pi08 ? n2722 : n2767;
  assign n2769 = pi07 ? n1703 : n2768;
  assign n2770 = pi06 ? n2707 : n2769;
  assign n2771 = pi16 ? n41 : n107;
  assign n2772 = pi16 ? n96 : n1143;
  assign n2773 = pi15 ? n2771 : n2772;
  assign n2774 = pi14 ? n115 : n2773;
  assign n2775 = pi14 ? n924 : n224;
  assign n2776 = pi13 ? n2774 : n2775;
  assign n2777 = pi12 ? n26 : n2776;
  assign n2778 = pi11 ? n26 : n2777;
  assign n2779 = pi14 ? n369 : n1653;
  assign n2780 = pi13 ? n2779 : n785;
  assign n2781 = pi12 ? n26 : n2780;
  assign n2782 = pi15 ? n41 : n936;
  assign n2783 = pi14 ? n369 : n2782;
  assign n2784 = pi13 ? n2783 : n797;
  assign n2785 = pi12 ? n26 : n2784;
  assign n2786 = pi11 ? n2781 : n2785;
  assign n2787 = pi10 ? n2778 : n2786;
  assign n2788 = pi09 ? n26 : n2787;
  assign n2789 = pi08 ? n26 : n2788;
  assign n2790 = pi07 ? n26 : n2789;
  assign n2791 = pi15 ? n26 : n229;
  assign n2792 = pi14 ? n2791 : n1927;
  assign n2793 = pi13 ? n2792 : n803;
  assign n2794 = pi12 ? n26 : n2793;
  assign n2795 = pi11 ? n2794 : n26;
  assign n2796 = pi10 ? n2795 : n26;
  assign n2797 = pi09 ? n2796 : n26;
  assign n2798 = pi08 ? n2797 : n26;
  assign n2799 = pi07 ? n2798 : n26;
  assign n2800 = pi06 ? n2790 : n2799;
  assign n2801 = pi05 ? n2770 : n2800;
  assign n2802 = pi14 ? n427 : n547;
  assign n2803 = pi13 ? n1577 : n2802;
  assign n2804 = pi12 ? n26 : n2803;
  assign n2805 = pi11 ? n26 : n2804;
  assign n2806 = pi14 ? n369 : n958;
  assign n2807 = pi14 ? n101 : n546;
  assign n2808 = pi13 ? n2806 : n2807;
  assign n2809 = pi12 ? n26 : n2808;
  assign n2810 = pi15 ? n552 : n333;
  assign n2811 = pi14 ? n2810 : n958;
  assign n2812 = pi13 ? n2811 : n1899;
  assign n2813 = pi12 ? n26 : n2812;
  assign n2814 = pi11 ? n2809 : n2813;
  assign n2815 = pi10 ? n2805 : n2814;
  assign n2816 = pi09 ? n26 : n2815;
  assign n2817 = pi08 ? n26 : n2816;
  assign n2818 = pi07 ? n26 : n2817;
  assign n2819 = pi15 ? n552 : n96;
  assign n2820 = pi15 ? n1549 : n542;
  assign n2821 = pi14 ? n2819 : n2820;
  assign n2822 = pi16 ? n1167 : n300;
  assign n2823 = pi15 ? n224 : n2822;
  assign n2824 = pi14 ? n494 : n2823;
  assign n2825 = pi13 ? n2821 : n2824;
  assign n2826 = pi12 ? n26 : n2825;
  assign n2827 = pi11 ? n2826 : n26;
  assign n2828 = pi10 ? n2827 : n26;
  assign n2829 = pi09 ? n2828 : n26;
  assign n2830 = pi08 ? n2829 : n26;
  assign n2831 = pi07 ? n2830 : n26;
  assign n2832 = pi06 ? n2818 : n2831;
  assign n2833 = pi14 ? n1186 : n101;
  assign n2834 = pi13 ? n426 : n2833;
  assign n2835 = pi12 ? n26 : n2834;
  assign n2836 = pi10 ? n2364 : n2835;
  assign n2837 = pi09 ? n26 : n2836;
  assign n2838 = pi08 ? n26 : n2837;
  assign n2839 = pi14 ? n26 : n2381;
  assign n2840 = pi13 ? n2839 : n75;
  assign n2841 = pi12 ? n26 : n2840;
  assign n2842 = pi11 ? n2835 : n2841;
  assign n2843 = pi13 ? n2382 : n1194;
  assign n2844 = pi12 ? n26 : n2843;
  assign n2845 = pi14 ? n294 : n2316;
  assign n2846 = pi14 ? n1193 : n1662;
  assign n2847 = pi13 ? n2845 : n2846;
  assign n2848 = pi12 ? n26 : n2847;
  assign n2849 = pi11 ? n2844 : n2848;
  assign n2850 = pi10 ? n2842 : n2849;
  assign n2851 = pi15 ? n26 : n997;
  assign n2852 = pi14 ? n2851 : n1200;
  assign n2853 = pi14 ? n124 : n323;
  assign n2854 = pi13 ? n2852 : n2853;
  assign n2855 = pi12 ? n26 : n2854;
  assign n2856 = pi14 ? n88 : n1206;
  assign n2857 = pi14 ? n1125 : n1210;
  assign n2858 = pi13 ? n2856 : n2857;
  assign n2859 = pi12 ? n26 : n2858;
  assign n2860 = pi11 ? n2855 : n2859;
  assign n2861 = pi15 ? n87 : n114;
  assign n2862 = pi14 ? n2861 : n958;
  assign n2863 = pi14 ? n523 : n840;
  assign n2864 = pi13 ? n2862 : n2863;
  assign n2865 = pi12 ? n26 : n2864;
  assign n2866 = pi15 ? n598 : n333;
  assign n2867 = pi14 ? n2866 : n958;
  assign n2868 = pi13 ? n2867 : n1158;
  assign n2869 = pi12 ? n26 : n2868;
  assign n2870 = pi11 ? n2865 : n2869;
  assign n2871 = pi10 ? n2860 : n2870;
  assign n2872 = pi09 ? n2850 : n2871;
  assign n2873 = pi08 ? n2835 : n2872;
  assign n2874 = pi07 ? n2838 : n2873;
  assign n2875 = pi14 ? n1615 : n543;
  assign n2876 = pi15 ? n224 : n1168;
  assign n2877 = pi14 ? n494 : n2876;
  assign n2878 = pi13 ? n2875 : n2877;
  assign n2879 = pi12 ? n26 : n2878;
  assign n2880 = pi14 ? n838 : n1325;
  assign n2881 = pi15 ? n997 : n26;
  assign n2882 = pi14 ? n840 : n2881;
  assign n2883 = pi13 ? n2880 : n2882;
  assign n2884 = pi12 ? n26 : n2883;
  assign n2885 = pi11 ? n2879 : n2884;
  assign n2886 = pi15 ? n286 : n542;
  assign n2887 = pi14 ? n2886 : n494;
  assign n2888 = pi16 ? n677 : n452;
  assign n2889 = pi15 ? n464 : n2888;
  assign n2890 = pi14 ? n2889 : n26;
  assign n2891 = pi13 ? n2887 : n2890;
  assign n2892 = pi12 ? n26 : n2891;
  assign n2893 = pi12 ? n26 : n1946;
  assign n2894 = pi11 ? n2892 : n2893;
  assign n2895 = pi10 ? n2885 : n2894;
  assign n2896 = pi12 ? n1880 : n1949;
  assign n2897 = pi14 ? n1385 : n26;
  assign n2898 = pi13 ? n1936 : n2897;
  assign n2899 = pi12 ? n1921 : n2898;
  assign n2900 = pi11 ? n2896 : n2899;
  assign n2901 = pi10 ? n2900 : n1956;
  assign n2902 = pi09 ? n2895 : n2901;
  assign n2903 = pi08 ? n2902 : n1956;
  assign n2904 = pi07 ? n2903 : n1966;
  assign n2905 = pi06 ? n2874 : n2904;
  assign n2906 = pi05 ? n2832 : n2905;
  assign n2907 = pi04 ? n2801 : n2906;
  assign n2908 = pi14 ? n365 : n323;
  assign n2909 = pi13 ? n2472 : n2908;
  assign n2910 = pi12 ? n26 : n2909;
  assign n2911 = pi14 ? n376 : n323;
  assign n2912 = pi13 ? n2476 : n2911;
  assign n2913 = pi12 ? n26 : n2912;
  assign n2914 = pi11 ? n2910 : n2913;
  assign n2915 = pi15 ? n41 : n136;
  assign n2916 = pi14 ? n2915 : n323;
  assign n2917 = pi13 ? n2479 : n2916;
  assign n2918 = pi12 ? n26 : n2917;
  assign n2919 = pi14 ? n1480 : n2456;
  assign n2920 = pi14 ? n820 : n323;
  assign n2921 = pi13 ? n2919 : n2920;
  assign n2922 = pi12 ? n26 : n2921;
  assign n2923 = pi11 ? n2918 : n2922;
  assign n2924 = pi10 ? n2914 : n2923;
  assign n2925 = pi14 ? n115 : n2341;
  assign n2926 = pi14 ? n124 : n1202;
  assign n2927 = pi13 ? n2925 : n2926;
  assign n2928 = pi12 ? n26 : n2927;
  assign n2929 = pi11 ? n2928 : n2859;
  assign n2930 = pi14 ? n88 : n1374;
  assign n2931 = pi15 ? n493 : n1814;
  assign n2932 = pi14 ? n348 : n2931;
  assign n2933 = pi13 ? n2930 : n2932;
  assign n2934 = pi12 ? n26 : n2933;
  assign n2935 = pi15 ? n81 : n554;
  assign n2936 = pi14 ? n2935 : n1374;
  assign n2937 = pi17 ? n107 : n224;
  assign n2938 = pi16 ? n2937 : n274;
  assign n2939 = pi15 ? n464 : n2938;
  assign n2940 = pi14 ? n899 : n2939;
  assign n2941 = pi13 ? n2936 : n2940;
  assign n2942 = pi12 ? n26 : n2941;
  assign n2943 = pi11 ? n2934 : n2942;
  assign n2944 = pi10 ? n2929 : n2943;
  assign n2945 = pi09 ? n2924 : n2944;
  assign n2946 = pi08 ? n2459 : n2945;
  assign n2947 = pi07 ? n2462 : n2946;
  assign n2948 = pi15 ? n591 : n96;
  assign n2949 = pi14 ? n2948 : n543;
  assign n2950 = pi13 ? n2949 : n1386;
  assign n2951 = pi12 ? n26 : n2950;
  assign n2952 = pi15 ? n643 : n96;
  assign n2953 = pi15 ? n542 : n377;
  assign n2954 = pi14 ? n2952 : n2953;
  assign n2955 = pi16 ? n1589 : n300;
  assign n2956 = pi15 ? n2955 : n26;
  assign n2957 = pi14 ? n224 : n2956;
  assign n2958 = pi13 ? n2954 : n2957;
  assign n2959 = pi12 ? n26 : n2958;
  assign n2960 = pi11 ? n2951 : n2959;
  assign n2961 = pi15 ? n519 : n122;
  assign n2962 = pi15 ? n542 : n771;
  assign n2963 = pi14 ? n2961 : n2962;
  assign n2964 = pi13 ? n2963 : n2018;
  assign n2965 = pi12 ? n26 : n2964;
  assign n2966 = pi15 ? n229 : n122;
  assign n2967 = pi14 ? n2966 : n899;
  assign n2968 = pi13 ? n2967 : n2025;
  assign n2969 = pi12 ? n26 : n2968;
  assign n2970 = pi11 ? n2965 : n2969;
  assign n2971 = pi10 ? n2960 : n2970;
  assign n2972 = pi13 ? n2037 : n2031;
  assign n2973 = pi12 ? n1880 : n2972;
  assign n2974 = pi12 ? n1921 : n2039;
  assign n2975 = pi11 ? n2973 : n2974;
  assign n2976 = pi10 ? n2975 : n2043;
  assign n2977 = pi09 ? n2971 : n2976;
  assign n2978 = pi08 ? n2977 : n2043;
  assign n2979 = pi14 ? n1374 : n910;
  assign n2980 = pi13 ? n2979 : n2041;
  assign n2981 = pi12 ? n1926 : n2980;
  assign n2982 = pi11 ? n2043 : n2981;
  assign n2983 = pi10 ? n2043 : n2982;
  assign n2984 = pi09 ? n2043 : n2983;
  assign n2985 = pi08 ? n2043 : n2984;
  assign n2986 = pi07 ? n2978 : n2985;
  assign n2987 = pi06 ? n2947 : n2986;
  assign n2988 = pi13 ? n2548 : n2588;
  assign n2989 = pi12 ? n26 : n2988;
  assign n2990 = pi11 ? n26 : n2989;
  assign n2991 = pi13 ? n2554 : n2588;
  assign n2992 = pi12 ? n26 : n2991;
  assign n2993 = pi10 ? n2990 : n2992;
  assign n2994 = pi09 ? n26 : n2993;
  assign n2995 = pi08 ? n26 : n2994;
  assign n2996 = pi11 ? n2992 : n2556;
  assign n2997 = pi10 ? n2992 : n2996;
  assign n2998 = pi09 ? n2992 : n2997;
  assign n2999 = pi15 ? n122 : n2491;
  assign n3000 = pi14 ? n2999 : n2549;
  assign n3001 = pi13 ? n2587 : n3000;
  assign n3002 = pi12 ? n26 : n3001;
  assign n3003 = pi16 ? n128 : n255;
  assign n3004 = pi15 ? n26 : n3003;
  assign n3005 = pi14 ? n3004 : n1400;
  assign n3006 = pi15 ? n122 : n53;
  assign n3007 = pi14 ? n3006 : n2699;
  assign n3008 = pi13 ? n3005 : n3007;
  assign n3009 = pi12 ? n26 : n3008;
  assign n3010 = pi11 ? n3002 : n3009;
  assign n3011 = pi15 ? n26 : n280;
  assign n3012 = pi14 ? n3011 : n1400;
  assign n3013 = pi14 ? n232 : n899;
  assign n3014 = pi13 ? n3012 : n3013;
  assign n3015 = pi12 ? n26 : n3014;
  assign n3016 = pi15 ? n26 : n186;
  assign n3017 = pi14 ? n3016 : n1481;
  assign n3018 = pi13 ? n3017 : n3013;
  assign n3019 = pi12 ? n26 : n3018;
  assign n3020 = pi11 ? n3015 : n3019;
  assign n3021 = pi10 ? n3010 : n3020;
  assign n3022 = pi14 ? n88 : n1533;
  assign n3023 = pi15 ? n979 : n377;
  assign n3024 = pi14 ? n3023 : n840;
  assign n3025 = pi13 ? n3022 : n3024;
  assign n3026 = pi12 ? n26 : n3025;
  assign n3027 = pi14 ? n82 : n1102;
  assign n3028 = pi14 ? n802 : n890;
  assign n3029 = pi13 ? n3027 : n3028;
  assign n3030 = pi12 ? n26 : n3029;
  assign n3031 = pi11 ? n3026 : n3030;
  assign n3032 = pi14 ? n82 : n1607;
  assign n3033 = pi15 ? n60 : n493;
  assign n3034 = pi15 ? n224 : n1216;
  assign n3035 = pi14 ? n3033 : n3034;
  assign n3036 = pi13 ? n3032 : n3035;
  assign n3037 = pi12 ? n26 : n3036;
  assign n3038 = pi16 ? n238 : n26;
  assign n3039 = pi15 ? n224 : n3038;
  assign n3040 = pi14 ? n899 : n3039;
  assign n3041 = pi13 ? n1906 : n3040;
  assign n3042 = pi12 ? n26 : n3041;
  assign n3043 = pi11 ? n3037 : n3042;
  assign n3044 = pi10 ? n3031 : n3043;
  assign n3045 = pi09 ? n3021 : n3044;
  assign n3046 = pi08 ? n2998 : n3045;
  assign n3047 = pi07 ? n2995 : n3046;
  assign n3048 = pi15 ? n1980 : n96;
  assign n3049 = pi16 ? n541 : n60;
  assign n3050 = pi15 ? n122 : n3049;
  assign n3051 = pi14 ? n3048 : n3050;
  assign n3052 = pi13 ? n3051 : n1386;
  assign n3053 = pi12 ? n26 : n3052;
  assign n3054 = pi15 ? n554 : n133;
  assign n3055 = pi14 ? n3054 : n770;
  assign n3056 = pi15 ? n464 : n26;
  assign n3057 = pi14 ? n494 : n3056;
  assign n3058 = pi13 ? n3055 : n3057;
  assign n3059 = pi12 ? n26 : n3058;
  assign n3060 = pi11 ? n3053 : n3059;
  assign n3061 = pi14 ? n1927 : n728;
  assign n3062 = pi15 ? n1064 : n475;
  assign n3063 = pi14 ? n3062 : n2017;
  assign n3064 = pi13 ? n3061 : n3063;
  assign n3065 = pi12 ? n26 : n3064;
  assign n3066 = pi15 ? n722 : n347;
  assign n3067 = pi14 ? n958 : n3066;
  assign n3068 = pi13 ? n3067 : n2119;
  assign n3069 = pi12 ? n1880 : n3068;
  assign n3070 = pi11 ? n3065 : n3069;
  assign n3071 = pi10 ? n3060 : n3070;
  assign n3072 = pi14 ? n1374 : n348;
  assign n3073 = pi13 ? n3072 : n2124;
  assign n3074 = pi12 ? n2088 : n3073;
  assign n3075 = pi14 ? n1607 : n323;
  assign n3076 = pi15 ? n1064 : n1983;
  assign n3077 = pi14 ? n3076 : n26;
  assign n3078 = pi13 ? n3075 : n3077;
  assign n3079 = pi12 ? n1770 : n3078;
  assign n3080 = pi11 ? n3074 : n3079;
  assign n3081 = pi14 ? n1820 : n348;
  assign n3082 = pi13 ? n3081 : n2140;
  assign n3083 = pi12 ? n2099 : n3082;
  assign n3084 = pi13 ? n3081 : n2145;
  assign n3085 = pi12 ? n1101 : n3084;
  assign n3086 = pi11 ? n3083 : n3085;
  assign n3087 = pi10 ? n3080 : n3086;
  assign n3088 = pi09 ? n3071 : n3087;
  assign n3089 = pi08 ? n3088 : n3085;
  assign n3090 = pi12 ? n2153 : n3084;
  assign n3091 = pi13 ? n3081 : n2038;
  assign n3092 = pi12 ? n2153 : n3091;
  assign n3093 = pi11 ? n3090 : n3092;
  assign n3094 = pi14 ? n1820 : n910;
  assign n3095 = pi13 ? n3094 : n2038;
  assign n3096 = pi12 ? n2153 : n3095;
  assign n3097 = pi10 ? n3093 : n3096;
  assign n3098 = pi09 ? n3085 : n3097;
  assign n3099 = pi08 ? n3085 : n3098;
  assign n3100 = pi07 ? n3089 : n3099;
  assign n3101 = pi06 ? n3047 : n3100;
  assign n3102 = pi05 ? n2987 : n3101;
  assign n3103 = pi14 ? n130 : n603;
  assign n3104 = pi13 ? n3103 : n1691;
  assign n3105 = pi12 ? n26 : n3104;
  assign n3106 = pi11 ? n26 : n3105;
  assign n3107 = pi14 ? n130 : n1653;
  assign n3108 = pi13 ? n3107 : n1698;
  assign n3109 = pi12 ? n26 : n3108;
  assign n3110 = pi10 ? n3106 : n3109;
  assign n3111 = pi09 ? n26 : n3110;
  assign n3112 = pi08 ? n26 : n3111;
  assign n3113 = pi14 ? n624 : n1653;
  assign n3114 = pi13 ? n3113 : n1646;
  assign n3115 = pi12 ? n26 : n3114;
  assign n3116 = pi13 ? n1710 : n1646;
  assign n3117 = pi12 ? n26 : n3116;
  assign n3118 = pi11 ? n3115 : n3117;
  assign n3119 = pi13 ? n1710 : n1655;
  assign n3120 = pi12 ? n26 : n3119;
  assign n3121 = pi16 ? n212 : n186;
  assign n3122 = pi15 ? n87 : n3121;
  assign n3123 = pi14 ? n3122 : n2730;
  assign n3124 = pi13 ? n3123 : n1650;
  assign n3125 = pi12 ? n26 : n3124;
  assign n3126 = pi11 ? n3120 : n3125;
  assign n3127 = pi10 ? n3118 : n3126;
  assign n3128 = pi14 ? n1719 : n958;
  assign n3129 = pi14 ? n67 : n2259;
  assign n3130 = pi13 ? n3128 : n3129;
  assign n3131 = pi12 ? n26 : n3130;
  assign n3132 = pi14 ? n101 : n2259;
  assign n3133 = pi13 ? n1856 : n3132;
  assign n3134 = pi12 ? n26 : n3133;
  assign n3135 = pi11 ? n3131 : n3134;
  assign n3136 = pi14 ? n82 : n1820;
  assign n3137 = pi15 ? n224 : n2518;
  assign n3138 = pi14 ? n910 : n3137;
  assign n3139 = pi13 ? n3136 : n3138;
  assign n3140 = pi12 ? n26 : n3139;
  assign n3141 = pi15 ? n34 : n480;
  assign n3142 = pi14 ? n3141 : n1374;
  assign n3143 = pi13 ? n3142 : n1677;
  assign n3144 = pi12 ? n26 : n3143;
  assign n3145 = pi11 ? n3140 : n3144;
  assign n3146 = pi10 ? n3135 : n3145;
  assign n3147 = pi09 ? n3127 : n3146;
  assign n3148 = pi08 ? n3109 : n3147;
  assign n3149 = pi07 ? n3112 : n3148;
  assign n3150 = pi15 ? n34 : n229;
  assign n3151 = pi14 ? n3150 : n3050;
  assign n3152 = pi13 ? n3151 : n2190;
  assign n3153 = pi12 ? n26 : n3152;
  assign n3154 = pi14 ? n3150 : n770;
  assign n3155 = pi15 ? n60 : n741;
  assign n3156 = pi14 ? n3155 : n2198;
  assign n3157 = pi13 ? n3154 : n3156;
  assign n3158 = pi12 ? n26 : n3157;
  assign n3159 = pi11 ? n3153 : n3158;
  assign n3160 = pi14 ? n2197 : n2204;
  assign n3161 = pi13 ? n2209 : n3160;
  assign n3162 = pi12 ? n26 : n3161;
  assign n3163 = pi13 ? n2224 : n2213;
  assign n3164 = pi12 ? n26 : n3163;
  assign n3165 = pi11 ? n3162 : n3164;
  assign n3166 = pi10 ? n3159 : n3165;
  assign n3167 = pi16 ? n1510 : n2210;
  assign n3168 = pi15 ? n60 : n3167;
  assign n3169 = pi14 ? n3168 : n2118;
  assign n3170 = pi13 ? n2224 : n3169;
  assign n3171 = pi12 ? n2088 : n3170;
  assign n3172 = pi12 ? n1770 : n2229;
  assign n3173 = pi11 ? n3171 : n3172;
  assign n3174 = pi14 ? n1206 : n101;
  assign n3175 = pi13 ? n3174 : n2231;
  assign n3176 = pi12 ? n2099 : n3175;
  assign n3177 = pi14 ? n1206 : n2130;
  assign n3178 = pi13 ? n3177 : n2237;
  assign n3179 = pi12 ? n1101 : n3178;
  assign n3180 = pi11 ? n3176 : n3179;
  assign n3181 = pi10 ? n3173 : n3180;
  assign n3182 = pi09 ? n3166 : n3181;
  assign n3183 = pi13 ? n3174 : n2237;
  assign n3184 = pi12 ? n1101 : n3183;
  assign n3185 = pi08 ? n3182 : n3184;
  assign n3186 = pi14 ? n1206 : n1125;
  assign n3187 = pi13 ? n3186 : n2247;
  assign n3188 = pi12 ? n1101 : n3187;
  assign n3189 = pi14 ? n2100 : n1125;
  assign n3190 = pi13 ? n3189 : n2254;
  assign n3191 = pi12 ? n2153 : n3190;
  assign n3192 = pi11 ? n3188 : n3191;
  assign n3193 = pi14 ? n2100 : n101;
  assign n3194 = pi13 ? n3193 : n2260;
  assign n3195 = pi12 ? n1101 : n3194;
  assign n3196 = pi14 ? n2250 : n101;
  assign n3197 = pi13 ? n3196 : n2263;
  assign n3198 = pi12 ? n1101 : n3197;
  assign n3199 = pi11 ? n3195 : n3198;
  assign n3200 = pi10 ? n3192 : n3199;
  assign n3201 = pi09 ? n3184 : n3200;
  assign n3202 = pi08 ? n3184 : n3201;
  assign n3203 = pi07 ? n3185 : n3202;
  assign n3204 = pi06 ? n3149 : n3203;
  assign n3205 = pi16 ? n97 : n41;
  assign n3206 = pi15 ? n32 : n3205;
  assign n3207 = pi14 ? n3206 : n2290;
  assign n3208 = pi13 ? n3207 : n2294;
  assign n3209 = pi12 ? n1101 : n3208;
  assign n3210 = pi11 ? n2289 : n3209;
  assign n3211 = pi14 ? n205 : n980;
  assign n3212 = pi13 ? n3211 : n2302;
  assign n3213 = pi12 ? n1101 : n3212;
  assign n3214 = pi15 ? n1560 : n41;
  assign n3215 = pi14 ? n3214 : n101;
  assign n3216 = pi13 ? n3215 : n2302;
  assign n3217 = pi12 ? n1101 : n3216;
  assign n3218 = pi11 ? n3213 : n3217;
  assign n3219 = pi10 ? n3210 : n3218;
  assign n3220 = pi09 ? n2285 : n3219;
  assign n3221 = pi08 ? n26 : n3220;
  assign n3222 = pi07 ? n26 : n3221;
  assign n3223 = pi06 ? n26 : n3222;
  assign n3224 = pi05 ? n3204 : n3223;
  assign n3225 = pi04 ? n3102 : n3224;
  assign n3226 = pi03 ? n2907 : n3225;
  assign n3227 = pi14 ? n1175 : n2317;
  assign n3228 = pi13 ? n3227 : n2321;
  assign n3229 = pi12 ? n1308 : n3228;
  assign n3230 = pi11 ? n26 : n3229;
  assign n3231 = pi10 ? n26 : n3230;
  assign n3232 = pi14 ? n1763 : n2328;
  assign n3233 = pi13 ? n3232 : n2331;
  assign n3234 = pi12 ? n1315 : n3233;
  assign n3235 = pi11 ? n3234 : n2339;
  assign n3236 = pi10 ? n3235 : n2355;
  assign n3237 = pi09 ? n3231 : n3236;
  assign n3238 = pi08 ? n26 : n3237;
  assign n3239 = pi07 ? n26 : n3238;
  assign n3240 = pi06 ? n26 : n3239;
  assign n3241 = pi13 ? n1176 : n2361;
  assign n3242 = pi12 ? n26 : n3241;
  assign n3243 = pi11 ? n26 : n3242;
  assign n3244 = pi10 ? n3243 : n2367;
  assign n3245 = pi09 ? n26 : n3244;
  assign n3246 = pi08 ? n26 : n3245;
  assign n3247 = pi07 ? n3246 : n2367;
  assign n3248 = pi06 ? n3247 : n2449;
  assign n3249 = pi05 ? n3240 : n3248;
  assign n3250 = pi10 ? n2455 : n2454;
  assign n3251 = pi09 ? n26 : n3250;
  assign n3252 = pi08 ? n26 : n3251;
  assign n3253 = pi07 ? n3252 : n2459;
  assign n3254 = pi06 ? n3253 : n2545;
  assign n3255 = pi14 ? n144 : n1034;
  assign n3256 = pi13 ? n3255 : n1394;
  assign n3257 = pi12 ? n26 : n3256;
  assign n3258 = pi11 ? n26 : n3257;
  assign n3259 = pi16 ? n32 : n563;
  assign n3260 = pi15 ? n32 : n3259;
  assign n3261 = pi14 ? n144 : n3260;
  assign n3262 = pi14 ? n315 : n2656;
  assign n3263 = pi13 ? n3261 : n3262;
  assign n3264 = pi12 ? n26 : n3263;
  assign n3265 = pi14 ? n144 : n2082;
  assign n3266 = pi13 ? n3265 : n2577;
  assign n3267 = pi12 ? n26 : n3266;
  assign n3268 = pi11 ? n3264 : n3267;
  assign n3269 = pi10 ? n3258 : n3268;
  assign n3270 = pi09 ? n26 : n3269;
  assign n3271 = pi08 ? n26 : n3270;
  assign n3272 = pi07 ? n3271 : n2556;
  assign n3273 = pi06 ? n3272 : n2674;
  assign n3274 = pi05 ? n3254 : n3273;
  assign n3275 = pi04 ? n3249 : n3274;
  assign n3276 = pi11 ? n26 : n2696;
  assign n3277 = pi14 ? n130 : n2697;
  assign n3278 = pi14 ? n124 : n1264;
  assign n3279 = pi13 ? n3277 : n3278;
  assign n3280 = pi12 ? n26 : n3279;
  assign n3281 = pi14 ? n124 : n2699;
  assign n3282 = pi13 ? n2698 : n3281;
  assign n3283 = pi12 ? n26 : n3282;
  assign n3284 = pi11 ? n3280 : n3283;
  assign n3285 = pi10 ? n3276 : n3284;
  assign n3286 = pi09 ? n26 : n3285;
  assign n3287 = pi08 ? n26 : n3286;
  assign n3288 = pi14 ? n130 : n386;
  assign n3289 = pi13 ? n3288 : n1698;
  assign n3290 = pi12 ? n26 : n3289;
  assign n3291 = pi10 ? n3290 : n1703;
  assign n3292 = pi09 ? n3291 : n1703;
  assign n3293 = pi08 ? n3292 : n1703;
  assign n3294 = pi07 ? n3287 : n3293;
  assign n3295 = pi06 ? n3294 : n2769;
  assign n3296 = pi14 ? n115 : n685;
  assign n3297 = pi14 ? n924 : n547;
  assign n3298 = pi13 ? n3296 : n3297;
  assign n3299 = pi12 ? n26 : n3298;
  assign n3300 = pi11 ? n26 : n3299;
  assign n3301 = pi15 ? n41 : n2772;
  assign n3302 = pi14 ? n115 : n3301;
  assign n3303 = pi14 ? n124 : n840;
  assign n3304 = pi13 ? n3302 : n3303;
  assign n3305 = pi12 ? n26 : n3304;
  assign n3306 = pi14 ? n115 : n1653;
  assign n3307 = pi14 ? n124 : n224;
  assign n3308 = pi13 ? n3306 : n3307;
  assign n3309 = pi12 ? n26 : n3308;
  assign n3310 = pi11 ? n3305 : n3309;
  assign n3311 = pi10 ? n3300 : n3310;
  assign n3312 = pi09 ? n26 : n3311;
  assign n3313 = pi08 ? n26 : n3312;
  assign n3314 = pi13 ? n2792 : n797;
  assign n3315 = pi12 ? n26 : n3314;
  assign n3316 = pi11 ? n3315 : n2794;
  assign n3317 = pi10 ? n3316 : n26;
  assign n3318 = pi09 ? n3317 : n26;
  assign n3319 = pi08 ? n3318 : n26;
  assign n3320 = pi07 ? n3313 : n3319;
  assign n3321 = pi06 ? n3320 : n26;
  assign n3322 = pi05 ? n3295 : n3321;
  assign n3323 = pi14 ? n105 : n937;
  assign n3324 = pi14 ? n770 : n926;
  assign n3325 = pi13 ? n3323 : n3324;
  assign n3326 = pi12 ? n26 : n3325;
  assign n3327 = pi11 ? n26 : n3326;
  assign n3328 = pi14 ? n105 : n958;
  assign n3329 = pi15 ? n58 : n377;
  assign n3330 = pi14 ? n3329 : n840;
  assign n3331 = pi13 ? n3328 : n3330;
  assign n3332 = pi12 ? n26 : n3331;
  assign n3333 = pi15 ? n58 : n493;
  assign n3334 = pi15 ? n224 : n546;
  assign n3335 = pi14 ? n3333 : n3334;
  assign n3336 = pi13 ? n1588 : n3335;
  assign n3337 = pi12 ? n26 : n3336;
  assign n3338 = pi11 ? n3332 : n3337;
  assign n3339 = pi10 ? n3327 : n3338;
  assign n3340 = pi09 ? n26 : n3339;
  assign n3341 = pi08 ? n26 : n3340;
  assign n3342 = pi14 ? n2819 : n958;
  assign n3343 = pi13 ? n3342 : n1899;
  assign n3344 = pi12 ? n26 : n3343;
  assign n3345 = pi15 ? n934 : n96;
  assign n3346 = pi14 ? n3345 : n2820;
  assign n3347 = pi13 ? n3346 : n2824;
  assign n3348 = pi12 ? n26 : n3347;
  assign n3349 = pi11 ? n3344 : n3348;
  assign n3350 = pi10 ? n3349 : n26;
  assign n3351 = pi09 ? n3350 : n26;
  assign n3352 = pi08 ? n3351 : n26;
  assign n3353 = pi07 ? n3341 : n3352;
  assign n3354 = pi06 ? n3353 : n26;
  assign n3355 = pi15 ? n108 : n122;
  assign n3356 = pi14 ? n88 : n3355;
  assign n3357 = pi14 ? n101 : n1118;
  assign n3358 = pi13 ? n3356 : n3357;
  assign n3359 = pi12 ? n26 : n3358;
  assign n3360 = pi11 ? n26 : n3359;
  assign n3361 = pi15 ? n58 : n66;
  assign n3362 = pi14 ? n3361 : n1852;
  assign n3363 = pi13 ? n1797 : n3362;
  assign n3364 = pi12 ? n26 : n3363;
  assign n3365 = pi15 ? n934 : n32;
  assign n3366 = pi14 ? n3365 : n958;
  assign n3367 = pi15 ? n58 : n771;
  assign n3368 = pi15 ? n464 : n1117;
  assign n3369 = pi14 ? n3367 : n3368;
  assign n3370 = pi13 ? n3366 : n3369;
  assign n3371 = pi12 ? n26 : n3370;
  assign n3372 = pi11 ? n3364 : n3371;
  assign n3373 = pi10 ? n3360 : n3372;
  assign n3374 = pi09 ? n26 : n3373;
  assign n3375 = pi08 ? n26 : n3374;
  assign n3376 = pi14 ? n3345 : n958;
  assign n3377 = pi14 ? n1155 : n1992;
  assign n3378 = pi13 ? n3376 : n3377;
  assign n3379 = pi12 ? n26 : n3378;
  assign n3380 = pi15 ? n1130 : n96;
  assign n3381 = pi14 ? n3380 : n543;
  assign n3382 = pi14 ? n1165 : n2876;
  assign n3383 = pi13 ? n3381 : n3382;
  assign n3384 = pi12 ? n26 : n3383;
  assign n3385 = pi11 ? n3379 : n3384;
  assign n3386 = pi14 ? n1852 : n2881;
  assign n3387 = pi13 ? n2880 : n3386;
  assign n3388 = pi12 ? n26 : n3387;
  assign n3389 = pi15 ? n464 : n678;
  assign n3390 = pi14 ? n3389 : n26;
  assign n3391 = pi13 ? n1936 : n3390;
  assign n3392 = pi12 ? n26 : n3391;
  assign n3393 = pi11 ? n3388 : n3392;
  assign n3394 = pi10 ? n3385 : n3393;
  assign n3395 = pi12 ? n1880 : n1946;
  assign n3396 = pi12 ? n1921 : n1949;
  assign n3397 = pi11 ? n3395 : n3396;
  assign n3398 = pi10 ? n3397 : n1956;
  assign n3399 = pi09 ? n3394 : n3398;
  assign n3400 = pi08 ? n3399 : n1956;
  assign n3401 = pi07 ? n3375 : n3400;
  assign n3402 = pi10 ? n1956 : n1959;
  assign n3403 = pi09 ? n1956 : n3402;
  assign n3404 = pi10 ? n1959 : n1956;
  assign n3405 = pi09 ? n3404 : n1956;
  assign n3406 = pi08 ? n3403 : n3405;
  assign n3407 = pi12 ? n1926 : n1961;
  assign n3408 = pi11 ? n1956 : n3407;
  assign n3409 = pi10 ? n1956 : n3408;
  assign n3410 = pi09 ? n1956 : n3409;
  assign n3411 = pi08 ? n1956 : n3410;
  assign n3412 = pi07 ? n3406 : n3411;
  assign n3413 = pi06 ? n3401 : n3412;
  assign n3414 = pi05 ? n3354 : n3413;
  assign n3415 = pi04 ? n3322 : n3414;
  assign n3416 = pi03 ? n3275 : n3415;
  assign n3417 = pi02 ? n3226 : n3416;
  assign n3418 = pi14 ? n101 : n1348;
  assign n3419 = pi13 ? n1797 : n3418;
  assign n3420 = pi12 ? n26 : n3419;
  assign n3421 = pi16 ? n545 : n1813;
  assign n3422 = pi15 ? n224 : n3421;
  assign n3423 = pi14 ? n1155 : n3422;
  assign n3424 = pi13 ? n3366 : n3423;
  assign n3425 = pi12 ? n26 : n3424;
  assign n3426 = pi11 ? n3420 : n3425;
  assign n3427 = pi10 ? n1796 : n3426;
  assign n3428 = pi09 ? n26 : n3427;
  assign n3429 = pi08 ? n26 : n3428;
  assign n3430 = pi14 ? n2948 : n1616;
  assign n3431 = pi14 ? n899 : n1157;
  assign n3432 = pi13 ? n3430 : n3431;
  assign n3433 = pi12 ? n26 : n3432;
  assign n3434 = pi15 ? n519 : n96;
  assign n3435 = pi14 ? n3434 : n543;
  assign n3436 = pi13 ? n3435 : n1386;
  assign n3437 = pi12 ? n26 : n3436;
  assign n3438 = pi11 ? n3433 : n3437;
  assign n3439 = pi15 ? n643 : n1622;
  assign n3440 = pi14 ? n3439 : n2953;
  assign n3441 = pi13 ? n3440 : n2013;
  assign n3442 = pi12 ? n26 : n3441;
  assign n3443 = pi14 ? n2966 : n2962;
  assign n3444 = pi13 ? n3443 : n2018;
  assign n3445 = pi12 ? n26 : n3444;
  assign n3446 = pi11 ? n3442 : n3445;
  assign n3447 = pi10 ? n3438 : n3446;
  assign n3448 = pi13 ? n2979 : n2025;
  assign n3449 = pi12 ? n1880 : n3448;
  assign n3450 = pi12 ? n1921 : n2972;
  assign n3451 = pi11 ? n3449 : n3450;
  assign n3452 = pi10 ? n3451 : n2044;
  assign n3453 = pi09 ? n3447 : n3452;
  assign n3454 = pi08 ? n3453 : n2043;
  assign n3455 = pi07 ? n3429 : n3454;
  assign n3456 = pi07 ? n2043 : n2985;
  assign n3457 = pi06 ? n3455 : n3456;
  assign n3458 = pi14 ? n523 : n1210;
  assign n3459 = pi13 ? n1890 : n3458;
  assign n3460 = pi12 ? n26 : n3459;
  assign n3461 = pi11 ? n26 : n3460;
  assign n3462 = pi14 ? n316 : n1583;
  assign n3463 = pi13 ? n1856 : n3462;
  assign n3464 = pi12 ? n26 : n3463;
  assign n3465 = pi15 ? n41 : n1162;
  assign n3466 = pi14 ? n1896 : n3465;
  assign n3467 = pi16 ? n1589 : n1215;
  assign n3468 = pi15 ? n464 : n3467;
  assign n3469 = pi14 ? n1155 : n3468;
  assign n3470 = pi13 ? n3466 : n3469;
  assign n3471 = pi12 ? n26 : n3470;
  assign n3472 = pi11 ? n3464 : n3471;
  assign n3473 = pi10 ? n3461 : n3472;
  assign n3474 = pi09 ? n26 : n3473;
  assign n3475 = pi08 ? n26 : n3474;
  assign n3476 = pi15 ? n579 : n705;
  assign n3477 = pi14 ? n3476 : n1616;
  assign n3478 = pi13 ? n3477 : n2000;
  assign n3479 = pi12 ? n26 : n3478;
  assign n3480 = pi15 ? n573 : n229;
  assign n3481 = pi14 ? n3480 : n543;
  assign n3482 = pi13 ? n3481 : n1386;
  assign n3483 = pi12 ? n26 : n3482;
  assign n3484 = pi11 ? n3479 : n3483;
  assign n3485 = pi15 ? n229 : n41;
  assign n3486 = pi14 ? n3485 : n433;
  assign n3487 = pi14 ? n1583 : n1565;
  assign n3488 = pi13 ? n3486 : n3487;
  assign n3489 = pi12 ? n26 : n3488;
  assign n3490 = pi15 ? n229 : n258;
  assign n3491 = pi14 ? n3490 : n728;
  assign n3492 = pi13 ? n3491 : n2109;
  assign n3493 = pi12 ? n1880 : n3492;
  assign n3494 = pi11 ? n3489 : n3493;
  assign n3495 = pi10 ? n3484 : n3494;
  assign n3496 = pi16 ? n224 : n212;
  assign n3497 = pi15 ? n1064 : n3496;
  assign n3498 = pi14 ? n3497 : n2118;
  assign n3499 = pi13 ? n3067 : n3498;
  assign n3500 = pi12 ? n2088 : n3499;
  assign n3501 = pi15 ? n503 : n347;
  assign n3502 = pi14 ? n958 : n3501;
  assign n3503 = pi13 ? n3502 : n2124;
  assign n3504 = pi12 ? n1770 : n3503;
  assign n3505 = pi11 ? n3500 : n3504;
  assign n3506 = pi12 ? n2099 : n3078;
  assign n3507 = pi12 ? n1101 : n3082;
  assign n3508 = pi11 ? n3506 : n3507;
  assign n3509 = pi10 ? n3505 : n3508;
  assign n3510 = pi09 ? n3495 : n3509;
  assign n3511 = pi08 ? n3510 : n3085;
  assign n3512 = pi07 ? n3475 : n3511;
  assign n3513 = pi11 ? n3085 : n3090;
  assign n3514 = pi10 ? n3085 : n3513;
  assign n3515 = pi15 ? n60 : n2655;
  assign n3516 = pi14 ? n1820 : n3515;
  assign n3517 = pi13 ? n3516 : n2038;
  assign n3518 = pi12 ? n2153 : n3517;
  assign n3519 = pi11 ? n3092 : n3518;
  assign n3520 = pi15 ? n546 : n1156;
  assign n3521 = pi14 ? n3520 : n26;
  assign n3522 = pi13 ? n3081 : n3521;
  assign n3523 = pi12 ? n1101 : n3522;
  assign n3524 = pi11 ? n3523 : n3085;
  assign n3525 = pi10 ? n3519 : n3524;
  assign n3526 = pi09 ? n3514 : n3525;
  assign n3527 = pi08 ? n3526 : n3085;
  assign n3528 = pi07 ? n3527 : n3085;
  assign n3529 = pi06 ? n3512 : n3528;
  assign n3530 = pi05 ? n3457 : n3529;
  assign n3531 = pi14 ? n82 : n2166;
  assign n3532 = pi15 ? n1633 : n226;
  assign n3533 = pi14 ? n523 : n3532;
  assign n3534 = pi13 ? n3531 : n3533;
  assign n3535 = pi12 ? n26 : n3534;
  assign n3536 = pi11 ? n26 : n3535;
  assign n3537 = pi15 ? n546 : n1814;
  assign n3538 = pi14 ? n316 : n3537;
  assign n3539 = pi13 ? n1863 : n3538;
  assign n3540 = pi12 ? n26 : n3539;
  assign n3541 = pi14 ? n35 : n1820;
  assign n3542 = pi14 ? n2656 : n1992;
  assign n3543 = pi13 ? n3541 : n3542;
  assign n3544 = pi12 ? n26 : n3543;
  assign n3545 = pi11 ? n3540 : n3544;
  assign n3546 = pi10 ? n3536 : n3545;
  assign n3547 = pi09 ? n26 : n3546;
  assign n3548 = pi08 ? n26 : n3547;
  assign n3549 = pi15 ? n34 : n705;
  assign n3550 = pi14 ? n3549 : n1616;
  assign n3551 = pi14 ? n910 : n1999;
  assign n3552 = pi13 ? n3550 : n3551;
  assign n3553 = pi12 ? n26 : n3552;
  assign n3554 = pi15 ? n34 : n2089;
  assign n3555 = pi14 ? n3554 : n543;
  assign n3556 = pi13 ? n3555 : n1772;
  assign n3557 = pi12 ? n26 : n3556;
  assign n3558 = pi11 ? n3553 : n3557;
  assign n3559 = pi14 ? n3155 : n3056;
  assign n3560 = pi13 ? n2195 : n3559;
  assign n3561 = pi12 ? n26 : n3560;
  assign n3562 = pi14 ? n190 : n427;
  assign n3563 = pi14 ? n2197 : n1932;
  assign n3564 = pi13 ? n3562 : n3563;
  assign n3565 = pi12 ? n26 : n3564;
  assign n3566 = pi11 ? n3561 : n3565;
  assign n3567 = pi10 ? n3558 : n3566;
  assign n3568 = pi12 ? n2088 : n3163;
  assign n3569 = pi12 ? n1770 : n3170;
  assign n3570 = pi11 ? n3568 : n3569;
  assign n3571 = pi12 ? n2099 : n2229;
  assign n3572 = pi11 ? n3571 : n2233;
  assign n3573 = pi10 ? n3570 : n3572;
  assign n3574 = pi09 ? n3567 : n3573;
  assign n3575 = pi11 ? n3179 : n3184;
  assign n3576 = pi10 ? n3575 : n3184;
  assign n3577 = pi09 ? n3576 : n3184;
  assign n3578 = pi08 ? n3574 : n3577;
  assign n3579 = pi07 ? n3548 : n3578;
  assign n3580 = pi13 ? n3186 : n2237;
  assign n3581 = pi12 ? n1101 : n3580;
  assign n3582 = pi11 ? n3581 : n3188;
  assign n3583 = pi10 ? n3184 : n3582;
  assign n3584 = pi15 ? n1064 : n2252;
  assign n3585 = pi14 ? n3584 : n26;
  assign n3586 = pi13 ? n3189 : n3585;
  assign n3587 = pi12 ? n2153 : n3586;
  assign n3588 = pi13 ? n3189 : n2260;
  assign n3589 = pi12 ? n1101 : n3588;
  assign n3590 = pi11 ? n3587 : n3589;
  assign n3591 = pi16 ? n1510 : n224;
  assign n3592 = pi15 ? n3591 : n1758;
  assign n3593 = pi14 ? n3592 : n26;
  assign n3594 = pi13 ? n3193 : n3593;
  assign n3595 = pi12 ? n1101 : n3594;
  assign n3596 = pi11 ? n3595 : n3184;
  assign n3597 = pi10 ? n3590 : n3596;
  assign n3598 = pi09 ? n3583 : n3597;
  assign n3599 = pi16 ? n1510 : n1813;
  assign n3600 = pi15 ? n60 : n3599;
  assign n3601 = pi14 ? n3600 : n26;
  assign n3602 = pi13 ? n3174 : n3601;
  assign n3603 = pi12 ? n1101 : n3602;
  assign n3604 = pi11 ? n3603 : n3184;
  assign n3605 = pi10 ? n3604 : n3184;
  assign n3606 = pi09 ? n3605 : n3184;
  assign n3607 = pi08 ? n3598 : n3606;
  assign n3608 = pi13 ? n3174 : n2247;
  assign n3609 = pi12 ? n1101 : n3608;
  assign n3610 = pi14 ? n2166 : n101;
  assign n3611 = pi16 ? n225 : n1366;
  assign n3612 = pi15 ? n1633 : n3611;
  assign n3613 = pi14 ? n3612 : n26;
  assign n3614 = pi13 ? n3610 : n3613;
  assign n3615 = pi12 ? n1101 : n3614;
  assign n3616 = pi11 ? n3609 : n3615;
  assign n3617 = pi10 ? n3184 : n3616;
  assign n3618 = pi09 ? n3184 : n3617;
  assign n3619 = pi08 ? n3184 : n3618;
  assign n3620 = pi07 ? n3607 : n3619;
  assign n3621 = pi06 ? n3579 : n3620;
  assign n3622 = pi14 ? n323 : n2227;
  assign n3623 = pi13 ? n2286 : n3622;
  assign n3624 = pi12 ? n1101 : n3623;
  assign n3625 = pi11 ? n2283 : n3624;
  assign n3626 = pi10 ? n26 : n3625;
  assign n3627 = pi15 ? n979 : n60;
  assign n3628 = pi14 ? n3206 : n3627;
  assign n3629 = pi14 ? n3584 : n2227;
  assign n3630 = pi13 ? n3628 : n3629;
  assign n3631 = pi12 ? n1101 : n3630;
  assign n3632 = pi16 ? n72 : n41;
  assign n3633 = pi15 ? n32 : n3632;
  assign n3634 = pi14 ? n3633 : n3627;
  assign n3635 = pi13 ? n3634 : n3629;
  assign n3636 = pi12 ? n1101 : n3635;
  assign n3637 = pi11 ? n3631 : n3636;
  assign n3638 = pi10 ? n3637 : n26;
  assign n3639 = pi09 ? n3626 : n3638;
  assign n3640 = pi08 ? n3639 : n26;
  assign n3641 = pi07 ? n3640 : n26;
  assign n3642 = pi06 ? n26 : n3641;
  assign n3643 = pi05 ? n3621 : n3642;
  assign n3644 = pi04 ? n3530 : n3643;
  assign n3645 = pi14 ? n1662 : n2330;
  assign n3646 = pi13 ? n3227 : n3645;
  assign n3647 = pi12 ? n1308 : n3646;
  assign n3648 = pi11 ? n3647 : n3234;
  assign n3649 = pi10 ? n26 : n3648;
  assign n3650 = pi15 ? n477 : n133;
  assign n3651 = pi14 ? n3650 : n2335;
  assign n3652 = pi14 ? n899 : n2347;
  assign n3653 = pi13 ? n3651 : n3652;
  assign n3654 = pi12 ? n1101 : n3653;
  assign n3655 = pi14 ? n1561 : n2276;
  assign n3656 = pi13 ? n3655 : n2348;
  assign n3657 = pi12 ? n1101 : n3656;
  assign n3658 = pi11 ? n3654 : n3657;
  assign n3659 = pi10 ? n3658 : n26;
  assign n3660 = pi09 ? n3649 : n3659;
  assign n3661 = pi08 ? n3660 : n26;
  assign n3662 = pi07 ? n3661 : n26;
  assign n3663 = pi06 ? n26 : n3662;
  assign n3664 = pi10 ? n3243 : n2835;
  assign n3665 = pi09 ? n26 : n3664;
  assign n3666 = pi08 ? n26 : n3665;
  assign n3667 = pi14 ? n1186 : n2383;
  assign n3668 = pi13 ? n426 : n3667;
  assign n3669 = pi12 ? n26 : n3668;
  assign n3670 = pi11 ? n2835 : n3669;
  assign n3671 = pi14 ? n74 : n292;
  assign n3672 = pi13 ? n2382 : n3671;
  assign n3673 = pi12 ? n26 : n3672;
  assign n3674 = pi13 ? n2393 : n2400;
  assign n3675 = pi12 ? n26 : n3674;
  assign n3676 = pi11 ? n3673 : n3675;
  assign n3677 = pi10 ? n3670 : n3676;
  assign n3678 = pi09 ? n2835 : n3677;
  assign n3679 = pi08 ? n2835 : n3678;
  assign n3680 = pi07 ? n3666 : n3679;
  assign n3681 = pi15 ? n62 : n26;
  assign n3682 = pi14 ? n1193 : n3681;
  assign n3683 = pi13 ? n2398 : n3682;
  assign n3684 = pi12 ? n26 : n3683;
  assign n3685 = pi15 ? n250 : n157;
  assign n3686 = pi14 ? n3685 : n1200;
  assign n3687 = pi13 ? n3686 : n2408;
  assign n3688 = pi12 ? n26 : n3687;
  assign n3689 = pi11 ? n3684 : n3688;
  assign n3690 = pi14 ? n425 : n2317;
  assign n3691 = pi15 ? n62 : n347;
  assign n3692 = pi14 ? n3691 : n2320;
  assign n3693 = pi13 ? n3690 : n3692;
  assign n3694 = pi12 ? n1539 : n3693;
  assign n3695 = pi15 ? n456 : n32;
  assign n3696 = pi16 ? n32 : n148;
  assign n3697 = pi15 ? n3696 : n2418;
  assign n3698 = pi14 ? n3695 : n3697;
  assign n3699 = pi14 ? n66 : n2320;
  assign n3700 = pi13 ? n3698 : n3699;
  assign n3701 = pi12 ? n1770 : n3700;
  assign n3702 = pi11 ? n3694 : n3701;
  assign n3703 = pi10 ? n3689 : n3702;
  assign n3704 = pi14 ? n117 : n2335;
  assign n3705 = pi15 ? n66 : n224;
  assign n3706 = pi14 ? n3705 : n2437;
  assign n3707 = pi13 ? n3704 : n3706;
  assign n3708 = pi12 ? n1315 : n3707;
  assign n3709 = pi14 ? n1653 : n2335;
  assign n3710 = pi13 ? n3709 : n2438;
  assign n3711 = pi12 ? n2441 : n3710;
  assign n3712 = pi11 ? n3708 : n3711;
  assign n3713 = pi16 ? n2274 : n135;
  assign n3714 = pi15 ? n3713 : n493;
  assign n3715 = pi14 ? n1927 : n3714;
  assign n3716 = pi14 ? n840 : n2118;
  assign n3717 = pi13 ? n3715 : n3716;
  assign n3718 = pi12 ? n522 : n3717;
  assign n3719 = pi14 ? n2820 : n494;
  assign n3720 = pi15 ? n464 : n2822;
  assign n3721 = pi14 ? n3720 : n26;
  assign n3722 = pi13 ? n3719 : n3721;
  assign n3723 = pi12 ? n522 : n3722;
  assign n3724 = pi11 ? n3718 : n3723;
  assign n3725 = pi10 ? n3712 : n3724;
  assign n3726 = pi09 ? n3703 : n3725;
  assign n3727 = pi12 ? n1926 : n2898;
  assign n3728 = pi11 ? n1950 : n3727;
  assign n3729 = pi10 ? n3728 : n1956;
  assign n3730 = pi09 ? n3729 : n1956;
  assign n3731 = pi08 ? n3726 : n3730;
  assign n3732 = pi07 ? n3731 : n3411;
  assign n3733 = pi06 ? n3680 : n3732;
  assign n3734 = pi05 ? n3663 : n3733;
  assign n3735 = pi13 ? n2476 : n2481;
  assign n3736 = pi12 ? n26 : n3735;
  assign n3737 = pi11 ? n2474 : n3736;
  assign n3738 = pi15 ? n60 : n291;
  assign n3739 = pi14 ? n2492 : n3738;
  assign n3740 = pi13 ? n2479 : n3739;
  assign n3741 = pi12 ? n26 : n3740;
  assign n3742 = pi14 ? n1411 : n2499;
  assign n3743 = pi13 ? n2490 : n3742;
  assign n3744 = pi12 ? n26 : n3743;
  assign n3745 = pi11 ? n3741 : n3744;
  assign n3746 = pi10 ? n3737 : n3745;
  assign n3747 = pi09 ? n2459 : n3746;
  assign n3748 = pi08 ? n2459 : n3747;
  assign n3749 = pi07 ? n3252 : n3748;
  assign n3750 = pi15 ? n405 : n178;
  assign n3751 = pi14 ? n3750 : n2456;
  assign n3752 = pi15 ? n60 : n26;
  assign n3753 = pi14 ? n820 : n3752;
  assign n3754 = pi13 ? n3751 : n3753;
  assign n3755 = pi12 ? n26 : n3754;
  assign n3756 = pi15 ? n701 : n997;
  assign n3757 = pi14 ? n3756 : n2341;
  assign n3758 = pi14 ? n124 : n3752;
  assign n3759 = pi13 ? n3757 : n3758;
  assign n3760 = pi12 ? n26 : n3759;
  assign n3761 = pi11 ? n3755 : n3760;
  assign n3762 = pi15 ? n62 : n60;
  assign n3763 = pi14 ? n3762 : n2320;
  assign n3764 = pi13 ? n2510 : n3763;
  assign n3765 = pi12 ? n26 : n3764;
  assign n3766 = pi16 ? n1589 : n452;
  assign n3767 = pi15 ? n3766 : n32;
  assign n3768 = pi15 ? n705 : n122;
  assign n3769 = pi14 ? n3767 : n3768;
  assign n3770 = pi15 ? n1661 : n60;
  assign n3771 = pi16 ? n60 : n274;
  assign n3772 = pi15 ? n3771 : n26;
  assign n3773 = pi14 ? n3770 : n3772;
  assign n3774 = pi13 ? n3769 : n3773;
  assign n3775 = pi12 ? n1770 : n3774;
  assign n3776 = pi11 ? n3765 : n3775;
  assign n3777 = pi10 ? n3761 : n3776;
  assign n3778 = pi14 ? n2697 : n723;
  assign n3779 = pi14 ? n910 : n2437;
  assign n3780 = pi13 ? n3778 : n3779;
  assign n3781 = pi12 ? n2526 : n3780;
  assign n3782 = pi11 ? n3781 : n2540;
  assign n3783 = pi15 ? n41 : n1622;
  assign n3784 = pi14 ? n3783 : n2953;
  assign n3785 = pi13 ? n3784 : n2302;
  assign n3786 = pi12 ? n1926 : n3785;
  assign n3787 = pi14 ? n958 : n2962;
  assign n3788 = pi14 ? n890 : n2118;
  assign n3789 = pi13 ? n3787 : n3788;
  assign n3790 = pi12 ? n1926 : n3789;
  assign n3791 = pi11 ? n3786 : n3790;
  assign n3792 = pi10 ? n3782 : n3791;
  assign n3793 = pi09 ? n3777 : n3792;
  assign n3794 = pi14 ? n958 : n899;
  assign n3795 = pi15 ? n224 : n2138;
  assign n3796 = pi14 ? n3795 : n26;
  assign n3797 = pi13 ? n3794 : n3796;
  assign n3798 = pi12 ? n1926 : n3797;
  assign n3799 = pi11 ? n3798 : n2040;
  assign n3800 = pi10 ? n3799 : n2043;
  assign n3801 = pi09 ? n3800 : n2043;
  assign n3802 = pi08 ? n3793 : n3801;
  assign n3803 = pi07 ? n3802 : n2985;
  assign n3804 = pi06 ? n3749 : n3803;
  assign n3805 = pi14 ? n365 : n1393;
  assign n3806 = pi13 ? n852 : n3805;
  assign n3807 = pi12 ? n26 : n3806;
  assign n3808 = pi11 ? n26 : n3807;
  assign n3809 = pi14 ? n365 : n2656;
  assign n3810 = pi13 ? n3265 : n3809;
  assign n3811 = pi12 ? n26 : n3810;
  assign n3812 = pi14 ? n365 : n2576;
  assign n3813 = pi13 ? n3265 : n3812;
  assign n3814 = pi12 ? n26 : n3813;
  assign n3815 = pi11 ? n3811 : n3814;
  assign n3816 = pi10 ? n3808 : n3815;
  assign n3817 = pi09 ? n26 : n3816;
  assign n3818 = pi08 ? n26 : n3817;
  assign n3819 = pi15 ? n123 : n2593;
  assign n3820 = pi14 ? n315 : n3819;
  assign n3821 = pi13 ? n2587 : n3820;
  assign n3822 = pi12 ? n26 : n3821;
  assign n3823 = pi15 ? n123 : n2601;
  assign n3824 = pi14 ? n365 : n3823;
  assign n3825 = pi13 ? n2592 : n3824;
  assign n3826 = pi12 ? n26 : n3825;
  assign n3827 = pi11 ? n3822 : n3826;
  assign n3828 = pi14 ? n2999 : n2613;
  assign n3829 = pi13 ? n2600 : n3828;
  assign n3830 = pi12 ? n26 : n3829;
  assign n3831 = pi13 ? n2611 : n2622;
  assign n3832 = pi12 ? n26 : n3831;
  assign n3833 = pi11 ? n3830 : n3832;
  assign n3834 = pi10 ? n3827 : n3833;
  assign n3835 = pi09 ? n2992 : n3834;
  assign n3836 = pi08 ? n2992 : n3835;
  assign n3837 = pi07 ? n3818 : n3836;
  assign n3838 = pi16 ? n32 : n156;
  assign n3839 = pi15 ? n405 : n3838;
  assign n3840 = pi15 ? n73 : n1836;
  assign n3841 = pi14 ? n3839 : n3840;
  assign n3842 = pi15 ? n60 : n2346;
  assign n3843 = pi14 ? n124 : n3842;
  assign n3844 = pi13 ? n3841 : n3843;
  assign n3845 = pi12 ? n26 : n3844;
  assign n3846 = pi15 ? n2737 : n32;
  assign n3847 = pi14 ? n3846 : n190;
  assign n3848 = pi15 ? n122 : n992;
  assign n3849 = pi14 ? n3848 : n2499;
  assign n3850 = pi13 ? n3847 : n3849;
  assign n3851 = pi12 ? n26 : n3850;
  assign n3852 = pi11 ? n3845 : n3851;
  assign n3853 = pi15 ? n493 : n26;
  assign n3854 = pi14 ? n1125 : n3853;
  assign n3855 = pi13 ? n2634 : n3854;
  assign n3856 = pi12 ? n26 : n3855;
  assign n3857 = pi15 ? n705 : n231;
  assign n3858 = pi14 ? n32 : n3857;
  assign n3859 = pi15 ? n123 : n60;
  assign n3860 = pi14 ? n3859 : n2198;
  assign n3861 = pi13 ? n3858 : n3860;
  assign n3862 = pi12 ? n1539 : n3861;
  assign n3863 = pi11 ? n3856 : n3862;
  assign n3864 = pi10 ? n3852 : n3863;
  assign n3865 = pi15 ? n573 : n32;
  assign n3866 = pi16 ? n502 : n121;
  assign n3867 = pi15 ? n122 : n3866;
  assign n3868 = pi14 ? n3865 : n3867;
  assign n3869 = pi15 ? n123 : n3591;
  assign n3870 = pi14 ? n3869 : n2204;
  assign n3871 = pi13 ? n3868 : n3870;
  assign n3872 = pi12 ? n2651 : n3871;
  assign n3873 = pi15 ? n573 : n705;
  assign n3874 = pi14 ? n3873 : n723;
  assign n3875 = pi17 ? n224 : n60;
  assign n3876 = pi16 ? n60 : n3875;
  assign n3877 = pi15 ? n3876 : n224;
  assign n3878 = pi14 ? n3877 : n2204;
  assign n3879 = pi13 ? n3874 : n3878;
  assign n3880 = pi12 ? n1315 : n3879;
  assign n3881 = pi11 ? n3872 : n3880;
  assign n3882 = pi14 ? n1997 : n433;
  assign n3883 = pi13 ? n3882 : n2438;
  assign n3884 = pi12 ? n1101 : n3883;
  assign n3885 = pi15 ? n573 : n936;
  assign n3886 = pi14 ? n3885 : n728;
  assign n3887 = pi14 ? n1165 : n2227;
  assign n3888 = pi13 ? n3886 : n3887;
  assign n3889 = pi12 ? n1101 : n3888;
  assign n3890 = pi11 ? n3884 : n3889;
  assign n3891 = pi10 ? n3881 : n3890;
  assign n3892 = pi09 ? n3864 : n3891;
  assign n3893 = pi14 ? n3062 : n2118;
  assign n3894 = pi13 ? n3067 : n3893;
  assign n3895 = pi12 ? n1101 : n3894;
  assign n3896 = pi15 ? n923 : n347;
  assign n3897 = pi14 ? n958 : n3896;
  assign n3898 = pi17 ? n32 : n355;
  assign n3899 = pi16 ? n224 : n3898;
  assign n3900 = pi15 ? n1064 : n3899;
  assign n3901 = pi14 ? n3900 : n26;
  assign n3902 = pi13 ? n3897 : n3901;
  assign n3903 = pi12 ? n1101 : n3902;
  assign n3904 = pi11 ? n3895 : n3903;
  assign n3905 = pi13 ? n3075 : n2140;
  assign n3906 = pi12 ? n1101 : n3905;
  assign n3907 = pi11 ? n3906 : n3085;
  assign n3908 = pi10 ? n3904 : n3907;
  assign n3909 = pi09 ? n3908 : n3085;
  assign n3910 = pi08 ? n3892 : n3909;
  assign n3911 = pi07 ? n3910 : n3085;
  assign n3912 = pi06 ? n3837 : n3911;
  assign n3913 = pi05 ? n3804 : n3912;
  assign n3914 = pi04 ? n3734 : n3913;
  assign n3915 = pi03 ? n3644 : n3914;
  assign n3916 = pi14 ? n130 : n134;
  assign n3917 = pi13 ? n3916 : n1036;
  assign n3918 = pi12 ? n26 : n3917;
  assign n3919 = pi11 ? n26 : n3918;
  assign n3920 = pi14 ? n130 : n783;
  assign n3921 = pi13 ? n3920 : n2694;
  assign n3922 = pi12 ? n26 : n3921;
  assign n3923 = pi14 ? n1044 : n783;
  assign n3924 = pi13 ? n3923 : n2700;
  assign n3925 = pi12 ? n26 : n3924;
  assign n3926 = pi11 ? n3922 : n3925;
  assign n3927 = pi10 ? n3919 : n3926;
  assign n3928 = pi09 ? n26 : n3927;
  assign n3929 = pi08 ? n26 : n3928;
  assign n3930 = pi14 ? n130 : n41;
  assign n3931 = pi13 ? n3930 : n1698;
  assign n3932 = pi12 ? n26 : n3931;
  assign n3933 = pi10 ? n3932 : n3109;
  assign n3934 = pi09 ? n3933 : n3109;
  assign n3935 = pi14 ? n383 : n1653;
  assign n3936 = pi14 ? n387 : n2253;
  assign n3937 = pi13 ? n3935 : n3936;
  assign n3938 = pi12 ? n26 : n3937;
  assign n3939 = pi14 ? n137 : n1668;
  assign n3940 = pi13 ? n2713 : n3939;
  assign n3941 = pi12 ? n26 : n3940;
  assign n3942 = pi11 ? n3938 : n3941;
  assign n3943 = pi13 ? n1710 : n2726;
  assign n3944 = pi12 ? n26 : n3943;
  assign n3945 = pi13 ? n2724 : n2733;
  assign n3946 = pi12 ? n26 : n3945;
  assign n3947 = pi11 ? n3944 : n3946;
  assign n3948 = pi10 ? n3942 : n3947;
  assign n3949 = pi09 ? n3109 : n3948;
  assign n3950 = pi08 ? n3934 : n3949;
  assign n3951 = pi07 ? n3929 : n3950;
  assign n3952 = pi15 ? n81 : n187;
  assign n3953 = pi15 ? n41 : n1836;
  assign n3954 = pi14 ? n3952 : n3953;
  assign n3955 = pi14 ? n770 : n2732;
  assign n3956 = pi13 ? n3954 : n3955;
  assign n3957 = pi12 ? n26 : n3956;
  assign n3958 = pi15 ? n34 : n808;
  assign n3959 = pi14 ? n3958 : n41;
  assign n3960 = pi14 ? n770 : n3853;
  assign n3961 = pi13 ? n3959 : n3960;
  assign n3962 = pi12 ? n26 : n3961;
  assign n3963 = pi11 ? n3957 : n3962;
  assign n3964 = pi14 ? n1175 : n958;
  assign n3965 = pi14 ? n101 : n2198;
  assign n3966 = pi13 ? n3964 : n3965;
  assign n3967 = pi12 ? n26 : n3966;
  assign n3968 = pi14 ? n2136 : n2198;
  assign n3969 = pi13 ? n2753 : n3968;
  assign n3970 = pi12 ? n2088 : n3969;
  assign n3971 = pi11 ? n3967 : n3970;
  assign n3972 = pi10 ? n3963 : n3971;
  assign n3973 = pi15 ? n477 : n554;
  assign n3974 = pi14 ? n3973 : n958;
  assign n3975 = pi14 ? n1393 : n2204;
  assign n3976 = pi13 ? n3974 : n3975;
  assign n3977 = pi12 ? n1770 : n3976;
  assign n3978 = pi12 ? n2099 : n2759;
  assign n3979 = pi11 ? n3977 : n3978;
  assign n3980 = pi14 ? n685 : n770;
  assign n3981 = pi14 ? n3155 : n2437;
  assign n3982 = pi13 ? n3980 : n3981;
  assign n3983 = pi12 ? n1101 : n3982;
  assign n3984 = pi16 ? n788 : n58;
  assign n3985 = pi15 ? n3984 : n66;
  assign n3986 = pi14 ? n685 : n3985;
  assign n3987 = pi14 ? n2197 : n2437;
  assign n3988 = pi13 ? n3986 : n3987;
  assign n3989 = pi12 ? n1101 : n3988;
  assign n3990 = pi11 ? n3983 : n3989;
  assign n3991 = pi10 ? n3979 : n3990;
  assign n3992 = pi09 ? n3972 : n3991;
  assign n3993 = pi15 ? n542 : n66;
  assign n3994 = pi14 ? n1206 : n3993;
  assign n3995 = pi13 ? n3994 : n2213;
  assign n3996 = pi12 ? n1101 : n3995;
  assign n3997 = pi13 ? n3994 : n3169;
  assign n3998 = pi12 ? n1101 : n3997;
  assign n3999 = pi11 ? n3996 : n3998;
  assign n4000 = pi13 ? n3994 : n2231;
  assign n4001 = pi12 ? n1101 : n4000;
  assign n4002 = pi11 ? n4001 : n2239;
  assign n4003 = pi10 ? n3999 : n4002;
  assign n4004 = pi09 ? n4003 : n3576;
  assign n4005 = pi08 ? n3992 : n4004;
  assign n4006 = pi07 ? n4005 : n3619;
  assign n4007 = pi06 ? n3951 : n4006;
  assign n4008 = pi14 ? n115 : n117;
  assign n4009 = pi13 ? n4008 : n834;
  assign n4010 = pi12 ? n26 : n4009;
  assign n4011 = pi11 ? n26 : n4010;
  assign n4012 = pi14 ? n115 : n783;
  assign n4013 = pi13 ? n4012 : n931;
  assign n4014 = pi12 ? n26 : n4013;
  assign n4015 = pi14 ? n115 : n41;
  assign n4016 = pi13 ? n4015 : n776;
  assign n4017 = pi12 ? n26 : n4016;
  assign n4018 = pi11 ? n4014 : n4017;
  assign n4019 = pi10 ? n4011 : n4018;
  assign n4020 = pi09 ? n26 : n4019;
  assign n4021 = pi08 ? n26 : n4020;
  assign n4022 = pi07 ? n4021 : n3319;
  assign n4023 = pi06 ? n4022 : n26;
  assign n4024 = pi05 ? n4007 : n4023;
  assign n4025 = pi14 ? n124 : n926;
  assign n4026 = pi13 ? n3323 : n4025;
  assign n4027 = pi12 ? n26 : n4026;
  assign n4028 = pi11 ? n26 : n4027;
  assign n4029 = pi14 ? n105 : n948;
  assign n4030 = pi13 ? n4029 : n3330;
  assign n4031 = pi12 ? n26 : n4030;
  assign n4032 = pi14 ? n1587 : n41;
  assign n4033 = pi14 ? n3333 : n939;
  assign n4034 = pi13 ? n4032 : n4033;
  assign n4035 = pi12 ? n26 : n4034;
  assign n4036 = pi11 ? n4031 : n4035;
  assign n4037 = pi10 ? n4028 : n4036;
  assign n4038 = pi09 ? n26 : n4037;
  assign n4039 = pi08 ? n26 : n4038;
  assign n4040 = pi15 ? n43 : n133;
  assign n4041 = pi14 ? n4040 : n958;
  assign n4042 = pi13 ? n4041 : n1899;
  assign n4043 = pi12 ? n26 : n4042;
  assign n4044 = pi14 ? n1605 : n2820;
  assign n4045 = pi13 ? n4044 : n2824;
  assign n4046 = pi12 ? n26 : n4045;
  assign n4047 = pi11 ? n4043 : n4046;
  assign n4048 = pi10 ? n4047 : n26;
  assign n4049 = pi09 ? n4048 : n26;
  assign n4050 = pi08 ? n4049 : n26;
  assign n4051 = pi07 ? n4039 : n4050;
  assign n4052 = pi06 ? n4051 : n26;
  assign n4053 = pi14 ? n3361 : n1348;
  assign n4054 = pi13 ? n1797 : n4053;
  assign n4055 = pi12 ? n26 : n4054;
  assign n4056 = pi13 ? n1802 : n3369;
  assign n4057 = pi12 ? n26 : n4056;
  assign n4058 = pi11 ? n4055 : n4057;
  assign n4059 = pi10 ? n3360 : n4058;
  assign n4060 = pi09 ? n26 : n4059;
  assign n4061 = pi08 ? n26 : n4060;
  assign n4062 = pi14 ? n1605 : n958;
  assign n4063 = pi13 ? n4062 : n1158;
  assign n4064 = pi12 ? n26 : n4063;
  assign n4065 = pi15 ? n475 : n1168;
  assign n4066 = pi14 ? n1165 : n4065;
  assign n4067 = pi13 ? n3381 : n4066;
  assign n4068 = pi12 ? n26 : n4067;
  assign n4069 = pi11 ? n4064 : n4068;
  assign n4070 = pi10 ? n4069 : n3393;
  assign n4071 = pi14 ? n26 : n1153;
  assign n4072 = pi13 ? n26 : n4071;
  assign n4073 = pi16 ? n175 : n300;
  assign n4074 = pi15 ? n475 : n4073;
  assign n4075 = pi14 ? n4074 : n26;
  assign n4076 = pi13 ? n1936 : n4075;
  assign n4077 = pi12 ? n4072 : n4076;
  assign n4078 = pi15 ? n26 : n643;
  assign n4079 = pi14 ? n26 : n4078;
  assign n4080 = pi13 ? n26 : n4079;
  assign n4081 = pi12 ? n4080 : n1949;
  assign n4082 = pi11 ? n4077 : n4081;
  assign n4083 = pi12 ? n909 : n1955;
  assign n4084 = pi15 ? n464 : n1384;
  assign n4085 = pi14 ? n4084 : n26;
  assign n4086 = pi13 ? n1936 : n4085;
  assign n4087 = pi12 ? n909 : n4086;
  assign n4088 = pi11 ? n4083 : n4087;
  assign n4089 = pi10 ? n4082 : n4088;
  assign n4090 = pi09 ? n4070 : n4089;
  assign n4091 = pi12 ? n909 : n2898;
  assign n4092 = pi10 ? n4091 : n4083;
  assign n4093 = pi09 ? n4092 : n4083;
  assign n4094 = pi08 ? n4090 : n4093;
  assign n4095 = pi07 ? n4061 : n4094;
  assign n4096 = pi12 ? n909 : n1961;
  assign n4097 = pi11 ? n4083 : n4096;
  assign n4098 = pi10 ? n4083 : n4097;
  assign n4099 = pi09 ? n4083 : n4098;
  assign n4100 = pi08 ? n4083 : n4099;
  assign n4101 = pi07 ? n4083 : n4100;
  assign n4102 = pi06 ? n4095 : n4101;
  assign n4103 = pi05 ? n4052 : n4102;
  assign n4104 = pi04 ? n4024 : n4103;
  assign n4105 = pi16 ? n1589 : n1813;
  assign n4106 = pi15 ? n224 : n4105;
  assign n4107 = pi14 ? n1155 : n4106;
  assign n4108 = pi13 ? n1856 : n4107;
  assign n4109 = pi12 ? n26 : n4108;
  assign n4110 = pi11 ? n3420 : n4109;
  assign n4111 = pi10 ? n1796 : n4110;
  assign n4112 = pi09 ? n26 : n4111;
  assign n4113 = pi08 ? n26 : n4112;
  assign n4114 = pi14 ? n3345 : n1374;
  assign n4115 = pi13 ? n4114 : n3431;
  assign n4116 = pi12 ? n26 : n4115;
  assign n4117 = pi13 ? n3381 : n1386;
  assign n4118 = pi12 ? n26 : n4117;
  assign n4119 = pi11 ? n4116 : n4118;
  assign n4120 = pi15 ? n789 : n1622;
  assign n4121 = pi14 ? n4120 : n2953;
  assign n4122 = pi13 ? n4121 : n2013;
  assign n4123 = pi12 ? n26 : n4122;
  assign n4124 = pi15 ? n464 : n475;
  assign n4125 = pi14 ? n4124 : n2017;
  assign n4126 = pi13 ? n3443 : n4125;
  assign n4127 = pi12 ? n1880 : n4126;
  assign n4128 = pi11 ? n4123 : n4127;
  assign n4129 = pi10 ? n4119 : n4128;
  assign n4130 = pi16 ? n42 : n96;
  assign n4131 = pi15 ? n26 : n4130;
  assign n4132 = pi14 ? n26 : n4131;
  assign n4133 = pi13 ? n26 : n4132;
  assign n4134 = pi14 ? n1607 : n899;
  assign n4135 = pi14 ? n475 : n26;
  assign n4136 = pi13 ? n4134 : n4135;
  assign n4137 = pi12 ? n4133 : n4136;
  assign n4138 = pi14 ? n1820 : n899;
  assign n4139 = pi15 ? n475 : n2138;
  assign n4140 = pi14 ? n4139 : n26;
  assign n4141 = pi13 ? n4138 : n4140;
  assign n4142 = pi12 ? n1926 : n4141;
  assign n4143 = pi11 ? n4137 : n4142;
  assign n4144 = pi14 ? n1912 : n26;
  assign n4145 = pi13 ? n4138 : n4144;
  assign n4146 = pi12 ? n1926 : n4145;
  assign n4147 = pi13 ? n4138 : n2041;
  assign n4148 = pi12 ? n1926 : n4147;
  assign n4149 = pi11 ? n4146 : n4148;
  assign n4150 = pi10 ? n4143 : n4149;
  assign n4151 = pi09 ? n4129 : n4150;
  assign n4152 = pi08 ? n4151 : n4148;
  assign n4153 = pi07 ? n4113 : n4152;
  assign n4154 = pi13 ? n3094 : n2041;
  assign n4155 = pi12 ? n1926 : n4154;
  assign n4156 = pi11 ? n4148 : n4155;
  assign n4157 = pi10 ? n4148 : n4156;
  assign n4158 = pi09 ? n4148 : n4157;
  assign n4159 = pi08 ? n4148 : n4158;
  assign n4160 = pi07 ? n4148 : n4159;
  assign n4161 = pi06 ? n4153 : n4160;
  assign n4162 = pi14 ? n3380 : n1616;
  assign n4163 = pi13 ? n4162 : n2000;
  assign n4164 = pi12 ? n26 : n4163;
  assign n4165 = pi14 ? n96 : n543;
  assign n4166 = pi13 ? n4165 : n1386;
  assign n4167 = pi12 ? n26 : n4166;
  assign n4168 = pi11 ? n4164 : n4167;
  assign n4169 = pi15 ? n1606 : n60;
  assign n4170 = pi14 ? n41 : n4169;
  assign n4171 = pi15 ? n771 : n475;
  assign n4172 = pi14 ? n4171 : n1565;
  assign n4173 = pi13 ? n4170 : n4172;
  assign n4174 = pi12 ? n1880 : n4173;
  assign n4175 = pi14 ? n958 : n1325;
  assign n4176 = pi14 ? n1852 : n2017;
  assign n4177 = pi13 ? n4175 : n4176;
  assign n4178 = pi12 ? n1921 : n4177;
  assign n4179 = pi11 ? n4174 : n4178;
  assign n4180 = pi10 ? n4168 : n4179;
  assign n4181 = pi16 ? n518 : n563;
  assign n4182 = pi15 ? n26 : n4181;
  assign n4183 = pi14 ? n26 : n4182;
  assign n4184 = pi13 ? n26 : n4183;
  assign n4185 = pi16 ? n251 : n2210;
  assign n4186 = pi15 ? n224 : n4185;
  assign n4187 = pi14 ? n4186 : n2118;
  assign n4188 = pi13 ? n3787 : n4187;
  assign n4189 = pi12 ? n4184 : n4188;
  assign n4190 = pi15 ? n923 : n771;
  assign n4191 = pi14 ? n958 : n4190;
  assign n4192 = pi16 ? n251 : n276;
  assign n4193 = pi15 ? n224 : n4192;
  assign n4194 = pi14 ? n4193 : n26;
  assign n4195 = pi13 ? n4191 : n4194;
  assign n4196 = pi12 ? n1926 : n4195;
  assign n4197 = pi11 ? n4189 : n4196;
  assign n4198 = pi17 ? n297 : n355;
  assign n4199 = pi16 ? n224 : n4198;
  assign n4200 = pi15 ? n224 : n4199;
  assign n4201 = pi14 ? n4200 : n26;
  assign n4202 = pi13 ? n2979 : n4201;
  assign n4203 = pi12 ? n2153 : n4202;
  assign n4204 = pi12 ? n2153 : n2039;
  assign n4205 = pi11 ? n4203 : n4204;
  assign n4206 = pi10 ? n4197 : n4205;
  assign n4207 = pi09 ? n4180 : n4206;
  assign n4208 = pi08 ? n4207 : n4204;
  assign n4209 = pi07 ? n3475 : n4208;
  assign n4210 = pi13 ? n2979 : n2038;
  assign n4211 = pi12 ? n2153 : n4210;
  assign n4212 = pi11 ? n4204 : n4211;
  assign n4213 = pi10 ? n4204 : n4212;
  assign n4214 = pi09 ? n4204 : n4213;
  assign n4215 = pi08 ? n4204 : n4214;
  assign n4216 = pi07 ? n4204 : n4215;
  assign n4217 = pi06 ? n4209 : n4216;
  assign n4218 = pi05 ? n4161 : n4217;
  assign n4219 = pi14 ? n323 : n3537;
  assign n4220 = pi13 ? n1863 : n4219;
  assign n4221 = pi12 ? n26 : n4220;
  assign n4222 = pi14 ? n1896 : n1820;
  assign n4223 = pi14 ? n2293 : n1992;
  assign n4224 = pi13 ? n4222 : n4223;
  assign n4225 = pi12 ? n26 : n4224;
  assign n4226 = pi11 ? n4221 : n4225;
  assign n4227 = pi10 ? n3461 : n4226;
  assign n4228 = pi09 ? n26 : n4227;
  assign n4229 = pi08 ? n26 : n4228;
  assign n4230 = pi15 ? n554 : n2089;
  assign n4231 = pi14 ? n4230 : n543;
  assign n4232 = pi13 ? n4231 : n1386;
  assign n4233 = pi12 ? n26 : n4232;
  assign n4234 = pi11 ? n3479 : n4233;
  assign n4235 = pi14 ? n41 : n770;
  assign n4236 = pi14 ? n1165 : n3056;
  assign n4237 = pi13 ? n4235 : n4236;
  assign n4238 = pi12 ? n1880 : n4237;
  assign n4239 = pi14 ? n2351 : n1562;
  assign n4240 = pi14 ? n1583 : n1932;
  assign n4241 = pi13 ? n4239 : n4240;
  assign n4242 = pi12 ? n1921 : n4241;
  assign n4243 = pi11 ? n4238 : n4242;
  assign n4244 = pi10 ? n4234 : n4243;
  assign n4245 = pi15 ? n493 : n3496;
  assign n4246 = pi14 ? n4245 : n2118;
  assign n4247 = pi13 ? n2108 : n4246;
  assign n4248 = pi12 ? n2099 : n4247;
  assign n4249 = pi14 ? n2100 : n728;
  assign n4250 = pi13 ? n4249 : n4246;
  assign n4251 = pi12 ? n2099 : n4250;
  assign n4252 = pi11 ? n4248 : n4251;
  assign n4253 = pi15 ? n493 : n2114;
  assign n4254 = pi14 ? n4253 : n2227;
  assign n4255 = pi13 ? n2108 : n4254;
  assign n4256 = pi12 ? n1101 : n4255;
  assign n4257 = pi15 ? n503 : n66;
  assign n4258 = pi14 ? n958 : n4257;
  assign n4259 = pi14 ? n1165 : n26;
  assign n4260 = pi13 ? n4258 : n4259;
  assign n4261 = pi12 ? n1101 : n4260;
  assign n4262 = pi11 ? n4256 : n4261;
  assign n4263 = pi10 ? n4252 : n4262;
  assign n4264 = pi09 ? n4244 : n4263;
  assign n4265 = pi14 ? n958 : n3859;
  assign n4266 = pi15 ? n493 : n1983;
  assign n4267 = pi14 ? n4266 : n26;
  assign n4268 = pi13 ? n4265 : n4267;
  assign n4269 = pi12 ? n1101 : n4268;
  assign n4270 = pi15 ? n493 : n1758;
  assign n4271 = pi14 ? n4270 : n26;
  assign n4272 = pi13 ? n4265 : n4271;
  assign n4273 = pi12 ? n1101 : n4272;
  assign n4274 = pi11 ? n4269 : n4273;
  assign n4275 = pi15 ? n923 : n60;
  assign n4276 = pi14 ? n958 : n4275;
  assign n4277 = pi13 ? n4276 : n4271;
  assign n4278 = pi12 ? n1101 : n4277;
  assign n4279 = pi10 ? n4274 : n4278;
  assign n4280 = pi09 ? n4279 : n4278;
  assign n4281 = pi08 ? n4264 : n4280;
  assign n4282 = pi07 ? n4229 : n4281;
  assign n4283 = pi06 ? n4282 : n4278;
  assign n4284 = pi14 ? n101 : n3532;
  assign n4285 = pi13 ? n2167 : n4284;
  assign n4286 = pi12 ? n26 : n4285;
  assign n4287 = pi11 ? n26 : n4286;
  assign n4288 = pi14 ? n35 : n1374;
  assign n4289 = pi14 ? n323 : n4266;
  assign n4290 = pi13 ? n4288 : n4289;
  assign n4291 = pi12 ? n26 : n4290;
  assign n4292 = pi15 ? n224 : n2601;
  assign n4293 = pi14 ? n910 : n4292;
  assign n4294 = pi13 ? n3541 : n4293;
  assign n4295 = pi12 ? n26 : n4294;
  assign n4296 = pi11 ? n4291 : n4295;
  assign n4297 = pi10 ? n4287 : n4296;
  assign n4298 = pi09 ? n26 : n4297;
  assign n4299 = pi08 ? n26 : n4298;
  assign n4300 = pi14 ? n706 : n1616;
  assign n4301 = pi13 ? n4300 : n1677;
  assign n4302 = pi12 ? n26 : n4301;
  assign n4303 = pi14 ? n2185 : n543;
  assign n4304 = pi13 ? n4303 : n2190;
  assign n4305 = pi12 ? n26 : n4304;
  assign n4306 = pi11 ? n4302 : n4305;
  assign n4307 = pi14 ? n2197 : n1782;
  assign n4308 = pi13 ? n2195 : n4307;
  assign n4309 = pi12 ? n2088 : n4308;
  assign n4310 = pi15 ? n1870 : n26;
  assign n4311 = pi14 ? n2203 : n4310;
  assign n4312 = pi13 ? n2195 : n4311;
  assign n4313 = pi12 ? n1770 : n4312;
  assign n4314 = pi11 ? n4309 : n4313;
  assign n4315 = pi10 ? n4306 : n4314;
  assign n4316 = pi14 ? n2298 : n728;
  assign n4317 = pi14 ? n2212 : n2017;
  assign n4318 = pi13 ? n4316 : n4317;
  assign n4319 = pi12 ? n2099 : n4318;
  assign n4320 = pi16 ? n740 : n238;
  assign n4321 = pi15 ? n60 : n4320;
  assign n4322 = pi14 ? n4321 : n2118;
  assign n4323 = pi13 ? n2224 : n4322;
  assign n4324 = pi12 ? n1101 : n4323;
  assign n4325 = pi11 ? n4319 : n4324;
  assign n4326 = pi12 ? n1101 : n3170;
  assign n4327 = pi14 ? n2203 : n2118;
  assign n4328 = pi13 ? n2224 : n4327;
  assign n4329 = pi12 ? n1101 : n4328;
  assign n4330 = pi11 ? n4326 : n4329;
  assign n4331 = pi10 ? n4325 : n4330;
  assign n4332 = pi09 ? n4315 : n4331;
  assign n4333 = pi13 ? n3186 : n2228;
  assign n4334 = pi12 ? n1101 : n4333;
  assign n4335 = pi15 ? n60 : n3591;
  assign n4336 = pi14 ? n4335 : n2227;
  assign n4337 = pi13 ? n2244 : n4336;
  assign n4338 = pi12 ? n1101 : n4337;
  assign n4339 = pi10 ? n4334 : n4338;
  assign n4340 = pi09 ? n4339 : n4338;
  assign n4341 = pi08 ? n4332 : n4340;
  assign n4342 = pi07 ? n4299 : n4341;
  assign n4343 = pi14 ? n910 : n2227;
  assign n4344 = pi13 ? n2244 : n4343;
  assign n4345 = pi12 ? n1101 : n4344;
  assign n4346 = pi14 ? n2166 : n2101;
  assign n4347 = pi14 ? n1634 : n2227;
  assign n4348 = pi13 ? n4346 : n4347;
  assign n4349 = pi12 ? n1101 : n4348;
  assign n4350 = pi11 ? n4345 : n4349;
  assign n4351 = pi10 ? n4338 : n4350;
  assign n4352 = pi09 ? n4338 : n4351;
  assign n4353 = pi08 ? n4338 : n4352;
  assign n4354 = pi07 ? n4338 : n4353;
  assign n4355 = pi06 ? n4342 : n4354;
  assign n4356 = pi05 ? n4283 : n4355;
  assign n4357 = pi04 ? n4218 : n4356;
  assign n4358 = pi03 ? n4104 : n4357;
  assign n4359 = pi02 ? n3915 : n4358;
  assign n4360 = pi01 ? n3417 : n4359;
  assign n4361 = pi00 ? n2680 : n4360;
  assign po0 = ~n4361;
endmodule


