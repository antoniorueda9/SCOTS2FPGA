// Benchmark "DD" written by ABC on Wed May 22 13:40:20 2019

module DD ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15,
    po0, po1  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15;
  output po0, po1;
  wire n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
    n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
    n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
    n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601;
  assign n19 = 1'b1;
  assign n20 = pi14 ? n19 : ~n19;
  assign n21 = pi13 ? n19 : n20;
  assign n22 = pi12 ? n19 : n21;
  assign n23 = pi11 ? n22 : ~n19;
  assign n24 = pi10 ? n23 : ~n19;
  assign n25 = pi09 ? n19 : n24;
  assign n26 = pi08 ? n25 : ~n19;
  assign n27 = pi07 ? n19 : n26;
  assign n28 = pi06 ? n19 : n27;
  assign n29 = pi05 ? n19 : n28;
  assign n30 = pi15 ? n19 : ~n19;
  assign n31 = pi14 ? n30 : ~n19;
  assign n32 = pi13 ? n19 : n31;
  assign n33 = pi12 ? n19 : n32;
  assign n34 = pi11 ? n33 : ~n19;
  assign n35 = pi10 ? n34 : ~n19;
  assign n36 = pi09 ? n19 : n35;
  assign n37 = pi08 ? n36 : ~n19;
  assign n38 = pi07 ? n26 : n37;
  assign n39 = pi13 ? n19 : ~n19;
  assign n40 = pi12 ? n19 : n39;
  assign n41 = pi11 ? n40 : ~n19;
  assign n42 = pi10 ? n41 : ~n19;
  assign n43 = pi09 ? n19 : n42;
  assign n44 = pi08 ? n43 : ~n19;
  assign n45 = pi07 ? n37 : n44;
  assign n46 = pi06 ? n38 : n45;
  assign n47 = pi14 ? n19 : n30;
  assign n48 = pi13 ? n47 : ~n19;
  assign n49 = pi12 ? n19 : n48;
  assign n50 = pi11 ? n49 : ~n19;
  assign n51 = pi10 ? n50 : ~n19;
  assign n52 = pi09 ? n19 : n51;
  assign n53 = pi08 ? n52 : ~n19;
  assign n54 = pi13 ? n20 : ~n19;
  assign n55 = pi12 ? n19 : n54;
  assign n56 = pi11 ? n55 : ~n19;
  assign n57 = pi10 ? n56 : ~n19;
  assign n58 = pi09 ? n19 : n57;
  assign n59 = pi08 ? n58 : ~n19;
  assign n60 = pi07 ? n53 : n59;
  assign n61 = pi06 ? n53 : n60;
  assign n62 = pi05 ? n46 : n61;
  assign n63 = pi04 ? n29 : n62;
  assign n64 = pi03 ? n19 : n63;
  assign n65 = pi02 ? n19 : n64;
  assign n66 = pi13 ? n31 : ~n19;
  assign n67 = pi12 ? n19 : n66;
  assign n68 = pi11 ? n67 : ~n19;
  assign n69 = pi10 ? n68 : ~n19;
  assign n70 = pi09 ? n19 : n69;
  assign n71 = pi08 ? n70 : ~n19;
  assign n72 = pi07 ? n59 : n71;
  assign n73 = pi12 ? n19 : ~n19;
  assign n74 = pi11 ? n73 : ~n19;
  assign n75 = pi10 ? n74 : ~n19;
  assign n76 = pi09 ? n19 : n75;
  assign n77 = pi08 ? n76 : ~n19;
  assign n78 = pi07 ? n71 : n77;
  assign n79 = pi06 ? n72 : n78;
  assign n80 = pi13 ? n19 : n47;
  assign n81 = pi12 ? n80 : ~n19;
  assign n82 = pi11 ? n81 : ~n19;
  assign n83 = pi10 ? n82 : ~n19;
  assign n84 = pi09 ? n19 : n83;
  assign n85 = pi08 ? n84 : ~n19;
  assign n86 = pi05 ? n79 : n85;
  assign n87 = pi12 ? n21 : ~n19;
  assign n88 = pi11 ? n87 : ~n19;
  assign n89 = pi10 ? n88 : ~n19;
  assign n90 = pi09 ? n19 : n89;
  assign n91 = pi08 ? n90 : ~n19;
  assign n92 = pi07 ? n85 : n91;
  assign n93 = pi12 ? n32 : ~n19;
  assign n94 = pi11 ? n93 : ~n19;
  assign n95 = pi10 ? n94 : ~n19;
  assign n96 = pi09 ? n19 : n95;
  assign n97 = pi08 ? n96 : ~n19;
  assign n98 = pi07 ? n91 : n97;
  assign n99 = pi06 ? n92 : n98;
  assign n100 = pi12 ? n39 : ~n19;
  assign n101 = pi11 ? n100 : ~n19;
  assign n102 = pi10 ? n101 : ~n19;
  assign n103 = pi09 ? n19 : n102;
  assign n104 = pi08 ? n103 : ~n19;
  assign n105 = pi05 ? n99 : n104;
  assign n106 = pi04 ? n86 : n105;
  assign n107 = pi12 ? n48 : ~n19;
  assign n108 = pi11 ? n107 : ~n19;
  assign n109 = pi10 ? n108 : ~n19;
  assign n110 = pi09 ? n19 : n109;
  assign n111 = pi08 ? n110 : ~n19;
  assign n112 = pi07 ? n104 : n111;
  assign n113 = pi12 ? n54 : ~n19;
  assign n114 = pi11 ? n113 : ~n19;
  assign n115 = pi10 ? n114 : ~n19;
  assign n116 = pi09 ? n19 : n115;
  assign n117 = pi08 ? n116 : ~n19;
  assign n118 = pi07 ? n111 : n117;
  assign n119 = pi06 ? n112 : n118;
  assign n120 = pi12 ? n66 : ~n19;
  assign n121 = pi11 ? n120 : ~n19;
  assign n122 = pi10 ? n121 : ~n19;
  assign n123 = pi09 ? n19 : n122;
  assign n124 = pi08 ? n123 : ~n19;
  assign n125 = pi10 ? n19 : n56;
  assign n126 = pi11 ? n19 : n73;
  assign n127 = pi10 ? n19 : n126;
  assign n128 = pi09 ? n125 : ~n127;
  assign n129 = pi08 ? n123 : ~n128;
  assign n130 = pi06 ? n124 : n129;
  assign n131 = pi05 ? n119 : n130;
  assign n132 = pi09 ? n19 : ~n19;
  assign n133 = pi08 ? n132 : ~n128;
  assign n134 = pi07 ? n129 : n133;
  assign n135 = pi12 ? n19 : n80;
  assign n136 = pi11 ? n19 : n135;
  assign n137 = pi10 ? n19 : n136;
  assign n138 = pi09 ? n137 : ~n19;
  assign n139 = pi08 ? n138 : ~n128;
  assign n140 = pi07 ? n133 : n139;
  assign n141 = pi06 ? n134 : n140;
  assign n142 = pi11 ? n19 : n22;
  assign n143 = pi10 ? n19 : n142;
  assign n144 = pi09 ? n143 : ~n19;
  assign n145 = pi10 ? n19 : n74;
  assign n146 = pi09 ? n145 : ~n127;
  assign n147 = pi08 ? n144 : ~n146;
  assign n148 = pi08 ? n144 : ~n128;
  assign n149 = pi07 ? n148 : n147;
  assign n150 = pi06 ? n147 : n149;
  assign n151 = pi05 ? n141 : n150;
  assign n152 = pi04 ? n131 : n151;
  assign n153 = pi03 ? n106 : n152;
  assign n154 = pi10 ? n19 : n82;
  assign n155 = pi09 ? n154 : ~n127;
  assign n156 = pi08 ? n144 : ~n155;
  assign n157 = pi07 ? n147 : n156;
  assign n158 = pi11 ? n19 : n33;
  assign n159 = pi10 ? n19 : n158;
  assign n160 = pi09 ? n159 : ~n19;
  assign n161 = pi08 ? n160 : ~n155;
  assign n162 = pi07 ? n156 : n161;
  assign n163 = pi06 ? n157 : n162;
  assign n164 = pi11 ? n19 : n40;
  assign n165 = pi10 ? n19 : n164;
  assign n166 = pi09 ? n165 : ~n19;
  assign n167 = pi08 ? n166 : ~n155;
  assign n168 = pi12 ? n21 : n54;
  assign n169 = pi11 ? n168 : ~n19;
  assign n170 = pi10 ? n19 : n169;
  assign n171 = pi09 ? n170 : ~n127;
  assign n172 = pi08 ? n166 : ~n171;
  assign n173 = pi07 ? n167 : n172;
  assign n174 = pi06 ? n173 : n172;
  assign n175 = pi05 ? n163 : n174;
  assign n176 = pi10 ? n19 : n101;
  assign n177 = pi09 ? n176 : ~n127;
  assign n178 = pi08 ? n166 : ~n177;
  assign n179 = pi12 ? n21 : n19;
  assign n180 = pi11 ? n179 : n19;
  assign n181 = pi10 ? n180 : n126;
  assign n182 = pi09 ? n176 : ~n181;
  assign n183 = pi08 ? n166 : ~n182;
  assign n184 = pi07 ? n178 : n183;
  assign n185 = pi11 ? n19 : n49;
  assign n186 = pi10 ? n19 : n185;
  assign n187 = pi09 ? n186 : ~n19;
  assign n188 = pi13 ? n47 : ~n20;
  assign n189 = pi12 ? n188 : ~n19;
  assign n190 = pi11 ? n189 : ~n19;
  assign n191 = pi10 ? n19 : n190;
  assign n192 = pi09 ? n191 : ~n127;
  assign n193 = pi08 ? n187 : ~n192;
  assign n194 = pi07 ? n178 : n193;
  assign n195 = pi06 ? n184 : n194;
  assign n196 = pi11 ? n19 : n55;
  assign n197 = pi10 ? n19 : n196;
  assign n198 = pi09 ? n197 : ~n19;
  assign n199 = pi13 ? n47 : n19;
  assign n200 = pi12 ? n199 : ~n19;
  assign n201 = pi11 ? n200 : ~n19;
  assign n202 = pi10 ? n19 : n201;
  assign n203 = pi09 ? n202 : ~n127;
  assign n204 = pi08 ? n198 : ~n203;
  assign n205 = pi13 ? n31 : n19;
  assign n206 = pi12 ? n205 : ~n19;
  assign n207 = pi11 ? n206 : ~n19;
  assign n208 = pi10 ? n19 : n207;
  assign n209 = pi09 ? n208 : ~n127;
  assign n210 = pi08 ? n198 : ~n209;
  assign n211 = pi07 ? n204 : n210;
  assign n212 = pi10 ? n19 : ~n19;
  assign n213 = pi09 ? n212 : ~n127;
  assign n214 = pi08 ? n198 : ~n213;
  assign n215 = pi06 ? n211 : n214;
  assign n216 = pi05 ? n195 : n215;
  assign n217 = pi04 ? n175 : n216;
  assign n218 = pi10 ? n74 : n19;
  assign n219 = pi09 ? n197 : ~n218;
  assign n220 = pi13 ? n19 : ~n20;
  assign n221 = pi12 ? n220 : n19;
  assign n222 = pi11 ? n221 : n19;
  assign n223 = pi10 ? n126 : n222;
  assign n224 = pi09 ? n223 : n127;
  assign n225 = pi08 ? n219 : n224;
  assign n226 = pi13 ? n20 : ~n20;
  assign n227 = pi12 ? n226 : n19;
  assign n228 = pi11 ? n227 : n19;
  assign n229 = pi10 ? n126 : n228;
  assign n230 = pi09 ? n229 : n127;
  assign n231 = pi08 ? n219 : n230;
  assign n232 = pi07 ? n225 : n231;
  assign n233 = pi12 ? n188 : n19;
  assign n234 = pi11 ? n233 : n19;
  assign n235 = pi10 ? n126 : n234;
  assign n236 = pi09 ? n235 : n127;
  assign n237 = pi08 ? n219 : n236;
  assign n238 = pi10 ? n126 : ~n88;
  assign n239 = pi09 ? n238 : n127;
  assign n240 = pi08 ? n219 : n239;
  assign n241 = pi07 ? n237 : n240;
  assign n242 = pi06 ? n232 : n241;
  assign n243 = pi09 ? n127 : ~n218;
  assign n244 = pi10 ? n164 : ~n88;
  assign n245 = pi09 ? n244 : n127;
  assign n246 = pi08 ? n243 : n245;
  assign n247 = pi13 ? n20 : n19;
  assign n248 = pi12 ? n247 : ~n19;
  assign n249 = pi11 ? n248 : ~n19;
  assign n250 = pi10 ? n249 : n19;
  assign n251 = pi09 ? n127 : ~n250;
  assign n252 = pi12 ? n19 : n220;
  assign n253 = pi11 ? n19 : n252;
  assign n254 = pi10 ? n253 : ~n101;
  assign n255 = pi09 ? n254 : n127;
  assign n256 = pi08 ? n251 : n255;
  assign n257 = pi07 ? n246 : n256;
  assign n258 = pi08 ? n243 : n255;
  assign n259 = pi13 ? n19 : ~n31;
  assign n260 = pi12 ? n259 : ~n19;
  assign n261 = pi11 ? n19 : n260;
  assign n262 = pi10 ? n19 : n261;
  assign n263 = pi09 ? n254 : n262;
  assign n264 = pi08 ? n243 : n263;
  assign n265 = pi07 ? n258 : n264;
  assign n266 = pi06 ? n257 : n265;
  assign n267 = pi05 ? n242 : n266;
  assign n268 = pi10 ? n101 : n19;
  assign n269 = pi09 ? n127 : ~n268;
  assign n270 = pi12 ? n247 : n19;
  assign n271 = pi11 ? n270 : n19;
  assign n272 = pi10 ? n253 : n271;
  assign n273 = pi09 ? n272 : n127;
  assign n274 = pi08 ? n269 : n273;
  assign n275 = pi10 ? n253 : n19;
  assign n276 = pi09 ? n275 : n127;
  assign n277 = pi08 ? n269 : n276;
  assign n278 = pi07 ? n274 : n277;
  assign n279 = pi09 ? n19 : n127;
  assign n280 = pi08 ? n269 : n279;
  assign n281 = pi10 ? n114 : n19;
  assign n282 = pi09 ? n127 : ~n281;
  assign n283 = pi08 ? n282 : n279;
  assign n284 = pi07 ? n280 : n283;
  assign n285 = pi06 ? n278 : n284;
  assign n286 = pi09 ? n127 : n212;
  assign n287 = pi08 ? n286 : n279;
  assign n288 = pi10 ? n19 : n222;
  assign n289 = pi09 ? n288 : n127;
  assign n290 = pi08 ? n286 : n289;
  assign n291 = pi07 ? n287 : n290;
  assign n292 = pi06 ? n283 : n291;
  assign n293 = pi05 ? n285 : n292;
  assign n294 = pi04 ? n267 : n293;
  assign n295 = pi03 ? n217 : n294;
  assign n296 = pi02 ? n153 : n295;
  assign n297 = pi01 ? n65 : n296;
  assign n298 = pi09 ? n127 : n19;
  assign n299 = pi08 ? n298 : n289;
  assign n300 = pi08 ? n298 : n279;
  assign n301 = pi14 ? n30 : n19;
  assign n302 = pi13 ? n301 : n19;
  assign n303 = pi12 ? n302 : n19;
  assign n304 = pi11 ? n303 : n19;
  assign n305 = pi10 ? n19 : n304;
  assign n306 = pi09 ? n305 : n127;
  assign n307 = pi08 ? n298 : n306;
  assign n308 = pi07 ? n300 : n307;
  assign n309 = pi12 ? n19 : ~n21;
  assign n310 = pi11 ? n19 : n309;
  assign n311 = pi10 ? n19 : n310;
  assign n312 = pi09 ? n311 : n19;
  assign n313 = pi10 ? n136 : n271;
  assign n314 = pi09 ? n313 : n127;
  assign n315 = pi08 ? n312 : n314;
  assign n316 = pi10 ? n19 : n271;
  assign n317 = pi09 ? n316 : n127;
  assign n318 = pi08 ? n312 : n317;
  assign n319 = pi07 ? n315 : n318;
  assign n320 = pi06 ? n308 : n319;
  assign n321 = pi05 ? n299 : n320;
  assign n322 = pi08 ? n312 : n279;
  assign n323 = pi12 ? n19 : ~n39;
  assign n324 = pi11 ? n19 : n323;
  assign n325 = pi10 ? n19 : n324;
  assign n326 = pi09 ? n325 : n19;
  assign n327 = pi08 ? n326 : n279;
  assign n328 = pi12 ? n19 : ~n80;
  assign n329 = pi11 ? n19 : n328;
  assign n330 = pi10 ? n19 : n329;
  assign n331 = pi09 ? n19 : n330;
  assign n332 = pi08 ? n326 : n331;
  assign n333 = pi07 ? n327 : n332;
  assign n334 = pi06 ? n322 : n333;
  assign n335 = pi05 ? n322 : n334;
  assign n336 = pi04 ? n321 : n335;
  assign n337 = pi12 ? n80 : ~n39;
  assign n338 = pi11 ? n19 : n337;
  assign n339 = pi10 ? n19 : n338;
  assign n340 = pi09 ? n339 : n19;
  assign n341 = pi08 ? n340 : n331;
  assign n342 = pi09 ? n19 : n311;
  assign n343 = pi08 ? n340 : n342;
  assign n344 = pi07 ? n341 : n343;
  assign n345 = pi12 ? n19 : ~n32;
  assign n346 = pi11 ? n19 : n345;
  assign n347 = pi10 ? n19 : n346;
  assign n348 = pi09 ? n19 : n347;
  assign n349 = pi08 ? n340 : n348;
  assign n350 = pi07 ? n343 : n349;
  assign n351 = pi06 ? n344 : n350;
  assign n352 = pi09 ? n19 : n325;
  assign n353 = pi08 ? n340 : n352;
  assign n354 = pi07 ? n349 : n353;
  assign n355 = pi12 ? n80 : ~n54;
  assign n356 = pi11 ? n19 : n355;
  assign n357 = pi10 ? n19 : n356;
  assign n358 = pi09 ? n357 : n19;
  assign n359 = pi08 ? n358 : n352;
  assign n360 = pi12 ? n19 : ~n48;
  assign n361 = pi11 ? n19 : n360;
  assign n362 = pi10 ? n19 : n361;
  assign n363 = pi09 ? n19 : n362;
  assign n364 = pi08 ? n358 : n363;
  assign n365 = pi07 ? n359 : n364;
  assign n366 = pi06 ? n354 : n365;
  assign n367 = pi05 ? n351 : n366;
  assign n368 = pi12 ? n19 : ~n54;
  assign n369 = pi11 ? n19 : n368;
  assign n370 = pi10 ? n19 : n369;
  assign n371 = pi09 ? n19 : n370;
  assign n372 = pi08 ? n358 : n371;
  assign n373 = pi07 ? n364 : n372;
  assign n374 = pi13 ? n19 : n301;
  assign n375 = pi12 ? n374 : ~n54;
  assign n376 = pi11 ? n19 : n375;
  assign n377 = pi10 ? n19 : n376;
  assign n378 = pi09 ? n19 : n377;
  assign n379 = pi08 ? n358 : n378;
  assign n380 = pi12 ? n19 : ~n66;
  assign n381 = pi11 ? n19 : n380;
  assign n382 = pi10 ? n19 : n381;
  assign n383 = pi09 ? n19 : n382;
  assign n384 = pi08 ? n358 : n383;
  assign n385 = pi07 ? n379 : n384;
  assign n386 = pi06 ? n373 : n385;
  assign n387 = pi08 ? n358 : n19;
  assign n388 = pi07 ? n384 : n387;
  assign n389 = pi12 ? n80 : n19;
  assign n390 = pi11 ? n19 : n389;
  assign n391 = pi10 ? n19 : n390;
  assign n392 = pi09 ? n391 : n19;
  assign n393 = pi08 ? n392 : n19;
  assign n394 = pi06 ? n388 : n393;
  assign n395 = pi05 ? n386 : n394;
  assign n396 = pi04 ? n367 : n395;
  assign n397 = pi03 ? n336 : n396;
  assign n398 = pi07 ? n393 : n19;
  assign n399 = pi06 ? n393 : n398;
  assign n400 = pi05 ? n399 : n19;
  assign n401 = pi04 ? n400 : n19;
  assign n402 = pi03 ? n401 : n19;
  assign n403 = pi02 ? n397 : n402;
  assign n404 = pi01 ? n403 : n19;
  assign n405 = pi00 ? n297 : n404;
  assign n406 = pi05 ? n119 : n124;
  assign n407 = pi08 ? n132 : ~n19;
  assign n408 = pi07 ? n124 : n407;
  assign n409 = pi08 ? n138 : ~n19;
  assign n410 = pi07 ? n407 : n409;
  assign n411 = pi06 ? n408 : n410;
  assign n412 = pi08 ? n144 : ~n19;
  assign n413 = pi05 ? n411 : n412;
  assign n414 = pi04 ? n406 : n413;
  assign n415 = pi03 ? n106 : n414;
  assign n416 = pi08 ? n160 : ~n19;
  assign n417 = pi07 ? n412 : n416;
  assign n418 = pi06 ? n412 : n417;
  assign n419 = pi08 ? n166 : ~n19;
  assign n420 = pi05 ? n418 : n419;
  assign n421 = pi08 ? n187 : ~n19;
  assign n422 = pi07 ? n419 : n421;
  assign n423 = pi06 ? n419 : n422;
  assign n424 = pi08 ? n198 : ~n19;
  assign n425 = pi05 ? n423 : n424;
  assign n426 = pi04 ? n420 : n425;
  assign n427 = pi11 ? n19 : n67;
  assign n428 = pi10 ? n19 : n427;
  assign n429 = pi09 ? n428 : ~n19;
  assign n430 = pi08 ? n429 : ~n19;
  assign n431 = pi07 ? n424 : n430;
  assign n432 = pi06 ? n424 : n431;
  assign n433 = pi09 ? n127 : ~n19;
  assign n434 = pi08 ? n433 : ~n19;
  assign n435 = pi05 ? n432 : n434;
  assign n436 = pi11 ? n19 : n81;
  assign n437 = pi10 ? n19 : n436;
  assign n438 = pi09 ? n437 : ~n19;
  assign n439 = pi08 ? n438 : ~n19;
  assign n440 = pi07 ? n434 : n439;
  assign n441 = pi06 ? n434 : n440;
  assign n442 = pi05 ? n441 : n439;
  assign n443 = pi04 ? n435 : n442;
  assign n444 = pi03 ? n426 : n443;
  assign n445 = pi02 ? n415 : n444;
  assign n446 = pi01 ? n65 : n445;
  assign n447 = pi09 ? n19 : n137;
  assign n448 = pi08 ? n438 : ~n447;
  assign n449 = pi07 ? n439 : n448;
  assign n450 = pi06 ? n439 : n449;
  assign n451 = pi05 ? n439 : n450;
  assign n452 = pi04 ? n439 : n451;
  assign n453 = pi09 ? n19 : n143;
  assign n454 = pi08 ? n438 : ~n453;
  assign n455 = pi07 ? n448 : n454;
  assign n456 = pi09 ? n19 : n159;
  assign n457 = pi08 ? n438 : ~n456;
  assign n458 = pi07 ? n454 : n457;
  assign n459 = pi06 ? n455 : n458;
  assign n460 = pi09 ? n19 : n165;
  assign n461 = pi08 ? n438 : ~n460;
  assign n462 = pi07 ? n457 : n461;
  assign n463 = pi09 ? n19 : n186;
  assign n464 = pi08 ? n438 : ~n463;
  assign n465 = pi07 ? n461 : n464;
  assign n466 = pi06 ? n462 : n465;
  assign n467 = pi05 ? n459 : n466;
  assign n468 = pi09 ? n19 : n197;
  assign n469 = pi08 ? n438 : ~n468;
  assign n470 = pi07 ? n464 : n469;
  assign n471 = pi09 ? n19 : n428;
  assign n472 = pi08 ? n438 : ~n471;
  assign n473 = pi07 ? n469 : n472;
  assign n474 = pi06 ? n470 : n473;
  assign n475 = pi08 ? n438 : ~n279;
  assign n476 = pi07 ? n472 : n475;
  assign n477 = pi06 ? n476 : n475;
  assign n478 = pi05 ? n474 : n477;
  assign n479 = pi04 ? n467 : n478;
  assign n480 = pi03 ? n452 : n479;
  assign n481 = pi09 ? n19 : n437;
  assign n482 = pi08 ? n438 : ~n481;
  assign n483 = pi06 ? n475 : n482;
  assign n484 = pi05 ? n475 : n483;
  assign n485 = pi04 ? n475 : n484;
  assign n486 = pi11 ? n19 : n87;
  assign n487 = pi10 ? n19 : n486;
  assign n488 = pi09 ? n19 : n487;
  assign n489 = pi08 ? n438 : ~n488;
  assign n490 = pi11 ? n19 : n93;
  assign n491 = pi10 ? n19 : n490;
  assign n492 = pi09 ? n19 : n491;
  assign n493 = pi08 ? n438 : ~n492;
  assign n494 = pi06 ? n489 : n493;
  assign n495 = pi11 ? n19 : n100;
  assign n496 = pi10 ? n19 : n495;
  assign n497 = pi09 ? n19 : n496;
  assign n498 = pi08 ? n438 : ~n497;
  assign n499 = pi11 ? n19 : n107;
  assign n500 = pi10 ? n19 : n499;
  assign n501 = pi09 ? n19 : n500;
  assign n502 = pi08 ? n438 : ~n501;
  assign n503 = pi06 ? n498 : n502;
  assign n504 = pi05 ? n494 : n503;
  assign n505 = pi11 ? n19 : n113;
  assign n506 = pi10 ? n19 : n505;
  assign n507 = pi09 ? n19 : n506;
  assign n508 = pi08 ? n438 : ~n507;
  assign n509 = pi11 ? n19 : n120;
  assign n510 = pi10 ? n19 : n509;
  assign n511 = pi09 ? n19 : n510;
  assign n512 = pi08 ? n438 : ~n511;
  assign n513 = pi06 ? n508 : n512;
  assign n514 = pi11 ? n19 : ~n19;
  assign n515 = pi10 ? n19 : n514;
  assign n516 = pi09 ? n19 : n515;
  assign n517 = pi08 ? n438 : ~n516;
  assign n518 = pi05 ? n513 : n517;
  assign n519 = pi04 ? n504 : n518;
  assign n520 = pi03 ? n485 : n519;
  assign n521 = pi02 ? n480 : n520;
  assign n522 = pi11 ? n135 : ~n19;
  assign n523 = pi10 ? n19 : n522;
  assign n524 = pi09 ? n19 : n523;
  assign n525 = pi08 ? n438 : ~n524;
  assign n526 = pi07 ? n517 : n525;
  assign n527 = pi10 ? n19 : n23;
  assign n528 = pi09 ? n19 : n527;
  assign n529 = pi08 ? n438 : ~n528;
  assign n530 = pi07 ? n525 : n529;
  assign n531 = pi06 ? n526 : n530;
  assign n532 = pi05 ? n517 : n531;
  assign n533 = pi04 ? n517 : n532;
  assign n534 = pi10 ? n19 : n34;
  assign n535 = pi09 ? n19 : n534;
  assign n536 = pi08 ? n438 : ~n535;
  assign n537 = pi07 ? n529 : n536;
  assign n538 = pi10 ? n19 : n41;
  assign n539 = pi09 ? n19 : n538;
  assign n540 = pi08 ? n438 : ~n539;
  assign n541 = pi07 ? n536 : n540;
  assign n542 = pi06 ? n537 : n541;
  assign n543 = pi10 ? n19 : n50;
  assign n544 = pi09 ? n19 : n543;
  assign n545 = pi08 ? n438 : ~n544;
  assign n546 = pi07 ? n540 : n545;
  assign n547 = pi09 ? n19 : n125;
  assign n548 = pi08 ? n438 : ~n547;
  assign n549 = pi07 ? n545 : n548;
  assign n550 = pi06 ? n546 : n549;
  assign n551 = pi05 ? n542 : n550;
  assign n552 = pi10 ? n19 : n68;
  assign n553 = pi09 ? n19 : n552;
  assign n554 = pi08 ? n438 : ~n553;
  assign n555 = pi07 ? n548 : n554;
  assign n556 = pi09 ? n19 : n145;
  assign n557 = pi08 ? n438 : ~n556;
  assign n558 = pi07 ? n554 : n557;
  assign n559 = pi06 ? n555 : n558;
  assign n560 = pi05 ? n559 : n557;
  assign n561 = pi04 ? n551 : n560;
  assign n562 = pi03 ? n533 : n561;
  assign n563 = pi09 ? n19 : n154;
  assign n564 = pi08 ? n438 : ~n563;
  assign n565 = pi10 ? n19 : n88;
  assign n566 = pi09 ? n19 : n565;
  assign n567 = pi08 ? n438 : ~n566;
  assign n568 = pi06 ? n564 : n567;
  assign n569 = pi05 ? n557 : n568;
  assign n570 = pi04 ? n557 : n569;
  assign n571 = pi10 ? n19 : n94;
  assign n572 = pi09 ? n19 : n571;
  assign n573 = pi08 ? n438 : ~n572;
  assign n574 = pi09 ? n19 : n176;
  assign n575 = pi08 ? n438 : ~n574;
  assign n576 = pi07 ? n573 : n575;
  assign n577 = pi06 ? n573 : n576;
  assign n578 = pi10 ? n19 : n108;
  assign n579 = pi09 ? n19 : n578;
  assign n580 = pi08 ? n438 : ~n579;
  assign n581 = pi07 ? n575 : n580;
  assign n582 = pi10 ? n19 : n114;
  assign n583 = pi09 ? n19 : n582;
  assign n584 = pi08 ? n438 : ~n583;
  assign n585 = pi07 ? n580 : n584;
  assign n586 = pi06 ? n581 : n585;
  assign n587 = pi05 ? n577 : n586;
  assign n588 = pi10 ? n19 : n121;
  assign n589 = pi09 ? n19 : n588;
  assign n590 = pi08 ? n438 : ~n589;
  assign n591 = pi07 ? n584 : n590;
  assign n592 = pi09 ? n19 : n212;
  assign n593 = pi08 ? n438 : ~n592;
  assign n594 = pi07 ? n590 : n593;
  assign n595 = pi06 ? n591 : n594;
  assign n596 = pi05 ? n595 : n593;
  assign n597 = pi04 ? n587 : n596;
  assign n598 = pi03 ? n570 : n597;
  assign n599 = pi02 ? n562 : n598;
  assign n600 = pi01 ? n521 : n599;
  assign n601 = pi00 ? n446 : n600;
  assign po0 = ~n405;
  assign po1 = ~n601;
endmodule


