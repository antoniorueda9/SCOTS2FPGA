// Benchmark "DD" written by ABC on Tue May 28 18:25:14 2019

module DD ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16,
    po0  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0;
  wire n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
    n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
    n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
    n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632;
  assign n19 = 1'b1;
  assign n20 = pi16 ? n19 : ~n19;
  assign n21 = pi14 ? n19 : ~n20;
  assign n22 = pi13 ? n19 : n21;
  assign n23 = pi12 ? n19 : n22;
  assign n24 = pi11 ? n23 : ~n20;
  assign n25 = pi10 ? n24 : ~n20;
  assign n26 = pi09 ? n19 : n25;
  assign n27 = pi08 ? n26 : ~n20;
  assign n28 = pi07 ? n19 : n27;
  assign n29 = pi06 ? n19 : n28;
  assign n30 = pi05 ? n19 : n29;
  assign n31 = pi15 ? n19 : ~n20;
  assign n32 = pi14 ? n31 : ~n20;
  assign n33 = pi13 ? n19 : n32;
  assign n34 = pi12 ? n19 : n33;
  assign n35 = pi11 ? n34 : ~n20;
  assign n36 = pi10 ? n35 : ~n20;
  assign n37 = pi09 ? n19 : n36;
  assign n38 = pi08 ? n37 : ~n20;
  assign n39 = pi07 ? n27 : n38;
  assign n40 = pi13 ? n19 : ~n20;
  assign n41 = pi12 ? n19 : n40;
  assign n42 = pi11 ? n41 : ~n20;
  assign n43 = pi10 ? n42 : ~n20;
  assign n44 = pi09 ? n19 : n43;
  assign n45 = pi08 ? n44 : ~n20;
  assign n46 = pi07 ? n38 : n45;
  assign n47 = pi06 ? n39 : n46;
  assign n48 = pi14 ? n19 : n31;
  assign n49 = pi13 ? n48 : ~n20;
  assign n50 = pi12 ? n19 : n49;
  assign n51 = pi11 ? n50 : ~n20;
  assign n52 = pi10 ? n51 : ~n20;
  assign n53 = pi09 ? n19 : n52;
  assign n54 = pi08 ? n53 : ~n20;
  assign n55 = pi13 ? n21 : ~n20;
  assign n56 = pi12 ? n19 : n55;
  assign n57 = pi11 ? n56 : ~n20;
  assign n58 = pi10 ? n57 : ~n20;
  assign n59 = pi09 ? n19 : n58;
  assign n60 = pi08 ? n59 : ~n20;
  assign n61 = pi07 ? n54 : n60;
  assign n62 = pi06 ? n54 : n61;
  assign n63 = pi05 ? n47 : n62;
  assign n64 = pi04 ? n30 : n63;
  assign n65 = pi03 ? n19 : n64;
  assign n66 = pi02 ? n19 : n65;
  assign n67 = pi13 ? n32 : ~n20;
  assign n68 = pi12 ? n19 : n67;
  assign n69 = pi11 ? n68 : ~n20;
  assign n70 = pi10 ? n69 : ~n20;
  assign n71 = pi09 ? n19 : n70;
  assign n72 = pi08 ? n71 : ~n20;
  assign n73 = pi07 ? n60 : n72;
  assign n74 = pi12 ? n19 : ~n20;
  assign n75 = pi11 ? n74 : ~n20;
  assign n76 = pi10 ? n75 : ~n20;
  assign n77 = pi09 ? n19 : n76;
  assign n78 = pi08 ? n77 : ~n20;
  assign n79 = pi07 ? n72 : n78;
  assign n80 = pi06 ? n73 : n79;
  assign n81 = pi13 ? n19 : n48;
  assign n82 = pi12 ? n81 : ~n20;
  assign n83 = pi11 ? n82 : ~n20;
  assign n84 = pi10 ? n83 : ~n20;
  assign n85 = pi09 ? n19 : n84;
  assign n86 = pi08 ? n85 : ~n20;
  assign n87 = pi05 ? n80 : n86;
  assign n88 = pi12 ? n22 : ~n20;
  assign n89 = pi11 ? n88 : ~n20;
  assign n90 = pi10 ? n89 : ~n20;
  assign n91 = pi09 ? n19 : n90;
  assign n92 = pi08 ? n91 : ~n20;
  assign n93 = pi07 ? n86 : n92;
  assign n94 = pi12 ? n33 : ~n20;
  assign n95 = pi11 ? n94 : ~n20;
  assign n96 = pi10 ? n95 : ~n20;
  assign n97 = pi09 ? n19 : n96;
  assign n98 = pi08 ? n97 : ~n20;
  assign n99 = pi07 ? n92 : n98;
  assign n100 = pi06 ? n93 : n99;
  assign n101 = pi12 ? n40 : ~n20;
  assign n102 = pi11 ? n101 : ~n20;
  assign n103 = pi10 ? n102 : ~n20;
  assign n104 = pi09 ? n19 : n103;
  assign n105 = pi08 ? n104 : ~n20;
  assign n106 = pi05 ? n100 : n105;
  assign n107 = pi04 ? n87 : n106;
  assign n108 = pi12 ? n49 : ~n20;
  assign n109 = pi11 ? n108 : ~n20;
  assign n110 = pi10 ? n109 : ~n20;
  assign n111 = pi09 ? n19 : n110;
  assign n112 = pi08 ? n111 : ~n20;
  assign n113 = pi07 ? n105 : n112;
  assign n114 = pi12 ? n55 : ~n20;
  assign n115 = pi11 ? n114 : ~n20;
  assign n116 = pi10 ? n115 : ~n20;
  assign n117 = pi09 ? n19 : n116;
  assign n118 = pi08 ? n117 : ~n20;
  assign n119 = pi07 ? n112 : n118;
  assign n120 = pi06 ? n113 : n119;
  assign n121 = pi12 ? n67 : ~n20;
  assign n122 = pi11 ? n121 : ~n20;
  assign n123 = pi10 ? n122 : ~n20;
  assign n124 = pi09 ? n19 : n123;
  assign n125 = pi08 ? n124 : ~n20;
  assign n126 = pi14 ? n20 : ~n20;
  assign n127 = pi13 ? n126 : ~n20;
  assign n128 = pi12 ? n20 : n127;
  assign n129 = pi11 ? n128 : ~n20;
  assign n130 = pi10 ? n20 : n129;
  assign n131 = pi12 ? n20 : ~n20;
  assign n132 = pi11 ? n20 : n131;
  assign n133 = pi10 ? n20 : n132;
  assign n134 = pi09 ? n130 : ~n133;
  assign n135 = pi08 ? n124 : ~n134;
  assign n136 = pi06 ? n125 : n135;
  assign n137 = pi05 ? n120 : n136;
  assign n138 = pi09 ? n19 : ~n20;
  assign n139 = pi08 ? n138 : ~n134;
  assign n140 = pi07 ? n135 : n139;
  assign n141 = pi12 ? n19 : n81;
  assign n142 = pi11 ? n19 : n141;
  assign n143 = pi10 ? n19 : n142;
  assign n144 = pi09 ? n143 : ~n20;
  assign n145 = pi08 ? n144 : ~n134;
  assign n146 = pi07 ? n139 : n145;
  assign n147 = pi06 ? n140 : n146;
  assign n148 = pi11 ? n19 : n23;
  assign n149 = pi10 ? n19 : n148;
  assign n150 = pi09 ? n149 : ~n20;
  assign n151 = pi11 ? n131 : ~n20;
  assign n152 = pi10 ? n20 : n151;
  assign n153 = pi09 ? n152 : ~n133;
  assign n154 = pi08 ? n150 : ~n153;
  assign n155 = pi08 ? n150 : ~n134;
  assign n156 = pi07 ? n155 : n154;
  assign n157 = pi06 ? n154 : n156;
  assign n158 = pi05 ? n147 : n157;
  assign n159 = pi04 ? n137 : n158;
  assign n160 = pi03 ? n107 : n159;
  assign n161 = pi15 ? n20 : ~n20;
  assign n162 = pi14 ? n20 : n161;
  assign n163 = pi13 ? n20 : n162;
  assign n164 = pi12 ? n163 : ~n20;
  assign n165 = pi11 ? n164 : ~n20;
  assign n166 = pi10 ? n20 : n165;
  assign n167 = pi09 ? n166 : ~n133;
  assign n168 = pi08 ? n150 : ~n167;
  assign n169 = pi07 ? n154 : n168;
  assign n170 = pi11 ? n19 : n34;
  assign n171 = pi10 ? n19 : n170;
  assign n172 = pi09 ? n171 : ~n20;
  assign n173 = pi08 ? n172 : ~n167;
  assign n174 = pi07 ? n168 : n173;
  assign n175 = pi06 ? n169 : n174;
  assign n176 = pi11 ? n19 : n41;
  assign n177 = pi10 ? n19 : n176;
  assign n178 = pi09 ? n177 : ~n20;
  assign n179 = pi08 ? n178 : ~n167;
  assign n180 = pi13 ? n20 : n126;
  assign n181 = pi12 ? n180 : n127;
  assign n182 = pi11 ? n181 : ~n20;
  assign n183 = pi10 ? n20 : n182;
  assign n184 = pi09 ? n183 : ~n133;
  assign n185 = pi08 ? n178 : ~n184;
  assign n186 = pi07 ? n179 : n185;
  assign n187 = pi06 ? n186 : n185;
  assign n188 = pi05 ? n175 : n187;
  assign n189 = pi13 ? n20 : ~n20;
  assign n190 = pi12 ? n189 : ~n20;
  assign n191 = pi11 ? n190 : ~n20;
  assign n192 = pi10 ? n20 : n191;
  assign n193 = pi09 ? n192 : ~n133;
  assign n194 = pi08 ? n178 : ~n193;
  assign n195 = pi12 ? n180 : n20;
  assign n196 = pi11 ? n195 : n20;
  assign n197 = pi10 ? n196 : n132;
  assign n198 = pi09 ? n192 : ~n197;
  assign n199 = pi08 ? n178 : ~n198;
  assign n200 = pi07 ? n194 : n199;
  assign n201 = pi11 ? n19 : n50;
  assign n202 = pi10 ? n19 : n201;
  assign n203 = pi09 ? n202 : ~n20;
  assign n204 = pi13 ? n162 : ~n126;
  assign n205 = pi12 ? n204 : ~n20;
  assign n206 = pi11 ? n205 : ~n20;
  assign n207 = pi10 ? n20 : n206;
  assign n208 = pi09 ? n207 : ~n133;
  assign n209 = pi08 ? n203 : ~n208;
  assign n210 = pi07 ? n194 : n209;
  assign n211 = pi06 ? n200 : n210;
  assign n212 = pi11 ? n19 : n56;
  assign n213 = pi10 ? n19 : n212;
  assign n214 = pi09 ? n213 : ~n20;
  assign n215 = pi13 ? n162 : n20;
  assign n216 = pi12 ? n215 : ~n20;
  assign n217 = pi11 ? n216 : ~n20;
  assign n218 = pi10 ? n20 : n217;
  assign n219 = pi09 ? n218 : ~n133;
  assign n220 = pi08 ? n214 : ~n219;
  assign n221 = pi14 ? n161 : ~n20;
  assign n222 = pi13 ? n221 : n20;
  assign n223 = pi12 ? n222 : ~n20;
  assign n224 = pi11 ? n223 : ~n20;
  assign n225 = pi10 ? n20 : n224;
  assign n226 = pi09 ? n225 : ~n133;
  assign n227 = pi08 ? n214 : ~n226;
  assign n228 = pi07 ? n220 : n227;
  assign n229 = pi10 ? n20 : ~n20;
  assign n230 = pi09 ? n229 : ~n133;
  assign n231 = pi08 ? n214 : ~n230;
  assign n232 = pi06 ? n228 : n231;
  assign n233 = pi05 ? n211 : n232;
  assign n234 = pi04 ? n188 : n233;
  assign n235 = pi10 ? n151 : n20;
  assign n236 = pi09 ? n213 : ~n235;
  assign n237 = pi13 ? n20 : ~n126;
  assign n238 = pi12 ? n237 : n20;
  assign n239 = pi11 ? n238 : n20;
  assign n240 = pi10 ? n132 : n239;
  assign n241 = pi09 ? n240 : n133;
  assign n242 = pi08 ? n236 : n241;
  assign n243 = pi13 ? n126 : ~n126;
  assign n244 = pi12 ? n243 : n20;
  assign n245 = pi11 ? n244 : n20;
  assign n246 = pi10 ? n132 : n245;
  assign n247 = pi09 ? n246 : n133;
  assign n248 = pi08 ? n236 : n247;
  assign n249 = pi07 ? n242 : n248;
  assign n250 = pi12 ? n204 : n20;
  assign n251 = pi11 ? n250 : n20;
  assign n252 = pi10 ? n132 : n251;
  assign n253 = pi09 ? n252 : n133;
  assign n254 = pi08 ? n236 : n253;
  assign n255 = pi15 ? n19 : n20;
  assign n256 = pi14 ? n255 : ~n20;
  assign n257 = pi13 ? n256 : ~n20;
  assign n258 = pi12 ? n19 : n257;
  assign n259 = pi11 ? n19 : n258;
  assign n260 = pi10 ? n19 : n259;
  assign n261 = pi09 ? n260 : ~n235;
  assign n262 = pi12 ? n180 : ~n20;
  assign n263 = pi11 ? n262 : ~n20;
  assign n264 = pi10 ? n132 : ~n263;
  assign n265 = pi09 ? n264 : n133;
  assign n266 = pi08 ? n261 : n265;
  assign n267 = pi07 ? n254 : n266;
  assign n268 = pi06 ? n249 : n267;
  assign n269 = pi11 ? n19 : n74;
  assign n270 = pi10 ? n19 : n269;
  assign n271 = pi09 ? n270 : ~n235;
  assign n272 = pi12 ? n20 : n189;
  assign n273 = pi11 ? n20 : n272;
  assign n274 = pi10 ? n273 : ~n263;
  assign n275 = pi09 ? n274 : n133;
  assign n276 = pi08 ? n271 : n275;
  assign n277 = pi13 ? n126 : n20;
  assign n278 = pi12 ? n277 : ~n20;
  assign n279 = pi11 ? n278 : ~n20;
  assign n280 = pi10 ? n279 : n20;
  assign n281 = pi09 ? n270 : ~n280;
  assign n282 = pi12 ? n20 : n237;
  assign n283 = pi11 ? n20 : n282;
  assign n284 = pi10 ? n283 : ~n191;
  assign n285 = pi09 ? n284 : n133;
  assign n286 = pi08 ? n281 : n285;
  assign n287 = pi07 ? n276 : n286;
  assign n288 = pi08 ? n271 : n285;
  assign n289 = pi13 ? n20 : ~n221;
  assign n290 = pi12 ? n289 : ~n20;
  assign n291 = pi11 ? n20 : n290;
  assign n292 = pi10 ? n20 : n291;
  assign n293 = pi09 ? n284 : n292;
  assign n294 = pi08 ? n271 : n293;
  assign n295 = pi07 ? n288 : n294;
  assign n296 = pi06 ? n287 : n295;
  assign n297 = pi05 ? n268 : n296;
  assign n298 = pi10 ? n191 : n20;
  assign n299 = pi09 ? n270 : ~n298;
  assign n300 = pi12 ? n277 : n20;
  assign n301 = pi11 ? n300 : n20;
  assign n302 = pi10 ? n283 : n301;
  assign n303 = pi09 ? n302 : n133;
  assign n304 = pi08 ? n299 : n303;
  assign n305 = pi10 ? n283 : n20;
  assign n306 = pi09 ? n305 : n133;
  assign n307 = pi08 ? n299 : n306;
  assign n308 = pi07 ? n304 : n307;
  assign n309 = pi09 ? n20 : n133;
  assign n310 = pi08 ? n299 : n309;
  assign n311 = pi14 ? n19 : n255;
  assign n312 = pi13 ? n19 : n311;
  assign n313 = pi12 ? n312 : ~n20;
  assign n314 = pi11 ? n19 : n313;
  assign n315 = pi10 ? n19 : n314;
  assign n316 = pi12 ? n127 : ~n20;
  assign n317 = pi11 ? n316 : ~n20;
  assign n318 = pi10 ? n317 : n20;
  assign n319 = pi09 ? n315 : ~n318;
  assign n320 = pi08 ? n319 : n309;
  assign n321 = pi07 ? n310 : n320;
  assign n322 = pi06 ? n308 : n321;
  assign n323 = pi09 ? n315 : n229;
  assign n324 = pi08 ? n323 : n309;
  assign n325 = pi10 ? n20 : n239;
  assign n326 = pi09 ? n325 : n133;
  assign n327 = pi08 ? n323 : n326;
  assign n328 = pi07 ? n324 : n327;
  assign n329 = pi06 ? n320 : n328;
  assign n330 = pi05 ? n322 : n329;
  assign n331 = pi04 ? n297 : n330;
  assign n332 = pi03 ? n234 : n331;
  assign n333 = pi02 ? n160 : n332;
  assign n334 = pi01 ? n66 : n333;
  assign n335 = pi09 ? n315 : n20;
  assign n336 = pi08 ? n335 : n326;
  assign n337 = pi08 ? n335 : n309;
  assign n338 = pi14 ? n161 : n20;
  assign n339 = pi13 ? n338 : n20;
  assign n340 = pi12 ? n339 : n20;
  assign n341 = pi11 ? n340 : n20;
  assign n342 = pi10 ? n20 : n341;
  assign n343 = pi09 ? n342 : n133;
  assign n344 = pi08 ? n335 : n343;
  assign n345 = pi07 ? n337 : n344;
  assign n346 = pi12 ? n312 : ~n180;
  assign n347 = pi11 ? n19 : n346;
  assign n348 = pi10 ? n19 : n347;
  assign n349 = pi09 ? n348 : n20;
  assign n350 = pi12 ? n20 : n163;
  assign n351 = pi11 ? n20 : n350;
  assign n352 = pi10 ? n351 : n301;
  assign n353 = pi09 ? n352 : n133;
  assign n354 = pi08 ? n349 : n353;
  assign n355 = pi10 ? n20 : n301;
  assign n356 = pi09 ? n355 : n133;
  assign n357 = pi08 ? n349 : n356;
  assign n358 = pi07 ? n354 : n357;
  assign n359 = pi06 ? n345 : n358;
  assign n360 = pi05 ? n336 : n359;
  assign n361 = pi08 ? n349 : n309;
  assign n362 = pi12 ? n312 : ~n189;
  assign n363 = pi11 ? n19 : n362;
  assign n364 = pi10 ? n19 : n363;
  assign n365 = pi09 ? n364 : n20;
  assign n366 = pi08 ? n365 : n309;
  assign n367 = pi15 ? n20 : ~n19;
  assign n368 = pi14 ? n20 : n367;
  assign n369 = pi13 ? n20 : n368;
  assign n370 = pi12 ? n20 : ~n369;
  assign n371 = pi11 ? n20 : n370;
  assign n372 = pi10 ? n20 : n371;
  assign n373 = pi09 ? n20 : n372;
  assign n374 = pi08 ? n365 : n373;
  assign n375 = pi07 ? n366 : n374;
  assign n376 = pi06 ? n361 : n375;
  assign n377 = pi05 ? n361 : n376;
  assign n378 = pi04 ? n360 : n377;
  assign n379 = pi12 ? n81 : ~n189;
  assign n380 = pi11 ? n19 : n379;
  assign n381 = pi10 ? n19 : n380;
  assign n382 = pi09 ? n381 : n20;
  assign n383 = pi08 ? n382 : n373;
  assign n384 = pi14 ? n20 : ~n19;
  assign n385 = pi13 ? n20 : n384;
  assign n386 = pi12 ? n20 : ~n385;
  assign n387 = pi11 ? n20 : n386;
  assign n388 = pi10 ? n20 : n387;
  assign n389 = pi09 ? n20 : n388;
  assign n390 = pi08 ? n382 : n389;
  assign n391 = pi07 ? n383 : n390;
  assign n392 = pi14 ? n367 : ~n19;
  assign n393 = pi13 ? n20 : n392;
  assign n394 = pi12 ? n20 : ~n393;
  assign n395 = pi11 ? n20 : n394;
  assign n396 = pi10 ? n20 : n395;
  assign n397 = pi09 ? n20 : n396;
  assign n398 = pi08 ? n382 : n397;
  assign n399 = pi07 ? n390 : n398;
  assign n400 = pi06 ? n391 : n399;
  assign n401 = pi13 ? n20 : ~n19;
  assign n402 = pi12 ? n20 : ~n401;
  assign n403 = pi11 ? n20 : n402;
  assign n404 = pi10 ? n20 : n403;
  assign n405 = pi09 ? n20 : n404;
  assign n406 = pi08 ? n382 : n405;
  assign n407 = pi07 ? n398 : n406;
  assign n408 = pi12 ? n81 : ~n127;
  assign n409 = pi11 ? n19 : n408;
  assign n410 = pi10 ? n19 : n409;
  assign n411 = pi09 ? n410 : n20;
  assign n412 = pi08 ? n411 : n405;
  assign n413 = pi13 ? n368 : ~n19;
  assign n414 = pi12 ? n20 : ~n413;
  assign n415 = pi11 ? n20 : n414;
  assign n416 = pi10 ? n20 : n415;
  assign n417 = pi09 ? n20 : n416;
  assign n418 = pi08 ? n411 : n417;
  assign n419 = pi07 ? n412 : n418;
  assign n420 = pi06 ? n407 : n419;
  assign n421 = pi05 ? n400 : n420;
  assign n422 = pi13 ? n384 : ~n19;
  assign n423 = pi12 ? n20 : ~n422;
  assign n424 = pi11 ? n20 : n423;
  assign n425 = pi10 ? n20 : n424;
  assign n426 = pi09 ? n20 : n425;
  assign n427 = pi08 ? n411 : n426;
  assign n428 = pi07 ? n418 : n427;
  assign n429 = pi13 ? n20 : n338;
  assign n430 = pi12 ? n429 : ~n422;
  assign n431 = pi11 ? n20 : n430;
  assign n432 = pi10 ? n20 : n431;
  assign n433 = pi09 ? n20 : n432;
  assign n434 = pi08 ? n411 : n433;
  assign n435 = pi13 ? n392 : ~n19;
  assign n436 = pi12 ? n20 : ~n435;
  assign n437 = pi11 ? n20 : n436;
  assign n438 = pi10 ? n20 : n437;
  assign n439 = pi09 ? n20 : n438;
  assign n440 = pi08 ? n411 : n439;
  assign n441 = pi07 ? n434 : n440;
  assign n442 = pi06 ? n428 : n441;
  assign n443 = pi12 ? n20 : n19;
  assign n444 = pi11 ? n20 : n443;
  assign n445 = pi10 ? n20 : n444;
  assign n446 = pi09 ? n20 : n445;
  assign n447 = pi08 ? n411 : n446;
  assign n448 = pi07 ? n440 : n447;
  assign n449 = pi12 ? n81 : n20;
  assign n450 = pi11 ? n19 : n449;
  assign n451 = pi10 ? n19 : n450;
  assign n452 = pi09 ? n451 : n20;
  assign n453 = pi08 ? n452 : n446;
  assign n454 = pi06 ? n448 : n453;
  assign n455 = pi05 ? n442 : n454;
  assign n456 = pi04 ? n421 : n455;
  assign n457 = pi03 ? n378 : n456;
  assign n458 = pi12 ? n312 : n20;
  assign n459 = pi11 ? n19 : n458;
  assign n460 = pi10 ? n19 : n459;
  assign n461 = pi09 ? n460 : n20;
  assign n462 = pi08 ? n461 : n446;
  assign n463 = pi07 ? n453 : n462;
  assign n464 = pi06 ? n453 : n463;
  assign n465 = pi05 ? n464 : n462;
  assign n466 = pi15 ? n20 : n19;
  assign n467 = pi14 ? n20 : n466;
  assign n468 = pi13 ? n20 : n467;
  assign n469 = pi12 ? n468 : n19;
  assign n470 = pi11 ? n20 : n469;
  assign n471 = pi10 ? n20 : n470;
  assign n472 = pi09 ? n20 : n471;
  assign n473 = pi08 ? n461 : n472;
  assign n474 = pi06 ? n462 : n473;
  assign n475 = pi05 ? n462 : n474;
  assign n476 = pi04 ? n465 : n475;
  assign n477 = pi14 ? n20 : n19;
  assign n478 = pi13 ? n20 : n477;
  assign n479 = pi12 ? n478 : n19;
  assign n480 = pi11 ? n20 : n479;
  assign n481 = pi10 ? n20 : n480;
  assign n482 = pi09 ? n20 : n481;
  assign n483 = pi08 ? n461 : n482;
  assign n484 = pi14 ? n466 : n19;
  assign n485 = pi13 ? n20 : n484;
  assign n486 = pi12 ? n485 : n19;
  assign n487 = pi11 ? n20 : n486;
  assign n488 = pi10 ? n20 : n487;
  assign n489 = pi09 ? n20 : n488;
  assign n490 = pi08 ? n461 : n489;
  assign n491 = pi06 ? n483 : n490;
  assign n492 = pi13 ? n20 : n19;
  assign n493 = pi12 ? n492 : n19;
  assign n494 = pi11 ? n20 : n493;
  assign n495 = pi10 ? n20 : n494;
  assign n496 = pi09 ? n20 : n495;
  assign n497 = pi08 ? n461 : n496;
  assign n498 = pi13 ? n467 : n19;
  assign n499 = pi12 ? n498 : n19;
  assign n500 = pi11 ? n20 : n499;
  assign n501 = pi10 ? n20 : n500;
  assign n502 = pi09 ? n20 : n501;
  assign n503 = pi08 ? n461 : n502;
  assign n504 = pi06 ? n497 : n503;
  assign n505 = pi05 ? n491 : n504;
  assign n506 = pi13 ? n477 : n19;
  assign n507 = pi12 ? n506 : n19;
  assign n508 = pi11 ? n20 : n507;
  assign n509 = pi10 ? n20 : n508;
  assign n510 = pi09 ? n20 : n509;
  assign n511 = pi08 ? n461 : n510;
  assign n512 = pi13 ? n484 : n19;
  assign n513 = pi12 ? n512 : n19;
  assign n514 = pi11 ? n20 : n513;
  assign n515 = pi10 ? n20 : n514;
  assign n516 = pi09 ? n20 : n515;
  assign n517 = pi08 ? n461 : n516;
  assign n518 = pi06 ? n511 : n517;
  assign n519 = pi11 ? n20 : n19;
  assign n520 = pi10 ? n20 : n519;
  assign n521 = pi09 ? n20 : n520;
  assign n522 = pi08 ? n461 : n521;
  assign n523 = pi05 ? n518 : n522;
  assign n524 = pi04 ? n505 : n523;
  assign n525 = pi03 ? n476 : n524;
  assign n526 = pi02 ? n457 : n525;
  assign n527 = pi12 ? n20 : n468;
  assign n528 = pi11 ? n527 : n19;
  assign n529 = pi10 ? n20 : n528;
  assign n530 = pi09 ? n20 : n529;
  assign n531 = pi08 ? n461 : n530;
  assign n532 = pi07 ? n522 : n531;
  assign n533 = pi12 ? n20 : n478;
  assign n534 = pi11 ? n533 : n19;
  assign n535 = pi10 ? n20 : n534;
  assign n536 = pi09 ? n20 : n535;
  assign n537 = pi08 ? n461 : n536;
  assign n538 = pi07 ? n531 : n537;
  assign n539 = pi06 ? n532 : n538;
  assign n540 = pi05 ? n522 : n539;
  assign n541 = pi04 ? n522 : n540;
  assign n542 = pi12 ? n20 : n485;
  assign n543 = pi11 ? n542 : n19;
  assign n544 = pi10 ? n20 : n543;
  assign n545 = pi09 ? n20 : n544;
  assign n546 = pi08 ? n461 : n545;
  assign n547 = pi07 ? n537 : n546;
  assign n548 = pi12 ? n20 : n492;
  assign n549 = pi11 ? n548 : n19;
  assign n550 = pi10 ? n20 : n549;
  assign n551 = pi09 ? n20 : n550;
  assign n552 = pi08 ? n461 : n551;
  assign n553 = pi07 ? n546 : n552;
  assign n554 = pi06 ? n547 : n553;
  assign n555 = pi12 ? n20 : n498;
  assign n556 = pi11 ? n555 : n19;
  assign n557 = pi10 ? n20 : n556;
  assign n558 = pi09 ? n20 : n557;
  assign n559 = pi08 ? n461 : n558;
  assign n560 = pi07 ? n552 : n559;
  assign n561 = pi12 ? n20 : n506;
  assign n562 = pi11 ? n561 : n19;
  assign n563 = pi10 ? n20 : n562;
  assign n564 = pi09 ? n20 : n563;
  assign n565 = pi08 ? n461 : n564;
  assign n566 = pi07 ? n559 : n565;
  assign n567 = pi06 ? n560 : n566;
  assign n568 = pi05 ? n554 : n567;
  assign n569 = pi12 ? n20 : n512;
  assign n570 = pi11 ? n569 : n19;
  assign n571 = pi10 ? n20 : n570;
  assign n572 = pi09 ? n20 : n571;
  assign n573 = pi08 ? n461 : n572;
  assign n574 = pi07 ? n565 : n573;
  assign n575 = pi11 ? n443 : n19;
  assign n576 = pi10 ? n20 : n575;
  assign n577 = pi09 ? n20 : n576;
  assign n578 = pi08 ? n461 : n577;
  assign n579 = pi07 ? n573 : n578;
  assign n580 = pi06 ? n574 : n579;
  assign n581 = pi05 ? n580 : n578;
  assign n582 = pi04 ? n568 : n581;
  assign n583 = pi03 ? n541 : n582;
  assign n584 = pi11 ? n469 : n19;
  assign n585 = pi10 ? n20 : n584;
  assign n586 = pi09 ? n20 : n585;
  assign n587 = pi08 ? n461 : n586;
  assign n588 = pi11 ? n479 : n19;
  assign n589 = pi10 ? n20 : n588;
  assign n590 = pi09 ? n20 : n589;
  assign n591 = pi08 ? n461 : n590;
  assign n592 = pi06 ? n587 : n591;
  assign n593 = pi05 ? n578 : n592;
  assign n594 = pi04 ? n578 : n593;
  assign n595 = pi11 ? n486 : n19;
  assign n596 = pi10 ? n20 : n595;
  assign n597 = pi09 ? n20 : n596;
  assign n598 = pi08 ? n461 : n597;
  assign n599 = pi11 ? n493 : n19;
  assign n600 = pi10 ? n20 : n599;
  assign n601 = pi09 ? n20 : n600;
  assign n602 = pi08 ? n461 : n601;
  assign n603 = pi07 ? n598 : n602;
  assign n604 = pi06 ? n598 : n603;
  assign n605 = pi11 ? n499 : n19;
  assign n606 = pi10 ? n20 : n605;
  assign n607 = pi09 ? n20 : n606;
  assign n608 = pi08 ? n461 : n607;
  assign n609 = pi07 ? n602 : n608;
  assign n610 = pi11 ? n507 : n19;
  assign n611 = pi10 ? n20 : n610;
  assign n612 = pi09 ? n20 : n611;
  assign n613 = pi08 ? n461 : n612;
  assign n614 = pi07 ? n608 : n613;
  assign n615 = pi06 ? n609 : n614;
  assign n616 = pi05 ? n604 : n615;
  assign n617 = pi11 ? n513 : n19;
  assign n618 = pi10 ? n20 : n617;
  assign n619 = pi09 ? n20 : n618;
  assign n620 = pi08 ? n461 : n619;
  assign n621 = pi07 ? n613 : n620;
  assign n622 = pi10 ? n20 : n19;
  assign n623 = pi09 ? n20 : n622;
  assign n624 = pi08 ? n461 : n623;
  assign n625 = pi07 ? n620 : n624;
  assign n626 = pi06 ? n621 : n625;
  assign n627 = pi05 ? n626 : n624;
  assign n628 = pi04 ? n616 : n627;
  assign n629 = pi03 ? n594 : n628;
  assign n630 = pi02 ? n583 : n629;
  assign n631 = pi01 ? n526 : n630;
  assign n632 = pi00 ? n334 : n631;
  assign po0 = ~n632;
endmodule


